// Latch-mapped netlist written by map_latches.py, 2017-08-22 08:02:33
// Written ISPD/ICCAD/TAU contest Verilog format. 
//    Input file:  cordic_ispd/cordic_ispd_remapped.v
//    Latch cell:  ms00f80
//    Clock port:  clk
//    Output file: cordic_ispd/cordic_ispd_remapped.v

module cordic_ispd (
clk,
beta_0,
beta_1,
beta_10,
beta_11,
beta_12,
beta_13,
beta_14,
beta_15,
beta_16,
beta_17,
beta_18,
beta_19,
beta_2,
beta_20,
beta_21,
beta_22,
beta_23,
beta_24,
beta_25,
beta_26,
beta_27,
beta_28,
beta_29,
beta_3,
beta_30,
beta_31,
beta_4,
beta_5,
beta_6,
beta_7,
beta_8,
beta_9,
rst,
tau_clk,
cos_out_0,
cos_out_1,
cos_out_10,
cos_out_11,
cos_out_12,
cos_out_13,
cos_out_14,
cos_out_15,
cos_out_16,
cos_out_17,
cos_out_18,
cos_out_19,
cos_out_2,
cos_out_20,
cos_out_21,
cos_out_22,
cos_out_23,
cos_out_24,
cos_out_25,
cos_out_26,
cos_out_27,
cos_out_28,
cos_out_29,
cos_out_3,
cos_out_30,
cos_out_31,
cos_out_4,
cos_out_5,
cos_out_6,
cos_out_7,
cos_out_8,
cos_out_9,
sin_out_0,
sin_out_1,
sin_out_10,
sin_out_11,
sin_out_12,
sin_out_13,
sin_out_14,
sin_out_15,
sin_out_16,
sin_out_17,
sin_out_18,
sin_out_19,
sin_out_2,
sin_out_20,
sin_out_21,
sin_out_22,
sin_out_23,
sin_out_24,
sin_out_25,
sin_out_26,
sin_out_27,
sin_out_28,
sin_out_29,
sin_out_3,
sin_out_30,
sin_out_31,
sin_out_4,
sin_out_5,
sin_out_6,
sin_out_7,
sin_out_8,
sin_out_9
);

// Start PIs
input clk;
input beta_0;
input beta_1;
input beta_10;
input beta_11;
input beta_12;
input beta_13;
input beta_14;
input beta_15;
input beta_16;
input beta_17;
input beta_18;
input beta_19;
input beta_2;
input beta_20;
input beta_21;
input beta_22;
input beta_23;
input beta_24;
input beta_25;
input beta_26;
input beta_27;
input beta_28;
input beta_29;
input beta_3;
input beta_30;
input beta_31;
input beta_4;
input beta_5;
input beta_6;
input beta_7;
input beta_8;
input beta_9;
input rst;
input tau_clk;

// Start POs
output cos_out_0;
output cos_out_1;
output cos_out_10;
output cos_out_11;
output cos_out_12;
output cos_out_13;
output cos_out_14;
output cos_out_15;
output cos_out_16;
output cos_out_17;
output cos_out_18;
output cos_out_19;
output cos_out_2;
output cos_out_20;
output cos_out_21;
output cos_out_22;
output cos_out_23;
output cos_out_24;
output cos_out_25;
output cos_out_26;
output cos_out_27;
output cos_out_28;
output cos_out_29;
output cos_out_3;
output cos_out_30;
output cos_out_31;
output cos_out_4;
output cos_out_5;
output cos_out_6;
output cos_out_7;
output cos_out_8;
output cos_out_9;
output sin_out_0;
output sin_out_1;
output sin_out_10;
output sin_out_11;
output sin_out_12;
output sin_out_13;
output sin_out_14;
output sin_out_15;
output sin_out_16;
output sin_out_17;
output sin_out_18;
output sin_out_19;
output sin_out_2;
output sin_out_20;
output sin_out_21;
output sin_out_22;
output sin_out_23;
output sin_out_24;
output sin_out_25;
output sin_out_26;
output sin_out_27;
output sin_out_28;
output sin_out_29;
output sin_out_3;
output sin_out_30;
output sin_out_31;
output sin_out_4;
output sin_out_5;
output sin_out_6;
output sin_out_7;
output sin_out_8;
output sin_out_9;

// Start wires
wire clk;
wire beta_0;
wire beta_1;
wire beta_10;
wire beta_11;
wire beta_12;
wire beta_13;
wire beta_14;
wire beta_15;
wire beta_16;
wire beta_17;
wire beta_18;
wire beta_19;
wire beta_2;
wire beta_20;
wire beta_21;
wire beta_22;
wire beta_23;
wire beta_24;
wire beta_25;
wire beta_26;
wire beta_27;
wire beta_28;
wire beta_29;
wire beta_3;
wire beta_30;
wire beta_31;
wire beta_4;
wire beta_5;
wire beta_6;
wire beta_7;
wire beta_8;
wire beta_9;
wire rst;
wire tau_clk;
wire cos_out_0;
wire cos_out_1;
wire cos_out_10;
wire cos_out_11;
wire cos_out_12;
wire cos_out_13;
wire cos_out_14;
wire cos_out_15;
wire cos_out_16;
wire cos_out_17;
wire cos_out_18;
wire cos_out_19;
wire cos_out_2;
wire cos_out_20;
wire cos_out_21;
wire cos_out_22;
wire cos_out_23;
wire cos_out_24;
wire cos_out_25;
wire cos_out_26;
wire cos_out_27;
wire cos_out_28;
wire cos_out_29;
wire cos_out_3;
wire cos_out_30;
wire cos_out_31;
wire cos_out_4;
wire cos_out_5;
wire cos_out_6;
wire cos_out_7;
wire cos_out_8;
wire cos_out_9;
wire sin_out_0;
wire sin_out_1;
wire sin_out_10;
wire sin_out_11;
wire sin_out_12;
wire sin_out_13;
wire sin_out_14;
wire sin_out_15;
wire sin_out_16;
wire sin_out_17;
wire sin_out_18;
wire sin_out_19;
wire sin_out_2;
wire sin_out_20;
wire sin_out_21;
wire sin_out_22;
wire sin_out_23;
wire sin_out_24;
wire sin_out_25;
wire sin_out_26;
wire sin_out_27;
wire sin_out_28;
wire sin_out_29;
wire sin_out_3;
wire sin_out_30;
wire sin_out_31;
wire sin_out_4;
wire sin_out_5;
wire sin_out_6;
wire sin_out_7;
wire sin_out_8;
wire sin_out_9;
wire cordic_combinational_sub_ln23_0_unr12_z_0_;
wire cordic_combinational_sub_ln23_0_unr16_z_0_;
wire cordic_combinational_sub_ln23_0_unr20_z_0_;
wire delay_add_ln22_unr11_stage5_stallmux_q_0_;
wire delay_add_ln22_unr11_stage5_stallmux_q_10_;
wire delay_add_ln22_unr11_stage5_stallmux_q_11_;
wire delay_add_ln22_unr11_stage5_stallmux_q_12_;
wire delay_add_ln22_unr11_stage5_stallmux_q_13_;
wire delay_add_ln22_unr11_stage5_stallmux_q_14_;
wire delay_add_ln22_unr11_stage5_stallmux_q_15_;
wire delay_add_ln22_unr11_stage5_stallmux_q_16_;
wire delay_add_ln22_unr11_stage5_stallmux_q_17_;
wire delay_add_ln22_unr11_stage5_stallmux_q_18_;
wire delay_add_ln22_unr11_stage5_stallmux_q_19_;
wire delay_add_ln22_unr11_stage5_stallmux_q_1_;
wire delay_add_ln22_unr11_stage5_stallmux_q_20_;
wire delay_add_ln22_unr11_stage5_stallmux_q_21_;
wire delay_add_ln22_unr11_stage5_stallmux_q_22_;
wire delay_add_ln22_unr11_stage5_stallmux_q_23_;
wire delay_add_ln22_unr11_stage5_stallmux_q_24_;
wire delay_add_ln22_unr11_stage5_stallmux_q_25_;
wire delay_add_ln22_unr11_stage5_stallmux_q_26_;
wire delay_add_ln22_unr11_stage5_stallmux_q_27_;
wire delay_add_ln22_unr11_stage5_stallmux_q_28_;
wire delay_add_ln22_unr11_stage5_stallmux_q_29_;
wire delay_add_ln22_unr11_stage5_stallmux_q_2_;
wire delay_add_ln22_unr11_stage5_stallmux_q_30_;
wire delay_add_ln22_unr11_stage5_stallmux_q_31_;
wire delay_add_ln22_unr11_stage5_stallmux_q_3_;
wire delay_add_ln22_unr11_stage5_stallmux_q_4_;
wire delay_add_ln22_unr11_stage5_stallmux_q_5_;
wire delay_add_ln22_unr11_stage5_stallmux_q_6_;
wire delay_add_ln22_unr11_stage5_stallmux_q_7_;
wire delay_add_ln22_unr11_stage5_stallmux_q_8_;
wire delay_add_ln22_unr11_stage5_stallmux_q_9_;
wire delay_add_ln22_unr14_stage6_stallmux_q_0_;
wire delay_add_ln22_unr14_stage6_stallmux_q_10_;
wire delay_add_ln22_unr14_stage6_stallmux_q_11_;
wire delay_add_ln22_unr14_stage6_stallmux_q_12_;
wire delay_add_ln22_unr14_stage6_stallmux_q_13_;
wire delay_add_ln22_unr14_stage6_stallmux_q_14_;
wire delay_add_ln22_unr14_stage6_stallmux_q_15_;
wire delay_add_ln22_unr14_stage6_stallmux_q_16_;
wire delay_add_ln22_unr14_stage6_stallmux_q_17_;
wire delay_add_ln22_unr14_stage6_stallmux_q_18_;
wire delay_add_ln22_unr14_stage6_stallmux_q_19_;
wire delay_add_ln22_unr14_stage6_stallmux_q_1_;
wire delay_add_ln22_unr14_stage6_stallmux_q_20_;
wire delay_add_ln22_unr14_stage6_stallmux_q_21_;
wire delay_add_ln22_unr14_stage6_stallmux_q_22_;
wire delay_add_ln22_unr14_stage6_stallmux_q_23_;
wire delay_add_ln22_unr14_stage6_stallmux_q_24_;
wire delay_add_ln22_unr14_stage6_stallmux_q_25_;
wire delay_add_ln22_unr14_stage6_stallmux_q_26_;
wire delay_add_ln22_unr14_stage6_stallmux_q_27_;
wire delay_add_ln22_unr14_stage6_stallmux_q_28_;
wire delay_add_ln22_unr14_stage6_stallmux_q_29_;
wire delay_add_ln22_unr14_stage6_stallmux_q_2_;
wire delay_add_ln22_unr14_stage6_stallmux_q_30_;
wire delay_add_ln22_unr14_stage6_stallmux_q_31_;
wire delay_add_ln22_unr14_stage6_stallmux_q_3_;
wire delay_add_ln22_unr14_stage6_stallmux_q_4_;
wire delay_add_ln22_unr14_stage6_stallmux_q_5_;
wire delay_add_ln22_unr14_stage6_stallmux_q_6_;
wire delay_add_ln22_unr14_stage6_stallmux_q_7_;
wire delay_add_ln22_unr14_stage6_stallmux_q_8_;
wire delay_add_ln22_unr14_stage6_stallmux_q_9_;
wire delay_add_ln22_unr17_stage7_stallmux_q_0_;
wire delay_add_ln22_unr17_stage7_stallmux_q_10_;
wire delay_add_ln22_unr17_stage7_stallmux_q_11_;
wire delay_add_ln22_unr17_stage7_stallmux_q_12_;
wire delay_add_ln22_unr17_stage7_stallmux_q_13_;
wire delay_add_ln22_unr17_stage7_stallmux_q_14_;
wire delay_add_ln22_unr17_stage7_stallmux_q_15_;
wire delay_add_ln22_unr17_stage7_stallmux_q_16_;
wire delay_add_ln22_unr17_stage7_stallmux_q_17_;
wire delay_add_ln22_unr17_stage7_stallmux_q_18_;
wire delay_add_ln22_unr17_stage7_stallmux_q_19_;
wire delay_add_ln22_unr17_stage7_stallmux_q_1_;
wire delay_add_ln22_unr17_stage7_stallmux_q_20_;
wire delay_add_ln22_unr17_stage7_stallmux_q_21_;
wire delay_add_ln22_unr17_stage7_stallmux_q_22_;
wire delay_add_ln22_unr17_stage7_stallmux_q_23_;
wire delay_add_ln22_unr17_stage7_stallmux_q_24_;
wire delay_add_ln22_unr17_stage7_stallmux_q_25_;
wire delay_add_ln22_unr17_stage7_stallmux_q_26_;
wire delay_add_ln22_unr17_stage7_stallmux_q_27_;
wire delay_add_ln22_unr17_stage7_stallmux_q_28_;
wire delay_add_ln22_unr17_stage7_stallmux_q_29_;
wire delay_add_ln22_unr17_stage7_stallmux_q_2_;
wire delay_add_ln22_unr17_stage7_stallmux_q_30_;
wire delay_add_ln22_unr17_stage7_stallmux_q_31_;
wire delay_add_ln22_unr17_stage7_stallmux_q_3_;
wire delay_add_ln22_unr17_stage7_stallmux_q_4_;
wire delay_add_ln22_unr17_stage7_stallmux_q_5_;
wire delay_add_ln22_unr17_stage7_stallmux_q_6_;
wire delay_add_ln22_unr17_stage7_stallmux_q_7_;
wire delay_add_ln22_unr17_stage7_stallmux_q_8_;
wire delay_add_ln22_unr17_stage7_stallmux_q_9_;
wire delay_add_ln22_unr20_stage8_stallmux_q_0_;
wire delay_add_ln22_unr20_stage8_stallmux_q_10_;
wire delay_add_ln22_unr20_stage8_stallmux_q_11_;
wire delay_add_ln22_unr20_stage8_stallmux_q_12_;
wire delay_add_ln22_unr20_stage8_stallmux_q_13_;
wire delay_add_ln22_unr20_stage8_stallmux_q_14_;
wire delay_add_ln22_unr20_stage8_stallmux_q_15_;
wire delay_add_ln22_unr20_stage8_stallmux_q_16_;
wire delay_add_ln22_unr20_stage8_stallmux_q_17_;
wire delay_add_ln22_unr20_stage8_stallmux_q_18_;
wire delay_add_ln22_unr20_stage8_stallmux_q_19_;
wire delay_add_ln22_unr20_stage8_stallmux_q_1_;
wire delay_add_ln22_unr20_stage8_stallmux_q_20_;
wire delay_add_ln22_unr20_stage8_stallmux_q_21_;
wire delay_add_ln22_unr20_stage8_stallmux_q_22_;
wire delay_add_ln22_unr20_stage8_stallmux_q_23_;
wire delay_add_ln22_unr20_stage8_stallmux_q_24_;
wire delay_add_ln22_unr20_stage8_stallmux_q_25_;
wire delay_add_ln22_unr20_stage8_stallmux_q_26_;
wire delay_add_ln22_unr20_stage8_stallmux_q_27_;
wire delay_add_ln22_unr20_stage8_stallmux_q_28_;
wire delay_add_ln22_unr20_stage8_stallmux_q_29_;
wire delay_add_ln22_unr20_stage8_stallmux_q_2_;
wire delay_add_ln22_unr20_stage8_stallmux_q_30_;
wire delay_add_ln22_unr20_stage8_stallmux_q_31_;
wire delay_add_ln22_unr20_stage8_stallmux_q_3_;
wire delay_add_ln22_unr20_stage8_stallmux_q_4_;
wire delay_add_ln22_unr20_stage8_stallmux_q_5_;
wire delay_add_ln22_unr20_stage8_stallmux_q_6_;
wire delay_add_ln22_unr20_stage8_stallmux_q_7_;
wire delay_add_ln22_unr20_stage8_stallmux_q_8_;
wire delay_add_ln22_unr20_stage8_stallmux_q_9_;
wire delay_add_ln22_unr23_stage9_stallmux_q_0_;
wire delay_add_ln22_unr23_stage9_stallmux_q_10_;
wire delay_add_ln22_unr23_stage9_stallmux_q_11_;
wire delay_add_ln22_unr23_stage9_stallmux_q_12_;
wire delay_add_ln22_unr23_stage9_stallmux_q_13_;
wire delay_add_ln22_unr23_stage9_stallmux_q_14_;
wire delay_add_ln22_unr23_stage9_stallmux_q_15_;
wire delay_add_ln22_unr23_stage9_stallmux_q_16_;
wire delay_add_ln22_unr23_stage9_stallmux_q_17_;
wire delay_add_ln22_unr23_stage9_stallmux_q_18_;
wire delay_add_ln22_unr23_stage9_stallmux_q_19_;
wire delay_add_ln22_unr23_stage9_stallmux_q_1_;
wire delay_add_ln22_unr23_stage9_stallmux_q_20_;
wire delay_add_ln22_unr23_stage9_stallmux_q_21_;
wire delay_add_ln22_unr23_stage9_stallmux_q_22_;
wire delay_add_ln22_unr23_stage9_stallmux_q_23_;
wire delay_add_ln22_unr23_stage9_stallmux_q_24_;
wire delay_add_ln22_unr23_stage9_stallmux_q_25_;
wire delay_add_ln22_unr23_stage9_stallmux_q_26_;
wire delay_add_ln22_unr23_stage9_stallmux_q_27_;
wire delay_add_ln22_unr23_stage9_stallmux_q_28_;
wire delay_add_ln22_unr23_stage9_stallmux_q_29_;
wire delay_add_ln22_unr23_stage9_stallmux_q_2_;
wire delay_add_ln22_unr23_stage9_stallmux_q_30_;
wire delay_add_ln22_unr23_stage9_stallmux_q_31_;
wire delay_add_ln22_unr23_stage9_stallmux_q_3_;
wire delay_add_ln22_unr23_stage9_stallmux_q_4_;
wire delay_add_ln22_unr23_stage9_stallmux_q_5_;
wire delay_add_ln22_unr23_stage9_stallmux_q_6_;
wire delay_add_ln22_unr23_stage9_stallmux_q_7_;
wire delay_add_ln22_unr23_stage9_stallmux_q_8_;
wire delay_add_ln22_unr23_stage9_stallmux_q_9_;
wire delay_add_ln22_unr27_stage10_stallmux_q_0_;
wire delay_add_ln22_unr27_stage10_stallmux_q_10_;
wire delay_add_ln22_unr27_stage10_stallmux_q_11_;
wire delay_add_ln22_unr27_stage10_stallmux_q_12_;
wire delay_add_ln22_unr27_stage10_stallmux_q_13_;
wire delay_add_ln22_unr27_stage10_stallmux_q_14_;
wire delay_add_ln22_unr27_stage10_stallmux_q_15_;
wire delay_add_ln22_unr27_stage10_stallmux_q_16_;
wire delay_add_ln22_unr27_stage10_stallmux_q_17_;
wire delay_add_ln22_unr27_stage10_stallmux_q_18_;
wire delay_add_ln22_unr27_stage10_stallmux_q_19_;
wire delay_add_ln22_unr27_stage10_stallmux_q_1_;
wire delay_add_ln22_unr27_stage10_stallmux_q_20_;
wire delay_add_ln22_unr27_stage10_stallmux_q_21_;
wire delay_add_ln22_unr27_stage10_stallmux_q_22_;
wire delay_add_ln22_unr27_stage10_stallmux_q_23_;
wire delay_add_ln22_unr27_stage10_stallmux_q_24_;
wire delay_add_ln22_unr27_stage10_stallmux_q_25_;
wire delay_add_ln22_unr27_stage10_stallmux_q_26_;
wire delay_add_ln22_unr27_stage10_stallmux_q_27_;
wire delay_add_ln22_unr27_stage10_stallmux_q_28_;
wire delay_add_ln22_unr27_stage10_stallmux_q_29_;
wire delay_add_ln22_unr27_stage10_stallmux_q_2_;
wire delay_add_ln22_unr27_stage10_stallmux_q_30_;
wire delay_add_ln22_unr27_stage10_stallmux_q_31_;
wire delay_add_ln22_unr27_stage10_stallmux_q_3_;
wire delay_add_ln22_unr27_stage10_stallmux_q_4_;
wire delay_add_ln22_unr27_stage10_stallmux_q_5_;
wire delay_add_ln22_unr27_stage10_stallmux_q_6_;
wire delay_add_ln22_unr27_stage10_stallmux_q_7_;
wire delay_add_ln22_unr27_stage10_stallmux_q_8_;
wire delay_add_ln22_unr27_stage10_stallmux_q_9_;
wire delay_add_ln22_unr2_stage2_stallmux_q_10_;
wire delay_add_ln22_unr2_stage2_stallmux_q_11_;
wire delay_add_ln22_unr2_stage2_stallmux_q_12_;
wire delay_add_ln22_unr2_stage2_stallmux_q_13_;
wire delay_add_ln22_unr2_stage2_stallmux_q_14_;
wire delay_add_ln22_unr2_stage2_stallmux_q_15_;
wire delay_add_ln22_unr2_stage2_stallmux_q_16_;
wire delay_add_ln22_unr2_stage2_stallmux_q_17_;
wire delay_add_ln22_unr2_stage2_stallmux_q_18_;
wire delay_add_ln22_unr2_stage2_stallmux_q_19_;
wire delay_add_ln22_unr2_stage2_stallmux_q_1_;
wire delay_add_ln22_unr2_stage2_stallmux_q_20_;
wire delay_add_ln22_unr2_stage2_stallmux_q_21_;
wire delay_add_ln22_unr2_stage2_stallmux_q_22_;
wire delay_add_ln22_unr2_stage2_stallmux_q_23_;
wire delay_add_ln22_unr2_stage2_stallmux_q_24_;
wire delay_add_ln22_unr2_stage2_stallmux_q_25_;
wire delay_add_ln22_unr2_stage2_stallmux_q_26_;
wire delay_add_ln22_unr2_stage2_stallmux_q_27_;
wire delay_add_ln22_unr2_stage2_stallmux_q_28_;
wire delay_add_ln22_unr2_stage2_stallmux_q_29_;
wire delay_add_ln22_unr2_stage2_stallmux_q_2_;
wire delay_add_ln22_unr2_stage2_stallmux_q_30_;
wire delay_add_ln22_unr2_stage2_stallmux_q_31_;
wire delay_add_ln22_unr2_stage2_stallmux_q_3_;
wire delay_add_ln22_unr2_stage2_stallmux_q_4_;
wire delay_add_ln22_unr2_stage2_stallmux_q_5_;
wire delay_add_ln22_unr2_stage2_stallmux_q_6_;
wire delay_add_ln22_unr2_stage2_stallmux_q_7_;
wire delay_add_ln22_unr2_stage2_stallmux_q_8_;
wire delay_add_ln22_unr2_stage2_stallmux_q_9_;
wire delay_add_ln22_unr5_stage3_stallmux_q_0_;
wire delay_add_ln22_unr5_stage3_stallmux_q_10_;
wire delay_add_ln22_unr5_stage3_stallmux_q_11_;
wire delay_add_ln22_unr5_stage3_stallmux_q_12_;
wire delay_add_ln22_unr5_stage3_stallmux_q_13_;
wire delay_add_ln22_unr5_stage3_stallmux_q_14_;
wire delay_add_ln22_unr5_stage3_stallmux_q_15_;
wire delay_add_ln22_unr5_stage3_stallmux_q_16_;
wire delay_add_ln22_unr5_stage3_stallmux_q_17_;
wire delay_add_ln22_unr5_stage3_stallmux_q_18_;
wire delay_add_ln22_unr5_stage3_stallmux_q_19_;
wire delay_add_ln22_unr5_stage3_stallmux_q_1_;
wire delay_add_ln22_unr5_stage3_stallmux_q_20_;
wire delay_add_ln22_unr5_stage3_stallmux_q_21_;
wire delay_add_ln22_unr5_stage3_stallmux_q_22_;
wire delay_add_ln22_unr5_stage3_stallmux_q_23_;
wire delay_add_ln22_unr5_stage3_stallmux_q_24_;
wire delay_add_ln22_unr5_stage3_stallmux_q_25_;
wire delay_add_ln22_unr5_stage3_stallmux_q_26_;
wire delay_add_ln22_unr5_stage3_stallmux_q_27_;
wire delay_add_ln22_unr5_stage3_stallmux_q_28_;
wire delay_add_ln22_unr5_stage3_stallmux_q_29_;
wire delay_add_ln22_unr5_stage3_stallmux_q_2_;
wire delay_add_ln22_unr5_stage3_stallmux_q_30_;
wire delay_add_ln22_unr5_stage3_stallmux_q_31_;
wire delay_add_ln22_unr5_stage3_stallmux_q_3_;
wire delay_add_ln22_unr5_stage3_stallmux_q_4_;
wire delay_add_ln22_unr5_stage3_stallmux_q_5_;
wire delay_add_ln22_unr5_stage3_stallmux_q_6_;
wire delay_add_ln22_unr5_stage3_stallmux_q_7_;
wire delay_add_ln22_unr5_stage3_stallmux_q_8_;
wire delay_add_ln22_unr5_stage3_stallmux_q_9_;
wire delay_add_ln22_unr8_stage4_stallmux_q_0_;
wire delay_add_ln22_unr8_stage4_stallmux_q_10_;
wire delay_add_ln22_unr8_stage4_stallmux_q_11_;
wire delay_add_ln22_unr8_stage4_stallmux_q_12_;
wire delay_add_ln22_unr8_stage4_stallmux_q_13_;
wire delay_add_ln22_unr8_stage4_stallmux_q_14_;
wire delay_add_ln22_unr8_stage4_stallmux_q_15_;
wire delay_add_ln22_unr8_stage4_stallmux_q_16_;
wire delay_add_ln22_unr8_stage4_stallmux_q_17_;
wire delay_add_ln22_unr8_stage4_stallmux_q_18_;
wire delay_add_ln22_unr8_stage4_stallmux_q_19_;
wire delay_add_ln22_unr8_stage4_stallmux_q_1_;
wire delay_add_ln22_unr8_stage4_stallmux_q_20_;
wire delay_add_ln22_unr8_stage4_stallmux_q_21_;
wire delay_add_ln22_unr8_stage4_stallmux_q_22_;
wire delay_add_ln22_unr8_stage4_stallmux_q_23_;
wire delay_add_ln22_unr8_stage4_stallmux_q_24_;
wire delay_add_ln22_unr8_stage4_stallmux_q_25_;
wire delay_add_ln22_unr8_stage4_stallmux_q_26_;
wire delay_add_ln22_unr8_stage4_stallmux_q_27_;
wire delay_add_ln22_unr8_stage4_stallmux_q_28_;
wire delay_add_ln22_unr8_stage4_stallmux_q_29_;
wire delay_add_ln22_unr8_stage4_stallmux_q_2_;
wire delay_add_ln22_unr8_stage4_stallmux_q_30_;
wire delay_add_ln22_unr8_stage4_stallmux_q_31_;
wire delay_add_ln22_unr8_stage4_stallmux_q_3_;
wire delay_add_ln22_unr8_stage4_stallmux_q_4_;
wire delay_add_ln22_unr8_stage4_stallmux_q_5_;
wire delay_add_ln22_unr8_stage4_stallmux_q_6_;
wire delay_add_ln22_unr8_stage4_stallmux_q_7_;
wire delay_add_ln22_unr8_stage4_stallmux_q_8_;
wire delay_add_ln22_unr8_stage4_stallmux_q_9_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_0_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_10_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_11_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_12_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_13_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_14_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_15_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_16_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_17_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_18_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_19_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_1_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_20_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_21_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_22_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_23_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_24_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_25_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_26_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_27_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_28_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_29_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_2_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_30_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_31_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_3_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_4_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_5_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_6_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_7_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_8_;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_9_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_0_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_10_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_11_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_12_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_13_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_14_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_15_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_16_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_17_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_18_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_19_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_1_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_20_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_21_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_22_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_23_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_24_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_25_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_26_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_27_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_28_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_29_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_2_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_30_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_31_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_3_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_4_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_5_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_6_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_7_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_8_;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_9_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_0_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_10_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_11_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_12_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_13_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_14_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_15_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_16_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_17_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_18_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_19_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_1_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_20_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_21_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_22_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_23_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_24_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_25_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_26_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_27_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_28_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_29_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_2_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_30_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_31_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_3_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_4_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_5_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_6_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_7_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_8_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_9_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_0_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_10_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_11_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_12_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_13_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_14_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_15_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_16_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_17_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_18_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_19_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_1_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_20_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_21_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_22_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_23_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_24_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_25_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_26_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_27_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_28_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_29_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_2_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_30_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_31_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_3_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_4_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_5_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_6_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_7_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_8_;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_9_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_0_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_10_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_11_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_12_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_13_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_14_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_15_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_16_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_17_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_18_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_19_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_1_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_20_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_21_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_22_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_23_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_24_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_25_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_26_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_27_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_28_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_29_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_2_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_30_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_31_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_3_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_4_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_5_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_6_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_7_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_8_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_9_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_0_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_10_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_11_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_12_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_13_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_14_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_15_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_16_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_17_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_18_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_19_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_1_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_20_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_21_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_22_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_23_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_24_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_25_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_26_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_27_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_28_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_29_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_2_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_30_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_31_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_3_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_4_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_5_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_6_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_7_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_8_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_9_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_0_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_10_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_12_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_13_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_15_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_16_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_17_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_18_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_19_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_1_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_20_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_21_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_22_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_23_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_24_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_25_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_26_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_27_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_28_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_29_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_2_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_3_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_4_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_5_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_6_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_7_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_8_;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_9_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_0_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_10_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_11_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_12_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_13_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_14_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_15_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_16_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_17_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_18_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_19_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_1_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_20_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_21_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_22_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_23_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_24_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_25_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_26_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_27_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_28_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_29_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_2_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_30_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_31_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_3_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_4_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_5_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_6_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_7_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_8_;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_9_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_0_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_10_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_11_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_12_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_13_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_14_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_15_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_16_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_17_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_18_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_19_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_1_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_20_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_21_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_22_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_23_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_24_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_25_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_26_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_27_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_28_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_29_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_2_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_30_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_31_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_3_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_4_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_5_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_6_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_7_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_8_;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_9_;
wire delay_sub_ln21_unr24_stage9_stallmux_q_1_;
wire delay_sub_ln21_unr24_stage9_stallmux_q_2_;
wire delay_sub_ln21_unr24_stage9_stallmux_q_3_;
wire delay_sub_ln21_unr24_stage9_stallmux_q_4_;
wire delay_sub_ln21_unr24_stage9_stallmux_q_5_;
wire delay_sub_ln21_unr24_stage9_stallmux_q_6_;
wire delay_sub_ln21_unr24_stage9_stallmux_q_7_;
wire delay_sub_ln21_unr24_stage9_stallmux_q_8_;
wire delay_sub_ln22_unr24_stage9_stallmux_q_0_;
wire delay_sub_ln22_unr24_stage9_stallmux_q_1_;
wire delay_sub_ln22_unr24_stage9_stallmux_q_2_;
wire delay_sub_ln22_unr24_stage9_stallmux_q_3_;
wire delay_sub_ln22_unr24_stage9_stallmux_q_4_;
wire delay_sub_ln22_unr24_stage9_stallmux_q_5_;
wire delay_sub_ln22_unr24_stage9_stallmux_q_6_;
wire delay_sub_ln22_unr24_stage9_stallmux_q_7_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_10_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_11_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_12_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_13_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_14_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_15_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_16_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_17_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_18_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_19_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_1_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_20_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_21_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_22_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_23_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_24_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_25_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_26_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_27_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_28_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_29_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_2_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_30_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_3_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_4_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_5_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_6_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_7_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_8_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_9_;
wire delay_sub_ln23_0_unr15_stage6_stallmux_q;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_10_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_11_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_12_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_13_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_14_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_15_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_16_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_17_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_18_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_19_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_1_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_20_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_21_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_22_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_23_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_24_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_25_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_26_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_27_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_28_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_29_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_2_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_30_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_3_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_4_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_5_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_6_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_7_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_8_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_9_;
wire delay_sub_ln23_0_unr1_stage2_stallmux_q_0_;
wire delay_sub_ln23_0_unr1_stage2_stallmux_q_1_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_10_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_11_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_12_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_13_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_14_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_15_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_16_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_17_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_18_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_19_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_1_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_20_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_21_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_22_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_23_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_24_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_25_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_26_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_27_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_28_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_29_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_2_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_30_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_3_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_4_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_5_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_6_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_7_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_8_;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_9_;
wire delay_sub_ln23_0_unr21_stage8_stallmux_q;
wire delay_sub_ln23_0_unr22_stage8_stallmux_q;
wire delay_sub_ln23_0_unr23_stage8_stallmux_q;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_0_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_10_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_11_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_12_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_13_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_14_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_15_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_16_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_17_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_18_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_19_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_1_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_20_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_21_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_22_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_23_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_24_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_25_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_26_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_27_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_28_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_29_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_2_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_30_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_3_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_4_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_5_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_6_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_7_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_8_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_9_;
wire delay_sub_ln23_0_unr24_stage9_stallmux_q;
wire delay_sub_ln23_0_unr25_stage9_stallmux_q;
wire delay_sub_ln23_0_unr26_stage9_stallmux_q_0_;
wire delay_sub_ln23_0_unr26_stage9_stallmux_q_1_;
wire delay_sub_ln23_0_unr26_stage9_stallmux_q_2_;
wire delay_sub_ln23_0_unr27_stage10_stallmux_z;
wire delay_sub_ln23_0_unr28_stage10_stallmux_q;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_0_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_10_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_11_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_12_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_13_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_14_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_15_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_16_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_17_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_18_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_19_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_1_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_20_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_21_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_22_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_23_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_24_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_25_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_26_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_27_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_28_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_2_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_3_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_4_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_5_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_6_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_7_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_8_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_9_;
wire delay_sub_ln23_0_unr29_stage10_stallmux_q;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_0_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_10_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_11_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_12_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_13_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_14_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_15_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_16_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_17_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_18_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_19_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_1_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_20_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_21_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_22_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_23_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_24_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_25_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_26_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_27_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_28_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_29_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_2_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_3_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_4_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_5_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_6_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_7_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_8_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_9_;
wire delay_sub_ln23_0_unr30_stage10_stallmux_q;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_0_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_10_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_11_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_12_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_13_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_14_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_15_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_16_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_17_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_18_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_19_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_1_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_20_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_21_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_22_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_23_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_24_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_25_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_26_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_27_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_28_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_29_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_2_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_30_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_31_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_3_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_4_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_5_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_6_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_7_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_8_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_9_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_0_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_10_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_11_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_12_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_13_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_14_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_15_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_16_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_17_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_18_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_19_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_1_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_20_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_21_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_22_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_23_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_24_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_25_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_26_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_27_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_28_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_29_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_2_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_3_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_4_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_5_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_6_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_7_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_8_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_9_;
wire delay_sub_ln23_unr13_stage5_stallmux_q_1_;
wire delay_sub_ln23_unr17_stage6_stallmux_q_1_;
wire delay_sub_ln23_unr21_stage7_stallmux_q_1_;
wire delay_sub_ln23_unr25_stage8_stallmux_q_1_;
wire delay_sub_ln23_unr25_stage8_stallmux_q_3_;
wire delay_sub_ln23_unr29_stage9_stallmux_q_2_;
wire delay_sub_ln23_unr9_stage4_stallmux_q_3_;
wire delay_xor_ln21_unr12_stage5_stallmux_q_10_;
wire delay_xor_ln21_unr12_stage5_stallmux_q_11_;
wire delay_xor_ln21_unr12_stage5_stallmux_q_12_;
wire delay_xor_ln21_unr12_stage5_stallmux_q_13_;
wire delay_xor_ln21_unr12_stage5_stallmux_q_14_;
wire delay_xor_ln21_unr12_stage5_stallmux_q_15_;
wire delay_xor_ln21_unr12_stage5_stallmux_q_16_;
wire delay_xor_ln21_unr12_stage5_stallmux_q_17_;
wire delay_xor_ln21_unr12_stage5_stallmux_q_18_;
wire delay_xor_ln21_unr12_stage5_stallmux_q_19_;
wire delay_xor_ln21_unr12_stage5_stallmux_q_2_;
wire delay_xor_ln21_unr12_stage5_stallmux_q_3_;
wire delay_xor_ln21_unr12_stage5_stallmux_q_4_;
wire delay_xor_ln21_unr12_stage5_stallmux_q_5_;
wire delay_xor_ln21_unr12_stage5_stallmux_q_6_;
wire delay_xor_ln21_unr12_stage5_stallmux_q_7_;
wire delay_xor_ln21_unr12_stage5_stallmux_q_8_;
wire delay_xor_ln21_unr12_stage5_stallmux_q_9_;
wire delay_xor_ln21_unr15_stage6_stallmux_q_0_;
wire delay_xor_ln21_unr15_stage6_stallmux_q_10_;
wire delay_xor_ln21_unr15_stage6_stallmux_q_11_;
wire delay_xor_ln21_unr15_stage6_stallmux_q_12_;
wire delay_xor_ln21_unr15_stage6_stallmux_q_13_;
wire delay_xor_ln21_unr15_stage6_stallmux_q_14_;
wire delay_xor_ln21_unr15_stage6_stallmux_q_15_;
wire delay_xor_ln21_unr15_stage6_stallmux_q_16_;
wire delay_xor_ln21_unr15_stage6_stallmux_q_1_;
wire delay_xor_ln21_unr15_stage6_stallmux_q_2_;
wire delay_xor_ln21_unr15_stage6_stallmux_q_3_;
wire delay_xor_ln21_unr15_stage6_stallmux_q_4_;
wire delay_xor_ln21_unr15_stage6_stallmux_q_5_;
wire delay_xor_ln21_unr15_stage6_stallmux_q_6_;
wire delay_xor_ln21_unr15_stage6_stallmux_q_7_;
wire delay_xor_ln21_unr15_stage6_stallmux_q_8_;
wire delay_xor_ln21_unr15_stage6_stallmux_q_9_;
wire delay_xor_ln21_unr18_stage7_stallmux_q_10_;
wire delay_xor_ln21_unr18_stage7_stallmux_q_11_;
wire delay_xor_ln21_unr18_stage7_stallmux_q_12_;
wire delay_xor_ln21_unr18_stage7_stallmux_q_13_;
wire delay_xor_ln21_unr18_stage7_stallmux_q_2_;
wire delay_xor_ln21_unr18_stage7_stallmux_q_3_;
wire delay_xor_ln21_unr18_stage7_stallmux_q_5_;
wire delay_xor_ln21_unr18_stage7_stallmux_q_6_;
wire delay_xor_ln21_unr18_stage7_stallmux_q_7_;
wire delay_xor_ln21_unr18_stage7_stallmux_q_8_;
wire delay_xor_ln21_unr18_stage7_stallmux_q_9_;
wire delay_xor_ln21_unr21_stage8_stallmux_q_0_;
wire delay_xor_ln21_unr21_stage8_stallmux_q_10_;
wire delay_xor_ln21_unr21_stage8_stallmux_q_1_;
wire delay_xor_ln21_unr21_stage8_stallmux_q_2_;
wire delay_xor_ln21_unr21_stage8_stallmux_q_3_;
wire delay_xor_ln21_unr21_stage8_stallmux_q_4_;
wire delay_xor_ln21_unr21_stage8_stallmux_q_5_;
wire delay_xor_ln21_unr21_stage8_stallmux_q_6_;
wire delay_xor_ln21_unr21_stage8_stallmux_q_7_;
wire delay_xor_ln21_unr21_stage8_stallmux_q_8_;
wire delay_xor_ln21_unr21_stage8_stallmux_q_9_;
wire delay_xor_ln21_unr28_stage10_stallmux_q_0_;
wire delay_xor_ln21_unr28_stage10_stallmux_q_1_;
wire delay_xor_ln21_unr28_stage10_stallmux_q_2_;
wire delay_xor_ln21_unr28_stage10_stallmux_q_3_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_0_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_10_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_11_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_12_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_13_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_14_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_15_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_16_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_17_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_18_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_19_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_1_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_20_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_21_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_22_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_23_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_24_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_25_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_26_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_27_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_28_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_2_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_3_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_4_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_5_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_6_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_7_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_8_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_9_;
wire delay_xor_ln21_unr6_stage3_stallmux_q_0_;
wire delay_xor_ln21_unr6_stage3_stallmux_q_10_;
wire delay_xor_ln21_unr6_stage3_stallmux_q_11_;
wire delay_xor_ln21_unr6_stage3_stallmux_q_12_;
wire delay_xor_ln21_unr6_stage3_stallmux_q_13_;
wire delay_xor_ln21_unr6_stage3_stallmux_q_14_;
wire delay_xor_ln21_unr6_stage3_stallmux_q_15_;
wire delay_xor_ln21_unr6_stage3_stallmux_q_16_;
wire delay_xor_ln21_unr6_stage3_stallmux_q_17_;
wire delay_xor_ln21_unr6_stage3_stallmux_q_18_;
wire delay_xor_ln21_unr6_stage3_stallmux_q_19_;
wire delay_xor_ln21_unr6_stage3_stallmux_q_1_;
wire delay_xor_ln21_unr6_stage3_stallmux_q_20_;
wire delay_xor_ln21_unr6_stage3_stallmux_q_21_;
wire delay_xor_ln21_unr6_stage3_stallmux_q_22_;
wire delay_xor_ln21_unr6_stage3_stallmux_q_23_;
wire delay_xor_ln21_unr6_stage3_stallmux_q_24_;
wire delay_xor_ln21_unr6_stage3_stallmux_q_25_;
wire delay_xor_ln21_unr6_stage3_stallmux_q_2_;
wire delay_xor_ln21_unr6_stage3_stallmux_q_3_;
wire delay_xor_ln21_unr6_stage3_stallmux_q_4_;
wire delay_xor_ln21_unr6_stage3_stallmux_q_5_;
wire delay_xor_ln21_unr6_stage3_stallmux_q_6_;
wire delay_xor_ln21_unr6_stage3_stallmux_q_7_;
wire delay_xor_ln21_unr6_stage3_stallmux_q_8_;
wire delay_xor_ln21_unr6_stage3_stallmux_q_9_;
wire delay_xor_ln21_unr9_stage4_stallmux_q_0_;
wire delay_xor_ln21_unr9_stage4_stallmux_q_10_;
wire delay_xor_ln21_unr9_stage4_stallmux_q_11_;
wire delay_xor_ln21_unr9_stage4_stallmux_q_12_;
wire delay_xor_ln21_unr9_stage4_stallmux_q_13_;
wire delay_xor_ln21_unr9_stage4_stallmux_q_14_;
wire delay_xor_ln21_unr9_stage4_stallmux_q_15_;
wire delay_xor_ln21_unr9_stage4_stallmux_q_16_;
wire delay_xor_ln21_unr9_stage4_stallmux_q_17_;
wire delay_xor_ln21_unr9_stage4_stallmux_q_18_;
wire delay_xor_ln21_unr9_stage4_stallmux_q_19_;
wire delay_xor_ln21_unr9_stage4_stallmux_q_1_;
wire delay_xor_ln21_unr9_stage4_stallmux_q_20_;
wire delay_xor_ln21_unr9_stage4_stallmux_q_21_;
wire delay_xor_ln21_unr9_stage4_stallmux_q_22_;
wire delay_xor_ln21_unr9_stage4_stallmux_q_2_;
wire delay_xor_ln21_unr9_stage4_stallmux_q_3_;
wire delay_xor_ln21_unr9_stage4_stallmux_q_4_;
wire delay_xor_ln21_unr9_stage4_stallmux_q_5_;
wire delay_xor_ln21_unr9_stage4_stallmux_q_6_;
wire delay_xor_ln21_unr9_stage4_stallmux_q_7_;
wire delay_xor_ln21_unr9_stage4_stallmux_q_8_;
wire delay_xor_ln21_unr9_stage4_stallmux_q_9_;
wire delay_xor_ln22_unr12_stage5_stallmux_q_0_;
wire delay_xor_ln22_unr12_stage5_stallmux_q_10_;
wire delay_xor_ln22_unr12_stage5_stallmux_q_11_;
wire delay_xor_ln22_unr12_stage5_stallmux_q_12_;
wire delay_xor_ln22_unr12_stage5_stallmux_q_13_;
wire delay_xor_ln22_unr12_stage5_stallmux_q_14_;
wire delay_xor_ln22_unr12_stage5_stallmux_q_15_;
wire delay_xor_ln22_unr12_stage5_stallmux_q_16_;
wire delay_xor_ln22_unr12_stage5_stallmux_q_17_;
wire delay_xor_ln22_unr12_stage5_stallmux_q_18_;
wire delay_xor_ln22_unr12_stage5_stallmux_q_19_;
wire delay_xor_ln22_unr12_stage5_stallmux_q_1_;
wire delay_xor_ln22_unr12_stage5_stallmux_q_2_;
wire delay_xor_ln22_unr12_stage5_stallmux_q_3_;
wire delay_xor_ln22_unr12_stage5_stallmux_q_4_;
wire delay_xor_ln22_unr12_stage5_stallmux_q_5_;
wire delay_xor_ln22_unr12_stage5_stallmux_q_6_;
wire delay_xor_ln22_unr12_stage5_stallmux_q_7_;
wire delay_xor_ln22_unr12_stage5_stallmux_q_8_;
wire delay_xor_ln22_unr12_stage5_stallmux_q_9_;
wire delay_xor_ln22_unr15_stage6_stallmux_q_0_;
wire delay_xor_ln22_unr15_stage6_stallmux_q_10_;
wire delay_xor_ln22_unr15_stage6_stallmux_q_11_;
wire delay_xor_ln22_unr15_stage6_stallmux_q_12_;
wire delay_xor_ln22_unr15_stage6_stallmux_q_13_;
wire delay_xor_ln22_unr15_stage6_stallmux_q_14_;
wire delay_xor_ln22_unr15_stage6_stallmux_q_15_;
wire delay_xor_ln22_unr15_stage6_stallmux_q_16_;
wire delay_xor_ln22_unr15_stage6_stallmux_q_2_;
wire delay_xor_ln22_unr15_stage6_stallmux_q_3_;
wire delay_xor_ln22_unr15_stage6_stallmux_q_4_;
wire delay_xor_ln22_unr15_stage6_stallmux_q_5_;
wire delay_xor_ln22_unr15_stage6_stallmux_q_6_;
wire delay_xor_ln22_unr15_stage6_stallmux_q_7_;
wire delay_xor_ln22_unr15_stage6_stallmux_q_8_;
wire delay_xor_ln22_unr15_stage6_stallmux_q_9_;
wire delay_xor_ln22_unr18_stage7_stallmux_q_0_;
wire delay_xor_ln22_unr18_stage7_stallmux_q_10_;
wire delay_xor_ln22_unr18_stage7_stallmux_q_11_;
wire delay_xor_ln22_unr18_stage7_stallmux_q_12_;
wire delay_xor_ln22_unr18_stage7_stallmux_q_13_;
wire delay_xor_ln22_unr18_stage7_stallmux_q_1_;
wire delay_xor_ln22_unr18_stage7_stallmux_q_2_;
wire delay_xor_ln22_unr18_stage7_stallmux_q_3_;
wire delay_xor_ln22_unr18_stage7_stallmux_q_4_;
wire delay_xor_ln22_unr18_stage7_stallmux_q_5_;
wire delay_xor_ln22_unr18_stage7_stallmux_q_6_;
wire delay_xor_ln22_unr18_stage7_stallmux_q_7_;
wire delay_xor_ln22_unr18_stage7_stallmux_q_8_;
wire delay_xor_ln22_unr18_stage7_stallmux_q_9_;
wire delay_xor_ln22_unr21_stage8_stallmux_q_0_;
wire delay_xor_ln22_unr21_stage8_stallmux_q_10_;
wire delay_xor_ln22_unr21_stage8_stallmux_q_1_;
wire delay_xor_ln22_unr21_stage8_stallmux_q_2_;
wire delay_xor_ln22_unr21_stage8_stallmux_q_3_;
wire delay_xor_ln22_unr21_stage8_stallmux_q_4_;
wire delay_xor_ln22_unr21_stage8_stallmux_q_5_;
wire delay_xor_ln22_unr21_stage8_stallmux_q_6_;
wire delay_xor_ln22_unr21_stage8_stallmux_q_7_;
wire delay_xor_ln22_unr21_stage8_stallmux_q_8_;
wire delay_xor_ln22_unr21_stage8_stallmux_q_9_;
wire delay_xor_ln22_unr28_stage10_stallmux_q_0_;
wire delay_xor_ln22_unr28_stage10_stallmux_q_1_;
wire delay_xor_ln22_unr28_stage10_stallmux_q_2_;
wire delay_xor_ln22_unr28_stage10_stallmux_q_3_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_0_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_10_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_11_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_12_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_13_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_14_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_15_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_16_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_17_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_18_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_19_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_1_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_20_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_21_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_22_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_23_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_24_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_25_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_26_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_27_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_28_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_2_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_3_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_4_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_5_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_6_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_7_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_8_;
wire delay_xor_ln22_unr3_stage2_stallmux_q_9_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_0_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_10_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_11_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_12_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_13_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_14_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_15_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_16_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_17_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_18_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_19_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_1_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_20_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_21_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_22_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_23_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_24_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_25_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_2_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_3_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_4_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_5_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_6_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_7_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_8_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_9_;
wire delay_xor_ln22_unr9_stage4_stallmux_q_10_;
wire delay_xor_ln22_unr9_stage4_stallmux_q_11_;
wire delay_xor_ln22_unr9_stage4_stallmux_q_12_;
wire delay_xor_ln22_unr9_stage4_stallmux_q_13_;
wire delay_xor_ln22_unr9_stage4_stallmux_q_14_;
wire delay_xor_ln22_unr9_stage4_stallmux_q_15_;
wire delay_xor_ln22_unr9_stage4_stallmux_q_16_;
wire delay_xor_ln22_unr9_stage4_stallmux_q_17_;
wire delay_xor_ln22_unr9_stage4_stallmux_q_18_;
wire delay_xor_ln22_unr9_stage4_stallmux_q_19_;
wire delay_xor_ln22_unr9_stage4_stallmux_q_20_;
wire delay_xor_ln22_unr9_stage4_stallmux_q_21_;
wire delay_xor_ln22_unr9_stage4_stallmux_q_22_;
wire delay_xor_ln22_unr9_stage4_stallmux_q_2_;
wire delay_xor_ln22_unr9_stage4_stallmux_q_3_;
wire delay_xor_ln22_unr9_stage4_stallmux_q_4_;
wire delay_xor_ln22_unr9_stage4_stallmux_q_5_;
wire delay_xor_ln22_unr9_stage4_stallmux_q_6_;
wire delay_xor_ln22_unr9_stage4_stallmux_q_7_;
wire delay_xor_ln22_unr9_stage4_stallmux_q_8_;
wire delay_xor_ln22_unr9_stage4_stallmux_q_9_;
wire delay_xor_ln23_unr3_stage2_stallmux_q;
wire delay_xor_ln23_unr6_stage3_stallmux_q;
wire mux_while_ln12_psv_q_1_;
wire mux_while_ln12_psv_q_2_;
wire mux_while_ln12_psv_q_3_;
wire mux_while_ln12_psv_q_4_;
wire mux_while_ln12_psv_q_5_;
wire mux_while_ln12_psv_q_6_;
wire mux_while_ln12_psv_q_7_;
wire mux_while_ln12_psv_q_8_;
wire n10000;
wire n10001;
wire n10002;
wire n10003;
wire n10004;
wire n10005;
wire n10006;
wire n10007;
wire n10008;
wire n10009;
wire n1001;
wire n10010;
wire n10011;
wire n10012;
wire n10013;
wire n10014;
wire n10015;
wire n10016;
wire n10017;
wire n10018;
wire n10019;
wire n10020;
wire n10021;
wire n10022;
wire n10023;
wire n10024;
wire n10025;
wire n10026;
wire n10027;
wire n10028;
wire n10030;
wire n10031;
wire n10032;
wire n10033;
wire n10034;
wire n10035;
wire n10036;
wire n10037;
wire n10038;
wire n10039;
wire n10040;
wire n10041;
wire n10042;
wire n10043;
wire n10044;
wire n10045;
wire n10046;
wire n10047;
wire n10048;
wire n10049;
wire n10050;
wire n10051;
wire n10052;
wire n10053;
wire n10054;
wire n10055;
wire n10056;
wire n10057;
wire n10058;
wire n10059;
wire n1006;
wire n10060;
wire n10061;
wire n10062;
wire n10063;
wire n10064;
wire n10065;
wire n10066;
wire n10067;
wire n10068;
wire n10069;
wire n10070;
wire n10071;
wire n10072;
wire n10073;
wire n10074;
wire n10075;
wire n10076;
wire n10077;
wire n10078;
wire n10079;
wire n10080;
wire n10081;
wire n10082;
wire n10083;
wire n10084;
wire n10085;
wire n10086;
wire n10087;
wire n10088;
wire n10089;
wire n10090;
wire n10091;
wire n10092;
wire n10093;
wire n10094;
wire n10095;
wire n10096;
wire n10097;
wire n10098;
wire n10099;
wire n10100;
wire n10101;
wire n10102;
wire n10103;
wire n10104;
wire n10105;
wire n10106;
wire n10107;
wire n10108;
wire n10109;
wire n1011;
wire n10110;
wire n10111;
wire n10112;
wire n10113;
wire n10114;
wire n10115;
wire n10116;
wire n10117;
wire n10118;
wire n10119;
wire n10120;
wire n10121;
wire n10122;
wire n10123;
wire n10124;
wire n10125;
wire n10126;
wire n10127;
wire n10128;
wire n10129;
wire n10130;
wire n10131;
wire n10132;
wire n10133;
wire n10134;
wire n10135;
wire n10136;
wire n10137;
wire n10138;
wire n10139;
wire n10140;
wire n10141;
wire n10142;
wire n10143;
wire n10144;
wire n10145;
wire n10146;
wire n10147;
wire n10148;
wire n10149;
wire n10150;
wire n10151;
wire n10152;
wire n10153;
wire n10154;
wire n10155;
wire n10156;
wire n10157;
wire n10158;
wire n10159;
wire n1016;
wire n10160;
wire n10161;
wire n10162;
wire n10163;
wire n10164;
wire n10165;
wire n10166;
wire n10167;
wire n10168;
wire n10169;
wire n10170;
wire n10171;
wire n10172;
wire n10173;
wire n10174;
wire n10175;
wire n10176;
wire n10177;
wire n10178;
wire n10179;
wire n10180;
wire n10181;
wire n10182;
wire n10183;
wire n10184;
wire n10185;
wire n10186;
wire n10187;
wire n10188;
wire n10189;
wire n10190;
wire n10191;
wire n10192;
wire n10193;
wire n10194;
wire n10195;
wire n10196;
wire n10197;
wire n10198;
wire n10199;
wire n10200;
wire n10201;
wire n10202;
wire n10203;
wire n10204;
wire n10205;
wire n10206;
wire n10207;
wire n10208;
wire n10209;
wire n1021;
wire n10210;
wire n10211;
wire n10212;
wire n10213;
wire n10214;
wire n10215;
wire n10216;
wire n10217;
wire n10218;
wire n10219;
wire n10220;
wire n10221;
wire n10222;
wire n10223;
wire n10224;
wire n10225;
wire n10226;
wire n10227;
wire n10228;
wire n10229;
wire n10230;
wire n10231;
wire n10232;
wire n10233;
wire n10234;
wire n10235;
wire n10236;
wire n10237;
wire n10238;
wire n10239;
wire n10240;
wire n10241;
wire n10242;
wire n10243;
wire n10244;
wire n10245;
wire n10246;
wire n10247;
wire n10248;
wire n10249;
wire n10250;
wire n10251;
wire n10252;
wire n10253;
wire n10254;
wire n10255;
wire n10256;
wire n10257;
wire n10258;
wire n10259;
wire n1026;
wire n10260;
wire n10261;
wire n10262;
wire n10263;
wire n10264;
wire n10265;
wire n10266;
wire n10267;
wire n10268;
wire n10269;
wire n10270;
wire n10271;
wire n10272;
wire n10273;
wire n10274;
wire n10275;
wire n10276;
wire n10277;
wire n10278;
wire n10279;
wire n10280;
wire n10281;
wire n10282;
wire n10283;
wire n10284;
wire n10285;
wire n10286;
wire n10287;
wire n10288;
wire n10289;
wire n10290;
wire n10291;
wire n10292;
wire n10293;
wire n10294;
wire n10295;
wire n10296;
wire n10297;
wire n10298;
wire n10299;
wire n10300;
wire n10301;
wire n10302;
wire n10303;
wire n10304;
wire n10305;
wire n10306;
wire n10307;
wire n10308;
wire n10309;
wire n1031;
wire n10310;
wire n10311;
wire n10312;
wire n10313;
wire n10314;
wire n10315;
wire n10316;
wire n10317;
wire n10318;
wire n10319;
wire n10320;
wire n10321;
wire n10322;
wire n10323;
wire n10324;
wire n10325;
wire n10326;
wire n10327;
wire n10328;
wire n10329;
wire n10330;
wire n10331;
wire n10332;
wire n10333;
wire n10334;
wire n10335;
wire n10336;
wire n10337;
wire n10338;
wire n10339;
wire n10340;
wire n10341;
wire n10342;
wire n10343;
wire n10344;
wire n10345;
wire n10346;
wire n10347;
wire n10348;
wire n10349;
wire n1035;
wire n10350;
wire n10351;
wire n10352;
wire n10353;
wire n10354;
wire n10355;
wire n10356;
wire n10357;
wire n10358;
wire n10359;
wire n10360;
wire n10361;
wire n10362;
wire n10363;
wire n10364;
wire n10365;
wire n10366;
wire n10367;
wire n10368;
wire n10369;
wire n10370;
wire n10371;
wire n10372;
wire n10373;
wire n10374;
wire n10375;
wire n10376;
wire n10377;
wire n10378;
wire n10379;
wire n10380;
wire n10381;
wire n10382;
wire n10383;
wire n10384;
wire n10385;
wire n10386;
wire n10387;
wire n10388;
wire n10389;
wire n10390;
wire n10391;
wire n10392;
wire n10393;
wire n10394;
wire n10395;
wire n10396;
wire n10397;
wire n10398;
wire n10399;
wire n1040;
wire n10400;
wire n10401;
wire n10402;
wire n10403;
wire n10404;
wire n10405;
wire n10406;
wire n10407;
wire n10408;
wire n10409;
wire n10410;
wire n10411;
wire n10412;
wire n10413;
wire n10414;
wire n10415;
wire n10416;
wire n10417;
wire n10418;
wire n10419;
wire n10420;
wire n10421;
wire n10422;
wire n10423;
wire n10424;
wire n10425;
wire n10426;
wire n10427;
wire n10429;
wire n10430;
wire n10431;
wire n10432;
wire n10433;
wire n10434;
wire n10435;
wire n10436;
wire n10437;
wire n10438;
wire n10439;
wire n10440;
wire n10441;
wire n10442;
wire n10443;
wire n10444;
wire n10445;
wire n10446;
wire n10447;
wire n10448;
wire n10449;
wire n1045;
wire n10450;
wire n10451;
wire n10452;
wire n10453;
wire n10454;
wire n10455;
wire n10456;
wire n10457;
wire n10458;
wire n10459;
wire n10460;
wire n10461;
wire n10462;
wire n10463;
wire n10464;
wire n10465;
wire n10466;
wire n10467;
wire n10468;
wire n10469;
wire n10470;
wire n10471;
wire n10472;
wire n10473;
wire n10474;
wire n10475;
wire n10476;
wire n10477;
wire n10478;
wire n10479;
wire n10480;
wire n10481;
wire n10482;
wire n10483;
wire n10484;
wire n10485;
wire n10486;
wire n10487;
wire n10488;
wire n10489;
wire n10490;
wire n10491;
wire n10492;
wire n10493;
wire n10494;
wire n10495;
wire n10496;
wire n10497;
wire n10498;
wire n10499;
wire n1050;
wire n10500;
wire n10501;
wire n10502;
wire n10503;
wire n10504;
wire n10505;
wire n10506;
wire n10507;
wire n10508;
wire n10509;
wire n10510;
wire n10511;
wire n10512;
wire n10513;
wire n10514;
wire n10515;
wire n10516;
wire n10517;
wire n10518;
wire n10519;
wire n10520;
wire n10521;
wire n10522;
wire n10523;
wire n10524;
wire n10525;
wire n10526;
wire n10527;
wire n10528;
wire n10529;
wire n10530;
wire n10531;
wire n10532;
wire n10533;
wire n10534;
wire n10535;
wire n10536;
wire n10537;
wire n10538;
wire n10539;
wire n10540;
wire n10541;
wire n10542;
wire n10543;
wire n10544;
wire n10545;
wire n10546;
wire n10547;
wire n10548;
wire n10549;
wire n1055;
wire n10550;
wire n10551;
wire n10552;
wire n10553;
wire n10554;
wire n10555;
wire n10556;
wire n10557;
wire n10558;
wire n10559;
wire n10560;
wire n10561;
wire n10562;
wire n10563;
wire n10564;
wire n10565;
wire n10566;
wire n10567;
wire n10568;
wire n10569;
wire n10570;
wire n10571;
wire n10572;
wire n10573;
wire n10574;
wire n10575;
wire n10576;
wire n10577;
wire n10578;
wire n10579;
wire n10580;
wire n10581;
wire n10582;
wire n10583;
wire n10584;
wire n10585;
wire n10586;
wire n10587;
wire n10588;
wire n10589;
wire n10590;
wire n10591;
wire n10592;
wire n10593;
wire n10594;
wire n10595;
wire n10596;
wire n10597;
wire n10598;
wire n10599;
wire n1060;
wire n10600;
wire n10601;
wire n10602;
wire n10603;
wire n10604;
wire n10605;
wire n10606;
wire n10607;
wire n10608;
wire n10609;
wire n10610;
wire n10611;
wire n10612;
wire n10613;
wire n10614;
wire n10615;
wire n10616;
wire n10617;
wire n10618;
wire n10619;
wire n10620;
wire n10621;
wire n10622;
wire n10623;
wire n10624;
wire n10625;
wire n10626;
wire n10627;
wire n10628;
wire n10629;
wire n10630;
wire n10631;
wire n10632;
wire n10633;
wire n10634;
wire n10635;
wire n10636;
wire n10637;
wire n10638;
wire n10639;
wire n10640;
wire n10641;
wire n10642;
wire n10643;
wire n10644;
wire n10645;
wire n10646;
wire n10647;
wire n10648;
wire n10649;
wire n1065;
wire n10650;
wire n10651;
wire n10652;
wire n10653;
wire n10654;
wire n10655;
wire n10656;
wire n10657;
wire n10658;
wire n10659;
wire n10660;
wire n10661;
wire n10662;
wire n10663;
wire n10664;
wire n10665;
wire n10666;
wire n10667;
wire n10668;
wire n10669;
wire n10670;
wire n10671;
wire n10672;
wire n10673;
wire n10674;
wire n10675;
wire n10676;
wire n10677;
wire n10678;
wire n10679;
wire n10680;
wire n10681;
wire n10682;
wire n10683;
wire n10684;
wire n10685;
wire n10686;
wire n10687;
wire n10688;
wire n10689;
wire n10690;
wire n10691;
wire n10692;
wire n10693;
wire n10694;
wire n10695;
wire n10696;
wire n10697;
wire n10698;
wire n10699;
wire n1070;
wire n10700;
wire n10701;
wire n10702;
wire n10703;
wire n10704;
wire n10705;
wire n10706;
wire n10707;
wire n10708;
wire n10709;
wire n10710;
wire n10711;
wire n10712;
wire n10713;
wire n10714;
wire n10715;
wire n10716;
wire n10717;
wire n10718;
wire n10719;
wire n10720;
wire n10721;
wire n10722;
wire n10723;
wire n10724;
wire n10725;
wire n10726;
wire n10727;
wire n10728;
wire n10729;
wire n10730;
wire n10731;
wire n10732;
wire n10733;
wire n10734;
wire n10735;
wire n10737;
wire n10738;
wire n10739;
wire n10740;
wire n10741;
wire n10742;
wire n10743;
wire n10744;
wire n10745;
wire n10746;
wire n10747;
wire n10748;
wire n10749;
wire n1075;
wire n10750;
wire n10751;
wire n10752;
wire n10753;
wire n10754;
wire n10755;
wire n10756;
wire n10757;
wire n10758;
wire n10759;
wire n10760;
wire n10761;
wire n10762;
wire n10763;
wire n10764;
wire n10765;
wire n10766;
wire n10767;
wire n10768;
wire n10769;
wire n10770;
wire n10771;
wire n10772;
wire n10773;
wire n10774;
wire n10775;
wire n10776;
wire n10777;
wire n10778;
wire n10779;
wire n10780;
wire n10781;
wire n10782;
wire n10783;
wire n10784;
wire n10785;
wire n10786;
wire n10787;
wire n10788;
wire n10789;
wire n10790;
wire n10791;
wire n10792;
wire n10793;
wire n10794;
wire n10795;
wire n10796;
wire n10797;
wire n10798;
wire n10799;
wire n1080;
wire n10800;
wire n10801;
wire n10802;
wire n10803;
wire n10804;
wire n10805;
wire n10806;
wire n10807;
wire n10808;
wire n10809;
wire n10810;
wire n10811;
wire n10812;
wire n10813;
wire n10814;
wire n10815;
wire n10816;
wire n10817;
wire n10818;
wire n10819;
wire n10820;
wire n10821;
wire n10822;
wire n10823;
wire n10824;
wire n10825;
wire n10826;
wire n10827;
wire n10828;
wire n10829;
wire n10830;
wire n10831;
wire n10833;
wire n10834;
wire n10835;
wire n10836;
wire n10837;
wire n10838;
wire n10839;
wire n10840;
wire n10841;
wire n10842;
wire n10843;
wire n10844;
wire n10845;
wire n10846;
wire n10847;
wire n10848;
wire n10849;
wire n1085;
wire n10850;
wire n10851;
wire n10852;
wire n10853;
wire n10854;
wire n10855;
wire n10856;
wire n10857;
wire n10858;
wire n10859;
wire n10860;
wire n10861;
wire n10862;
wire n10863;
wire n10864;
wire n10865;
wire n10866;
wire n10867;
wire n10868;
wire n10869;
wire n10870;
wire n10871;
wire n10872;
wire n10873;
wire n10874;
wire n10875;
wire n10876;
wire n10877;
wire n10878;
wire n10879;
wire n10880;
wire n10881;
wire n10882;
wire n10883;
wire n10884;
wire n10885;
wire n10886;
wire n10887;
wire n10888;
wire n10889;
wire n10890;
wire n10891;
wire n10892;
wire n10893;
wire n10894;
wire n10895;
wire n10896;
wire n10897;
wire n10898;
wire n10899;
wire n1090;
wire n10900;
wire n10901;
wire n10902;
wire n10903;
wire n10904;
wire n10905;
wire n10906;
wire n10907;
wire n10908;
wire n10909;
wire n10910;
wire n10911;
wire n10912;
wire n10913;
wire n10914;
wire n10915;
wire n10916;
wire n10917;
wire n10918;
wire n10919;
wire n10920;
wire n10921;
wire n10922;
wire n10923;
wire n10924;
wire n10925;
wire n10926;
wire n10927;
wire n10928;
wire n10929;
wire n10930;
wire n10931;
wire n10932;
wire n10933;
wire n10934;
wire n10935;
wire n10936;
wire n10937;
wire n10938;
wire n10939;
wire n10940;
wire n10941;
wire n10942;
wire n10943;
wire n10944;
wire n10945;
wire n10946;
wire n10947;
wire n10948;
wire n10949;
wire n1095;
wire n10950;
wire n10951;
wire n10952;
wire n10953;
wire n10954;
wire n10955;
wire n10956;
wire n10957;
wire n10958;
wire n10959;
wire n10960;
wire n10961;
wire n10962;
wire n10963;
wire n10964;
wire n10965;
wire n10966;
wire n10967;
wire n10968;
wire n10969;
wire n10970;
wire n10971;
wire n10972;
wire n10973;
wire n10974;
wire n10975;
wire n10976;
wire n10977;
wire n10978;
wire n10979;
wire n10980;
wire n10981;
wire n10982;
wire n10983;
wire n10984;
wire n10985;
wire n10986;
wire n10987;
wire n10988;
wire n10989;
wire n10990;
wire n10991;
wire n10992;
wire n10993;
wire n10994;
wire n10995;
wire n10996;
wire n10997;
wire n10998;
wire n10999;
wire n1100;
wire n11000;
wire n11001;
wire n11002;
wire n11003;
wire n11004;
wire n11005;
wire n11006;
wire n11007;
wire n11008;
wire n11009;
wire n11010;
wire n11011;
wire n11012;
wire n11013;
wire n11015;
wire n11016;
wire n11017;
wire n11018;
wire n11019;
wire n11020;
wire n11021;
wire n11022;
wire n11023;
wire n11024;
wire n11025;
wire n11026;
wire n11027;
wire n11028;
wire n11029;
wire n11030;
wire n11031;
wire n11032;
wire n11033;
wire n11034;
wire n11035;
wire n11036;
wire n11037;
wire n11038;
wire n11039;
wire n11040;
wire n11041;
wire n11042;
wire n11043;
wire n11044;
wire n11045;
wire n11046;
wire n11047;
wire n11048;
wire n11049;
wire n1105;
wire n11050;
wire n11051;
wire n11052;
wire n11053;
wire n11054;
wire n11055;
wire n11056;
wire n11057;
wire n11058;
wire n11059;
wire n11060;
wire n11061;
wire n11062;
wire n11063;
wire n11064;
wire n11065;
wire n11066;
wire n11067;
wire n11068;
wire n11069;
wire n11070;
wire n11071;
wire n11072;
wire n11073;
wire n11074;
wire n11075;
wire n11076;
wire n11077;
wire n11078;
wire n11079;
wire n11080;
wire n11081;
wire n11082;
wire n11083;
wire n11084;
wire n11085;
wire n11086;
wire n11087;
wire n11088;
wire n11089;
wire n11090;
wire n11091;
wire n11092;
wire n11093;
wire n11094;
wire n11095;
wire n11096;
wire n11097;
wire n11098;
wire n11099;
wire n1110;
wire n11100;
wire n11101;
wire n11102;
wire n11103;
wire n11104;
wire n11105;
wire n11106;
wire n11107;
wire n11108;
wire n11109;
wire n11110;
wire n11111;
wire n11112;
wire n11113;
wire n11114;
wire n11115;
wire n11116;
wire n11117;
wire n11118;
wire n11119;
wire n11120;
wire n11121;
wire n11122;
wire n11123;
wire n11124;
wire n11125;
wire n11126;
wire n11127;
wire n11128;
wire n11129;
wire n11130;
wire n11131;
wire n11132;
wire n11133;
wire n11134;
wire n11135;
wire n11136;
wire n11137;
wire n11138;
wire n11139;
wire n11140;
wire n11141;
wire n11142;
wire n11143;
wire n11144;
wire n11145;
wire n11146;
wire n11147;
wire n11148;
wire n11149;
wire n1115;
wire n11150;
wire n11151;
wire n11152;
wire n11153;
wire n11154;
wire n11155;
wire n11156;
wire n11157;
wire n11158;
wire n11159;
wire n11160;
wire n11161;
wire n11162;
wire n11163;
wire n11164;
wire n11165;
wire n11166;
wire n11167;
wire n11168;
wire n11169;
wire n11170;
wire n11171;
wire n11172;
wire n11173;
wire n11174;
wire n11175;
wire n11176;
wire n11177;
wire n11178;
wire n11179;
wire n11180;
wire n11181;
wire n11182;
wire n11183;
wire n11184;
wire n11185;
wire n11186;
wire n11187;
wire n11188;
wire n11189;
wire n11190;
wire n11191;
wire n11192;
wire n11193;
wire n11194;
wire n11195;
wire n11196;
wire n11197;
wire n11198;
wire n11199;
wire n1120;
wire n11200;
wire n11201;
wire n11202;
wire n11203;
wire n11204;
wire n11205;
wire n11206;
wire n11207;
wire n11208;
wire n11209;
wire n11210;
wire n11211;
wire n11212;
wire n11213;
wire n11214;
wire n11215;
wire n11216;
wire n11217;
wire n11218;
wire n11219;
wire n11220;
wire n11221;
wire n11222;
wire n11223;
wire n11224;
wire n11225;
wire n11226;
wire n11227;
wire n11228;
wire n11229;
wire n11230;
wire n11231;
wire n11232;
wire n11233;
wire n11234;
wire n11235;
wire n11236;
wire n11237;
wire n11238;
wire n11239;
wire n11240;
wire n11241;
wire n11242;
wire n11243;
wire n11244;
wire n11245;
wire n11246;
wire n11247;
wire n11248;
wire n11249;
wire n1125;
wire n11250;
wire n11251;
wire n11252;
wire n11253;
wire n11254;
wire n11255;
wire n11256;
wire n11257;
wire n11258;
wire n11259;
wire n11260;
wire n11261;
wire n11262;
wire n11263;
wire n11264;
wire n11265;
wire n11266;
wire n11267;
wire n11268;
wire n11269;
wire n11270;
wire n11271;
wire n11272;
wire n11273;
wire n11274;
wire n11275;
wire n11276;
wire n11277;
wire n11278;
wire n11279;
wire n11280;
wire n11281;
wire n11282;
wire n11283;
wire n11284;
wire n11285;
wire n11286;
wire n11287;
wire n11288;
wire n11289;
wire n11290;
wire n11291;
wire n11292;
wire n11293;
wire n11294;
wire n11295;
wire n11296;
wire n11297;
wire n11298;
wire n11299;
wire n1130;
wire n11300;
wire n11301;
wire n11302;
wire n11303;
wire n11304;
wire n11305;
wire n11306;
wire n11307;
wire n11308;
wire n11309;
wire n11310;
wire n11311;
wire n11312;
wire n11313;
wire n11314;
wire n11315;
wire n11316;
wire n11317;
wire n11318;
wire n11319;
wire n11320;
wire n11321;
wire n11322;
wire n11323;
wire n11324;
wire n11325;
wire n11326;
wire n11327;
wire n11328;
wire n11329;
wire n11330;
wire n11331;
wire n11332;
wire n11333;
wire n11334;
wire n11335;
wire n11336;
wire n11337;
wire n11338;
wire n11339;
wire n11340;
wire n11341;
wire n11342;
wire n11343;
wire n11344;
wire n11345;
wire n11346;
wire n11347;
wire n11348;
wire n11349;
wire n1135;
wire n11350;
wire n11351;
wire n11352;
wire n11353;
wire n11354;
wire n11355;
wire n11356;
wire n11357;
wire n11358;
wire n11359;
wire n11360;
wire n11361;
wire n11362;
wire n11363;
wire n11364;
wire n11365;
wire n11366;
wire n11367;
wire n11368;
wire n11369;
wire n11370;
wire n11371;
wire n11372;
wire n11373;
wire n11374;
wire n11375;
wire n11376;
wire n11377;
wire n11378;
wire n11379;
wire n11380;
wire n11381;
wire n11382;
wire n11383;
wire n11384;
wire n11385;
wire n11386;
wire n11387;
wire n11388;
wire n11389;
wire n11390;
wire n11391;
wire n11392;
wire n11393;
wire n11394;
wire n11395;
wire n11396;
wire n11397;
wire n11398;
wire n11399;
wire n1140;
wire n11400;
wire n11401;
wire n11402;
wire n11403;
wire n11404;
wire n11405;
wire n11406;
wire n11407;
wire n11408;
wire n11409;
wire n11410;
wire n11411;
wire n11412;
wire n11413;
wire n11414;
wire n11415;
wire n11416;
wire n11417;
wire n11418;
wire n11419;
wire n11420;
wire n11421;
wire n11422;
wire n11423;
wire n11424;
wire n11425;
wire n11426;
wire n11427;
wire n11428;
wire n11429;
wire n11430;
wire n11431;
wire n11432;
wire n11433;
wire n11434;
wire n11435;
wire n11436;
wire n11437;
wire n11438;
wire n11439;
wire n11440;
wire n11441;
wire n11442;
wire n11443;
wire n11444;
wire n11445;
wire n11446;
wire n11447;
wire n11448;
wire n11449;
wire n1145;
wire n11450;
wire n11451;
wire n11452;
wire n11453;
wire n11454;
wire n11455;
wire n11456;
wire n11457;
wire n11458;
wire n11459;
wire n11460;
wire n11461;
wire n11462;
wire n11463;
wire n11464;
wire n11465;
wire n11466;
wire n11467;
wire n11468;
wire n11469;
wire n11470;
wire n11471;
wire n11472;
wire n11473;
wire n11474;
wire n11475;
wire n11476;
wire n11477;
wire n11478;
wire n11479;
wire n11480;
wire n11481;
wire n11482;
wire n11483;
wire n11484;
wire n11485;
wire n11486;
wire n11487;
wire n11488;
wire n11489;
wire n11490;
wire n11491;
wire n11492;
wire n11493;
wire n11494;
wire n11495;
wire n11496;
wire n11497;
wire n11498;
wire n11499;
wire n1150;
wire n11500;
wire n11501;
wire n11502;
wire n11503;
wire n11504;
wire n11505;
wire n11506;
wire n11507;
wire n11508;
wire n11509;
wire n11510;
wire n11511;
wire n11512;
wire n11513;
wire n11514;
wire n11515;
wire n11516;
wire n11517;
wire n11518;
wire n11519;
wire n11520;
wire n11521;
wire n11522;
wire n11523;
wire n11524;
wire n11525;
wire n11526;
wire n11527;
wire n11528;
wire n11529;
wire n11530;
wire n11531;
wire n11532;
wire n11533;
wire n11534;
wire n11535;
wire n11536;
wire n11537;
wire n11538;
wire n11539;
wire n11540;
wire n11541;
wire n11542;
wire n11543;
wire n11544;
wire n11545;
wire n11546;
wire n11547;
wire n11548;
wire n11549;
wire n1155;
wire n11550;
wire n11551;
wire n11552;
wire n11553;
wire n11554;
wire n11555;
wire n11556;
wire n11557;
wire n11558;
wire n11559;
wire n11560;
wire n11561;
wire n11562;
wire n11563;
wire n11564;
wire n11565;
wire n11566;
wire n11567;
wire n11568;
wire n11569;
wire n11570;
wire n11571;
wire n11572;
wire n11573;
wire n11574;
wire n11575;
wire n11576;
wire n11577;
wire n11578;
wire n11579;
wire n11580;
wire n11581;
wire n11582;
wire n11583;
wire n11584;
wire n11585;
wire n11586;
wire n11587;
wire n11588;
wire n11589;
wire n11590;
wire n11591;
wire n11592;
wire n11593;
wire n11594;
wire n11595;
wire n11596;
wire n11597;
wire n11598;
wire n11599;
wire n1160;
wire n11600;
wire n11601;
wire n11602;
wire n11603;
wire n11604;
wire n11605;
wire n11606;
wire n11607;
wire n11608;
wire n11609;
wire n11610;
wire n11611;
wire n11612;
wire n11613;
wire n11614;
wire n11615;
wire n11616;
wire n11617;
wire n11618;
wire n11619;
wire n11620;
wire n11621;
wire n11622;
wire n11623;
wire n11624;
wire n11625;
wire n11626;
wire n11627;
wire n11628;
wire n11629;
wire n11630;
wire n11631;
wire n11632;
wire n11633;
wire n11634;
wire n11635;
wire n11636;
wire n11637;
wire n11638;
wire n11639;
wire n11640;
wire n11641;
wire n11642;
wire n11643;
wire n11644;
wire n11645;
wire n11646;
wire n11647;
wire n11648;
wire n11649;
wire n1165;
wire n11650;
wire n11651;
wire n11652;
wire n11653;
wire n11654;
wire n11655;
wire n11656;
wire n11657;
wire n11658;
wire n11659;
wire n11660;
wire n11661;
wire n11662;
wire n11663;
wire n11664;
wire n11665;
wire n11666;
wire n11667;
wire n11668;
wire n11669;
wire n11670;
wire n11671;
wire n11672;
wire n11673;
wire n11674;
wire n11675;
wire n11676;
wire n11677;
wire n11678;
wire n11679;
wire n11680;
wire n11681;
wire n11682;
wire n11683;
wire n11684;
wire n11685;
wire n11686;
wire n11687;
wire n11688;
wire n11689;
wire n11690;
wire n11691;
wire n11692;
wire n11693;
wire n11694;
wire n11695;
wire n11696;
wire n11697;
wire n11698;
wire n11699;
wire n1170;
wire n11700;
wire n11701;
wire n11702;
wire n11703;
wire n11704;
wire n11705;
wire n11706;
wire n11707;
wire n11708;
wire n11709;
wire n11710;
wire n11711;
wire n11712;
wire n11713;
wire n11714;
wire n11715;
wire n11716;
wire n11717;
wire n11718;
wire n11719;
wire n11720;
wire n11721;
wire n11722;
wire n11723;
wire n11724;
wire n11725;
wire n11726;
wire n11727;
wire n11728;
wire n11729;
wire n11730;
wire n11731;
wire n11732;
wire n11733;
wire n11734;
wire n11735;
wire n11736;
wire n11737;
wire n11738;
wire n11739;
wire n11740;
wire n11741;
wire n11742;
wire n11743;
wire n11744;
wire n11745;
wire n11746;
wire n11747;
wire n11748;
wire n11749;
wire n1175;
wire n11750;
wire n11751;
wire n11752;
wire n11753;
wire n11754;
wire n11755;
wire n11756;
wire n11757;
wire n11758;
wire n11759;
wire n11760;
wire n11761;
wire n11762;
wire n11763;
wire n11764;
wire n11765;
wire n11766;
wire n11767;
wire n11768;
wire n11769;
wire n11770;
wire n11771;
wire n11772;
wire n11773;
wire n11774;
wire n11775;
wire n11776;
wire n11777;
wire n11778;
wire n11779;
wire n11780;
wire n11781;
wire n11782;
wire n11783;
wire n11784;
wire n11785;
wire n11786;
wire n11787;
wire n11788;
wire n11789;
wire n11790;
wire n11791;
wire n11792;
wire n11793;
wire n11794;
wire n11795;
wire n11796;
wire n11797;
wire n11798;
wire n11799;
wire n1180;
wire n11800;
wire n11801;
wire n11802;
wire n11803;
wire n11804;
wire n11805;
wire n11806;
wire n11807;
wire n11808;
wire n11809;
wire n11810;
wire n11811;
wire n11812;
wire n11813;
wire n11814;
wire n11815;
wire n11816;
wire n11817;
wire n11818;
wire n11819;
wire n11820;
wire n11821;
wire n11822;
wire n11823;
wire n11824;
wire n11825;
wire n11826;
wire n11827;
wire n11828;
wire n11829;
wire n11830;
wire n11831;
wire n11832;
wire n11833;
wire n11834;
wire n11835;
wire n11836;
wire n11837;
wire n11838;
wire n11839;
wire n11840;
wire n11841;
wire n11842;
wire n11843;
wire n11844;
wire n11845;
wire n11846;
wire n11847;
wire n11848;
wire n11849;
wire n1185;
wire n11850;
wire n11851;
wire n11852;
wire n11853;
wire n11854;
wire n11855;
wire n11856;
wire n11857;
wire n11858;
wire n11859;
wire n11860;
wire n11861;
wire n11862;
wire n11863;
wire n11864;
wire n11865;
wire n11866;
wire n11867;
wire n11868;
wire n11870;
wire n11871;
wire n11872;
wire n11873;
wire n11874;
wire n11875;
wire n11876;
wire n11877;
wire n11878;
wire n11879;
wire n11880;
wire n11881;
wire n11882;
wire n11883;
wire n11884;
wire n11885;
wire n11886;
wire n11887;
wire n11888;
wire n11889;
wire n11890;
wire n11891;
wire n11892;
wire n11893;
wire n11894;
wire n11895;
wire n11896;
wire n11897;
wire n11898;
wire n11899;
wire n1190;
wire n11900;
wire n11901;
wire n11902;
wire n11903;
wire n11904;
wire n11905;
wire n11906;
wire n11907;
wire n11908;
wire n11909;
wire n11910;
wire n11911;
wire n11912;
wire n11913;
wire n11914;
wire n11915;
wire n11916;
wire n11917;
wire n11918;
wire n11919;
wire n11920;
wire n11921;
wire n11922;
wire n11923;
wire n11924;
wire n11925;
wire n11926;
wire n11927;
wire n11928;
wire n11929;
wire n11930;
wire n11931;
wire n11932;
wire n11933;
wire n11934;
wire n11935;
wire n11936;
wire n11937;
wire n11938;
wire n11939;
wire n11940;
wire n11941;
wire n11942;
wire n11943;
wire n11944;
wire n11945;
wire n11946;
wire n11947;
wire n11948;
wire n11949;
wire n1195;
wire n11950;
wire n11951;
wire n11952;
wire n11953;
wire n11954;
wire n11955;
wire n11956;
wire n11957;
wire n11958;
wire n11959;
wire n11960;
wire n11961;
wire n11962;
wire n11963;
wire n11964;
wire n11965;
wire n11966;
wire n11967;
wire n11968;
wire n11969;
wire n11970;
wire n11971;
wire n11972;
wire n11973;
wire n11974;
wire n11975;
wire n11976;
wire n11977;
wire n11978;
wire n11979;
wire n11980;
wire n11981;
wire n11982;
wire n11983;
wire n11984;
wire n11985;
wire n11986;
wire n11987;
wire n11988;
wire n11989;
wire n11990;
wire n11991;
wire n11992;
wire n11993;
wire n11994;
wire n11995;
wire n11996;
wire n11997;
wire n11998;
wire n11999;
wire n1200;
wire n12000;
wire n12001;
wire n12002;
wire n12003;
wire n12004;
wire n12005;
wire n12006;
wire n12007;
wire n12008;
wire n12009;
wire n12010;
wire n12011;
wire n12012;
wire n12013;
wire n12014;
wire n12015;
wire n12016;
wire n12017;
wire n12018;
wire n12019;
wire n12020;
wire n12021;
wire n12022;
wire n12023;
wire n12024;
wire n12025;
wire n12026;
wire n12027;
wire n12028;
wire n12029;
wire n12030;
wire n12031;
wire n12032;
wire n12033;
wire n12034;
wire n12035;
wire n12036;
wire n12037;
wire n12038;
wire n12039;
wire n12040;
wire n12041;
wire n12042;
wire n12043;
wire n12044;
wire n12045;
wire n12046;
wire n12047;
wire n12048;
wire n12049;
wire n1205;
wire n12050;
wire n12051;
wire n12052;
wire n12053;
wire n12054;
wire n12055;
wire n12056;
wire n12057;
wire n12058;
wire n12059;
wire n12060;
wire n12061;
wire n12062;
wire n12063;
wire n12064;
wire n12065;
wire n12066;
wire n12067;
wire n12068;
wire n12069;
wire n12070;
wire n12071;
wire n12072;
wire n12073;
wire n12074;
wire n12075;
wire n12076;
wire n12077;
wire n12078;
wire n12079;
wire n12080;
wire n12081;
wire n12082;
wire n12083;
wire n12084;
wire n12085;
wire n12086;
wire n12087;
wire n12088;
wire n12089;
wire n12090;
wire n12091;
wire n12092;
wire n12093;
wire n12094;
wire n12095;
wire n12096;
wire n12097;
wire n12098;
wire n12099;
wire n1210;
wire n12100;
wire n12101;
wire n12102;
wire n12103;
wire n12104;
wire n12105;
wire n12106;
wire n12107;
wire n12108;
wire n12109;
wire n12110;
wire n12111;
wire n12112;
wire n12113;
wire n12114;
wire n12115;
wire n12116;
wire n12117;
wire n12118;
wire n12119;
wire n12120;
wire n12121;
wire n12122;
wire n12123;
wire n12124;
wire n12125;
wire n12126;
wire n12127;
wire n12128;
wire n12129;
wire n12130;
wire n12131;
wire n12132;
wire n12133;
wire n12134;
wire n12135;
wire n12136;
wire n12137;
wire n12138;
wire n12139;
wire n12140;
wire n12141;
wire n12142;
wire n12143;
wire n12144;
wire n12145;
wire n12146;
wire n12147;
wire n12148;
wire n12149;
wire n1215;
wire n12150;
wire n12151;
wire n12152;
wire n12153;
wire n12154;
wire n12155;
wire n12156;
wire n12157;
wire n12158;
wire n12159;
wire n12160;
wire n12161;
wire n12162;
wire n12163;
wire n12164;
wire n12165;
wire n12166;
wire n12167;
wire n12168;
wire n12169;
wire n12170;
wire n12171;
wire n12172;
wire n12173;
wire n12174;
wire n12175;
wire n12176;
wire n12177;
wire n12178;
wire n12179;
wire n12180;
wire n12181;
wire n12182;
wire n12183;
wire n12184;
wire n12185;
wire n12186;
wire n12187;
wire n12188;
wire n12189;
wire n12190;
wire n12191;
wire n12192;
wire n12193;
wire n12194;
wire n12195;
wire n12196;
wire n12197;
wire n12198;
wire n12199;
wire n1220;
wire n12200;
wire n12201;
wire n12202;
wire n12203;
wire n12204;
wire n12205;
wire n12206;
wire n12207;
wire n12208;
wire n12209;
wire n12210;
wire n12211;
wire n12212;
wire n12213;
wire n12214;
wire n12215;
wire n12216;
wire n12217;
wire n12218;
wire n12219;
wire n12220;
wire n12221;
wire n12222;
wire n12223;
wire n12224;
wire n12225;
wire n12226;
wire n12227;
wire n12228;
wire n12229;
wire n12230;
wire n12231;
wire n12232;
wire n12233;
wire n12234;
wire n12235;
wire n12236;
wire n12237;
wire n12238;
wire n12239;
wire n12240;
wire n12241;
wire n12242;
wire n12243;
wire n12244;
wire n12245;
wire n12246;
wire n12247;
wire n12248;
wire n12249;
wire n1225;
wire n12250;
wire n12251;
wire n12252;
wire n12253;
wire n12254;
wire n12255;
wire n12256;
wire n12257;
wire n12258;
wire n12259;
wire n12260;
wire n12261;
wire n12262;
wire n12263;
wire n12264;
wire n12265;
wire n12266;
wire n12267;
wire n12268;
wire n12269;
wire n12270;
wire n12271;
wire n12272;
wire n12273;
wire n12274;
wire n12275;
wire n12276;
wire n12277;
wire n12278;
wire n12279;
wire n12280;
wire n12281;
wire n12282;
wire n12283;
wire n12284;
wire n12285;
wire n12286;
wire n12287;
wire n12288;
wire n12289;
wire n12290;
wire n12291;
wire n12292;
wire n12293;
wire n12294;
wire n12295;
wire n12296;
wire n12297;
wire n12298;
wire n12299;
wire n1230;
wire n12300;
wire n12301;
wire n12302;
wire n12303;
wire n12304;
wire n12305;
wire n12306;
wire n12307;
wire n12308;
wire n12309;
wire n12310;
wire n12311;
wire n12312;
wire n12313;
wire n12314;
wire n12315;
wire n12316;
wire n12317;
wire n12318;
wire n12319;
wire n12320;
wire n12321;
wire n12322;
wire n12323;
wire n12324;
wire n12325;
wire n12326;
wire n12327;
wire n12328;
wire n12329;
wire n12330;
wire n12331;
wire n12332;
wire n12333;
wire n12334;
wire n12335;
wire n12336;
wire n12337;
wire n12338;
wire n12339;
wire n12340;
wire n12341;
wire n12342;
wire n12343;
wire n12344;
wire n12345;
wire n12346;
wire n12347;
wire n12348;
wire n12349;
wire n1235;
wire n12350;
wire n12351;
wire n12352;
wire n12353;
wire n12354;
wire n12355;
wire n12356;
wire n12357;
wire n12358;
wire n12359;
wire n12360;
wire n12361;
wire n12362;
wire n12363;
wire n12364;
wire n12365;
wire n12366;
wire n12367;
wire n12368;
wire n12369;
wire n12370;
wire n12371;
wire n12372;
wire n12373;
wire n12374;
wire n12375;
wire n12376;
wire n12377;
wire n12378;
wire n12379;
wire n12380;
wire n12381;
wire n12382;
wire n12383;
wire n12384;
wire n12385;
wire n12386;
wire n12387;
wire n12388;
wire n12389;
wire n12390;
wire n12391;
wire n12392;
wire n12393;
wire n12394;
wire n12395;
wire n12396;
wire n12397;
wire n12398;
wire n12399;
wire n1240;
wire n12400;
wire n12401;
wire n12402;
wire n12403;
wire n12404;
wire n12405;
wire n12406;
wire n12407;
wire n12408;
wire n12409;
wire n12410;
wire n12411;
wire n12412;
wire n12413;
wire n12414;
wire n12415;
wire n12416;
wire n12417;
wire n12418;
wire n12419;
wire n12420;
wire n12421;
wire n12422;
wire n12423;
wire n12424;
wire n12425;
wire n12426;
wire n12427;
wire n12428;
wire n12429;
wire n12430;
wire n12431;
wire n12432;
wire n12433;
wire n12434;
wire n12435;
wire n12436;
wire n12437;
wire n12438;
wire n12439;
wire n12440;
wire n12441;
wire n12442;
wire n12443;
wire n12444;
wire n12445;
wire n12446;
wire n12447;
wire n12448;
wire n12449;
wire n1245;
wire n12450;
wire n12451;
wire n12452;
wire n12453;
wire n12454;
wire n12455;
wire n12456;
wire n12457;
wire n12458;
wire n12459;
wire n12460;
wire n12461;
wire n12462;
wire n12463;
wire n12464;
wire n12465;
wire n12466;
wire n12467;
wire n12468;
wire n12469;
wire n12470;
wire n12471;
wire n12472;
wire n12473;
wire n12474;
wire n12475;
wire n12476;
wire n12477;
wire n12478;
wire n12479;
wire n12480;
wire n12481;
wire n12482;
wire n12483;
wire n12484;
wire n12485;
wire n12486;
wire n12487;
wire n12488;
wire n12489;
wire n12490;
wire n12491;
wire n12492;
wire n12493;
wire n12494;
wire n12495;
wire n12496;
wire n12497;
wire n12498;
wire n12499;
wire n1250;
wire n12500;
wire n12501;
wire n12502;
wire n12503;
wire n12504;
wire n12505;
wire n12506;
wire n12507;
wire n12508;
wire n12509;
wire n12510;
wire n12511;
wire n12512;
wire n12513;
wire n12514;
wire n12515;
wire n12516;
wire n12517;
wire n12518;
wire n12519;
wire n12520;
wire n12521;
wire n12522;
wire n12523;
wire n12524;
wire n12525;
wire n12526;
wire n12527;
wire n12528;
wire n12529;
wire n12530;
wire n12531;
wire n12532;
wire n12533;
wire n12534;
wire n12535;
wire n12536;
wire n12537;
wire n12538;
wire n12539;
wire n12540;
wire n12541;
wire n12542;
wire n12543;
wire n12544;
wire n12545;
wire n12546;
wire n12547;
wire n12548;
wire n12549;
wire n1255;
wire n12550;
wire n12551;
wire n12552;
wire n12553;
wire n12554;
wire n12555;
wire n12556;
wire n12557;
wire n12558;
wire n12559;
wire n12560;
wire n12561;
wire n12562;
wire n12563;
wire n12564;
wire n12565;
wire n12566;
wire n12567;
wire n12568;
wire n12569;
wire n12570;
wire n12571;
wire n12572;
wire n12573;
wire n12574;
wire n12575;
wire n12576;
wire n12577;
wire n12578;
wire n12579;
wire n12580;
wire n12581;
wire n12582;
wire n12583;
wire n12584;
wire n12585;
wire n12586;
wire n12587;
wire n12588;
wire n12589;
wire n12590;
wire n12591;
wire n12592;
wire n12593;
wire n12594;
wire n12595;
wire n12596;
wire n12597;
wire n12598;
wire n12599;
wire n1260;
wire n12600;
wire n12601;
wire n12602;
wire n12603;
wire n12604;
wire n12605;
wire n12606;
wire n12607;
wire n12608;
wire n12609;
wire n12610;
wire n12611;
wire n12612;
wire n12613;
wire n12614;
wire n12615;
wire n12616;
wire n12617;
wire n12618;
wire n12619;
wire n12620;
wire n12621;
wire n12622;
wire n12623;
wire n12624;
wire n12625;
wire n12626;
wire n12627;
wire n12628;
wire n12629;
wire n12630;
wire n12631;
wire n12632;
wire n12633;
wire n12634;
wire n12635;
wire n12636;
wire n12637;
wire n12638;
wire n12639;
wire n12640;
wire n12641;
wire n12642;
wire n12643;
wire n12644;
wire n12645;
wire n12646;
wire n12647;
wire n12648;
wire n12649;
wire n1265;
wire n12650;
wire n12651;
wire n12652;
wire n12653;
wire n12654;
wire n12655;
wire n12656;
wire n12657;
wire n12658;
wire n12659;
wire n12660;
wire n12661;
wire n12662;
wire n12663;
wire n12664;
wire n12665;
wire n12666;
wire n12667;
wire n12668;
wire n12669;
wire n12670;
wire n12671;
wire n12672;
wire n12673;
wire n12674;
wire n12675;
wire n12676;
wire n12677;
wire n12678;
wire n12679;
wire n12680;
wire n12681;
wire n12682;
wire n12683;
wire n12684;
wire n12685;
wire n12686;
wire n12687;
wire n12688;
wire n12689;
wire n12690;
wire n12691;
wire n12692;
wire n12693;
wire n12694;
wire n12695;
wire n12696;
wire n12697;
wire n12698;
wire n12699;
wire n1270;
wire n12700;
wire n12701;
wire n12702;
wire n12703;
wire n12704;
wire n12705;
wire n12706;
wire n12707;
wire n12708;
wire n12709;
wire n12710;
wire n12711;
wire n12712;
wire n12713;
wire n12714;
wire n12715;
wire n12716;
wire n12717;
wire n12718;
wire n12719;
wire n12720;
wire n12721;
wire n12722;
wire n12723;
wire n12724;
wire n12725;
wire n12726;
wire n12727;
wire n12728;
wire n12729;
wire n12730;
wire n12731;
wire n12732;
wire n12733;
wire n12734;
wire n12735;
wire n12736;
wire n12737;
wire n12738;
wire n12739;
wire n12740;
wire n12741;
wire n12742;
wire n12743;
wire n12744;
wire n12745;
wire n12746;
wire n12747;
wire n12748;
wire n12749;
wire n1275;
wire n12750;
wire n12751;
wire n12752;
wire n12753;
wire n12754;
wire n12755;
wire n12756;
wire n12757;
wire n12758;
wire n12759;
wire n12760;
wire n12761;
wire n12762;
wire n12763;
wire n12764;
wire n12765;
wire n12766;
wire n12767;
wire n12768;
wire n12769;
wire n12770;
wire n12771;
wire n12772;
wire n12773;
wire n12774;
wire n12775;
wire n12776;
wire n12777;
wire n12778;
wire n12779;
wire n12780;
wire n12781;
wire n12782;
wire n12783;
wire n12784;
wire n12785;
wire n12786;
wire n12787;
wire n12788;
wire n12789;
wire n12790;
wire n12791;
wire n12792;
wire n12793;
wire n12794;
wire n12795;
wire n12796;
wire n12797;
wire n12798;
wire n12799;
wire n1280;
wire n12800;
wire n12801;
wire n12802;
wire n12803;
wire n12804;
wire n12805;
wire n12806;
wire n12807;
wire n12808;
wire n12809;
wire n12810;
wire n12811;
wire n12812;
wire n12813;
wire n12814;
wire n12815;
wire n12816;
wire n12817;
wire n12818;
wire n12819;
wire n12820;
wire n12821;
wire n12822;
wire n12823;
wire n12824;
wire n12825;
wire n12826;
wire n12827;
wire n12828;
wire n12829;
wire n12830;
wire n12831;
wire n12832;
wire n12833;
wire n12834;
wire n12835;
wire n12836;
wire n12837;
wire n12838;
wire n12839;
wire n12840;
wire n12841;
wire n12842;
wire n12843;
wire n12844;
wire n12845;
wire n12846;
wire n12847;
wire n12848;
wire n12849;
wire n1285;
wire n12850;
wire n12851;
wire n12852;
wire n12853;
wire n12854;
wire n12855;
wire n12856;
wire n12857;
wire n12858;
wire n12859;
wire n12860;
wire n12861;
wire n12862;
wire n12863;
wire n12864;
wire n12865;
wire n12866;
wire n12867;
wire n12868;
wire n12869;
wire n12870;
wire n12871;
wire n12872;
wire n12873;
wire n12874;
wire n12875;
wire n12876;
wire n12877;
wire n12878;
wire n12879;
wire n12880;
wire n12881;
wire n12882;
wire n12883;
wire n12884;
wire n12885;
wire n12886;
wire n12887;
wire n12888;
wire n12889;
wire n12890;
wire n12891;
wire n12892;
wire n12893;
wire n12894;
wire n12895;
wire n12896;
wire n12897;
wire n12898;
wire n12899;
wire n1290;
wire n12900;
wire n12901;
wire n12902;
wire n12903;
wire n12904;
wire n12905;
wire n12906;
wire n12907;
wire n12908;
wire n12909;
wire n12910;
wire n12911;
wire n12912;
wire n12913;
wire n12914;
wire n12915;
wire n12916;
wire n12917;
wire n12918;
wire n12919;
wire n12920;
wire n12921;
wire n12922;
wire n12923;
wire n12924;
wire n12925;
wire n12926;
wire n12927;
wire n12928;
wire n12929;
wire n12930;
wire n12931;
wire n12932;
wire n12933;
wire n12934;
wire n12935;
wire n12936;
wire n12937;
wire n12938;
wire n12939;
wire n12940;
wire n12941;
wire n12942;
wire n12943;
wire n12944;
wire n12945;
wire n12946;
wire n12947;
wire n12948;
wire n12949;
wire n1295;
wire n12950;
wire n12951;
wire n12952;
wire n12953;
wire n12954;
wire n12955;
wire n12956;
wire n12957;
wire n12958;
wire n12959;
wire n12960;
wire n12961;
wire n12962;
wire n12963;
wire n12964;
wire n12965;
wire n12966;
wire n12967;
wire n12968;
wire n12969;
wire n12970;
wire n12971;
wire n12972;
wire n12973;
wire n12974;
wire n12975;
wire n12976;
wire n12977;
wire n12978;
wire n12979;
wire n12980;
wire n12981;
wire n12982;
wire n12983;
wire n12984;
wire n12985;
wire n12986;
wire n12987;
wire n12988;
wire n12989;
wire n12990;
wire n12991;
wire n12992;
wire n12993;
wire n12994;
wire n12995;
wire n12996;
wire n12997;
wire n12998;
wire n12999;
wire n1300;
wire n13000;
wire n13001;
wire n13002;
wire n13003;
wire n13004;
wire n13005;
wire n13006;
wire n13007;
wire n13008;
wire n13009;
wire n13010;
wire n13011;
wire n13012;
wire n13013;
wire n13014;
wire n13015;
wire n13016;
wire n13017;
wire n13018;
wire n13019;
wire n13020;
wire n13021;
wire n13022;
wire n13023;
wire n13024;
wire n13025;
wire n13026;
wire n13027;
wire n13028;
wire n13029;
wire n13030;
wire n13031;
wire n13032;
wire n13033;
wire n13034;
wire n13035;
wire n13036;
wire n13037;
wire n13038;
wire n13039;
wire n13040;
wire n13041;
wire n13042;
wire n13043;
wire n13044;
wire n13045;
wire n13046;
wire n13047;
wire n13048;
wire n13049;
wire n1305;
wire n13050;
wire n13051;
wire n13052;
wire n13053;
wire n13054;
wire n13055;
wire n13056;
wire n13057;
wire n13058;
wire n13059;
wire n13060;
wire n13061;
wire n13062;
wire n13063;
wire n13064;
wire n13065;
wire n13066;
wire n13067;
wire n13068;
wire n13069;
wire n13070;
wire n13071;
wire n13072;
wire n13073;
wire n13074;
wire n13075;
wire n13076;
wire n13077;
wire n13078;
wire n13079;
wire n13080;
wire n13081;
wire n13082;
wire n13083;
wire n13084;
wire n13085;
wire n13086;
wire n13087;
wire n13088;
wire n13089;
wire n13090;
wire n13091;
wire n13092;
wire n13093;
wire n13094;
wire n13095;
wire n13096;
wire n13097;
wire n13098;
wire n13099;
wire n1310;
wire n13100;
wire n13101;
wire n13102;
wire n13103;
wire n13104;
wire n13105;
wire n13106;
wire n13107;
wire n13108;
wire n13109;
wire n13110;
wire n13111;
wire n13112;
wire n13113;
wire n13114;
wire n13115;
wire n13116;
wire n13117;
wire n13118;
wire n13119;
wire n13120;
wire n13121;
wire n13122;
wire n13123;
wire n13124;
wire n13125;
wire n13126;
wire n13127;
wire n13128;
wire n13129;
wire n13130;
wire n13131;
wire n13132;
wire n13133;
wire n13134;
wire n13135;
wire n13136;
wire n13137;
wire n13138;
wire n13139;
wire n13140;
wire n13141;
wire n13142;
wire n13143;
wire n13144;
wire n13145;
wire n13146;
wire n13147;
wire n13148;
wire n13149;
wire n1315;
wire n13150;
wire n13151;
wire n13152;
wire n13153;
wire n13154;
wire n13155;
wire n13156;
wire n13157;
wire n13158;
wire n13159;
wire n13160;
wire n13161;
wire n13162;
wire n13163;
wire n13164;
wire n13165;
wire n13166;
wire n13167;
wire n13168;
wire n13169;
wire n13170;
wire n13171;
wire n13172;
wire n13173;
wire n13174;
wire n13175;
wire n13176;
wire n13177;
wire n13178;
wire n13179;
wire n13180;
wire n13181;
wire n13182;
wire n13183;
wire n13184;
wire n13185;
wire n13186;
wire n13187;
wire n13188;
wire n13189;
wire n1319;
wire n13190;
wire n13191;
wire n13192;
wire n13193;
wire n13194;
wire n13195;
wire n13196;
wire n13197;
wire n13198;
wire n13199;
wire n13200;
wire n13201;
wire n13202;
wire n13203;
wire n13204;
wire n13205;
wire n13206;
wire n13207;
wire n13208;
wire n13209;
wire n13210;
wire n13211;
wire n13212;
wire n13213;
wire n13214;
wire n13215;
wire n13216;
wire n13217;
wire n13218;
wire n13219;
wire n13220;
wire n13221;
wire n13222;
wire n13223;
wire n13224;
wire n13225;
wire n13226;
wire n13227;
wire n13228;
wire n13229;
wire n13230;
wire n13231;
wire n13232;
wire n13233;
wire n13234;
wire n13235;
wire n13236;
wire n13237;
wire n13238;
wire n13239;
wire n1324;
wire n13240;
wire n13241;
wire n13242;
wire n13243;
wire n13244;
wire n13245;
wire n13246;
wire n13247;
wire n13248;
wire n13249;
wire n13250;
wire n13251;
wire n13252;
wire n13253;
wire n13254;
wire n13255;
wire n13256;
wire n13257;
wire n13258;
wire n13259;
wire n13260;
wire n13261;
wire n13262;
wire n13263;
wire n13264;
wire n13265;
wire n13266;
wire n13267;
wire n13268;
wire n13269;
wire n13270;
wire n13271;
wire n13272;
wire n13273;
wire n13274;
wire n13275;
wire n13276;
wire n13277;
wire n13278;
wire n13279;
wire n13280;
wire n13281;
wire n13282;
wire n13283;
wire n13284;
wire n13285;
wire n13286;
wire n13287;
wire n13288;
wire n13289;
wire n1329;
wire n13290;
wire n13291;
wire n13292;
wire n13293;
wire n13294;
wire n13295;
wire n13296;
wire n13297;
wire n13298;
wire n13299;
wire n13300;
wire n13301;
wire n13302;
wire n13303;
wire n13304;
wire n13305;
wire n13306;
wire n13307;
wire n13308;
wire n13309;
wire n13310;
wire n13311;
wire n13312;
wire n13313;
wire n13314;
wire n13315;
wire n13316;
wire n13317;
wire n13318;
wire n13319;
wire n13320;
wire n13321;
wire n13322;
wire n13323;
wire n13324;
wire n13325;
wire n13326;
wire n13327;
wire n13328;
wire n13329;
wire n13330;
wire n13331;
wire n13332;
wire n13333;
wire n13334;
wire n13335;
wire n13336;
wire n13337;
wire n13338;
wire n13339;
wire n1334;
wire n13340;
wire n13341;
wire n13342;
wire n13343;
wire n13344;
wire n13345;
wire n13346;
wire n13347;
wire n13348;
wire n13349;
wire n13350;
wire n13351;
wire n13352;
wire n13353;
wire n13354;
wire n13355;
wire n13356;
wire n13357;
wire n13358;
wire n13359;
wire n13360;
wire n13361;
wire n13362;
wire n13363;
wire n13364;
wire n13365;
wire n13366;
wire n13367;
wire n13368;
wire n13369;
wire n13370;
wire n13371;
wire n13372;
wire n13373;
wire n13374;
wire n13375;
wire n13376;
wire n13377;
wire n13378;
wire n13379;
wire n13380;
wire n13381;
wire n13382;
wire n13383;
wire n13384;
wire n13385;
wire n13386;
wire n13387;
wire n13388;
wire n13389;
wire n1339;
wire n13390;
wire n13391;
wire n13392;
wire n13393;
wire n13394;
wire n13395;
wire n13396;
wire n13397;
wire n13398;
wire n13399;
wire n13400;
wire n13401;
wire n13402;
wire n13403;
wire n13404;
wire n13405;
wire n13406;
wire n13407;
wire n13408;
wire n13409;
wire n13410;
wire n13411;
wire n13412;
wire n13413;
wire n13414;
wire n13415;
wire n13416;
wire n13417;
wire n13418;
wire n13419;
wire n13420;
wire n13421;
wire n13422;
wire n13423;
wire n13424;
wire n13425;
wire n13426;
wire n13427;
wire n13428;
wire n13429;
wire n13430;
wire n13431;
wire n13432;
wire n13433;
wire n13434;
wire n13435;
wire n13436;
wire n13437;
wire n13438;
wire n13439;
wire n1344;
wire n13440;
wire n13441;
wire n13442;
wire n13443;
wire n13444;
wire n13445;
wire n13446;
wire n13447;
wire n13448;
wire n13449;
wire n13450;
wire n13451;
wire n13452;
wire n13453;
wire n13454;
wire n13455;
wire n13456;
wire n13457;
wire n13458;
wire n13459;
wire n13460;
wire n13461;
wire n13462;
wire n13463;
wire n13464;
wire n13465;
wire n13466;
wire n13467;
wire n13468;
wire n13469;
wire n13470;
wire n13471;
wire n13472;
wire n13473;
wire n13474;
wire n13475;
wire n13476;
wire n13477;
wire n13478;
wire n13479;
wire n1348;
wire n13480;
wire n13481;
wire n13482;
wire n13483;
wire n13484;
wire n13485;
wire n13486;
wire n13487;
wire n13488;
wire n13489;
wire n13490;
wire n13491;
wire n13492;
wire n13493;
wire n13494;
wire n13495;
wire n13496;
wire n13497;
wire n13498;
wire n13499;
wire n13500;
wire n13501;
wire n13502;
wire n13503;
wire n13504;
wire n13505;
wire n13506;
wire n13507;
wire n13508;
wire n13509;
wire n13510;
wire n13511;
wire n13512;
wire n13513;
wire n13514;
wire n13515;
wire n13516;
wire n13517;
wire n13518;
wire n13519;
wire n13520;
wire n13521;
wire n13522;
wire n13523;
wire n13524;
wire n13525;
wire n13526;
wire n13527;
wire n13528;
wire n13529;
wire n1353;
wire n13530;
wire n13531;
wire n13532;
wire n13533;
wire n13534;
wire n13535;
wire n13536;
wire n13537;
wire n13538;
wire n13539;
wire n13540;
wire n13541;
wire n13542;
wire n13543;
wire n13544;
wire n13545;
wire n13546;
wire n13547;
wire n13548;
wire n13549;
wire n13550;
wire n13551;
wire n13552;
wire n13553;
wire n13554;
wire n13555;
wire n13556;
wire n13557;
wire n13558;
wire n13559;
wire n13560;
wire n13561;
wire n13562;
wire n13563;
wire n13564;
wire n13565;
wire n13566;
wire n13567;
wire n13568;
wire n13569;
wire n13570;
wire n13571;
wire n13572;
wire n13573;
wire n13574;
wire n13575;
wire n13576;
wire n13577;
wire n13578;
wire n13579;
wire n1358;
wire n13580;
wire n13581;
wire n13582;
wire n13583;
wire n13584;
wire n13585;
wire n13586;
wire n13587;
wire n13588;
wire n13589;
wire n13590;
wire n13591;
wire n13592;
wire n13593;
wire n13594;
wire n13595;
wire n13596;
wire n13597;
wire n13598;
wire n13599;
wire n13600;
wire n13601;
wire n13602;
wire n13603;
wire n13604;
wire n13605;
wire n13606;
wire n13607;
wire n13608;
wire n13609;
wire n13610;
wire n13611;
wire n13612;
wire n13613;
wire n13614;
wire n13615;
wire n13616;
wire n13617;
wire n13618;
wire n13619;
wire n13620;
wire n13621;
wire n13622;
wire n13623;
wire n13624;
wire n13625;
wire n13626;
wire n13627;
wire n13628;
wire n13629;
wire n1363;
wire n13630;
wire n13631;
wire n13632;
wire n13633;
wire n13634;
wire n13635;
wire n13636;
wire n13637;
wire n13638;
wire n13639;
wire n13640;
wire n13641;
wire n13642;
wire n13643;
wire n13644;
wire n13645;
wire n13646;
wire n13647;
wire n13648;
wire n13649;
wire n13650;
wire n13651;
wire n13652;
wire n13653;
wire n13654;
wire n13655;
wire n13656;
wire n13657;
wire n13658;
wire n13659;
wire n13660;
wire n13661;
wire n13662;
wire n13663;
wire n13664;
wire n13665;
wire n13666;
wire n13667;
wire n13668;
wire n13669;
wire n13670;
wire n13671;
wire n13672;
wire n13673;
wire n13674;
wire n13675;
wire n13676;
wire n13677;
wire n13678;
wire n13679;
wire n1368;
wire n13680;
wire n13681;
wire n13682;
wire n13683;
wire n13684;
wire n13685;
wire n13686;
wire n13687;
wire n13688;
wire n13689;
wire n13690;
wire n13691;
wire n13692;
wire n13693;
wire n13694;
wire n13695;
wire n13696;
wire n13697;
wire n13698;
wire n13699;
wire n13700;
wire n13701;
wire n13702;
wire n13703;
wire n13704;
wire n13705;
wire n13706;
wire n13707;
wire n13708;
wire n13709;
wire n13710;
wire n13711;
wire n13712;
wire n13713;
wire n13714;
wire n13715;
wire n13716;
wire n13717;
wire n13718;
wire n13719;
wire n13720;
wire n13721;
wire n13722;
wire n13723;
wire n13724;
wire n13725;
wire n13726;
wire n13727;
wire n13728;
wire n13729;
wire n1373;
wire n13730;
wire n13731;
wire n13732;
wire n13733;
wire n13734;
wire n13735;
wire n13736;
wire n13737;
wire n13738;
wire n13739;
wire n13740;
wire n13741;
wire n13742;
wire n13743;
wire n13744;
wire n13745;
wire n13746;
wire n13747;
wire n13748;
wire n13749;
wire n13750;
wire n13751;
wire n13752;
wire n13753;
wire n13754;
wire n13755;
wire n13756;
wire n13757;
wire n13758;
wire n13759;
wire n13760;
wire n13761;
wire n13762;
wire n13763;
wire n13764;
wire n13765;
wire n13766;
wire n13767;
wire n13768;
wire n13769;
wire n1377;
wire n13770;
wire n13771;
wire n13772;
wire n13773;
wire n13774;
wire n13775;
wire n13776;
wire n13777;
wire n13778;
wire n13779;
wire n13780;
wire n13781;
wire n13782;
wire n13783;
wire n13784;
wire n13785;
wire n13786;
wire n13787;
wire n13788;
wire n13789;
wire n13790;
wire n13791;
wire n13792;
wire n13793;
wire n13794;
wire n13795;
wire n13796;
wire n13797;
wire n13798;
wire n13799;
wire n13800;
wire n13801;
wire n13802;
wire n13803;
wire n13804;
wire n13805;
wire n13806;
wire n13807;
wire n13808;
wire n13809;
wire n13810;
wire n13811;
wire n13812;
wire n13813;
wire n13814;
wire n13815;
wire n13816;
wire n13817;
wire n13818;
wire n13819;
wire n1382;
wire n13820;
wire n13821;
wire n13822;
wire n13823;
wire n13824;
wire n13825;
wire n13826;
wire n13827;
wire n13828;
wire n13829;
wire n13830;
wire n13831;
wire n13832;
wire n13833;
wire n13834;
wire n13835;
wire n13836;
wire n13837;
wire n13838;
wire n13839;
wire n13840;
wire n13841;
wire n13842;
wire n13843;
wire n13844;
wire n13845;
wire n13846;
wire n13847;
wire n13848;
wire n13849;
wire n13850;
wire n13851;
wire n13852;
wire n13853;
wire n13854;
wire n13855;
wire n13856;
wire n13857;
wire n13858;
wire n13859;
wire n13860;
wire n13861;
wire n13862;
wire n13863;
wire n13864;
wire n13865;
wire n13866;
wire n13867;
wire n13868;
wire n13869;
wire n1387;
wire n13870;
wire n13871;
wire n13872;
wire n13873;
wire n13874;
wire n13875;
wire n13876;
wire n13877;
wire n13878;
wire n13879;
wire n13880;
wire n13881;
wire n13882;
wire n13883;
wire n13884;
wire n13885;
wire n13886;
wire n13887;
wire n13888;
wire n13889;
wire n13890;
wire n13891;
wire n13892;
wire n13893;
wire n13894;
wire n13895;
wire n13896;
wire n13897;
wire n13898;
wire n13899;
wire n13900;
wire n13901;
wire n13902;
wire n13903;
wire n13904;
wire n13905;
wire n13906;
wire n13907;
wire n13908;
wire n13909;
wire n13910;
wire n13911;
wire n13912;
wire n13913;
wire n13914;
wire n13915;
wire n13916;
wire n13917;
wire n13918;
wire n13919;
wire n1392;
wire n13920;
wire n13921;
wire n13922;
wire n13923;
wire n13924;
wire n13925;
wire n13926;
wire n13927;
wire n13928;
wire n13929;
wire n13930;
wire n13931;
wire n13932;
wire n13933;
wire n13934;
wire n13935;
wire n13936;
wire n13937;
wire n13938;
wire n13939;
wire n13940;
wire n13941;
wire n13942;
wire n13943;
wire n13944;
wire n13945;
wire n13946;
wire n13947;
wire n13948;
wire n13949;
wire n13950;
wire n13951;
wire n13952;
wire n13953;
wire n13954;
wire n13955;
wire n13956;
wire n13957;
wire n13958;
wire n13959;
wire n1396;
wire n13960;
wire n13961;
wire n13962;
wire n13963;
wire n13964;
wire n13965;
wire n13966;
wire n13967;
wire n13968;
wire n13969;
wire n13970;
wire n13971;
wire n13972;
wire n13973;
wire n13974;
wire n13975;
wire n13976;
wire n13977;
wire n13978;
wire n13979;
wire n13980;
wire n13981;
wire n13982;
wire n13983;
wire n13984;
wire n13985;
wire n13986;
wire n13987;
wire n13988;
wire n13989;
wire n13990;
wire n13991;
wire n13992;
wire n13993;
wire n13994;
wire n13995;
wire n13996;
wire n13997;
wire n13998;
wire n13999;
wire n14000;
wire n14001;
wire n14002;
wire n14003;
wire n14004;
wire n14005;
wire n14006;
wire n14007;
wire n14008;
wire n14009;
wire n1401;
wire n14010;
wire n14011;
wire n14012;
wire n14013;
wire n14014;
wire n14015;
wire n14016;
wire n14017;
wire n14018;
wire n14019;
wire n14020;
wire n14021;
wire n14022;
wire n14023;
wire n14024;
wire n14025;
wire n14026;
wire n14027;
wire n14028;
wire n14029;
wire n14030;
wire n14031;
wire n14032;
wire n14033;
wire n14034;
wire n14035;
wire n14036;
wire n14037;
wire n14038;
wire n14039;
wire n14040;
wire n14041;
wire n14042;
wire n14043;
wire n14044;
wire n14045;
wire n14046;
wire n14047;
wire n14048;
wire n14049;
wire n14050;
wire n14051;
wire n14052;
wire n14053;
wire n14054;
wire n14055;
wire n14056;
wire n14057;
wire n14058;
wire n14059;
wire n1406;
wire n14060;
wire n14061;
wire n14062;
wire n14063;
wire n14064;
wire n14065;
wire n14066;
wire n14067;
wire n14068;
wire n14069;
wire n14070;
wire n14071;
wire n14072;
wire n14073;
wire n14074;
wire n14075;
wire n14076;
wire n14077;
wire n14078;
wire n14079;
wire n14080;
wire n14081;
wire n14082;
wire n14083;
wire n14084;
wire n14085;
wire n14086;
wire n14087;
wire n14088;
wire n14089;
wire n14090;
wire n14091;
wire n14092;
wire n14093;
wire n14094;
wire n14095;
wire n14096;
wire n14097;
wire n14098;
wire n14099;
wire n14100;
wire n14101;
wire n14102;
wire n14103;
wire n14104;
wire n14105;
wire n14106;
wire n14107;
wire n14108;
wire n14109;
wire n1411;
wire n14110;
wire n14111;
wire n14112;
wire n14113;
wire n14114;
wire n14115;
wire n14116;
wire n14117;
wire n14118;
wire n14119;
wire n14120;
wire n14121;
wire n14122;
wire n14123;
wire n14124;
wire n14125;
wire n14126;
wire n14127;
wire n14128;
wire n14129;
wire n14130;
wire n14131;
wire n14132;
wire n14133;
wire n14134;
wire n14135;
wire n14136;
wire n14137;
wire n14138;
wire n14139;
wire n14140;
wire n14141;
wire n14142;
wire n14143;
wire n14144;
wire n14145;
wire n14146;
wire n14147;
wire n14148;
wire n14149;
wire n14150;
wire n14151;
wire n14152;
wire n14153;
wire n14154;
wire n14155;
wire n14156;
wire n14157;
wire n14158;
wire n14159;
wire n1416;
wire n14160;
wire n14161;
wire n14162;
wire n14163;
wire n14164;
wire n14165;
wire n14166;
wire n14167;
wire n14168;
wire n14169;
wire n14170;
wire n14171;
wire n14172;
wire n14173;
wire n14174;
wire n14175;
wire n14176;
wire n14177;
wire n14178;
wire n14179;
wire n14180;
wire n14181;
wire n14182;
wire n14183;
wire n14184;
wire n14185;
wire n14186;
wire n14187;
wire n14188;
wire n14189;
wire n14190;
wire n14191;
wire n14192;
wire n14193;
wire n14194;
wire n14195;
wire n14196;
wire n14197;
wire n14198;
wire n14199;
wire n14200;
wire n14201;
wire n14202;
wire n14203;
wire n14204;
wire n14205;
wire n14206;
wire n14207;
wire n14208;
wire n14209;
wire n1421;
wire n14210;
wire n14211;
wire n14212;
wire n14213;
wire n14214;
wire n14215;
wire n14216;
wire n14217;
wire n14218;
wire n14219;
wire n14220;
wire n14221;
wire n14222;
wire n14223;
wire n14224;
wire n14225;
wire n14226;
wire n14227;
wire n14228;
wire n14229;
wire n14230;
wire n14231;
wire n14232;
wire n14233;
wire n14234;
wire n14235;
wire n14236;
wire n14237;
wire n14238;
wire n14239;
wire n14240;
wire n14241;
wire n14242;
wire n14243;
wire n14244;
wire n14245;
wire n14246;
wire n14247;
wire n14248;
wire n14249;
wire n14250;
wire n14251;
wire n14252;
wire n14253;
wire n14254;
wire n14255;
wire n14256;
wire n14257;
wire n14258;
wire n14259;
wire n1426;
wire n14260;
wire n14261;
wire n14262;
wire n14263;
wire n14264;
wire n14265;
wire n14266;
wire n14267;
wire n14268;
wire n14269;
wire n14270;
wire n14271;
wire n14272;
wire n14273;
wire n14274;
wire n14275;
wire n14276;
wire n14277;
wire n14278;
wire n14279;
wire n14280;
wire n14281;
wire n14282;
wire n14283;
wire n14284;
wire n14285;
wire n14286;
wire n14287;
wire n14288;
wire n14289;
wire n14290;
wire n14291;
wire n14292;
wire n14293;
wire n14294;
wire n14295;
wire n14296;
wire n14297;
wire n14298;
wire n14299;
wire n14300;
wire n14301;
wire n14302;
wire n14303;
wire n14304;
wire n14305;
wire n14306;
wire n14307;
wire n14308;
wire n14309;
wire n1431;
wire n14310;
wire n14311;
wire n14312;
wire n14313;
wire n14314;
wire n14315;
wire n14316;
wire n14317;
wire n14318;
wire n14319;
wire n14320;
wire n14321;
wire n14322;
wire n14323;
wire n14324;
wire n14325;
wire n14326;
wire n14327;
wire n14328;
wire n14329;
wire n14330;
wire n14331;
wire n14332;
wire n14333;
wire n14334;
wire n14335;
wire n14336;
wire n14337;
wire n14338;
wire n14339;
wire n14340;
wire n14341;
wire n14343;
wire n14344;
wire n14345;
wire n14347;
wire n14349;
wire n14350;
wire n14351;
wire n14352;
wire n14353;
wire n14354;
wire n14355;
wire n14356;
wire n14357;
wire n14358;
wire n14359;
wire n1436;
wire n14360;
wire n14361;
wire n14362;
wire n14363;
wire n14364;
wire n14365;
wire n14366;
wire n14367;
wire n14368;
wire n14369;
wire n14370;
wire n14371;
wire n14372;
wire n14373;
wire n14374;
wire n14375;
wire n14376;
wire n14377;
wire n14378;
wire n14379;
wire n14380;
wire n14381;
wire n14382;
wire n14383;
wire n14384;
wire n14385;
wire n14386;
wire n14387;
wire n14388;
wire n14389;
wire n14390;
wire n14391;
wire n14392;
wire n14393;
wire n14394;
wire n14395;
wire n14396;
wire n14397;
wire n14398;
wire n14399;
wire n14400;
wire n14401;
wire n14402;
wire n14403;
wire n14404;
wire n14405;
wire n14406;
wire n14407;
wire n14408;
wire n14409;
wire n1441;
wire n14410;
wire n14411;
wire n14412;
wire n14413;
wire n14414;
wire n14415;
wire n14416;
wire n14417;
wire n14418;
wire n14419;
wire n14420;
wire n14421;
wire n14422;
wire n14423;
wire n14424;
wire n14425;
wire n14426;
wire n14427;
wire n14428;
wire n14429;
wire n14430;
wire n14431;
wire n14432;
wire n14433;
wire n14434;
wire n14435;
wire n14436;
wire n14437;
wire n14438;
wire n14439;
wire n14440;
wire n14441;
wire n14442;
wire n14443;
wire n14444;
wire n14445;
wire n14446;
wire n14447;
wire n14448;
wire n14449;
wire n14450;
wire n14451;
wire n14452;
wire n14453;
wire n14454;
wire n14455;
wire n14456;
wire n14457;
wire n14458;
wire n14459;
wire n1446;
wire n14460;
wire n14461;
wire n14462;
wire n14463;
wire n14464;
wire n14465;
wire n14466;
wire n14467;
wire n14468;
wire n14469;
wire n14470;
wire n14471;
wire n14472;
wire n14473;
wire n14474;
wire n14475;
wire n14476;
wire n14477;
wire n14478;
wire n14479;
wire n14480;
wire n14481;
wire n14482;
wire n14483;
wire n14484;
wire n14485;
wire n14486;
wire n14487;
wire n14488;
wire n14489;
wire n14490;
wire n14491;
wire n14492;
wire n14493;
wire n14494;
wire n14495;
wire n14496;
wire n14497;
wire n14498;
wire n14499;
wire n14500;
wire n14501;
wire n14502;
wire n14503;
wire n14504;
wire n14505;
wire n14506;
wire n14507;
wire n14508;
wire n14509;
wire n1451;
wire n14510;
wire n14511;
wire n14512;
wire n14513;
wire n14514;
wire n14515;
wire n14516;
wire n14517;
wire n14518;
wire n14519;
wire n14520;
wire n14521;
wire n14522;
wire n14523;
wire n14524;
wire n14525;
wire n14526;
wire n14527;
wire n14528;
wire n14529;
wire n14530;
wire n14531;
wire n14532;
wire n14533;
wire n14534;
wire n14535;
wire n14536;
wire n14537;
wire n14538;
wire n14539;
wire n14540;
wire n14541;
wire n14542;
wire n14543;
wire n14544;
wire n14545;
wire n14546;
wire n14547;
wire n14548;
wire n14549;
wire n14550;
wire n14551;
wire n14552;
wire n14553;
wire n14554;
wire n14555;
wire n14556;
wire n14557;
wire n14558;
wire n14559;
wire n1456;
wire n14560;
wire n14561;
wire n14562;
wire n14563;
wire n14564;
wire n14565;
wire n14566;
wire n14567;
wire n14568;
wire n14569;
wire n14570;
wire n14571;
wire n14572;
wire n14573;
wire n14574;
wire n14575;
wire n14576;
wire n14577;
wire n14578;
wire n14579;
wire n14580;
wire n14581;
wire n14582;
wire n14583;
wire n14584;
wire n14585;
wire n14586;
wire n14587;
wire n14588;
wire n14589;
wire n14590;
wire n14591;
wire n14592;
wire n14593;
wire n14594;
wire n14595;
wire n14596;
wire n14597;
wire n14598;
wire n14599;
wire n14600;
wire n14601;
wire n14602;
wire n14603;
wire n14604;
wire n14605;
wire n14606;
wire n14607;
wire n14608;
wire n14609;
wire n1461;
wire n14610;
wire n14611;
wire n14612;
wire n14613;
wire n14614;
wire n14615;
wire n14616;
wire n14617;
wire n14618;
wire n14619;
wire n14620;
wire n14621;
wire n14622;
wire n14623;
wire n14624;
wire n14625;
wire n14626;
wire n14627;
wire n14628;
wire n14629;
wire n14630;
wire n14631;
wire n14632;
wire n14633;
wire n14634;
wire n14635;
wire n14636;
wire n14637;
wire n14638;
wire n14639;
wire n14640;
wire n14641;
wire n14642;
wire n14643;
wire n14644;
wire n14645;
wire n14646;
wire n14647;
wire n14648;
wire n14649;
wire n14650;
wire n14651;
wire n14652;
wire n14653;
wire n14654;
wire n14655;
wire n14656;
wire n14657;
wire n14658;
wire n14659;
wire n1466;
wire n14660;
wire n14661;
wire n14662;
wire n14663;
wire n14664;
wire n14665;
wire n14666;
wire n14667;
wire n14668;
wire n14669;
wire n14670;
wire n14671;
wire n14672;
wire n14673;
wire n14674;
wire n14675;
wire n14676;
wire n14677;
wire n14678;
wire n14679;
wire n14680;
wire n14681;
wire n14682;
wire n14683;
wire n14684;
wire n14685;
wire n14686;
wire n14687;
wire n14688;
wire n14689;
wire n14690;
wire n14691;
wire n14692;
wire n14693;
wire n14694;
wire n14695;
wire n14696;
wire n14697;
wire n14698;
wire n14699;
wire n14700;
wire n14701;
wire n14702;
wire n14703;
wire n14704;
wire n14705;
wire n14706;
wire n14707;
wire n14708;
wire n14709;
wire n1471;
wire n14710;
wire n14711;
wire n14712;
wire n14713;
wire n14714;
wire n14715;
wire n14716;
wire n14717;
wire n14718;
wire n14719;
wire n14720;
wire n14721;
wire n14722;
wire n14723;
wire n14724;
wire n14725;
wire n14726;
wire n14727;
wire n14728;
wire n14729;
wire n14730;
wire n14731;
wire n14732;
wire n14733;
wire n14734;
wire n14735;
wire n14736;
wire n14737;
wire n14738;
wire n14739;
wire n14740;
wire n14741;
wire n14742;
wire n14743;
wire n14744;
wire n14745;
wire n14746;
wire n14747;
wire n14748;
wire n14749;
wire n14750;
wire n14751;
wire n14752;
wire n14753;
wire n14754;
wire n14755;
wire n14756;
wire n14757;
wire n14758;
wire n14759;
wire n1476;
wire n14760;
wire n14761;
wire n14762;
wire n14763;
wire n14764;
wire n14765;
wire n14766;
wire n14767;
wire n14768;
wire n14769;
wire n14770;
wire n14771;
wire n14772;
wire n14773;
wire n14774;
wire n14775;
wire n14776;
wire n14777;
wire n14778;
wire n14779;
wire n14780;
wire n14781;
wire n14782;
wire n14783;
wire n14784;
wire n14785;
wire n14786;
wire n14787;
wire n14788;
wire n14789;
wire n14790;
wire n14791;
wire n14792;
wire n14793;
wire n14794;
wire n14795;
wire n14796;
wire n14797;
wire n14798;
wire n14799;
wire n14800;
wire n14801;
wire n14802;
wire n14803;
wire n14804;
wire n14805;
wire n14806;
wire n14807;
wire n14808;
wire n14809;
wire n1481;
wire n14810;
wire n14811;
wire n14812;
wire n14813;
wire n14814;
wire n14815;
wire n14816;
wire n14817;
wire n14818;
wire n14819;
wire n14820;
wire n14821;
wire n14822;
wire n14823;
wire n14824;
wire n14825;
wire n14826;
wire n14827;
wire n14828;
wire n14829;
wire n14830;
wire n14831;
wire n14832;
wire n14833;
wire n14834;
wire n14835;
wire n14836;
wire n14837;
wire n14838;
wire n14839;
wire n14840;
wire n14841;
wire n14842;
wire n14843;
wire n14844;
wire n14845;
wire n14846;
wire n14847;
wire n14848;
wire n14849;
wire n14850;
wire n14851;
wire n14852;
wire n14853;
wire n14854;
wire n14855;
wire n14856;
wire n14857;
wire n14858;
wire n14859;
wire n1486;
wire n14860;
wire n14861;
wire n14862;
wire n14863;
wire n14864;
wire n14865;
wire n14866;
wire n14867;
wire n14868;
wire n14869;
wire n14870;
wire n14871;
wire n14872;
wire n14873;
wire n14874;
wire n14875;
wire n14876;
wire n14877;
wire n14878;
wire n14879;
wire n14880;
wire n14881;
wire n14882;
wire n14883;
wire n14884;
wire n14885;
wire n14886;
wire n14887;
wire n14888;
wire n14889;
wire n14890;
wire n14891;
wire n14892;
wire n14893;
wire n14894;
wire n14895;
wire n14896;
wire n14897;
wire n14898;
wire n14899;
wire n14900;
wire n14901;
wire n14902;
wire n14903;
wire n14904;
wire n14905;
wire n14906;
wire n14907;
wire n14908;
wire n14909;
wire n1491;
wire n14910;
wire n14911;
wire n14912;
wire n14913;
wire n14914;
wire n14915;
wire n14916;
wire n14917;
wire n14918;
wire n14919;
wire n14920;
wire n14921;
wire n14922;
wire n14923;
wire n14924;
wire n14925;
wire n14926;
wire n14927;
wire n14928;
wire n14929;
wire n14930;
wire n14931;
wire n14932;
wire n14933;
wire n14934;
wire n14935;
wire n14936;
wire n14937;
wire n14938;
wire n14939;
wire n14940;
wire n14941;
wire n14942;
wire n14943;
wire n14944;
wire n14945;
wire n14946;
wire n14947;
wire n14948;
wire n14949;
wire n14950;
wire n14951;
wire n14952;
wire n14953;
wire n14954;
wire n14955;
wire n14956;
wire n14957;
wire n14958;
wire n14959;
wire n1496;
wire n14960;
wire n14961;
wire n14962;
wire n14963;
wire n14964;
wire n14965;
wire n14966;
wire n14967;
wire n14968;
wire n14969;
wire n14970;
wire n14971;
wire n14972;
wire n14973;
wire n14974;
wire n14975;
wire n14976;
wire n14977;
wire n14978;
wire n14979;
wire n14980;
wire n14981;
wire n14982;
wire n14983;
wire n14984;
wire n14985;
wire n14986;
wire n14987;
wire n14988;
wire n14989;
wire n14990;
wire n14991;
wire n14992;
wire n14993;
wire n14994;
wire n14995;
wire n14996;
wire n14997;
wire n14998;
wire n14999;
wire n15000;
wire n15001;
wire n15002;
wire n15003;
wire n15004;
wire n15005;
wire n15006;
wire n15007;
wire n15008;
wire n15009;
wire n1501;
wire n15010;
wire n15011;
wire n15012;
wire n15013;
wire n15014;
wire n15015;
wire n15016;
wire n15017;
wire n15018;
wire n15019;
wire n15020;
wire n15021;
wire n15022;
wire n15023;
wire n15024;
wire n15025;
wire n15026;
wire n15027;
wire n15028;
wire n15029;
wire n15030;
wire n15031;
wire n15032;
wire n15033;
wire n15034;
wire n15035;
wire n15036;
wire n15037;
wire n15038;
wire n15039;
wire n15040;
wire n15041;
wire n15042;
wire n15043;
wire n15044;
wire n15045;
wire n15046;
wire n15047;
wire n15048;
wire n15049;
wire n15050;
wire n15051;
wire n15052;
wire n15053;
wire n15054;
wire n15055;
wire n15056;
wire n15057;
wire n15058;
wire n15059;
wire n1506;
wire n15060;
wire n15061;
wire n15062;
wire n15063;
wire n15064;
wire n15065;
wire n15066;
wire n15067;
wire n15068;
wire n15069;
wire n15070;
wire n15071;
wire n15072;
wire n15073;
wire n15074;
wire n15075;
wire n15076;
wire n15077;
wire n15078;
wire n15079;
wire n15080;
wire n15081;
wire n15082;
wire n15083;
wire n15084;
wire n15085;
wire n15086;
wire n15087;
wire n15088;
wire n15089;
wire n15090;
wire n15091;
wire n15092;
wire n15093;
wire n15094;
wire n15095;
wire n15096;
wire n15097;
wire n15098;
wire n15099;
wire n15100;
wire n15101;
wire n15102;
wire n15103;
wire n15104;
wire n15105;
wire n15106;
wire n15107;
wire n15108;
wire n15109;
wire n1511;
wire n15110;
wire n15111;
wire n15112;
wire n15113;
wire n15114;
wire n15115;
wire n15116;
wire n15117;
wire n15118;
wire n15119;
wire n15120;
wire n15121;
wire n15122;
wire n15123;
wire n15124;
wire n15125;
wire n15126;
wire n15127;
wire n15128;
wire n15129;
wire n15130;
wire n15131;
wire n15132;
wire n15133;
wire n15134;
wire n15135;
wire n15136;
wire n15137;
wire n15138;
wire n15139;
wire n15140;
wire n15141;
wire n15142;
wire n15143;
wire n15144;
wire n15145;
wire n15146;
wire n15147;
wire n15148;
wire n15149;
wire n15150;
wire n15151;
wire n15152;
wire n15153;
wire n15154;
wire n15155;
wire n15156;
wire n15157;
wire n15158;
wire n15159;
wire n1516;
wire n15160;
wire n15161;
wire n15162;
wire n15163;
wire n15164;
wire n15165;
wire n15166;
wire n15167;
wire n15168;
wire n15169;
wire n15170;
wire n15171;
wire n15172;
wire n15173;
wire n15174;
wire n15175;
wire n15176;
wire n15177;
wire n15178;
wire n15179;
wire n15180;
wire n15181;
wire n15182;
wire n15183;
wire n15184;
wire n15185;
wire n15186;
wire n15187;
wire n15188;
wire n15189;
wire n15190;
wire n15191;
wire n15192;
wire n15193;
wire n15194;
wire n15195;
wire n15196;
wire n15197;
wire n15198;
wire n15199;
wire n15200;
wire n15201;
wire n15202;
wire n15203;
wire n15204;
wire n15205;
wire n15206;
wire n15207;
wire n15208;
wire n15209;
wire n1521;
wire n15210;
wire n15211;
wire n15212;
wire n15213;
wire n15214;
wire n15215;
wire n15216;
wire n15217;
wire n15218;
wire n15219;
wire n15220;
wire n15221;
wire n15222;
wire n15223;
wire n15224;
wire n15225;
wire n15226;
wire n15227;
wire n15228;
wire n15229;
wire n15230;
wire n15231;
wire n15232;
wire n15233;
wire n15234;
wire n15235;
wire n15236;
wire n15237;
wire n15238;
wire n15239;
wire n15240;
wire n15241;
wire n15242;
wire n15243;
wire n15244;
wire n15245;
wire n15246;
wire n15247;
wire n15248;
wire n15249;
wire n15250;
wire n15251;
wire n15252;
wire n15253;
wire n15254;
wire n15255;
wire n15256;
wire n15257;
wire n15258;
wire n15259;
wire n1526;
wire n15260;
wire n15261;
wire n15262;
wire n15263;
wire n15264;
wire n15265;
wire n15266;
wire n15267;
wire n15268;
wire n15269;
wire n15270;
wire n15271;
wire n15272;
wire n15273;
wire n15274;
wire n15275;
wire n15276;
wire n15277;
wire n15278;
wire n15279;
wire n15280;
wire n15281;
wire n15282;
wire n15283;
wire n15284;
wire n15285;
wire n15286;
wire n15287;
wire n15288;
wire n15289;
wire n15290;
wire n15291;
wire n15292;
wire n15293;
wire n15294;
wire n15295;
wire n15296;
wire n15297;
wire n15298;
wire n15299;
wire n15300;
wire n15301;
wire n15302;
wire n15303;
wire n15304;
wire n15305;
wire n15306;
wire n15307;
wire n15308;
wire n15309;
wire n1531;
wire n15310;
wire n15311;
wire n15312;
wire n15313;
wire n15314;
wire n15315;
wire n15316;
wire n15317;
wire n15318;
wire n15319;
wire n15320;
wire n15321;
wire n15322;
wire n15323;
wire n15324;
wire n15325;
wire n15326;
wire n15327;
wire n15328;
wire n15329;
wire n15330;
wire n15331;
wire n15332;
wire n15333;
wire n15334;
wire n15335;
wire n15336;
wire n15337;
wire n15338;
wire n15339;
wire n15340;
wire n15341;
wire n15342;
wire n15343;
wire n15344;
wire n15345;
wire n15346;
wire n15347;
wire n15348;
wire n15349;
wire n15350;
wire n15351;
wire n15352;
wire n15353;
wire n15354;
wire n15355;
wire n15356;
wire n15357;
wire n15358;
wire n15359;
wire n1536;
wire n15360;
wire n15361;
wire n15362;
wire n15363;
wire n15364;
wire n15365;
wire n15366;
wire n15367;
wire n15368;
wire n15369;
wire n15370;
wire n15371;
wire n15372;
wire n15373;
wire n15374;
wire n15375;
wire n15376;
wire n15377;
wire n15378;
wire n15379;
wire n15380;
wire n15381;
wire n15382;
wire n15383;
wire n15384;
wire n15385;
wire n15386;
wire n15387;
wire n15388;
wire n15389;
wire n15390;
wire n15391;
wire n15392;
wire n15393;
wire n15394;
wire n15395;
wire n15396;
wire n15397;
wire n15398;
wire n15399;
wire n1540;
wire n15400;
wire n15401;
wire n15402;
wire n15403;
wire n15404;
wire n15405;
wire n15406;
wire n15407;
wire n15408;
wire n15409;
wire n15410;
wire n15411;
wire n15412;
wire n15413;
wire n15414;
wire n15415;
wire n15416;
wire n15417;
wire n15418;
wire n15419;
wire n15420;
wire n15421;
wire n15422;
wire n15423;
wire n15424;
wire n15425;
wire n15426;
wire n15427;
wire n15428;
wire n15429;
wire n15430;
wire n15431;
wire n15432;
wire n15433;
wire n15434;
wire n15435;
wire n15436;
wire n15437;
wire n15438;
wire n15439;
wire n15440;
wire n15441;
wire n15442;
wire n15443;
wire n15444;
wire n15445;
wire n15446;
wire n15447;
wire n15448;
wire n15449;
wire n1545;
wire n15450;
wire n15451;
wire n15452;
wire n15453;
wire n15454;
wire n15455;
wire n15456;
wire n15457;
wire n15458;
wire n15459;
wire n15460;
wire n15461;
wire n15462;
wire n15463;
wire n15464;
wire n15465;
wire n15466;
wire n15467;
wire n15468;
wire n15469;
wire n15470;
wire n15471;
wire n15472;
wire n15473;
wire n15474;
wire n15475;
wire n15476;
wire n15477;
wire n15478;
wire n15479;
wire n15480;
wire n15481;
wire n15482;
wire n15483;
wire n15484;
wire n15485;
wire n15486;
wire n15487;
wire n15488;
wire n15489;
wire n15490;
wire n15491;
wire n15492;
wire n15493;
wire n15494;
wire n15495;
wire n15496;
wire n15497;
wire n15498;
wire n15499;
wire n1550;
wire n15500;
wire n15501;
wire n15502;
wire n15503;
wire n15504;
wire n15505;
wire n15506;
wire n15507;
wire n15508;
wire n15509;
wire n15510;
wire n15511;
wire n15512;
wire n15513;
wire n15514;
wire n15515;
wire n15516;
wire n15517;
wire n15518;
wire n15519;
wire n15520;
wire n15521;
wire n15522;
wire n15523;
wire n15524;
wire n15525;
wire n15526;
wire n15527;
wire n15528;
wire n15529;
wire n15530;
wire n15531;
wire n15532;
wire n15533;
wire n15534;
wire n15535;
wire n15536;
wire n15537;
wire n15538;
wire n15539;
wire n15540;
wire n15541;
wire n15542;
wire n15543;
wire n15544;
wire n15545;
wire n15546;
wire n15547;
wire n15548;
wire n15549;
wire n1555;
wire n15550;
wire n15551;
wire n15552;
wire n15553;
wire n15554;
wire n15555;
wire n15556;
wire n15557;
wire n15558;
wire n15559;
wire n15560;
wire n15561;
wire n15562;
wire n15563;
wire n15564;
wire n15565;
wire n15566;
wire n15567;
wire n15568;
wire n15569;
wire n15570;
wire n15571;
wire n15572;
wire n15573;
wire n15574;
wire n15575;
wire n15576;
wire n15577;
wire n15578;
wire n15579;
wire n15580;
wire n15581;
wire n15582;
wire n15583;
wire n15584;
wire n15585;
wire n15586;
wire n15587;
wire n15588;
wire n15589;
wire n15590;
wire n15591;
wire n15592;
wire n15593;
wire n15594;
wire n15595;
wire n15596;
wire n15597;
wire n15598;
wire n15599;
wire n1560;
wire n15600;
wire n15601;
wire n15602;
wire n15603;
wire n15604;
wire n15605;
wire n15606;
wire n15607;
wire n15608;
wire n15609;
wire n15610;
wire n15611;
wire n15612;
wire n15613;
wire n15614;
wire n15615;
wire n15616;
wire n15617;
wire n15618;
wire n15619;
wire n15620;
wire n15621;
wire n15622;
wire n15623;
wire n15624;
wire n15625;
wire n15626;
wire n15627;
wire n15628;
wire n15629;
wire n15630;
wire n15631;
wire n15632;
wire n15633;
wire n15634;
wire n15635;
wire n15636;
wire n15637;
wire n15638;
wire n15639;
wire n15640;
wire n15641;
wire n15642;
wire n15643;
wire n15644;
wire n15645;
wire n15646;
wire n15647;
wire n15648;
wire n15649;
wire n1565;
wire n15650;
wire n15651;
wire n15652;
wire n15653;
wire n15654;
wire n15655;
wire n15656;
wire n15657;
wire n15658;
wire n15659;
wire n15660;
wire n15661;
wire n15662;
wire n15663;
wire n15664;
wire n15665;
wire n15666;
wire n15667;
wire n15668;
wire n15669;
wire n15670;
wire n15671;
wire n15672;
wire n15673;
wire n15674;
wire n15675;
wire n15676;
wire n15677;
wire n15678;
wire n15679;
wire n15680;
wire n15681;
wire n15682;
wire n15683;
wire n15684;
wire n15685;
wire n15686;
wire n15687;
wire n15688;
wire n15689;
wire n15690;
wire n15691;
wire n15692;
wire n15693;
wire n15694;
wire n15695;
wire n15696;
wire n15697;
wire n15698;
wire n15699;
wire n1570;
wire n15700;
wire n15701;
wire n15702;
wire n15703;
wire n15704;
wire n15705;
wire n15706;
wire n15707;
wire n15708;
wire n15709;
wire n15710;
wire n15711;
wire n15712;
wire n15713;
wire n15714;
wire n15715;
wire n15716;
wire n15717;
wire n15718;
wire n15719;
wire n15720;
wire n15721;
wire n15722;
wire n15723;
wire n15724;
wire n15725;
wire n15726;
wire n15727;
wire n15728;
wire n15729;
wire n15730;
wire n15731;
wire n15732;
wire n15733;
wire n15734;
wire n15735;
wire n15736;
wire n15737;
wire n15738;
wire n15739;
wire n15740;
wire n15741;
wire n15742;
wire n15743;
wire n15744;
wire n15745;
wire n15746;
wire n15747;
wire n15748;
wire n15749;
wire n1575;
wire n15750;
wire n15751;
wire n15752;
wire n15753;
wire n15754;
wire n15755;
wire n15756;
wire n15757;
wire n15758;
wire n15759;
wire n15760;
wire n15761;
wire n15762;
wire n15763;
wire n15764;
wire n15765;
wire n15766;
wire n15767;
wire n15768;
wire n15769;
wire n15770;
wire n15771;
wire n15772;
wire n15773;
wire n15774;
wire n15775;
wire n15776;
wire n15777;
wire n15778;
wire n15779;
wire n15780;
wire n15781;
wire n15782;
wire n15783;
wire n15784;
wire n15785;
wire n15786;
wire n15787;
wire n15788;
wire n15789;
wire n15790;
wire n15791;
wire n15792;
wire n15793;
wire n15794;
wire n15795;
wire n15796;
wire n15797;
wire n15798;
wire n15799;
wire n1580;
wire n15800;
wire n15801;
wire n15802;
wire n15803;
wire n15804;
wire n15805;
wire n15806;
wire n15807;
wire n15808;
wire n15809;
wire n15810;
wire n15811;
wire n15812;
wire n15813;
wire n15814;
wire n15815;
wire n15816;
wire n15817;
wire n15818;
wire n15819;
wire n15820;
wire n15821;
wire n15822;
wire n15823;
wire n15824;
wire n15825;
wire n15826;
wire n15827;
wire n15828;
wire n15829;
wire n15830;
wire n15831;
wire n15832;
wire n15833;
wire n15834;
wire n15835;
wire n15836;
wire n15837;
wire n15838;
wire n15839;
wire n15840;
wire n15841;
wire n15842;
wire n15843;
wire n15844;
wire n15845;
wire n15846;
wire n15847;
wire n15848;
wire n15849;
wire n1585;
wire n15850;
wire n15851;
wire n15852;
wire n15853;
wire n15854;
wire n15855;
wire n15856;
wire n15857;
wire n15858;
wire n15859;
wire n15860;
wire n15861;
wire n15862;
wire n15863;
wire n15864;
wire n15865;
wire n15866;
wire n15867;
wire n15868;
wire n15869;
wire n15870;
wire n15871;
wire n15872;
wire n15873;
wire n15874;
wire n15875;
wire n15876;
wire n15877;
wire n15878;
wire n15879;
wire n15880;
wire n15881;
wire n15882;
wire n15883;
wire n15884;
wire n15885;
wire n15886;
wire n15887;
wire n15888;
wire n15889;
wire n15890;
wire n15891;
wire n15892;
wire n15893;
wire n15894;
wire n15895;
wire n15896;
wire n15897;
wire n15898;
wire n15899;
wire n1590;
wire n15900;
wire n15901;
wire n15902;
wire n15903;
wire n15904;
wire n15905;
wire n15906;
wire n15907;
wire n15908;
wire n15909;
wire n15910;
wire n15911;
wire n15912;
wire n15913;
wire n15914;
wire n15915;
wire n15916;
wire n15917;
wire n15918;
wire n15919;
wire n15920;
wire n15921;
wire n15922;
wire n15923;
wire n15924;
wire n15925;
wire n15926;
wire n15927;
wire n15928;
wire n15929;
wire n15930;
wire n15931;
wire n15932;
wire n15933;
wire n15934;
wire n15935;
wire n15936;
wire n15937;
wire n15938;
wire n15939;
wire n15940;
wire n15941;
wire n15942;
wire n15943;
wire n15944;
wire n15945;
wire n15946;
wire n15947;
wire n15948;
wire n15949;
wire n1595;
wire n15950;
wire n15951;
wire n15952;
wire n15953;
wire n15954;
wire n15955;
wire n15956;
wire n15957;
wire n15958;
wire n15959;
wire n15960;
wire n15961;
wire n15962;
wire n15963;
wire n15964;
wire n15965;
wire n15966;
wire n15967;
wire n15968;
wire n15969;
wire n15970;
wire n15971;
wire n15972;
wire n15973;
wire n15974;
wire n15975;
wire n15976;
wire n15977;
wire n15978;
wire n15979;
wire n15980;
wire n15981;
wire n15982;
wire n15983;
wire n15984;
wire n15985;
wire n15986;
wire n15987;
wire n15988;
wire n15989;
wire n15990;
wire n15991;
wire n15992;
wire n15993;
wire n15994;
wire n15995;
wire n15996;
wire n15997;
wire n15998;
wire n15999;
wire n1600;
wire n16000;
wire n16001;
wire n16002;
wire n16003;
wire n16004;
wire n16005;
wire n16006;
wire n16007;
wire n16008;
wire n16009;
wire n16010;
wire n16011;
wire n16012;
wire n16013;
wire n16014;
wire n16015;
wire n16016;
wire n16017;
wire n16018;
wire n16019;
wire n16020;
wire n16021;
wire n16022;
wire n16023;
wire n16024;
wire n16025;
wire n16026;
wire n16027;
wire n16028;
wire n16029;
wire n16030;
wire n16031;
wire n16032;
wire n16033;
wire n16034;
wire n16035;
wire n16036;
wire n16037;
wire n16038;
wire n16039;
wire n16040;
wire n16041;
wire n16042;
wire n16043;
wire n16044;
wire n16045;
wire n16046;
wire n16047;
wire n16048;
wire n16049;
wire n1605;
wire n16050;
wire n16051;
wire n16052;
wire n16053;
wire n16054;
wire n16055;
wire n16056;
wire n16057;
wire n16058;
wire n16059;
wire n16060;
wire n16061;
wire n16062;
wire n16063;
wire n16064;
wire n16065;
wire n16066;
wire n16067;
wire n16068;
wire n16069;
wire n16070;
wire n16071;
wire n16072;
wire n16073;
wire n16074;
wire n16075;
wire n16076;
wire n16077;
wire n16078;
wire n16079;
wire n16080;
wire n16081;
wire n16082;
wire n16083;
wire n16084;
wire n16085;
wire n16086;
wire n16087;
wire n16088;
wire n16089;
wire n16090;
wire n16091;
wire n16092;
wire n16093;
wire n16094;
wire n16095;
wire n16096;
wire n16097;
wire n16098;
wire n16099;
wire n1610;
wire n16100;
wire n16101;
wire n16102;
wire n16103;
wire n16104;
wire n16105;
wire n16106;
wire n16107;
wire n16108;
wire n16109;
wire n16110;
wire n16111;
wire n16112;
wire n16113;
wire n16114;
wire n16115;
wire n16116;
wire n16117;
wire n16118;
wire n16119;
wire n16120;
wire n16121;
wire n16122;
wire n16123;
wire n16124;
wire n16125;
wire n16126;
wire n16127;
wire n16128;
wire n16129;
wire n16130;
wire n16131;
wire n16132;
wire n16133;
wire n16134;
wire n16135;
wire n16136;
wire n16137;
wire n16138;
wire n16139;
wire n16140;
wire n16141;
wire n16142;
wire n16143;
wire n16144;
wire n16145;
wire n16146;
wire n16147;
wire n16148;
wire n16149;
wire n1615;
wire n16150;
wire n16151;
wire n16152;
wire n16153;
wire n16154;
wire n16155;
wire n16156;
wire n16157;
wire n16158;
wire n16159;
wire n16160;
wire n16161;
wire n16162;
wire n16163;
wire n16164;
wire n16165;
wire n16166;
wire n16167;
wire n16168;
wire n16169;
wire n16170;
wire n16171;
wire n16172;
wire n16173;
wire n16174;
wire n16175;
wire n16176;
wire n16177;
wire n16178;
wire n16179;
wire n16180;
wire n16181;
wire n16182;
wire n16183;
wire n16184;
wire n16185;
wire n16186;
wire n16187;
wire n16188;
wire n16189;
wire n16190;
wire n16191;
wire n16192;
wire n16193;
wire n16194;
wire n16195;
wire n16196;
wire n16197;
wire n16198;
wire n16199;
wire n1620;
wire n16200;
wire n16201;
wire n16202;
wire n16203;
wire n16204;
wire n16205;
wire n16206;
wire n16207;
wire n16208;
wire n16209;
wire n16210;
wire n16211;
wire n16212;
wire n16213;
wire n16214;
wire n16215;
wire n16216;
wire n16217;
wire n16218;
wire n16219;
wire n16220;
wire n16221;
wire n16222;
wire n16223;
wire n16224;
wire n16225;
wire n16226;
wire n16227;
wire n16228;
wire n16229;
wire n16230;
wire n16231;
wire n16232;
wire n16233;
wire n16234;
wire n16235;
wire n16236;
wire n16237;
wire n16238;
wire n16239;
wire n16240;
wire n16241;
wire n16242;
wire n16243;
wire n16244;
wire n16245;
wire n16246;
wire n16247;
wire n16248;
wire n16249;
wire n1625;
wire n16250;
wire n16251;
wire n16252;
wire n16253;
wire n16254;
wire n16255;
wire n16256;
wire n16257;
wire n16258;
wire n16259;
wire n16260;
wire n16261;
wire n16262;
wire n16263;
wire n16264;
wire n16265;
wire n16266;
wire n16267;
wire n16268;
wire n16269;
wire n16270;
wire n16271;
wire n16272;
wire n16273;
wire n16274;
wire n16275;
wire n16276;
wire n16277;
wire n16278;
wire n16279;
wire n16280;
wire n16281;
wire n16282;
wire n16283;
wire n16284;
wire n16285;
wire n16286;
wire n16287;
wire n16288;
wire n16289;
wire n16290;
wire n16291;
wire n16292;
wire n16293;
wire n16294;
wire n16295;
wire n16296;
wire n16297;
wire n16298;
wire n16299;
wire n1630;
wire n16300;
wire n16301;
wire n16302;
wire n16303;
wire n16304;
wire n16305;
wire n16306;
wire n16307;
wire n16308;
wire n16309;
wire n16310;
wire n16311;
wire n16312;
wire n16313;
wire n16314;
wire n16315;
wire n16316;
wire n16317;
wire n16318;
wire n16319;
wire n16320;
wire n16321;
wire n16322;
wire n16323;
wire n16324;
wire n16325;
wire n16326;
wire n16327;
wire n16328;
wire n16329;
wire n16330;
wire n16331;
wire n16332;
wire n16333;
wire n16334;
wire n16335;
wire n16336;
wire n16337;
wire n16338;
wire n16339;
wire n16340;
wire n16341;
wire n16342;
wire n16343;
wire n16344;
wire n16345;
wire n16346;
wire n16347;
wire n16348;
wire n16349;
wire n1635;
wire n16350;
wire n16351;
wire n16352;
wire n16353;
wire n16354;
wire n16355;
wire n16356;
wire n16357;
wire n16358;
wire n16359;
wire n16360;
wire n16361;
wire n16362;
wire n16363;
wire n16364;
wire n16365;
wire n16366;
wire n16367;
wire n16368;
wire n16369;
wire n16370;
wire n16371;
wire n16372;
wire n16373;
wire n16374;
wire n16375;
wire n16376;
wire n16377;
wire n16378;
wire n16379;
wire n16380;
wire n16381;
wire n16382;
wire n16383;
wire n16384;
wire n16385;
wire n16386;
wire n16387;
wire n16388;
wire n16389;
wire n16390;
wire n16391;
wire n16392;
wire n16393;
wire n16394;
wire n16395;
wire n16396;
wire n16397;
wire n16398;
wire n16399;
wire n1640;
wire n16400;
wire n16401;
wire n16402;
wire n16403;
wire n16404;
wire n16405;
wire n16406;
wire n16407;
wire n16408;
wire n16409;
wire n16410;
wire n16411;
wire n16412;
wire n16413;
wire n16414;
wire n16415;
wire n16416;
wire n16417;
wire n16418;
wire n16419;
wire n16420;
wire n16421;
wire n16422;
wire n16423;
wire n16424;
wire n16425;
wire n16426;
wire n16427;
wire n16428;
wire n16429;
wire n16430;
wire n16431;
wire n16432;
wire n16433;
wire n16434;
wire n16435;
wire n16436;
wire n16437;
wire n16438;
wire n16439;
wire n16440;
wire n16441;
wire n16442;
wire n16443;
wire n16444;
wire n16445;
wire n16446;
wire n16447;
wire n16448;
wire n16449;
wire n1645;
wire n16450;
wire n16451;
wire n16452;
wire n16453;
wire n16454;
wire n16455;
wire n16456;
wire n16457;
wire n16458;
wire n16459;
wire n16460;
wire n16461;
wire n16462;
wire n16463;
wire n16464;
wire n16465;
wire n16466;
wire n16467;
wire n16468;
wire n16469;
wire n16470;
wire n16471;
wire n16472;
wire n16473;
wire n16474;
wire n16475;
wire n16476;
wire n16477;
wire n16478;
wire n16479;
wire n16480;
wire n16481;
wire n16482;
wire n16483;
wire n16484;
wire n16485;
wire n16486;
wire n16487;
wire n16488;
wire n16489;
wire n16490;
wire n16491;
wire n16492;
wire n16493;
wire n16494;
wire n16495;
wire n16496;
wire n16497;
wire n16498;
wire n16499;
wire n1650;
wire n16500;
wire n16501;
wire n16502;
wire n16503;
wire n16504;
wire n16505;
wire n16506;
wire n16507;
wire n16508;
wire n16509;
wire n16510;
wire n16511;
wire n16512;
wire n16513;
wire n16514;
wire n16515;
wire n16516;
wire n16517;
wire n16518;
wire n16519;
wire n16520;
wire n16521;
wire n16522;
wire n16523;
wire n16524;
wire n16525;
wire n16526;
wire n16527;
wire n16528;
wire n16529;
wire n16530;
wire n16531;
wire n16532;
wire n16533;
wire n16534;
wire n16535;
wire n16536;
wire n16537;
wire n16538;
wire n16539;
wire n16540;
wire n16541;
wire n16542;
wire n16543;
wire n16544;
wire n16545;
wire n16546;
wire n16547;
wire n16549;
wire n1655;
wire n16550;
wire n16551;
wire n16552;
wire n16553;
wire n16554;
wire n16555;
wire n16556;
wire n16557;
wire n16558;
wire n16559;
wire n16560;
wire n16561;
wire n16562;
wire n16563;
wire n16564;
wire n16565;
wire n16566;
wire n16567;
wire n16568;
wire n16569;
wire n16570;
wire n16571;
wire n16572;
wire n16573;
wire n16574;
wire n16575;
wire n16576;
wire n16577;
wire n16578;
wire n16579;
wire n16580;
wire n16581;
wire n16582;
wire n16583;
wire n16584;
wire n16585;
wire n16586;
wire n16587;
wire n16588;
wire n16589;
wire n16590;
wire n16591;
wire n16592;
wire n16593;
wire n16594;
wire n16595;
wire n16596;
wire n16597;
wire n16598;
wire n16599;
wire n1660;
wire n16600;
wire n16601;
wire n16602;
wire n16603;
wire n16604;
wire n16605;
wire n16606;
wire n16607;
wire n16608;
wire n16609;
wire n16610;
wire n16611;
wire n16612;
wire n16613;
wire n16614;
wire n16615;
wire n16616;
wire n16617;
wire n16618;
wire n16619;
wire n16620;
wire n16621;
wire n16622;
wire n16623;
wire n16624;
wire n16625;
wire n16626;
wire n16627;
wire n16628;
wire n16629;
wire n16630;
wire n16631;
wire n16632;
wire n16633;
wire n16634;
wire n16635;
wire n16636;
wire n16637;
wire n16638;
wire n16639;
wire n1664;
wire n16640;
wire n16641;
wire n16642;
wire n16643;
wire n16644;
wire n16645;
wire n16646;
wire n16647;
wire n16648;
wire n16649;
wire n16650;
wire n16651;
wire n16652;
wire n16653;
wire n16654;
wire n16655;
wire n16656;
wire n16657;
wire n16658;
wire n16659;
wire n16660;
wire n16661;
wire n16662;
wire n16663;
wire n16664;
wire n16665;
wire n16666;
wire n16667;
wire n16668;
wire n16669;
wire n16670;
wire n16671;
wire n16672;
wire n16673;
wire n16674;
wire n16675;
wire n16676;
wire n16677;
wire n16678;
wire n16679;
wire n16680;
wire n16681;
wire n16682;
wire n16683;
wire n16684;
wire n16685;
wire n16686;
wire n16687;
wire n16688;
wire n16689;
wire n1669;
wire n16690;
wire n16691;
wire n16692;
wire n16693;
wire n16694;
wire n16695;
wire n16696;
wire n16697;
wire n16698;
wire n16699;
wire n16700;
wire n16701;
wire n16702;
wire n16703;
wire n16704;
wire n16705;
wire n16706;
wire n16707;
wire n16708;
wire n16709;
wire n16710;
wire n16711;
wire n16712;
wire n16713;
wire n16714;
wire n16715;
wire n16716;
wire n16717;
wire n16718;
wire n16719;
wire n16720;
wire n16721;
wire n16722;
wire n16723;
wire n16724;
wire n16725;
wire n16726;
wire n16727;
wire n16728;
wire n16729;
wire n16730;
wire n16731;
wire n16732;
wire n16733;
wire n16734;
wire n16735;
wire n16736;
wire n16737;
wire n16738;
wire n16739;
wire n1674;
wire n16740;
wire n16741;
wire n16742;
wire n16743;
wire n16744;
wire n16745;
wire n16746;
wire n16747;
wire n16748;
wire n16749;
wire n16750;
wire n16751;
wire n16752;
wire n16753;
wire n16754;
wire n16755;
wire n16756;
wire n16757;
wire n16758;
wire n16759;
wire n16760;
wire n16761;
wire n16762;
wire n16763;
wire n16764;
wire n16765;
wire n16766;
wire n16767;
wire n16768;
wire n16769;
wire n16770;
wire n16771;
wire n16772;
wire n16773;
wire n16774;
wire n16775;
wire n16776;
wire n16777;
wire n16778;
wire n16779;
wire n16780;
wire n16781;
wire n16782;
wire n16783;
wire n16784;
wire n16785;
wire n16786;
wire n16787;
wire n16788;
wire n16789;
wire n1679;
wire n16790;
wire n16791;
wire n16792;
wire n16793;
wire n16794;
wire n16795;
wire n16796;
wire n16797;
wire n16798;
wire n16799;
wire n16800;
wire n16801;
wire n16802;
wire n16803;
wire n16804;
wire n16805;
wire n16806;
wire n16807;
wire n16808;
wire n16809;
wire n16810;
wire n16811;
wire n16812;
wire n16813;
wire n16814;
wire n16815;
wire n16816;
wire n16817;
wire n16818;
wire n16819;
wire n16820;
wire n16821;
wire n16822;
wire n16823;
wire n16824;
wire n16825;
wire n16826;
wire n16827;
wire n16828;
wire n16829;
wire n16830;
wire n16831;
wire n16832;
wire n16833;
wire n16834;
wire n16835;
wire n16836;
wire n16837;
wire n16838;
wire n16839;
wire n1684;
wire n16840;
wire n16841;
wire n16842;
wire n16843;
wire n16844;
wire n16845;
wire n16846;
wire n16847;
wire n16848;
wire n16849;
wire n16850;
wire n16851;
wire n16852;
wire n16853;
wire n16854;
wire n16855;
wire n16856;
wire n16857;
wire n16858;
wire n16859;
wire n16860;
wire n16861;
wire n16862;
wire n16863;
wire n16864;
wire n16865;
wire n16866;
wire n16867;
wire n16868;
wire n16869;
wire n16870;
wire n16871;
wire n16872;
wire n16873;
wire n16874;
wire n16875;
wire n16876;
wire n16877;
wire n16878;
wire n16879;
wire n16880;
wire n16881;
wire n16882;
wire n16883;
wire n16884;
wire n16885;
wire n16886;
wire n16887;
wire n16888;
wire n16889;
wire n1689;
wire n16890;
wire n16891;
wire n16892;
wire n16893;
wire n16894;
wire n16895;
wire n16896;
wire n16897;
wire n16898;
wire n16899;
wire n16900;
wire n16901;
wire n16902;
wire n16903;
wire n16904;
wire n16905;
wire n16906;
wire n16907;
wire n16908;
wire n16909;
wire n16910;
wire n16911;
wire n16912;
wire n16913;
wire n16914;
wire n16915;
wire n16916;
wire n16917;
wire n16918;
wire n16919;
wire n16920;
wire n16921;
wire n16922;
wire n16923;
wire n16924;
wire n16925;
wire n16926;
wire n16927;
wire n16928;
wire n16929;
wire n16930;
wire n16931;
wire n16932;
wire n16933;
wire n16934;
wire n16935;
wire n16936;
wire n16937;
wire n16938;
wire n16939;
wire n1694;
wire n16940;
wire n16941;
wire n16942;
wire n16943;
wire n16944;
wire n16945;
wire n16946;
wire n16947;
wire n16948;
wire n16949;
wire n16950;
wire n16951;
wire n16952;
wire n16953;
wire n16954;
wire n16955;
wire n16956;
wire n16957;
wire n16958;
wire n16959;
wire n16960;
wire n16961;
wire n16962;
wire n16963;
wire n16964;
wire n16965;
wire n16966;
wire n16967;
wire n16968;
wire n16969;
wire n16970;
wire n16971;
wire n16972;
wire n16973;
wire n16974;
wire n16975;
wire n16976;
wire n16977;
wire n16978;
wire n16979;
wire n16980;
wire n16981;
wire n16982;
wire n16983;
wire n16984;
wire n16985;
wire n16986;
wire n16987;
wire n16988;
wire n16989;
wire n1699;
wire n16990;
wire n16991;
wire n16992;
wire n16993;
wire n16994;
wire n16995;
wire n16996;
wire n16997;
wire n16998;
wire n16999;
wire n17000;
wire n17001;
wire n17002;
wire n17003;
wire n17004;
wire n17005;
wire n17006;
wire n17007;
wire n17008;
wire n17009;
wire n17010;
wire n17011;
wire n17012;
wire n17013;
wire n17014;
wire n17015;
wire n17016;
wire n17017;
wire n17018;
wire n17019;
wire n17020;
wire n17021;
wire n17022;
wire n17023;
wire n17024;
wire n17025;
wire n17026;
wire n17027;
wire n17028;
wire n17029;
wire n17030;
wire n17031;
wire n17032;
wire n17033;
wire n17034;
wire n17035;
wire n17036;
wire n17037;
wire n17038;
wire n17039;
wire n1704;
wire n17040;
wire n17041;
wire n17042;
wire n17043;
wire n17044;
wire n17045;
wire n17046;
wire n17047;
wire n17048;
wire n17049;
wire n17050;
wire n17051;
wire n17052;
wire n17053;
wire n17054;
wire n17055;
wire n17056;
wire n17057;
wire n17058;
wire n17059;
wire n17060;
wire n17061;
wire n17062;
wire n17063;
wire n17064;
wire n17065;
wire n17066;
wire n17067;
wire n17068;
wire n17069;
wire n17070;
wire n17071;
wire n17072;
wire n17073;
wire n17074;
wire n17075;
wire n17076;
wire n17077;
wire n17078;
wire n17079;
wire n17080;
wire n17081;
wire n17082;
wire n17083;
wire n17084;
wire n17085;
wire n17086;
wire n17087;
wire n17088;
wire n17089;
wire n1709;
wire n17090;
wire n17091;
wire n17092;
wire n17093;
wire n17094;
wire n17095;
wire n17096;
wire n17097;
wire n17098;
wire n17099;
wire n17100;
wire n17101;
wire n17102;
wire n17103;
wire n17104;
wire n17105;
wire n17106;
wire n17107;
wire n17108;
wire n17109;
wire n17110;
wire n17111;
wire n17112;
wire n17113;
wire n17114;
wire n17115;
wire n17116;
wire n17117;
wire n17118;
wire n17119;
wire n17120;
wire n17121;
wire n17122;
wire n17123;
wire n17124;
wire n17125;
wire n17126;
wire n17127;
wire n17128;
wire n17129;
wire n17130;
wire n17131;
wire n17132;
wire n17133;
wire n17134;
wire n17135;
wire n17136;
wire n17137;
wire n17138;
wire n17139;
wire n1714;
wire n17140;
wire n17141;
wire n17142;
wire n17143;
wire n17144;
wire n17145;
wire n17146;
wire n17147;
wire n17148;
wire n17149;
wire n17150;
wire n17151;
wire n17152;
wire n17153;
wire n17154;
wire n17155;
wire n17156;
wire n17157;
wire n17158;
wire n17159;
wire n17160;
wire n17161;
wire n17162;
wire n17163;
wire n17164;
wire n17165;
wire n17166;
wire n17167;
wire n17168;
wire n17169;
wire n17170;
wire n17171;
wire n17172;
wire n17173;
wire n17174;
wire n17175;
wire n17176;
wire n17177;
wire n17178;
wire n17179;
wire n17180;
wire n17181;
wire n17182;
wire n17183;
wire n17184;
wire n17185;
wire n17186;
wire n17187;
wire n17188;
wire n17189;
wire n1719;
wire n17190;
wire n17191;
wire n17192;
wire n17193;
wire n17194;
wire n17195;
wire n17196;
wire n17197;
wire n17198;
wire n17199;
wire n17200;
wire n17201;
wire n17202;
wire n17203;
wire n17204;
wire n17205;
wire n17206;
wire n17207;
wire n17208;
wire n17209;
wire n17210;
wire n17211;
wire n17212;
wire n17213;
wire n17214;
wire n17215;
wire n17216;
wire n17217;
wire n17218;
wire n17219;
wire n17220;
wire n17221;
wire n17222;
wire n17223;
wire n17224;
wire n17225;
wire n17226;
wire n17227;
wire n17228;
wire n17229;
wire n17230;
wire n17231;
wire n17232;
wire n17233;
wire n17234;
wire n17235;
wire n17236;
wire n17237;
wire n17238;
wire n17239;
wire n1724;
wire n17240;
wire n17241;
wire n17242;
wire n17243;
wire n17244;
wire n17245;
wire n17246;
wire n17247;
wire n17248;
wire n17249;
wire n17250;
wire n17251;
wire n17252;
wire n17253;
wire n17254;
wire n17255;
wire n17256;
wire n17257;
wire n17258;
wire n17259;
wire n17260;
wire n17261;
wire n17262;
wire n17263;
wire n17264;
wire n17265;
wire n17266;
wire n17267;
wire n17268;
wire n17269;
wire n17270;
wire n17271;
wire n17272;
wire n17273;
wire n17274;
wire n17275;
wire n17276;
wire n17277;
wire n17278;
wire n17279;
wire n17280;
wire n17281;
wire n17282;
wire n17283;
wire n17284;
wire n17285;
wire n17286;
wire n17287;
wire n17288;
wire n17289;
wire n1729;
wire n17290;
wire n17291;
wire n17292;
wire n17293;
wire n17294;
wire n17295;
wire n17296;
wire n17297;
wire n17298;
wire n17299;
wire n17300;
wire n17301;
wire n17302;
wire n17303;
wire n17304;
wire n17305;
wire n17306;
wire n17307;
wire n17308;
wire n17309;
wire n17310;
wire n17311;
wire n17312;
wire n17313;
wire n17314;
wire n17315;
wire n17316;
wire n17317;
wire n17318;
wire n17319;
wire n17320;
wire n17321;
wire n17322;
wire n17323;
wire n17324;
wire n17325;
wire n17326;
wire n17327;
wire n17328;
wire n17329;
wire n17330;
wire n17331;
wire n17332;
wire n17333;
wire n17334;
wire n17335;
wire n17336;
wire n17337;
wire n17338;
wire n17339;
wire n1734;
wire n17340;
wire n17341;
wire n17342;
wire n17343;
wire n17344;
wire n17345;
wire n17346;
wire n17347;
wire n17348;
wire n17349;
wire n17350;
wire n17351;
wire n17352;
wire n17353;
wire n17354;
wire n17355;
wire n17356;
wire n17357;
wire n17358;
wire n17359;
wire n17360;
wire n17361;
wire n17362;
wire n17363;
wire n17364;
wire n17365;
wire n17366;
wire n17367;
wire n17368;
wire n17369;
wire n17370;
wire n17371;
wire n17372;
wire n17373;
wire n17374;
wire n17375;
wire n17376;
wire n17377;
wire n17378;
wire n17379;
wire n17380;
wire n17381;
wire n17382;
wire n17383;
wire n17384;
wire n17385;
wire n17386;
wire n17387;
wire n17388;
wire n17389;
wire n1739;
wire n17390;
wire n17391;
wire n17392;
wire n17393;
wire n17394;
wire n17395;
wire n17396;
wire n17397;
wire n17398;
wire n17399;
wire n17400;
wire n17401;
wire n17402;
wire n17403;
wire n17404;
wire n17405;
wire n17406;
wire n17407;
wire n17408;
wire n17409;
wire n17410;
wire n17411;
wire n17412;
wire n17413;
wire n17414;
wire n17415;
wire n17416;
wire n17417;
wire n17418;
wire n17419;
wire n17420;
wire n17421;
wire n17422;
wire n17423;
wire n17424;
wire n17425;
wire n17426;
wire n17427;
wire n17428;
wire n17429;
wire n17430;
wire n17431;
wire n17432;
wire n17433;
wire n17434;
wire n17435;
wire n17436;
wire n17437;
wire n17438;
wire n17439;
wire n1744;
wire n17440;
wire n17441;
wire n17442;
wire n17443;
wire n17444;
wire n17445;
wire n17446;
wire n17447;
wire n17448;
wire n17449;
wire n17450;
wire n17451;
wire n17452;
wire n17453;
wire n17454;
wire n17455;
wire n17456;
wire n17457;
wire n17458;
wire n17459;
wire n17460;
wire n17461;
wire n17462;
wire n17463;
wire n17464;
wire n17465;
wire n17466;
wire n17467;
wire n17468;
wire n17469;
wire n17470;
wire n17471;
wire n17472;
wire n17473;
wire n17474;
wire n17475;
wire n17476;
wire n17477;
wire n17478;
wire n17479;
wire n17480;
wire n17481;
wire n17482;
wire n17483;
wire n17484;
wire n17485;
wire n17486;
wire n17487;
wire n17488;
wire n17489;
wire n1749;
wire n17490;
wire n17491;
wire n17492;
wire n17493;
wire n17494;
wire n17495;
wire n17496;
wire n17497;
wire n17498;
wire n17499;
wire n17500;
wire n17501;
wire n17502;
wire n17503;
wire n17504;
wire n17505;
wire n17506;
wire n17507;
wire n17508;
wire n17509;
wire n17510;
wire n17511;
wire n17512;
wire n17513;
wire n17514;
wire n17515;
wire n17516;
wire n17517;
wire n17518;
wire n17519;
wire n17520;
wire n17521;
wire n17522;
wire n17523;
wire n17524;
wire n17525;
wire n17526;
wire n17527;
wire n17528;
wire n17529;
wire n17530;
wire n17531;
wire n17532;
wire n17533;
wire n17534;
wire n17535;
wire n17536;
wire n17537;
wire n17538;
wire n17539;
wire n1754;
wire n17540;
wire n17541;
wire n17542;
wire n17543;
wire n17544;
wire n17545;
wire n17546;
wire n17547;
wire n17548;
wire n17549;
wire n17550;
wire n17551;
wire n17552;
wire n17553;
wire n17554;
wire n17555;
wire n17556;
wire n17557;
wire n17558;
wire n17559;
wire n17560;
wire n17561;
wire n17562;
wire n17563;
wire n17564;
wire n17565;
wire n17566;
wire n17567;
wire n17568;
wire n17569;
wire n17570;
wire n17571;
wire n17572;
wire n17573;
wire n17574;
wire n17575;
wire n17576;
wire n17577;
wire n17578;
wire n17579;
wire n17580;
wire n17581;
wire n17582;
wire n17583;
wire n17584;
wire n17585;
wire n17586;
wire n17587;
wire n17588;
wire n17589;
wire n1759;
wire n17590;
wire n17591;
wire n17592;
wire n17593;
wire n17594;
wire n17595;
wire n17596;
wire n17597;
wire n17598;
wire n17599;
wire n17600;
wire n17601;
wire n17602;
wire n17603;
wire n17604;
wire n17605;
wire n17606;
wire n17607;
wire n17608;
wire n17609;
wire n17610;
wire n17611;
wire n17612;
wire n17613;
wire n17614;
wire n17615;
wire n17616;
wire n17617;
wire n17618;
wire n17619;
wire n17620;
wire n17621;
wire n17622;
wire n17623;
wire n17624;
wire n17625;
wire n17626;
wire n17627;
wire n17628;
wire n17629;
wire n1763;
wire n17630;
wire n17631;
wire n17632;
wire n17633;
wire n17634;
wire n17635;
wire n17636;
wire n17637;
wire n17638;
wire n17639;
wire n17640;
wire n17641;
wire n17642;
wire n17643;
wire n17644;
wire n17645;
wire n17646;
wire n17647;
wire n17648;
wire n17649;
wire n17650;
wire n17651;
wire n17652;
wire n17653;
wire n17654;
wire n17655;
wire n17656;
wire n17657;
wire n17658;
wire n17659;
wire n17660;
wire n17661;
wire n17662;
wire n17663;
wire n17664;
wire n17665;
wire n17666;
wire n17667;
wire n17668;
wire n17669;
wire n1767;
wire n17670;
wire n17671;
wire n17672;
wire n17673;
wire n17674;
wire n17675;
wire n17676;
wire n17677;
wire n17678;
wire n17679;
wire n17680;
wire n17681;
wire n17682;
wire n17683;
wire n17684;
wire n17685;
wire n17686;
wire n17687;
wire n17688;
wire n17689;
wire n17690;
wire n17691;
wire n17692;
wire n17693;
wire n17694;
wire n17695;
wire n17696;
wire n17697;
wire n17698;
wire n17699;
wire n17700;
wire n17701;
wire n17702;
wire n17703;
wire n17704;
wire n17705;
wire n17706;
wire n17707;
wire n17708;
wire n17709;
wire n17710;
wire n17711;
wire n17712;
wire n17713;
wire n17714;
wire n17715;
wire n17716;
wire n17717;
wire n17718;
wire n17719;
wire n1772;
wire n17720;
wire n17721;
wire n17722;
wire n17723;
wire n17724;
wire n17725;
wire n17726;
wire n17727;
wire n17728;
wire n17729;
wire n17730;
wire n17731;
wire n17732;
wire n17733;
wire n17734;
wire n17735;
wire n17736;
wire n17737;
wire n17738;
wire n17739;
wire n17740;
wire n17741;
wire n17742;
wire n17743;
wire n17744;
wire n17745;
wire n17746;
wire n17747;
wire n17748;
wire n17749;
wire n17750;
wire n17751;
wire n17752;
wire n17753;
wire n17754;
wire n17755;
wire n17756;
wire n17757;
wire n17758;
wire n17759;
wire n17760;
wire n17761;
wire n17762;
wire n17763;
wire n17764;
wire n17765;
wire n17766;
wire n17767;
wire n17768;
wire n17769;
wire n1777;
wire n17770;
wire n17771;
wire n17772;
wire n17773;
wire n17774;
wire n17775;
wire n17776;
wire n17777;
wire n17778;
wire n17779;
wire n17780;
wire n17781;
wire n17782;
wire n17783;
wire n17784;
wire n17785;
wire n17786;
wire n17787;
wire n17788;
wire n17789;
wire n17790;
wire n17791;
wire n17792;
wire n17793;
wire n17794;
wire n17795;
wire n17796;
wire n17797;
wire n17798;
wire n17799;
wire n17800;
wire n17801;
wire n17802;
wire n17803;
wire n17804;
wire n17805;
wire n17806;
wire n17807;
wire n17808;
wire n17809;
wire n17810;
wire n17811;
wire n17812;
wire n17813;
wire n17814;
wire n17815;
wire n17816;
wire n17817;
wire n17818;
wire n17819;
wire n1782;
wire n17820;
wire n17821;
wire n17822;
wire n17823;
wire n17824;
wire n17825;
wire n17826;
wire n17827;
wire n17828;
wire n17829;
wire n17830;
wire n17831;
wire n17832;
wire n17833;
wire n17834;
wire n17835;
wire n17836;
wire n17837;
wire n17838;
wire n17839;
wire n17840;
wire n17841;
wire n17842;
wire n17843;
wire n17844;
wire n17845;
wire n17846;
wire n17847;
wire n17848;
wire n17849;
wire n17850;
wire n17851;
wire n17852;
wire n17853;
wire n17854;
wire n17855;
wire n17856;
wire n17857;
wire n17858;
wire n17859;
wire n17860;
wire n17861;
wire n17862;
wire n17863;
wire n17864;
wire n17865;
wire n17866;
wire n17867;
wire n17868;
wire n17869;
wire n1787;
wire n17870;
wire n17871;
wire n17872;
wire n17873;
wire n17874;
wire n17875;
wire n17876;
wire n17877;
wire n17878;
wire n17879;
wire n17880;
wire n17881;
wire n17882;
wire n17883;
wire n17884;
wire n17885;
wire n17886;
wire n17887;
wire n17888;
wire n17889;
wire n17890;
wire n17891;
wire n17892;
wire n17893;
wire n17894;
wire n17895;
wire n17896;
wire n17897;
wire n17898;
wire n17899;
wire n17900;
wire n17901;
wire n17902;
wire n17903;
wire n17904;
wire n17905;
wire n17906;
wire n17907;
wire n17908;
wire n17909;
wire n17910;
wire n17911;
wire n17912;
wire n17913;
wire n17914;
wire n17915;
wire n17916;
wire n17917;
wire n17918;
wire n17919;
wire n1792;
wire n17920;
wire n17921;
wire n17922;
wire n17923;
wire n17924;
wire n17925;
wire n17926;
wire n17927;
wire n17928;
wire n17929;
wire n17930;
wire n17931;
wire n17932;
wire n17933;
wire n17934;
wire n17935;
wire n17936;
wire n17937;
wire n17938;
wire n17939;
wire n17940;
wire n17941;
wire n17942;
wire n17943;
wire n17944;
wire n17945;
wire n17946;
wire n17947;
wire n17948;
wire n17949;
wire n17950;
wire n17951;
wire n17952;
wire n17953;
wire n17954;
wire n17955;
wire n17956;
wire n17957;
wire n17958;
wire n17959;
wire n1796;
wire n17961;
wire n17962;
wire n17964;
wire n17965;
wire n17966;
wire n17967;
wire n17968;
wire n17969;
wire n17970;
wire n17971;
wire n17972;
wire n17973;
wire n17974;
wire n17975;
wire n17976;
wire n17977;
wire n17978;
wire n17979;
wire n17980;
wire n17981;
wire n17982;
wire n17983;
wire n17984;
wire n17985;
wire n17986;
wire n17987;
wire n17988;
wire n17989;
wire n17990;
wire n17991;
wire n17992;
wire n17993;
wire n17994;
wire n17995;
wire n17996;
wire n17997;
wire n17998;
wire n17999;
wire n18000;
wire n18001;
wire n18002;
wire n18003;
wire n18004;
wire n18005;
wire n18006;
wire n18007;
wire n18008;
wire n18009;
wire n1801;
wire n18010;
wire n18011;
wire n18012;
wire n18013;
wire n18014;
wire n18015;
wire n18016;
wire n18017;
wire n18018;
wire n18019;
wire n18020;
wire n18021;
wire n18022;
wire n18023;
wire n18024;
wire n18025;
wire n18026;
wire n18027;
wire n18028;
wire n18029;
wire n18030;
wire n18031;
wire n18032;
wire n18033;
wire n18034;
wire n18035;
wire n18036;
wire n18037;
wire n18038;
wire n18039;
wire n18040;
wire n18041;
wire n18042;
wire n18043;
wire n18044;
wire n18045;
wire n18046;
wire n18047;
wire n18048;
wire n18049;
wire n18050;
wire n18051;
wire n18052;
wire n18053;
wire n18054;
wire n18055;
wire n18056;
wire n18057;
wire n18058;
wire n18059;
wire n1806;
wire n18060;
wire n18061;
wire n18062;
wire n18063;
wire n18064;
wire n18065;
wire n18066;
wire n18067;
wire n18068;
wire n18069;
wire n18070;
wire n18071;
wire n18072;
wire n18073;
wire n18074;
wire n18075;
wire n18076;
wire n18077;
wire n18078;
wire n18079;
wire n18080;
wire n18081;
wire n18082;
wire n18083;
wire n18084;
wire n18085;
wire n18086;
wire n18087;
wire n18088;
wire n18089;
wire n18090;
wire n18091;
wire n18092;
wire n18093;
wire n18094;
wire n18095;
wire n18096;
wire n18097;
wire n18098;
wire n18099;
wire n18100;
wire n18101;
wire n18102;
wire n18103;
wire n18104;
wire n18105;
wire n18106;
wire n18107;
wire n18108;
wire n18109;
wire n1811;
wire n18110;
wire n18111;
wire n18112;
wire n18113;
wire n18114;
wire n18115;
wire n18116;
wire n18117;
wire n18118;
wire n18119;
wire n18120;
wire n18121;
wire n18122;
wire n18123;
wire n18124;
wire n18125;
wire n18126;
wire n18127;
wire n18128;
wire n18129;
wire n18130;
wire n18131;
wire n18132;
wire n18133;
wire n18134;
wire n18135;
wire n18136;
wire n18137;
wire n18138;
wire n18139;
wire n18140;
wire n18141;
wire n18142;
wire n18143;
wire n18144;
wire n18145;
wire n18146;
wire n18147;
wire n18148;
wire n18149;
wire n18150;
wire n18151;
wire n18152;
wire n18153;
wire n18154;
wire n18155;
wire n18156;
wire n18157;
wire n18158;
wire n18159;
wire n1816;
wire n18160;
wire n18161;
wire n18162;
wire n18163;
wire n18164;
wire n18165;
wire n18166;
wire n18167;
wire n18168;
wire n18169;
wire n18170;
wire n18171;
wire n18172;
wire n18173;
wire n18174;
wire n18175;
wire n18176;
wire n18177;
wire n18178;
wire n18180;
wire n18181;
wire n18182;
wire n18183;
wire n18184;
wire n18185;
wire n18186;
wire n18187;
wire n18188;
wire n18189;
wire n18190;
wire n18191;
wire n18192;
wire n18193;
wire n18194;
wire n18195;
wire n18196;
wire n18197;
wire n18198;
wire n18199;
wire n18200;
wire n18201;
wire n18202;
wire n18203;
wire n18204;
wire n18205;
wire n18206;
wire n18207;
wire n18208;
wire n18209;
wire n1821;
wire n18210;
wire n18211;
wire n18212;
wire n18213;
wire n18214;
wire n18215;
wire n18216;
wire n18217;
wire n18218;
wire n18219;
wire n18220;
wire n18221;
wire n18222;
wire n18223;
wire n18224;
wire n18225;
wire n18226;
wire n18227;
wire n18228;
wire n18229;
wire n18230;
wire n18231;
wire n18232;
wire n18233;
wire n18234;
wire n18235;
wire n18236;
wire n18237;
wire n18238;
wire n18239;
wire n18240;
wire n18241;
wire n18242;
wire n18243;
wire n18244;
wire n18245;
wire n18246;
wire n18247;
wire n18248;
wire n18249;
wire n18250;
wire n18251;
wire n18252;
wire n18253;
wire n18254;
wire n18255;
wire n18256;
wire n18257;
wire n18258;
wire n18259;
wire n1826;
wire n18260;
wire n18261;
wire n18262;
wire n18263;
wire n18264;
wire n18265;
wire n18266;
wire n18267;
wire n18268;
wire n18269;
wire n18270;
wire n18271;
wire n18272;
wire n18273;
wire n18274;
wire n18275;
wire n18276;
wire n18277;
wire n18278;
wire n18279;
wire n18280;
wire n18281;
wire n18282;
wire n18283;
wire n18284;
wire n18285;
wire n18286;
wire n18287;
wire n18288;
wire n18289;
wire n18290;
wire n18291;
wire n18292;
wire n18293;
wire n18294;
wire n18295;
wire n18296;
wire n18297;
wire n18298;
wire n18299;
wire n18300;
wire n18301;
wire n18302;
wire n18303;
wire n18304;
wire n18305;
wire n18306;
wire n18307;
wire n18308;
wire n18309;
wire n1831;
wire n18310;
wire n18311;
wire n18312;
wire n18313;
wire n18314;
wire n18315;
wire n18316;
wire n18317;
wire n18318;
wire n18319;
wire n18320;
wire n18321;
wire n18322;
wire n18323;
wire n18324;
wire n18325;
wire n18326;
wire n18327;
wire n18328;
wire n18329;
wire n18330;
wire n18331;
wire n18332;
wire n18333;
wire n18334;
wire n18335;
wire n18336;
wire n18337;
wire n18338;
wire n18339;
wire n18340;
wire n18341;
wire n18342;
wire n18343;
wire n18344;
wire n18345;
wire n18346;
wire n18347;
wire n18348;
wire n18349;
wire n1835;
wire n18350;
wire n18351;
wire n18352;
wire n18353;
wire n18354;
wire n18355;
wire n18356;
wire n18357;
wire n18358;
wire n18359;
wire n18360;
wire n18361;
wire n18362;
wire n18363;
wire n18364;
wire n18365;
wire n18366;
wire n18367;
wire n18368;
wire n18369;
wire n18370;
wire n18371;
wire n18372;
wire n18373;
wire n18374;
wire n18375;
wire n18376;
wire n18377;
wire n18378;
wire n18379;
wire n18380;
wire n18381;
wire n18382;
wire n18383;
wire n18384;
wire n18385;
wire n18386;
wire n18387;
wire n18388;
wire n18389;
wire n18390;
wire n18391;
wire n18392;
wire n18393;
wire n18394;
wire n18395;
wire n18396;
wire n18397;
wire n18398;
wire n18399;
wire n1840;
wire n18400;
wire n18401;
wire n18402;
wire n18403;
wire n18404;
wire n18405;
wire n18406;
wire n18407;
wire n18408;
wire n18409;
wire n18410;
wire n18411;
wire n18412;
wire n18413;
wire n18414;
wire n18415;
wire n18416;
wire n18417;
wire n18418;
wire n18419;
wire n18420;
wire n18421;
wire n18422;
wire n18423;
wire n18424;
wire n18425;
wire n18426;
wire n18427;
wire n18428;
wire n18429;
wire n18430;
wire n18431;
wire n18432;
wire n18433;
wire n18434;
wire n18435;
wire n18436;
wire n18437;
wire n18438;
wire n18439;
wire n18440;
wire n18441;
wire n18442;
wire n18443;
wire n18444;
wire n18445;
wire n18446;
wire n18447;
wire n18448;
wire n18449;
wire n1845;
wire n18450;
wire n18451;
wire n18452;
wire n18453;
wire n18454;
wire n18455;
wire n18456;
wire n18457;
wire n18458;
wire n18459;
wire n18460;
wire n18461;
wire n18462;
wire n18463;
wire n18464;
wire n18465;
wire n18466;
wire n18467;
wire n18468;
wire n18469;
wire n18470;
wire n18471;
wire n18472;
wire n18473;
wire n18474;
wire n18475;
wire n18476;
wire n18477;
wire n18478;
wire n18479;
wire n18480;
wire n18481;
wire n18482;
wire n18483;
wire n18484;
wire n18485;
wire n18486;
wire n18487;
wire n18488;
wire n18489;
wire n18490;
wire n18491;
wire n18492;
wire n18493;
wire n18494;
wire n18495;
wire n18496;
wire n18497;
wire n18498;
wire n18499;
wire n1850;
wire n18500;
wire n18501;
wire n18502;
wire n18503;
wire n18504;
wire n18505;
wire n18506;
wire n18507;
wire n18508;
wire n18509;
wire n18510;
wire n18511;
wire n18512;
wire n18513;
wire n18514;
wire n18515;
wire n18516;
wire n18517;
wire n18518;
wire n18519;
wire n18520;
wire n18521;
wire n18522;
wire n18523;
wire n18524;
wire n18525;
wire n18526;
wire n18527;
wire n18528;
wire n18529;
wire n18530;
wire n18531;
wire n18532;
wire n18533;
wire n18534;
wire n18535;
wire n18536;
wire n18537;
wire n18538;
wire n18539;
wire n18540;
wire n18541;
wire n18542;
wire n18543;
wire n18544;
wire n18545;
wire n18546;
wire n18547;
wire n18548;
wire n18549;
wire n1855;
wire n18550;
wire n18551;
wire n18552;
wire n18553;
wire n18554;
wire n18555;
wire n18556;
wire n18557;
wire n18558;
wire n18559;
wire n18560;
wire n18561;
wire n18562;
wire n18563;
wire n18564;
wire n18565;
wire n18566;
wire n18567;
wire n18568;
wire n18569;
wire n18570;
wire n18571;
wire n18572;
wire n18573;
wire n18574;
wire n18575;
wire n18576;
wire n18577;
wire n18578;
wire n18579;
wire n18580;
wire n18581;
wire n18582;
wire n18583;
wire n18584;
wire n18585;
wire n18586;
wire n18587;
wire n18588;
wire n18589;
wire n18590;
wire n18591;
wire n18592;
wire n18593;
wire n18594;
wire n18595;
wire n18596;
wire n18597;
wire n18598;
wire n18599;
wire n1860;
wire n18600;
wire n18601;
wire n18602;
wire n18603;
wire n18604;
wire n18605;
wire n18606;
wire n18607;
wire n18608;
wire n18609;
wire n18610;
wire n18611;
wire n18612;
wire n18613;
wire n18614;
wire n18615;
wire n18616;
wire n18617;
wire n18618;
wire n18619;
wire n18620;
wire n18621;
wire n18622;
wire n18623;
wire n18624;
wire n18625;
wire n18626;
wire n18627;
wire n18628;
wire n18629;
wire n18630;
wire n18631;
wire n18632;
wire n18633;
wire n18634;
wire n18635;
wire n18636;
wire n18637;
wire n18638;
wire n18639;
wire n18640;
wire n18641;
wire n18642;
wire n18643;
wire n18644;
wire n18645;
wire n18646;
wire n18647;
wire n18648;
wire n18649;
wire n1865;
wire n18650;
wire n18651;
wire n18652;
wire n18653;
wire n18654;
wire n18655;
wire n18656;
wire n18657;
wire n18658;
wire n18659;
wire n18660;
wire n18661;
wire n18662;
wire n18663;
wire n18664;
wire n18665;
wire n18666;
wire n18667;
wire n18668;
wire n18669;
wire n18670;
wire n18671;
wire n18672;
wire n18673;
wire n18674;
wire n18675;
wire n18676;
wire n18677;
wire n18678;
wire n18679;
wire n18680;
wire n18681;
wire n18682;
wire n18683;
wire n18684;
wire n18685;
wire n18686;
wire n18687;
wire n18688;
wire n18689;
wire n1869;
wire n18690;
wire n18691;
wire n18692;
wire n18693;
wire n18694;
wire n18695;
wire n18696;
wire n18697;
wire n18698;
wire n18699;
wire n18700;
wire n18701;
wire n18702;
wire n18703;
wire n18704;
wire n18705;
wire n18706;
wire n18707;
wire n18708;
wire n18709;
wire n18710;
wire n18711;
wire n18712;
wire n18713;
wire n18714;
wire n18715;
wire n18716;
wire n18717;
wire n18718;
wire n18719;
wire n18720;
wire n18721;
wire n18722;
wire n18723;
wire n18724;
wire n18725;
wire n18726;
wire n18727;
wire n18728;
wire n18729;
wire n18730;
wire n18731;
wire n18732;
wire n18733;
wire n18734;
wire n18735;
wire n18736;
wire n18737;
wire n18738;
wire n18739;
wire n1874;
wire n18740;
wire n18741;
wire n18742;
wire n18743;
wire n18744;
wire n18745;
wire n18746;
wire n18747;
wire n18748;
wire n18749;
wire n18750;
wire n18751;
wire n18752;
wire n18753;
wire n18754;
wire n18755;
wire n18756;
wire n18757;
wire n18758;
wire n18759;
wire n18760;
wire n18761;
wire n18762;
wire n18763;
wire n18764;
wire n18765;
wire n18766;
wire n18767;
wire n18768;
wire n18769;
wire n18770;
wire n18771;
wire n18772;
wire n18773;
wire n18774;
wire n18775;
wire n18776;
wire n18777;
wire n18778;
wire n18779;
wire n18780;
wire n18781;
wire n18782;
wire n18783;
wire n18784;
wire n18785;
wire n18786;
wire n18787;
wire n18788;
wire n18789;
wire n1879;
wire n18790;
wire n18791;
wire n18792;
wire n18793;
wire n18794;
wire n18795;
wire n18796;
wire n18797;
wire n18798;
wire n18799;
wire n18800;
wire n18801;
wire n18802;
wire n18803;
wire n18804;
wire n18805;
wire n18806;
wire n18807;
wire n18808;
wire n18809;
wire n18810;
wire n18811;
wire n18812;
wire n18813;
wire n18814;
wire n18815;
wire n18816;
wire n18817;
wire n18818;
wire n18819;
wire n18820;
wire n18821;
wire n18822;
wire n18823;
wire n18824;
wire n18825;
wire n18826;
wire n18827;
wire n18828;
wire n18829;
wire n18830;
wire n18831;
wire n18832;
wire n18833;
wire n18834;
wire n18835;
wire n18836;
wire n18837;
wire n18838;
wire n18839;
wire n1884;
wire n18840;
wire n18841;
wire n18842;
wire n18843;
wire n18844;
wire n18845;
wire n18846;
wire n18847;
wire n18848;
wire n18849;
wire n18850;
wire n18851;
wire n18852;
wire n18853;
wire n18854;
wire n18855;
wire n18856;
wire n18857;
wire n18858;
wire n18859;
wire n18860;
wire n18861;
wire n18862;
wire n18863;
wire n18864;
wire n18865;
wire n18866;
wire n18867;
wire n18868;
wire n18869;
wire n18870;
wire n18871;
wire n18872;
wire n18873;
wire n18874;
wire n18875;
wire n18876;
wire n18877;
wire n18878;
wire n18879;
wire n18880;
wire n18881;
wire n18882;
wire n18883;
wire n18884;
wire n18885;
wire n18886;
wire n18887;
wire n18888;
wire n18889;
wire n1889;
wire n18890;
wire n18891;
wire n18892;
wire n18893;
wire n18894;
wire n18895;
wire n18896;
wire n18897;
wire n18898;
wire n18899;
wire n18900;
wire n18901;
wire n18902;
wire n18903;
wire n18904;
wire n18905;
wire n18906;
wire n18907;
wire n18908;
wire n18909;
wire n18910;
wire n18911;
wire n18912;
wire n18913;
wire n18914;
wire n18915;
wire n18916;
wire n18917;
wire n18918;
wire n18919;
wire n18920;
wire n18921;
wire n18922;
wire n18923;
wire n18924;
wire n18925;
wire n18926;
wire n18927;
wire n18928;
wire n18929;
wire n18930;
wire n18931;
wire n18932;
wire n18933;
wire n18934;
wire n18935;
wire n18936;
wire n18937;
wire n18938;
wire n18939;
wire n1894;
wire n18940;
wire n18941;
wire n18942;
wire n18943;
wire n18944;
wire n18945;
wire n18946;
wire n18947;
wire n18948;
wire n18949;
wire n18950;
wire n18951;
wire n18952;
wire n18953;
wire n18954;
wire n18955;
wire n18956;
wire n18957;
wire n18958;
wire n18959;
wire n18960;
wire n18961;
wire n18962;
wire n18963;
wire n18964;
wire n18965;
wire n18966;
wire n18967;
wire n18968;
wire n18969;
wire n18970;
wire n18971;
wire n18972;
wire n18973;
wire n18974;
wire n18975;
wire n18976;
wire n18977;
wire n18978;
wire n18979;
wire n18980;
wire n18981;
wire n18982;
wire n18983;
wire n18984;
wire n18985;
wire n18986;
wire n18987;
wire n18988;
wire n18989;
wire n1899;
wire n18990;
wire n18991;
wire n18992;
wire n18993;
wire n18994;
wire n18995;
wire n18996;
wire n18997;
wire n18998;
wire n18999;
wire n19000;
wire n19001;
wire n19002;
wire n19003;
wire n19004;
wire n19005;
wire n19006;
wire n19007;
wire n19008;
wire n19009;
wire n19010;
wire n19011;
wire n19012;
wire n19013;
wire n19014;
wire n19015;
wire n19016;
wire n19017;
wire n19018;
wire n19019;
wire n19020;
wire n19021;
wire n19022;
wire n19023;
wire n19024;
wire n19025;
wire n19026;
wire n19027;
wire n19028;
wire n19029;
wire n19030;
wire n19031;
wire n19032;
wire n19033;
wire n19034;
wire n19035;
wire n19036;
wire n19037;
wire n19038;
wire n19039;
wire n1904;
wire n19040;
wire n19041;
wire n19042;
wire n19043;
wire n19044;
wire n19045;
wire n19046;
wire n19047;
wire n19048;
wire n19049;
wire n19050;
wire n19051;
wire n19052;
wire n19053;
wire n19054;
wire n19055;
wire n19056;
wire n19057;
wire n19058;
wire n19059;
wire n19060;
wire n19061;
wire n19062;
wire n19063;
wire n19064;
wire n19065;
wire n19066;
wire n19067;
wire n19068;
wire n19069;
wire n19070;
wire n19071;
wire n19072;
wire n19073;
wire n19074;
wire n19075;
wire n19076;
wire n19077;
wire n19078;
wire n19079;
wire n19080;
wire n19081;
wire n19082;
wire n19083;
wire n19084;
wire n19085;
wire n19086;
wire n19087;
wire n19088;
wire n19089;
wire n1909;
wire n19090;
wire n19091;
wire n19092;
wire n19093;
wire n19094;
wire n19095;
wire n19096;
wire n19097;
wire n19098;
wire n19099;
wire n19100;
wire n19101;
wire n19102;
wire n19103;
wire n19104;
wire n19105;
wire n19106;
wire n19107;
wire n19108;
wire n19109;
wire n19110;
wire n19111;
wire n19112;
wire n19113;
wire n19114;
wire n19115;
wire n19116;
wire n19117;
wire n19118;
wire n19119;
wire n19120;
wire n19121;
wire n19122;
wire n19123;
wire n19124;
wire n19125;
wire n19126;
wire n19127;
wire n19128;
wire n19129;
wire n19130;
wire n19131;
wire n19132;
wire n19133;
wire n19134;
wire n19135;
wire n19136;
wire n19137;
wire n19138;
wire n19139;
wire n1914;
wire n19140;
wire n19141;
wire n19142;
wire n19143;
wire n19144;
wire n19145;
wire n19146;
wire n19147;
wire n19148;
wire n19149;
wire n19150;
wire n19151;
wire n19152;
wire n19153;
wire n19154;
wire n19155;
wire n19156;
wire n19157;
wire n19158;
wire n19159;
wire n19160;
wire n19161;
wire n19162;
wire n19163;
wire n19164;
wire n19165;
wire n19166;
wire n19167;
wire n19168;
wire n19169;
wire n19170;
wire n19171;
wire n19172;
wire n19173;
wire n19174;
wire n19175;
wire n19176;
wire n19177;
wire n19178;
wire n19179;
wire n19180;
wire n19181;
wire n19182;
wire n19183;
wire n19184;
wire n19185;
wire n19186;
wire n19187;
wire n19188;
wire n19189;
wire n1919;
wire n19190;
wire n19191;
wire n19192;
wire n19193;
wire n19194;
wire n19195;
wire n19196;
wire n19197;
wire n19198;
wire n19199;
wire n19200;
wire n19201;
wire n19202;
wire n19203;
wire n19204;
wire n19205;
wire n19206;
wire n19207;
wire n19208;
wire n19209;
wire n19210;
wire n19211;
wire n19212;
wire n19213;
wire n19214;
wire n19215;
wire n19216;
wire n19217;
wire n19218;
wire n19219;
wire n19220;
wire n19221;
wire n19222;
wire n19223;
wire n19224;
wire n19225;
wire n19226;
wire n19227;
wire n19228;
wire n19229;
wire n19230;
wire n19231;
wire n19232;
wire n19233;
wire n19234;
wire n19235;
wire n19236;
wire n19237;
wire n19238;
wire n19239;
wire n1924;
wire n19240;
wire n19241;
wire n19242;
wire n19243;
wire n19244;
wire n19245;
wire n19246;
wire n19247;
wire n19248;
wire n19249;
wire n19250;
wire n19251;
wire n19252;
wire n19253;
wire n19254;
wire n19255;
wire n19256;
wire n19257;
wire n19258;
wire n19259;
wire n19260;
wire n19261;
wire n19262;
wire n19263;
wire n19264;
wire n19265;
wire n19266;
wire n19267;
wire n19268;
wire n19269;
wire n19270;
wire n19271;
wire n19272;
wire n19273;
wire n19274;
wire n19275;
wire n19276;
wire n19277;
wire n19278;
wire n19279;
wire n19280;
wire n19281;
wire n19282;
wire n19283;
wire n19284;
wire n19285;
wire n19286;
wire n19287;
wire n19288;
wire n19289;
wire n1929;
wire n19290;
wire n19291;
wire n19292;
wire n19293;
wire n19294;
wire n19295;
wire n19296;
wire n19297;
wire n19298;
wire n19299;
wire n19300;
wire n19301;
wire n19302;
wire n19303;
wire n19304;
wire n19305;
wire n19306;
wire n19307;
wire n19308;
wire n19309;
wire n19310;
wire n19311;
wire n19312;
wire n19313;
wire n19314;
wire n19315;
wire n19316;
wire n19317;
wire n19318;
wire n19319;
wire n19320;
wire n19321;
wire n19322;
wire n19323;
wire n19324;
wire n19325;
wire n19326;
wire n19327;
wire n19328;
wire n19329;
wire n19330;
wire n19331;
wire n19332;
wire n19333;
wire n19334;
wire n19335;
wire n19336;
wire n19337;
wire n19338;
wire n19339;
wire n1934;
wire n19340;
wire n19341;
wire n19342;
wire n19343;
wire n19344;
wire n19345;
wire n19346;
wire n19347;
wire n19348;
wire n19349;
wire n19350;
wire n19351;
wire n19352;
wire n19353;
wire n19354;
wire n19355;
wire n19356;
wire n19357;
wire n19358;
wire n19359;
wire n19360;
wire n19361;
wire n19362;
wire n19363;
wire n19364;
wire n19365;
wire n19366;
wire n19367;
wire n19368;
wire n19369;
wire n19370;
wire n19371;
wire n19372;
wire n19373;
wire n19374;
wire n19375;
wire n19376;
wire n19377;
wire n19378;
wire n19379;
wire n19380;
wire n19381;
wire n19382;
wire n19383;
wire n19384;
wire n19385;
wire n19386;
wire n19387;
wire n19388;
wire n19389;
wire n1939;
wire n19390;
wire n19391;
wire n19392;
wire n19393;
wire n19394;
wire n19395;
wire n19396;
wire n19397;
wire n19398;
wire n19399;
wire n19400;
wire n19401;
wire n19402;
wire n19403;
wire n19404;
wire n19405;
wire n19406;
wire n19407;
wire n19408;
wire n19409;
wire n19410;
wire n19411;
wire n19412;
wire n19413;
wire n19414;
wire n19415;
wire n19416;
wire n19417;
wire n19418;
wire n19419;
wire n19420;
wire n19421;
wire n19422;
wire n19423;
wire n19424;
wire n19425;
wire n19426;
wire n19427;
wire n19428;
wire n19429;
wire n19430;
wire n19431;
wire n19432;
wire n19433;
wire n19434;
wire n19435;
wire n19436;
wire n19437;
wire n19438;
wire n19439;
wire n1944;
wire n19440;
wire n19441;
wire n19442;
wire n19443;
wire n19444;
wire n19445;
wire n19446;
wire n19447;
wire n19448;
wire n19449;
wire n19450;
wire n19451;
wire n19452;
wire n19453;
wire n19454;
wire n19455;
wire n19456;
wire n19457;
wire n19458;
wire n19459;
wire n19460;
wire n19461;
wire n19462;
wire n19463;
wire n19464;
wire n19465;
wire n19466;
wire n19467;
wire n19468;
wire n19469;
wire n19470;
wire n19471;
wire n19472;
wire n19473;
wire n19474;
wire n19475;
wire n19476;
wire n19477;
wire n19478;
wire n19479;
wire n19480;
wire n19481;
wire n19482;
wire n19483;
wire n19484;
wire n19485;
wire n19486;
wire n19487;
wire n19488;
wire n19489;
wire n1949;
wire n19490;
wire n19491;
wire n19492;
wire n19493;
wire n19494;
wire n19495;
wire n19496;
wire n19497;
wire n19498;
wire n19499;
wire n19500;
wire n19501;
wire n19502;
wire n19503;
wire n19504;
wire n19505;
wire n19506;
wire n19507;
wire n19508;
wire n19509;
wire n19510;
wire n19511;
wire n19512;
wire n19513;
wire n19514;
wire n19515;
wire n19516;
wire n19517;
wire n19518;
wire n19519;
wire n19520;
wire n19521;
wire n19522;
wire n19523;
wire n19524;
wire n19525;
wire n19526;
wire n19527;
wire n19528;
wire n19529;
wire n19530;
wire n19531;
wire n19532;
wire n19533;
wire n19534;
wire n19535;
wire n19536;
wire n19537;
wire n19538;
wire n19539;
wire n1954;
wire n19540;
wire n19541;
wire n19542;
wire n19543;
wire n19544;
wire n19545;
wire n19546;
wire n19547;
wire n19548;
wire n19549;
wire n19550;
wire n19551;
wire n19552;
wire n19553;
wire n19554;
wire n19555;
wire n19556;
wire n19557;
wire n19558;
wire n19559;
wire n19560;
wire n19561;
wire n19562;
wire n19563;
wire n19564;
wire n19565;
wire n19566;
wire n19567;
wire n19568;
wire n19569;
wire n19570;
wire n19571;
wire n19572;
wire n19573;
wire n19574;
wire n19575;
wire n19576;
wire n19577;
wire n19578;
wire n19579;
wire n19580;
wire n19581;
wire n19582;
wire n19583;
wire n19584;
wire n19585;
wire n19586;
wire n19587;
wire n19588;
wire n19589;
wire n1959;
wire n19590;
wire n19591;
wire n19592;
wire n19593;
wire n19594;
wire n19595;
wire n19596;
wire n19597;
wire n19598;
wire n19599;
wire n19600;
wire n19601;
wire n19602;
wire n19603;
wire n19604;
wire n19605;
wire n19606;
wire n19607;
wire n19608;
wire n19609;
wire n19610;
wire n19611;
wire n19612;
wire n19613;
wire n19614;
wire n19615;
wire n19616;
wire n19617;
wire n19618;
wire n19619;
wire n19620;
wire n19621;
wire n19622;
wire n19623;
wire n19624;
wire n19625;
wire n19626;
wire n19627;
wire n19628;
wire n19629;
wire n19630;
wire n19631;
wire n19632;
wire n19633;
wire n19634;
wire n19635;
wire n19636;
wire n19637;
wire n19638;
wire n19639;
wire n1964;
wire n19640;
wire n19641;
wire n19642;
wire n19643;
wire n19644;
wire n19645;
wire n19646;
wire n19647;
wire n19648;
wire n19649;
wire n19650;
wire n19651;
wire n19652;
wire n19653;
wire n19654;
wire n19655;
wire n19656;
wire n19657;
wire n19658;
wire n19659;
wire n19660;
wire n19661;
wire n19662;
wire n19663;
wire n19664;
wire n19665;
wire n19666;
wire n19667;
wire n19668;
wire n19669;
wire n19670;
wire n19671;
wire n19672;
wire n19673;
wire n19674;
wire n19675;
wire n19676;
wire n19677;
wire n19678;
wire n19679;
wire n19680;
wire n19681;
wire n19682;
wire n19683;
wire n19684;
wire n19685;
wire n19686;
wire n19687;
wire n19688;
wire n19689;
wire n1969;
wire n19690;
wire n19691;
wire n19692;
wire n19693;
wire n19694;
wire n19695;
wire n19696;
wire n19697;
wire n19698;
wire n19699;
wire n19700;
wire n19701;
wire n19702;
wire n19703;
wire n19704;
wire n19705;
wire n19706;
wire n19707;
wire n19708;
wire n19709;
wire n19710;
wire n19711;
wire n19712;
wire n19713;
wire n19714;
wire n19715;
wire n19716;
wire n19717;
wire n19718;
wire n19719;
wire n19720;
wire n19721;
wire n19722;
wire n19723;
wire n19724;
wire n19725;
wire n19726;
wire n19727;
wire n19728;
wire n19729;
wire n19730;
wire n19731;
wire n19732;
wire n19733;
wire n19734;
wire n19735;
wire n19736;
wire n19737;
wire n19738;
wire n19739;
wire n1974;
wire n19740;
wire n19741;
wire n19742;
wire n19743;
wire n19744;
wire n19745;
wire n19746;
wire n19747;
wire n19748;
wire n19749;
wire n19750;
wire n19751;
wire n19752;
wire n19753;
wire n19754;
wire n19755;
wire n19756;
wire n19757;
wire n19758;
wire n19759;
wire n19760;
wire n19761;
wire n19762;
wire n19763;
wire n19764;
wire n19765;
wire n19766;
wire n19767;
wire n19768;
wire n19769;
wire n19770;
wire n19771;
wire n19772;
wire n19773;
wire n19774;
wire n19775;
wire n19776;
wire n19777;
wire n19778;
wire n19779;
wire n19780;
wire n19781;
wire n19782;
wire n19783;
wire n19784;
wire n19785;
wire n19786;
wire n19787;
wire n19788;
wire n19789;
wire n1979;
wire n19790;
wire n19791;
wire n19792;
wire n19793;
wire n19794;
wire n19795;
wire n19796;
wire n19797;
wire n19798;
wire n19799;
wire n198;
wire n19800;
wire n19801;
wire n19802;
wire n19803;
wire n19804;
wire n19805;
wire n19806;
wire n19807;
wire n19808;
wire n19809;
wire n19810;
wire n19811;
wire n19812;
wire n19813;
wire n19814;
wire n19815;
wire n19816;
wire n19817;
wire n19818;
wire n19819;
wire n19820;
wire n19821;
wire n19822;
wire n19823;
wire n19824;
wire n19825;
wire n19826;
wire n19827;
wire n19828;
wire n19829;
wire n1983;
wire n19830;
wire n19831;
wire n19832;
wire n19833;
wire n19834;
wire n19835;
wire n19836;
wire n19837;
wire n19838;
wire n19839;
wire n19840;
wire n19841;
wire n19842;
wire n19843;
wire n19844;
wire n19845;
wire n19846;
wire n19847;
wire n19848;
wire n19849;
wire n19850;
wire n19851;
wire n19852;
wire n19853;
wire n19854;
wire n19855;
wire n19856;
wire n19857;
wire n19858;
wire n19859;
wire n19860;
wire n19861;
wire n19862;
wire n19863;
wire n19864;
wire n19865;
wire n19866;
wire n19867;
wire n19868;
wire n19869;
wire n19870;
wire n19871;
wire n19872;
wire n19873;
wire n19874;
wire n19875;
wire n19876;
wire n19877;
wire n19878;
wire n19879;
wire n1988;
wire n19880;
wire n19881;
wire n19882;
wire n19883;
wire n19884;
wire n19885;
wire n19886;
wire n19887;
wire n19888;
wire n19889;
wire n19890;
wire n19891;
wire n19892;
wire n19893;
wire n19894;
wire n19895;
wire n19896;
wire n19897;
wire n19898;
wire n19899;
wire n19900;
wire n19901;
wire n19902;
wire n19903;
wire n19904;
wire n19905;
wire n19906;
wire n19907;
wire n19908;
wire n19909;
wire n19910;
wire n19911;
wire n19912;
wire n19913;
wire n19914;
wire n19915;
wire n19916;
wire n19917;
wire n19918;
wire n19919;
wire n19920;
wire n19921;
wire n19922;
wire n19923;
wire n19924;
wire n19925;
wire n19926;
wire n19927;
wire n19928;
wire n19929;
wire n1993;
wire n19930;
wire n19931;
wire n19932;
wire n19933;
wire n19934;
wire n19935;
wire n19936;
wire n19937;
wire n19938;
wire n19939;
wire n19940;
wire n19941;
wire n19942;
wire n19943;
wire n19944;
wire n19945;
wire n19946;
wire n19947;
wire n19948;
wire n19949;
wire n19950;
wire n19951;
wire n19952;
wire n19953;
wire n19954;
wire n19955;
wire n19956;
wire n19957;
wire n19958;
wire n19959;
wire n19960;
wire n19961;
wire n19962;
wire n19963;
wire n19964;
wire n19965;
wire n19966;
wire n19967;
wire n19968;
wire n19969;
wire n19970;
wire n19971;
wire n19972;
wire n19973;
wire n19974;
wire n19975;
wire n19976;
wire n19977;
wire n19978;
wire n19979;
wire n1998;
wire n19980;
wire n19981;
wire n19982;
wire n19983;
wire n19984;
wire n19985;
wire n19986;
wire n19987;
wire n19988;
wire n19989;
wire n19990;
wire n19991;
wire n19992;
wire n19993;
wire n19994;
wire n19995;
wire n19996;
wire n19997;
wire n19998;
wire n19999;
wire n20000;
wire n20001;
wire n20002;
wire n20003;
wire n20004;
wire n20005;
wire n20006;
wire n20007;
wire n20008;
wire n20009;
wire n20010;
wire n20011;
wire n20012;
wire n20013;
wire n20014;
wire n20015;
wire n20016;
wire n20017;
wire n20018;
wire n20019;
wire n20020;
wire n20021;
wire n20022;
wire n20023;
wire n20024;
wire n20025;
wire n20026;
wire n20027;
wire n20028;
wire n20029;
wire n2003;
wire n20030;
wire n20031;
wire n20032;
wire n20033;
wire n20034;
wire n20035;
wire n20036;
wire n20037;
wire n20038;
wire n20039;
wire n20040;
wire n20041;
wire n20042;
wire n20043;
wire n20044;
wire n20045;
wire n20046;
wire n20047;
wire n20048;
wire n20049;
wire n20050;
wire n20051;
wire n20052;
wire n20053;
wire n20054;
wire n20055;
wire n20056;
wire n20057;
wire n20058;
wire n20059;
wire n20060;
wire n20061;
wire n20062;
wire n20063;
wire n20064;
wire n20065;
wire n20066;
wire n20067;
wire n20068;
wire n20069;
wire n20070;
wire n20071;
wire n20072;
wire n20073;
wire n20074;
wire n20075;
wire n20076;
wire n20077;
wire n20078;
wire n20079;
wire n2008;
wire n20080;
wire n20081;
wire n20082;
wire n20083;
wire n20084;
wire n20085;
wire n20086;
wire n20087;
wire n20088;
wire n20089;
wire n20090;
wire n20091;
wire n20092;
wire n20093;
wire n20094;
wire n20095;
wire n20096;
wire n20097;
wire n20098;
wire n20099;
wire n20100;
wire n20101;
wire n20102;
wire n20103;
wire n20104;
wire n20105;
wire n20106;
wire n20107;
wire n20108;
wire n20109;
wire n20110;
wire n20111;
wire n20112;
wire n20113;
wire n20114;
wire n20115;
wire n20116;
wire n20117;
wire n20118;
wire n20119;
wire n20120;
wire n20121;
wire n20122;
wire n20123;
wire n20124;
wire n20125;
wire n20126;
wire n20127;
wire n20128;
wire n20129;
wire n2013;
wire n20130;
wire n20131;
wire n20132;
wire n20133;
wire n20134;
wire n20135;
wire n20136;
wire n20137;
wire n20138;
wire n20139;
wire n20140;
wire n20141;
wire n20142;
wire n20143;
wire n20144;
wire n20145;
wire n20146;
wire n20147;
wire n20148;
wire n20149;
wire n20150;
wire n20151;
wire n20152;
wire n20153;
wire n20154;
wire n20155;
wire n20156;
wire n20157;
wire n20158;
wire n20159;
wire n20160;
wire n20161;
wire n20162;
wire n20163;
wire n20164;
wire n20165;
wire n20166;
wire n20167;
wire n20168;
wire n20169;
wire n20170;
wire n20171;
wire n20172;
wire n20173;
wire n20174;
wire n20175;
wire n20176;
wire n20177;
wire n20178;
wire n20179;
wire n2018;
wire n20180;
wire n20181;
wire n20182;
wire n20183;
wire n20184;
wire n20185;
wire n20186;
wire n20187;
wire n20188;
wire n20189;
wire n20190;
wire n20191;
wire n20192;
wire n20193;
wire n20194;
wire n20195;
wire n20196;
wire n20197;
wire n20198;
wire n20199;
wire n20200;
wire n20201;
wire n20202;
wire n20203;
wire n20204;
wire n20205;
wire n20206;
wire n20207;
wire n20208;
wire n20209;
wire n20210;
wire n20211;
wire n20212;
wire n20213;
wire n20214;
wire n20215;
wire n20216;
wire n20217;
wire n20218;
wire n20219;
wire n20220;
wire n20221;
wire n20222;
wire n20223;
wire n20224;
wire n20225;
wire n20226;
wire n20227;
wire n20228;
wire n20229;
wire n2023;
wire n20230;
wire n20231;
wire n20232;
wire n20233;
wire n20234;
wire n20235;
wire n20236;
wire n20237;
wire n20238;
wire n20239;
wire n20240;
wire n20241;
wire n20242;
wire n20243;
wire n20244;
wire n20245;
wire n20246;
wire n20247;
wire n20248;
wire n20249;
wire n20250;
wire n20251;
wire n20252;
wire n20253;
wire n20254;
wire n20255;
wire n20256;
wire n20257;
wire n20258;
wire n20259;
wire n20260;
wire n20261;
wire n20262;
wire n20263;
wire n20264;
wire n20265;
wire n20266;
wire n20267;
wire n20268;
wire n20269;
wire n20270;
wire n20271;
wire n20272;
wire n20273;
wire n20274;
wire n20275;
wire n20276;
wire n20277;
wire n20278;
wire n20279;
wire n2028;
wire n20280;
wire n20281;
wire n20282;
wire n20283;
wire n20284;
wire n20285;
wire n20286;
wire n20287;
wire n20288;
wire n20289;
wire n20290;
wire n20291;
wire n20292;
wire n20293;
wire n20294;
wire n20295;
wire n20296;
wire n20297;
wire n20298;
wire n20299;
wire n203;
wire n20300;
wire n20301;
wire n20302;
wire n20303;
wire n20304;
wire n20305;
wire n20306;
wire n20307;
wire n20308;
wire n20309;
wire n20310;
wire n20311;
wire n20312;
wire n20313;
wire n20314;
wire n20315;
wire n20316;
wire n20317;
wire n20318;
wire n20319;
wire n20320;
wire n20321;
wire n20322;
wire n20323;
wire n20324;
wire n20325;
wire n20326;
wire n20327;
wire n20328;
wire n20329;
wire n2033;
wire n20330;
wire n20331;
wire n20332;
wire n20333;
wire n20334;
wire n20335;
wire n20336;
wire n20337;
wire n20338;
wire n20339;
wire n20340;
wire n20341;
wire n20342;
wire n20343;
wire n20344;
wire n20345;
wire n20346;
wire n20347;
wire n20348;
wire n20349;
wire n20350;
wire n20351;
wire n20352;
wire n20353;
wire n20354;
wire n20355;
wire n20356;
wire n20357;
wire n20358;
wire n20359;
wire n20360;
wire n20361;
wire n20362;
wire n20363;
wire n20364;
wire n20365;
wire n20366;
wire n20367;
wire n20368;
wire n20369;
wire n20370;
wire n20371;
wire n20372;
wire n20373;
wire n20374;
wire n20375;
wire n20376;
wire n20377;
wire n20378;
wire n20379;
wire n2038;
wire n20380;
wire n20381;
wire n20382;
wire n20383;
wire n20384;
wire n20385;
wire n20386;
wire n20387;
wire n20388;
wire n20389;
wire n20390;
wire n20391;
wire n20392;
wire n20393;
wire n20394;
wire n20395;
wire n20396;
wire n20397;
wire n20398;
wire n20399;
wire n20400;
wire n20401;
wire n20402;
wire n20403;
wire n20404;
wire n20405;
wire n20406;
wire n20407;
wire n20408;
wire n20409;
wire n20410;
wire n20411;
wire n20412;
wire n20413;
wire n20414;
wire n20415;
wire n20416;
wire n20417;
wire n20418;
wire n20419;
wire n20420;
wire n20421;
wire n20422;
wire n20423;
wire n20424;
wire n20425;
wire n20426;
wire n20427;
wire n20428;
wire n20429;
wire n2043;
wire n20430;
wire n20431;
wire n20432;
wire n20433;
wire n20434;
wire n20435;
wire n20436;
wire n20437;
wire n20438;
wire n20439;
wire n20440;
wire n20441;
wire n20442;
wire n20443;
wire n20444;
wire n20445;
wire n20446;
wire n20447;
wire n20448;
wire n20449;
wire n20450;
wire n20451;
wire n20452;
wire n20453;
wire n20454;
wire n20455;
wire n20456;
wire n20457;
wire n20458;
wire n20459;
wire n20460;
wire n20461;
wire n20462;
wire n20463;
wire n20464;
wire n20465;
wire n20466;
wire n20467;
wire n20468;
wire n20469;
wire n20470;
wire n20471;
wire n20472;
wire n20473;
wire n20474;
wire n20475;
wire n20476;
wire n20477;
wire n20478;
wire n20479;
wire n2048;
wire n20480;
wire n20481;
wire n20482;
wire n20483;
wire n20484;
wire n20485;
wire n20486;
wire n20487;
wire n20488;
wire n20489;
wire n20490;
wire n20491;
wire n20492;
wire n20493;
wire n20494;
wire n20495;
wire n20496;
wire n20497;
wire n20498;
wire n20499;
wire n20500;
wire n20501;
wire n20502;
wire n20503;
wire n20504;
wire n20505;
wire n20506;
wire n20507;
wire n20508;
wire n20509;
wire n20510;
wire n20511;
wire n20512;
wire n20513;
wire n20514;
wire n20515;
wire n20516;
wire n20517;
wire n20518;
wire n20519;
wire n20520;
wire n20521;
wire n20522;
wire n20523;
wire n20524;
wire n20525;
wire n20526;
wire n20527;
wire n20528;
wire n20529;
wire n2053;
wire n20530;
wire n20531;
wire n20532;
wire n20533;
wire n20534;
wire n20535;
wire n20536;
wire n20537;
wire n20538;
wire n20539;
wire n20540;
wire n20541;
wire n20542;
wire n20543;
wire n20544;
wire n20545;
wire n20546;
wire n20547;
wire n20548;
wire n20549;
wire n20550;
wire n20551;
wire n20552;
wire n20553;
wire n20554;
wire n20555;
wire n20556;
wire n20557;
wire n20558;
wire n20559;
wire n20560;
wire n20561;
wire n20562;
wire n20563;
wire n20564;
wire n20565;
wire n20566;
wire n20567;
wire n20568;
wire n20569;
wire n20570;
wire n20571;
wire n20572;
wire n20573;
wire n20574;
wire n20575;
wire n20576;
wire n20577;
wire n20578;
wire n20579;
wire n2058;
wire n20580;
wire n20581;
wire n20582;
wire n20583;
wire n20584;
wire n20585;
wire n20586;
wire n20587;
wire n20588;
wire n20589;
wire n20590;
wire n20591;
wire n20592;
wire n20593;
wire n20594;
wire n20595;
wire n20596;
wire n20597;
wire n20598;
wire n20599;
wire n20600;
wire n20601;
wire n20602;
wire n20603;
wire n20604;
wire n20605;
wire n20606;
wire n20607;
wire n20608;
wire n20609;
wire n20610;
wire n20611;
wire n20612;
wire n20613;
wire n20614;
wire n20615;
wire n20616;
wire n20617;
wire n20618;
wire n20619;
wire n20620;
wire n20621;
wire n20622;
wire n20623;
wire n20624;
wire n20625;
wire n20626;
wire n20627;
wire n20628;
wire n20629;
wire n2063;
wire n20630;
wire n20631;
wire n20632;
wire n20633;
wire n20634;
wire n20635;
wire n20636;
wire n20637;
wire n20638;
wire n20639;
wire n20640;
wire n20641;
wire n20642;
wire n20643;
wire n20644;
wire n20645;
wire n20646;
wire n20647;
wire n20648;
wire n20649;
wire n20650;
wire n20651;
wire n20652;
wire n20653;
wire n20654;
wire n20655;
wire n20656;
wire n20657;
wire n20658;
wire n20659;
wire n20660;
wire n20661;
wire n20662;
wire n20663;
wire n20664;
wire n20665;
wire n20666;
wire n20667;
wire n20668;
wire n20669;
wire n20670;
wire n20671;
wire n20672;
wire n20673;
wire n20674;
wire n20675;
wire n20676;
wire n20677;
wire n20678;
wire n20679;
wire n2068;
wire n20680;
wire n20681;
wire n20682;
wire n20683;
wire n20684;
wire n20685;
wire n20686;
wire n20687;
wire n20688;
wire n20689;
wire n20690;
wire n20691;
wire n20692;
wire n20693;
wire n20694;
wire n20695;
wire n20696;
wire n20697;
wire n20698;
wire n20699;
wire n20700;
wire n20701;
wire n20702;
wire n20703;
wire n20704;
wire n20705;
wire n20706;
wire n20707;
wire n20708;
wire n20709;
wire n20710;
wire n20711;
wire n20712;
wire n20713;
wire n20714;
wire n20715;
wire n20716;
wire n20717;
wire n20718;
wire n20719;
wire n2072;
wire n20720;
wire n20721;
wire n20722;
wire n20723;
wire n20724;
wire n20725;
wire n20726;
wire n20727;
wire n20728;
wire n20729;
wire n20730;
wire n20731;
wire n20732;
wire n20733;
wire n20734;
wire n20735;
wire n20736;
wire n20737;
wire n20738;
wire n20739;
wire n20740;
wire n20741;
wire n20742;
wire n20743;
wire n20744;
wire n20745;
wire n20746;
wire n20747;
wire n20748;
wire n20749;
wire n20750;
wire n20751;
wire n20752;
wire n20753;
wire n20754;
wire n20755;
wire n20756;
wire n20757;
wire n20758;
wire n20759;
wire n20760;
wire n20761;
wire n20762;
wire n20763;
wire n20764;
wire n20765;
wire n20766;
wire n20767;
wire n20768;
wire n20769;
wire n2077;
wire n20770;
wire n20771;
wire n20772;
wire n20773;
wire n20774;
wire n20775;
wire n20776;
wire n20777;
wire n20778;
wire n20779;
wire n20780;
wire n20781;
wire n20782;
wire n20783;
wire n20784;
wire n20785;
wire n20786;
wire n20787;
wire n20788;
wire n20789;
wire n20790;
wire n20791;
wire n20792;
wire n20793;
wire n20794;
wire n20795;
wire n20796;
wire n20797;
wire n20798;
wire n20799;
wire n208;
wire n20800;
wire n20801;
wire n20802;
wire n20803;
wire n20804;
wire n20805;
wire n20806;
wire n20807;
wire n20808;
wire n20809;
wire n20810;
wire n20811;
wire n20812;
wire n20813;
wire n20814;
wire n20815;
wire n20816;
wire n20817;
wire n20818;
wire n20819;
wire n2082;
wire n20820;
wire n20821;
wire n20822;
wire n20823;
wire n20824;
wire n20825;
wire n20826;
wire n20827;
wire n20828;
wire n20829;
wire n20830;
wire n20831;
wire n20832;
wire n20833;
wire n20834;
wire n20835;
wire n20836;
wire n20837;
wire n20838;
wire n20839;
wire n20840;
wire n20841;
wire n20842;
wire n20843;
wire n20844;
wire n20845;
wire n20846;
wire n20847;
wire n20848;
wire n20849;
wire n20850;
wire n20851;
wire n20852;
wire n20853;
wire n20854;
wire n20855;
wire n20856;
wire n20857;
wire n20858;
wire n20859;
wire n20860;
wire n20861;
wire n20862;
wire n20863;
wire n20864;
wire n20865;
wire n20866;
wire n20867;
wire n20868;
wire n20869;
wire n2087;
wire n20870;
wire n20871;
wire n20872;
wire n20873;
wire n20874;
wire n20875;
wire n20876;
wire n20877;
wire n20878;
wire n20879;
wire n20880;
wire n20881;
wire n20882;
wire n20883;
wire n20884;
wire n20885;
wire n20886;
wire n20887;
wire n20888;
wire n20889;
wire n20890;
wire n20891;
wire n20892;
wire n20893;
wire n20894;
wire n20895;
wire n20896;
wire n20897;
wire n20898;
wire n20899;
wire n20900;
wire n20901;
wire n20902;
wire n20903;
wire n20904;
wire n20905;
wire n20906;
wire n20907;
wire n20908;
wire n20909;
wire n20910;
wire n20911;
wire n20912;
wire n20913;
wire n20914;
wire n20915;
wire n20916;
wire n20917;
wire n20918;
wire n20919;
wire n2092;
wire n20920;
wire n20921;
wire n20922;
wire n20923;
wire n20924;
wire n20925;
wire n20926;
wire n20927;
wire n20928;
wire n20929;
wire n20930;
wire n20931;
wire n20932;
wire n20933;
wire n20934;
wire n20935;
wire n20936;
wire n20937;
wire n20938;
wire n20939;
wire n20940;
wire n20941;
wire n20942;
wire n20943;
wire n20944;
wire n20945;
wire n20946;
wire n20947;
wire n20948;
wire n20949;
wire n20950;
wire n20951;
wire n20952;
wire n20953;
wire n20954;
wire n20955;
wire n20956;
wire n20957;
wire n20958;
wire n20959;
wire n20960;
wire n20961;
wire n20962;
wire n20963;
wire n20964;
wire n20965;
wire n20966;
wire n20967;
wire n20968;
wire n20969;
wire n2097;
wire n20970;
wire n20971;
wire n20972;
wire n20973;
wire n20974;
wire n20975;
wire n20976;
wire n20977;
wire n20978;
wire n20979;
wire n20980;
wire n20981;
wire n20982;
wire n20983;
wire n20984;
wire n20985;
wire n20986;
wire n20987;
wire n20988;
wire n20989;
wire n20990;
wire n20991;
wire n20992;
wire n20993;
wire n20994;
wire n20995;
wire n20996;
wire n20997;
wire n20998;
wire n20999;
wire n21000;
wire n21001;
wire n21002;
wire n21003;
wire n21004;
wire n21005;
wire n21006;
wire n21007;
wire n21008;
wire n21009;
wire n21010;
wire n21011;
wire n21012;
wire n21013;
wire n21014;
wire n21015;
wire n21016;
wire n21017;
wire n21018;
wire n21019;
wire n2102;
wire n21020;
wire n21021;
wire n21022;
wire n21023;
wire n21024;
wire n21025;
wire n21026;
wire n21027;
wire n21028;
wire n21029;
wire n21030;
wire n21031;
wire n21032;
wire n21033;
wire n21034;
wire n21035;
wire n21036;
wire n21037;
wire n21038;
wire n21039;
wire n21040;
wire n21041;
wire n21042;
wire n21043;
wire n21044;
wire n21045;
wire n21046;
wire n21047;
wire n21048;
wire n21049;
wire n21050;
wire n21051;
wire n21052;
wire n21053;
wire n21054;
wire n21055;
wire n21056;
wire n21057;
wire n21058;
wire n21059;
wire n21060;
wire n21061;
wire n21062;
wire n21063;
wire n21064;
wire n21065;
wire n21066;
wire n21067;
wire n21068;
wire n21069;
wire n2107;
wire n21070;
wire n21071;
wire n21072;
wire n21073;
wire n21074;
wire n21075;
wire n21076;
wire n21077;
wire n21078;
wire n21079;
wire n21080;
wire n21081;
wire n21082;
wire n21083;
wire n21084;
wire n21085;
wire n21086;
wire n21087;
wire n21088;
wire n21089;
wire n21090;
wire n21091;
wire n21092;
wire n21093;
wire n21094;
wire n21095;
wire n21096;
wire n21097;
wire n21098;
wire n21099;
wire n21100;
wire n21101;
wire n21102;
wire n21103;
wire n21104;
wire n21105;
wire n21106;
wire n21107;
wire n21108;
wire n21109;
wire n21110;
wire n21111;
wire n21112;
wire n21113;
wire n21114;
wire n21115;
wire n21116;
wire n21117;
wire n21118;
wire n21119;
wire n2112;
wire n21120;
wire n21121;
wire n21122;
wire n21123;
wire n21124;
wire n21125;
wire n21126;
wire n21127;
wire n21128;
wire n21129;
wire n21130;
wire n21131;
wire n21132;
wire n21133;
wire n21134;
wire n21135;
wire n21136;
wire n21137;
wire n21138;
wire n21139;
wire n21140;
wire n21141;
wire n21142;
wire n21143;
wire n21144;
wire n21145;
wire n21146;
wire n21147;
wire n21148;
wire n21149;
wire n21150;
wire n21151;
wire n21152;
wire n21153;
wire n21154;
wire n21155;
wire n21156;
wire n21157;
wire n21158;
wire n21159;
wire n21160;
wire n21161;
wire n21162;
wire n21163;
wire n21164;
wire n21165;
wire n21166;
wire n21167;
wire n21168;
wire n21169;
wire n2117;
wire n21170;
wire n21171;
wire n21172;
wire n21173;
wire n21174;
wire n21175;
wire n21176;
wire n21177;
wire n21178;
wire n21179;
wire n21180;
wire n21181;
wire n21182;
wire n21183;
wire n21184;
wire n21185;
wire n21186;
wire n21187;
wire n21188;
wire n21189;
wire n21190;
wire n21191;
wire n21192;
wire n21193;
wire n21194;
wire n21195;
wire n21196;
wire n21197;
wire n21198;
wire n21199;
wire n21200;
wire n21201;
wire n21202;
wire n21203;
wire n21204;
wire n21205;
wire n21206;
wire n21207;
wire n21208;
wire n21209;
wire n2121;
wire n21210;
wire n21211;
wire n21212;
wire n21213;
wire n21214;
wire n21215;
wire n21216;
wire n21217;
wire n21218;
wire n21219;
wire n21220;
wire n21221;
wire n21222;
wire n21223;
wire n21224;
wire n21225;
wire n21226;
wire n21227;
wire n21228;
wire n21229;
wire n21230;
wire n21231;
wire n21232;
wire n21233;
wire n21234;
wire n21235;
wire n21236;
wire n21237;
wire n21238;
wire n21239;
wire n21240;
wire n21241;
wire n21242;
wire n21243;
wire n21244;
wire n21245;
wire n21246;
wire n21247;
wire n21248;
wire n21249;
wire n21250;
wire n21251;
wire n21252;
wire n21253;
wire n21254;
wire n21255;
wire n21256;
wire n21257;
wire n21258;
wire n21259;
wire n2126;
wire n21260;
wire n21261;
wire n21262;
wire n21263;
wire n21264;
wire n21265;
wire n21266;
wire n21267;
wire n21268;
wire n21269;
wire n21270;
wire n21271;
wire n21272;
wire n21273;
wire n21274;
wire n21275;
wire n21276;
wire n21277;
wire n21278;
wire n21279;
wire n21280;
wire n21281;
wire n21282;
wire n21283;
wire n21284;
wire n21285;
wire n21286;
wire n21287;
wire n21288;
wire n21289;
wire n21290;
wire n21291;
wire n21292;
wire n21293;
wire n21294;
wire n21295;
wire n21296;
wire n21297;
wire n21298;
wire n21299;
wire n213;
wire n21300;
wire n21301;
wire n21302;
wire n21303;
wire n21304;
wire n21305;
wire n21306;
wire n21307;
wire n21308;
wire n21309;
wire n2131;
wire n21310;
wire n21311;
wire n21312;
wire n21313;
wire n21314;
wire n21315;
wire n21316;
wire n21317;
wire n21318;
wire n21319;
wire n21320;
wire n21321;
wire n21322;
wire n21323;
wire n21324;
wire n21325;
wire n21326;
wire n21327;
wire n21328;
wire n21329;
wire n21330;
wire n21331;
wire n21332;
wire n21333;
wire n21334;
wire n21335;
wire n21336;
wire n21337;
wire n21339;
wire n21340;
wire n21341;
wire n21342;
wire n21343;
wire n21344;
wire n21345;
wire n21347;
wire n21348;
wire n21349;
wire n21350;
wire n21351;
wire n21352;
wire n21353;
wire n21354;
wire n21355;
wire n21356;
wire n21357;
wire n21358;
wire n21359;
wire n2136;
wire n21360;
wire n21361;
wire n21362;
wire n21363;
wire n21364;
wire n21365;
wire n21366;
wire n21367;
wire n21368;
wire n21369;
wire n21370;
wire n21371;
wire n21372;
wire n21373;
wire n21374;
wire n21375;
wire n21376;
wire n21377;
wire n21378;
wire n21379;
wire n21380;
wire n21381;
wire n21382;
wire n21383;
wire n21384;
wire n21385;
wire n21386;
wire n21387;
wire n21388;
wire n21389;
wire n21390;
wire n21391;
wire n21392;
wire n21393;
wire n21394;
wire n21395;
wire n21396;
wire n21397;
wire n21398;
wire n21399;
wire n21400;
wire n21401;
wire n21402;
wire n21403;
wire n21404;
wire n21405;
wire n21406;
wire n21407;
wire n21408;
wire n21409;
wire n2141;
wire n21410;
wire n21411;
wire n21412;
wire n21413;
wire n21414;
wire n21415;
wire n21416;
wire n21417;
wire n21418;
wire n21419;
wire n21420;
wire n21421;
wire n21422;
wire n21423;
wire n21424;
wire n21425;
wire n21426;
wire n21427;
wire n21428;
wire n21429;
wire n21430;
wire n21431;
wire n21432;
wire n21433;
wire n21434;
wire n21435;
wire n21436;
wire n21437;
wire n21438;
wire n21439;
wire n21440;
wire n21441;
wire n21442;
wire n21443;
wire n21444;
wire n21445;
wire n21446;
wire n21447;
wire n21448;
wire n21449;
wire n21450;
wire n21451;
wire n21452;
wire n21453;
wire n21454;
wire n21455;
wire n21456;
wire n21457;
wire n21458;
wire n21459;
wire n2146;
wire n21460;
wire n21461;
wire n21462;
wire n21463;
wire n21464;
wire n21465;
wire n21466;
wire n21467;
wire n21468;
wire n21469;
wire n21470;
wire n21471;
wire n21472;
wire n21473;
wire n21474;
wire n21475;
wire n21476;
wire n21477;
wire n21478;
wire n21479;
wire n21480;
wire n21481;
wire n21482;
wire n21483;
wire n21484;
wire n21485;
wire n21486;
wire n21487;
wire n21488;
wire n21489;
wire n21490;
wire n21491;
wire n21492;
wire n21493;
wire n21494;
wire n21495;
wire n21496;
wire n21497;
wire n21498;
wire n21499;
wire n21500;
wire n21501;
wire n21502;
wire n21503;
wire n21504;
wire n21505;
wire n21506;
wire n21507;
wire n21508;
wire n21509;
wire n2151;
wire n21510;
wire n21511;
wire n21512;
wire n21513;
wire n21514;
wire n21515;
wire n21516;
wire n21517;
wire n21518;
wire n21519;
wire n21520;
wire n21521;
wire n21522;
wire n21523;
wire n21524;
wire n21525;
wire n21526;
wire n21527;
wire n21528;
wire n21529;
wire n21530;
wire n21531;
wire n21532;
wire n21533;
wire n21534;
wire n21535;
wire n21536;
wire n21537;
wire n21538;
wire n21539;
wire n21540;
wire n21541;
wire n21542;
wire n21543;
wire n21544;
wire n21545;
wire n21546;
wire n21547;
wire n21548;
wire n21549;
wire n2155;
wire n21550;
wire n21551;
wire n21552;
wire n21553;
wire n21554;
wire n21555;
wire n21556;
wire n21557;
wire n21558;
wire n21559;
wire n21560;
wire n21561;
wire n21562;
wire n21563;
wire n21564;
wire n21565;
wire n21566;
wire n21567;
wire n21568;
wire n21569;
wire n21570;
wire n21571;
wire n21572;
wire n21573;
wire n21574;
wire n21575;
wire n21576;
wire n21577;
wire n21578;
wire n21579;
wire n21580;
wire n21581;
wire n21582;
wire n21583;
wire n21584;
wire n21585;
wire n21586;
wire n21587;
wire n21588;
wire n21589;
wire n21590;
wire n21591;
wire n21592;
wire n21593;
wire n21594;
wire n21595;
wire n21596;
wire n21597;
wire n21598;
wire n21599;
wire n2160;
wire n21600;
wire n21601;
wire n21602;
wire n21603;
wire n21604;
wire n21605;
wire n21606;
wire n21607;
wire n21608;
wire n21609;
wire n21610;
wire n21611;
wire n21612;
wire n21613;
wire n21614;
wire n21615;
wire n21616;
wire n21617;
wire n21618;
wire n21619;
wire n21620;
wire n21621;
wire n21622;
wire n21623;
wire n21624;
wire n21626;
wire n21627;
wire n21628;
wire n21629;
wire n21630;
wire n21631;
wire n21632;
wire n21633;
wire n21634;
wire n21635;
wire n21636;
wire n21637;
wire n21638;
wire n21639;
wire n21640;
wire n21641;
wire n21642;
wire n21643;
wire n21644;
wire n21645;
wire n21646;
wire n21647;
wire n21648;
wire n21649;
wire n2165;
wire n21650;
wire n21651;
wire n21652;
wire n21653;
wire n21654;
wire n21655;
wire n21656;
wire n21657;
wire n21658;
wire n21659;
wire n21660;
wire n21661;
wire n21662;
wire n21663;
wire n21664;
wire n21665;
wire n21666;
wire n21667;
wire n21668;
wire n21669;
wire n21670;
wire n21671;
wire n21672;
wire n21673;
wire n21674;
wire n21675;
wire n21676;
wire n21677;
wire n21678;
wire n21679;
wire n21680;
wire n21681;
wire n21682;
wire n21683;
wire n21684;
wire n21685;
wire n21686;
wire n21687;
wire n21688;
wire n21689;
wire n2169;
wire n21690;
wire n21691;
wire n21692;
wire n21693;
wire n21694;
wire n21695;
wire n21696;
wire n21697;
wire n21698;
wire n21699;
wire n21700;
wire n21701;
wire n21702;
wire n21703;
wire n21704;
wire n21705;
wire n21706;
wire n21707;
wire n21708;
wire n21709;
wire n21710;
wire n21711;
wire n21712;
wire n21713;
wire n21714;
wire n21715;
wire n21716;
wire n21717;
wire n21718;
wire n21719;
wire n21720;
wire n21721;
wire n21722;
wire n21723;
wire n21724;
wire n21725;
wire n21726;
wire n21727;
wire n21728;
wire n21729;
wire n21730;
wire n21731;
wire n21732;
wire n21733;
wire n21734;
wire n21735;
wire n21736;
wire n21737;
wire n21738;
wire n21739;
wire n2174;
wire n21740;
wire n21741;
wire n21742;
wire n21743;
wire n21744;
wire n21745;
wire n21746;
wire n21747;
wire n21748;
wire n21749;
wire n21750;
wire n21751;
wire n21752;
wire n21753;
wire n21754;
wire n21755;
wire n21756;
wire n21757;
wire n21758;
wire n21759;
wire n21760;
wire n21761;
wire n21762;
wire n21763;
wire n21764;
wire n21765;
wire n21766;
wire n21767;
wire n21768;
wire n21769;
wire n21770;
wire n21771;
wire n21772;
wire n21773;
wire n21774;
wire n21775;
wire n21776;
wire n21777;
wire n21778;
wire n21779;
wire n21780;
wire n21781;
wire n21782;
wire n21783;
wire n21784;
wire n21785;
wire n21786;
wire n21787;
wire n21788;
wire n21789;
wire n2179;
wire n21790;
wire n21791;
wire n21792;
wire n21793;
wire n21794;
wire n21795;
wire n21796;
wire n21797;
wire n21798;
wire n21799;
wire n218;
wire n21800;
wire n21801;
wire n21802;
wire n21803;
wire n21804;
wire n21805;
wire n21806;
wire n21807;
wire n21808;
wire n21809;
wire n21810;
wire n21811;
wire n21812;
wire n21813;
wire n21814;
wire n21815;
wire n21816;
wire n21817;
wire n21818;
wire n21819;
wire n21820;
wire n21821;
wire n21822;
wire n21823;
wire n21824;
wire n21825;
wire n21826;
wire n21827;
wire n21828;
wire n21829;
wire n21830;
wire n21831;
wire n21832;
wire n21833;
wire n21834;
wire n21835;
wire n21836;
wire n21837;
wire n21838;
wire n21839;
wire n2184;
wire n21840;
wire n21841;
wire n21842;
wire n21843;
wire n21844;
wire n21845;
wire n21846;
wire n21847;
wire n21848;
wire n21849;
wire n21850;
wire n21851;
wire n21852;
wire n21853;
wire n21854;
wire n21855;
wire n21856;
wire n21857;
wire n21858;
wire n21859;
wire n21860;
wire n21861;
wire n21862;
wire n21863;
wire n21864;
wire n21865;
wire n21866;
wire n21867;
wire n21868;
wire n21869;
wire n21870;
wire n21871;
wire n21872;
wire n21873;
wire n21874;
wire n21875;
wire n21876;
wire n21877;
wire n21878;
wire n21879;
wire n21880;
wire n21881;
wire n21882;
wire n21883;
wire n21884;
wire n21885;
wire n21886;
wire n21887;
wire n21888;
wire n21889;
wire n2189;
wire n21890;
wire n21891;
wire n21892;
wire n21893;
wire n21894;
wire n21895;
wire n21896;
wire n21897;
wire n21898;
wire n21899;
wire n21900;
wire n21901;
wire n21902;
wire n21903;
wire n21904;
wire n21905;
wire n21906;
wire n21907;
wire n21908;
wire n21909;
wire n21910;
wire n21911;
wire n21912;
wire n21913;
wire n21914;
wire n21915;
wire n21916;
wire n21917;
wire n21918;
wire n21919;
wire n21920;
wire n21921;
wire n21922;
wire n21923;
wire n21924;
wire n21925;
wire n21926;
wire n21927;
wire n21928;
wire n21929;
wire n21930;
wire n21931;
wire n21932;
wire n21933;
wire n21934;
wire n21935;
wire n21936;
wire n21937;
wire n21938;
wire n21939;
wire n2194;
wire n21940;
wire n21941;
wire n21942;
wire n21943;
wire n21944;
wire n21945;
wire n21946;
wire n21947;
wire n21948;
wire n21949;
wire n21950;
wire n21951;
wire n21952;
wire n21953;
wire n21954;
wire n21955;
wire n21956;
wire n21957;
wire n21958;
wire n21959;
wire n21960;
wire n21961;
wire n21962;
wire n21963;
wire n21964;
wire n21965;
wire n21966;
wire n21967;
wire n21968;
wire n21969;
wire n21970;
wire n21971;
wire n21972;
wire n21973;
wire n21974;
wire n21975;
wire n21976;
wire n21977;
wire n21978;
wire n21979;
wire n2198;
wire n21980;
wire n21981;
wire n21982;
wire n21983;
wire n21984;
wire n21985;
wire n21986;
wire n21987;
wire n21988;
wire n21989;
wire n21990;
wire n21991;
wire n21992;
wire n21993;
wire n21994;
wire n21995;
wire n21996;
wire n21997;
wire n21998;
wire n21999;
wire n22000;
wire n22001;
wire n22002;
wire n22003;
wire n22004;
wire n22005;
wire n22006;
wire n22007;
wire n22008;
wire n22009;
wire n22010;
wire n22011;
wire n22012;
wire n22013;
wire n22014;
wire n22015;
wire n22016;
wire n22017;
wire n22018;
wire n22019;
wire n22020;
wire n22021;
wire n22022;
wire n22023;
wire n22024;
wire n22025;
wire n22026;
wire n22027;
wire n22028;
wire n22029;
wire n2203;
wire n22030;
wire n22031;
wire n22032;
wire n22033;
wire n22034;
wire n22035;
wire n22036;
wire n22037;
wire n22038;
wire n22039;
wire n22040;
wire n22041;
wire n22042;
wire n22043;
wire n22044;
wire n22045;
wire n22046;
wire n22047;
wire n22048;
wire n22049;
wire n22050;
wire n22051;
wire n22052;
wire n22053;
wire n22054;
wire n22055;
wire n22056;
wire n22057;
wire n22058;
wire n22059;
wire n22060;
wire n22061;
wire n22062;
wire n22063;
wire n22064;
wire n22065;
wire n22066;
wire n22067;
wire n22068;
wire n22069;
wire n22070;
wire n22071;
wire n22072;
wire n22073;
wire n22074;
wire n22075;
wire n22076;
wire n22077;
wire n22078;
wire n22079;
wire n2208;
wire n22080;
wire n22081;
wire n22082;
wire n22083;
wire n22084;
wire n22085;
wire n22086;
wire n22087;
wire n22088;
wire n22089;
wire n22090;
wire n22091;
wire n22092;
wire n22093;
wire n22094;
wire n22095;
wire n22096;
wire n22097;
wire n22098;
wire n22099;
wire n22100;
wire n22101;
wire n22102;
wire n22103;
wire n22104;
wire n22105;
wire n22106;
wire n22107;
wire n22108;
wire n22109;
wire n22110;
wire n22111;
wire n22112;
wire n22113;
wire n22114;
wire n22115;
wire n22116;
wire n22117;
wire n22118;
wire n22119;
wire n22120;
wire n22121;
wire n22122;
wire n22123;
wire n22124;
wire n22125;
wire n22126;
wire n22127;
wire n22128;
wire n22129;
wire n2213;
wire n22130;
wire n22131;
wire n22132;
wire n22133;
wire n22134;
wire n22135;
wire n22136;
wire n22137;
wire n22138;
wire n22139;
wire n22140;
wire n22141;
wire n22142;
wire n22143;
wire n22144;
wire n22145;
wire n22146;
wire n22147;
wire n22148;
wire n22149;
wire n22150;
wire n22151;
wire n22152;
wire n22153;
wire n22154;
wire n22155;
wire n22156;
wire n22157;
wire n22158;
wire n22159;
wire n22160;
wire n22161;
wire n22162;
wire n22163;
wire n22164;
wire n22165;
wire n22166;
wire n22167;
wire n22168;
wire n22169;
wire n22170;
wire n22171;
wire n22172;
wire n22173;
wire n22174;
wire n22175;
wire n22176;
wire n22177;
wire n22178;
wire n22179;
wire n2218;
wire n22180;
wire n22181;
wire n22182;
wire n22183;
wire n22184;
wire n22185;
wire n22186;
wire n22187;
wire n22188;
wire n22189;
wire n22190;
wire n22191;
wire n22192;
wire n22193;
wire n22194;
wire n22195;
wire n22196;
wire n22197;
wire n22198;
wire n22199;
wire n22200;
wire n22201;
wire n22202;
wire n22203;
wire n22204;
wire n22205;
wire n22206;
wire n22207;
wire n22208;
wire n22209;
wire n22210;
wire n22211;
wire n22212;
wire n22213;
wire n22214;
wire n22215;
wire n22216;
wire n22217;
wire n22218;
wire n22219;
wire n22220;
wire n22221;
wire n22222;
wire n22223;
wire n22224;
wire n22225;
wire n22226;
wire n22227;
wire n22228;
wire n22229;
wire n2223;
wire n22230;
wire n22231;
wire n22232;
wire n22233;
wire n22234;
wire n22235;
wire n22236;
wire n22237;
wire n22238;
wire n22239;
wire n22240;
wire n22241;
wire n22242;
wire n22243;
wire n22244;
wire n22245;
wire n22246;
wire n22247;
wire n22248;
wire n22249;
wire n22250;
wire n22251;
wire n22252;
wire n22253;
wire n22254;
wire n22255;
wire n22256;
wire n22257;
wire n22258;
wire n22259;
wire n22260;
wire n22261;
wire n22262;
wire n22263;
wire n22264;
wire n22265;
wire n22266;
wire n22267;
wire n22268;
wire n22269;
wire n2227;
wire n22270;
wire n22271;
wire n22272;
wire n22273;
wire n22274;
wire n22275;
wire n22276;
wire n22277;
wire n22278;
wire n22279;
wire n22280;
wire n22281;
wire n22282;
wire n22283;
wire n22284;
wire n22285;
wire n22286;
wire n22287;
wire n22288;
wire n22289;
wire n22290;
wire n22291;
wire n22292;
wire n22293;
wire n22294;
wire n22295;
wire n22296;
wire n22297;
wire n22298;
wire n22299;
wire n223;
wire n22300;
wire n22301;
wire n22302;
wire n22303;
wire n22304;
wire n22305;
wire n22306;
wire n22307;
wire n22308;
wire n22309;
wire n22310;
wire n22311;
wire n22312;
wire n22313;
wire n22314;
wire n22315;
wire n22316;
wire n22317;
wire n22318;
wire n22319;
wire n2232;
wire n22320;
wire n22321;
wire n22322;
wire n22323;
wire n22324;
wire n22325;
wire n22326;
wire n22327;
wire n22328;
wire n22329;
wire n22330;
wire n22331;
wire n22332;
wire n22333;
wire n22334;
wire n22335;
wire n22336;
wire n22337;
wire n22338;
wire n22339;
wire n22340;
wire n22341;
wire n22342;
wire n22343;
wire n22344;
wire n22345;
wire n22346;
wire n22347;
wire n22348;
wire n22349;
wire n22350;
wire n22351;
wire n22352;
wire n22353;
wire n22354;
wire n22355;
wire n22356;
wire n22357;
wire n22358;
wire n22359;
wire n22360;
wire n22361;
wire n22362;
wire n22363;
wire n22364;
wire n22365;
wire n22366;
wire n22367;
wire n22368;
wire n22369;
wire n2237;
wire n22370;
wire n22371;
wire n22372;
wire n22373;
wire n22374;
wire n22375;
wire n22376;
wire n22377;
wire n22378;
wire n22379;
wire n22380;
wire n22381;
wire n22382;
wire n22383;
wire n22384;
wire n22385;
wire n22386;
wire n22387;
wire n22388;
wire n22389;
wire n22390;
wire n22391;
wire n22392;
wire n22393;
wire n22394;
wire n22395;
wire n22396;
wire n22397;
wire n22398;
wire n22399;
wire n22400;
wire n22401;
wire n22402;
wire n22403;
wire n22404;
wire n22405;
wire n22406;
wire n22407;
wire n22408;
wire n22409;
wire n22410;
wire n22411;
wire n22412;
wire n22413;
wire n22414;
wire n22415;
wire n22416;
wire n22417;
wire n22418;
wire n22419;
wire n2242;
wire n22420;
wire n22421;
wire n22422;
wire n22423;
wire n22424;
wire n22425;
wire n22426;
wire n22427;
wire n22428;
wire n22429;
wire n22430;
wire n22431;
wire n22432;
wire n22433;
wire n22434;
wire n22435;
wire n22436;
wire n22437;
wire n22438;
wire n22439;
wire n22440;
wire n22441;
wire n22442;
wire n22443;
wire n22444;
wire n22445;
wire n22446;
wire n22447;
wire n22448;
wire n22449;
wire n22450;
wire n22451;
wire n22452;
wire n22453;
wire n22454;
wire n22455;
wire n22456;
wire n22457;
wire n22458;
wire n22459;
wire n22460;
wire n22461;
wire n22462;
wire n22463;
wire n22464;
wire n22465;
wire n22466;
wire n22467;
wire n22468;
wire n22469;
wire n2247;
wire n22470;
wire n22471;
wire n22472;
wire n22473;
wire n22474;
wire n22475;
wire n22476;
wire n22477;
wire n22478;
wire n22479;
wire n22480;
wire n22481;
wire n22482;
wire n22483;
wire n22484;
wire n22485;
wire n22486;
wire n22487;
wire n22488;
wire n22489;
wire n22490;
wire n22492;
wire n22493;
wire n22494;
wire n22495;
wire n22496;
wire n22497;
wire n22498;
wire n22499;
wire n22500;
wire n22501;
wire n22502;
wire n22503;
wire n22504;
wire n22505;
wire n22506;
wire n22507;
wire n22508;
wire n22509;
wire n22510;
wire n22511;
wire n22512;
wire n22513;
wire n22514;
wire n22515;
wire n22516;
wire n22517;
wire n22518;
wire n22519;
wire n2252;
wire n22520;
wire n22521;
wire n22522;
wire n22523;
wire n22524;
wire n22525;
wire n22526;
wire n22527;
wire n22528;
wire n22529;
wire n22530;
wire n22531;
wire n22532;
wire n22533;
wire n22534;
wire n22535;
wire n22536;
wire n22537;
wire n22538;
wire n22539;
wire n22540;
wire n22541;
wire n22542;
wire n22543;
wire n22544;
wire n22545;
wire n22546;
wire n22547;
wire n22548;
wire n22549;
wire n22550;
wire n22551;
wire n22552;
wire n22553;
wire n22554;
wire n22555;
wire n22556;
wire n22557;
wire n22558;
wire n22559;
wire n22560;
wire n22561;
wire n22562;
wire n22563;
wire n22565;
wire n22566;
wire n22567;
wire n22568;
wire n22569;
wire n2257;
wire n22570;
wire n22571;
wire n22572;
wire n22573;
wire n22574;
wire n22575;
wire n22576;
wire n22577;
wire n22578;
wire n22579;
wire n22580;
wire n22581;
wire n22582;
wire n22583;
wire n22584;
wire n22585;
wire n22586;
wire n22587;
wire n22588;
wire n22589;
wire n22590;
wire n22591;
wire n22592;
wire n22593;
wire n22594;
wire n22595;
wire n22596;
wire n22597;
wire n22598;
wire n22599;
wire n22600;
wire n22601;
wire n22602;
wire n22603;
wire n22604;
wire n22605;
wire n22606;
wire n22607;
wire n22608;
wire n22609;
wire n22610;
wire n22611;
wire n22612;
wire n22613;
wire n22614;
wire n22615;
wire n22616;
wire n22617;
wire n22618;
wire n22619;
wire n2262;
wire n22620;
wire n22621;
wire n22622;
wire n22623;
wire n22624;
wire n22625;
wire n22626;
wire n22627;
wire n22628;
wire n22629;
wire n22630;
wire n22631;
wire n22632;
wire n22633;
wire n22634;
wire n22635;
wire n22636;
wire n22637;
wire n22638;
wire n22639;
wire n22640;
wire n22641;
wire n22642;
wire n22643;
wire n22644;
wire n22645;
wire n22646;
wire n22647;
wire n22648;
wire n22649;
wire n22650;
wire n22651;
wire n22652;
wire n22653;
wire n22654;
wire n22655;
wire n22656;
wire n22657;
wire n22658;
wire n22659;
wire n22660;
wire n22661;
wire n22662;
wire n22663;
wire n22664;
wire n22665;
wire n22666;
wire n22667;
wire n22668;
wire n22669;
wire n2267;
wire n22670;
wire n22671;
wire n22672;
wire n22673;
wire n22674;
wire n22675;
wire n22676;
wire n22677;
wire n22678;
wire n22679;
wire n22680;
wire n22681;
wire n22682;
wire n22683;
wire n22684;
wire n22685;
wire n22686;
wire n22687;
wire n22688;
wire n22689;
wire n22690;
wire n22691;
wire n22692;
wire n22693;
wire n22694;
wire n22695;
wire n22696;
wire n22697;
wire n22698;
wire n22699;
wire n22700;
wire n22701;
wire n22702;
wire n22703;
wire n22704;
wire n22705;
wire n22706;
wire n22707;
wire n22708;
wire n22709;
wire n22710;
wire n22711;
wire n22712;
wire n22713;
wire n22714;
wire n22715;
wire n22716;
wire n22717;
wire n22718;
wire n22719;
wire n2272;
wire n22720;
wire n22721;
wire n22722;
wire n22723;
wire n22724;
wire n22725;
wire n22726;
wire n22727;
wire n22728;
wire n22729;
wire n22730;
wire n22731;
wire n22732;
wire n22733;
wire n22734;
wire n22735;
wire n22736;
wire n22737;
wire n22738;
wire n22739;
wire n22740;
wire n22741;
wire n22742;
wire n22743;
wire n22744;
wire n22745;
wire n22746;
wire n22747;
wire n22748;
wire n22749;
wire n22750;
wire n22751;
wire n22752;
wire n22753;
wire n22754;
wire n22755;
wire n22756;
wire n22758;
wire n22759;
wire n22760;
wire n22761;
wire n22762;
wire n22763;
wire n22764;
wire n22765;
wire n22767;
wire n22768;
wire n22769;
wire n2277;
wire n22770;
wire n22771;
wire n22772;
wire n22773;
wire n22774;
wire n22775;
wire n22776;
wire n22777;
wire n22778;
wire n22779;
wire n22780;
wire n22781;
wire n22782;
wire n22783;
wire n22784;
wire n22785;
wire n22786;
wire n22787;
wire n22788;
wire n22789;
wire n22790;
wire n22791;
wire n22792;
wire n22793;
wire n22794;
wire n22795;
wire n22796;
wire n22797;
wire n22798;
wire n22799;
wire n228;
wire n22800;
wire n22801;
wire n22802;
wire n22803;
wire n22804;
wire n22805;
wire n22806;
wire n22807;
wire n22808;
wire n22809;
wire n22810;
wire n22811;
wire n22812;
wire n22813;
wire n22814;
wire n22815;
wire n22816;
wire n22817;
wire n22818;
wire n22819;
wire n2282;
wire n22820;
wire n22821;
wire n22822;
wire n22823;
wire n22824;
wire n22825;
wire n22826;
wire n22827;
wire n22828;
wire n22829;
wire n22830;
wire n22831;
wire n22832;
wire n22833;
wire n22834;
wire n22835;
wire n22836;
wire n22837;
wire n22838;
wire n22839;
wire n22840;
wire n22841;
wire n22842;
wire n22843;
wire n22844;
wire n22845;
wire n22846;
wire n22847;
wire n22848;
wire n22849;
wire n22850;
wire n22851;
wire n22852;
wire n22853;
wire n22854;
wire n22855;
wire n22856;
wire n22857;
wire n22858;
wire n22859;
wire n22860;
wire n22861;
wire n22862;
wire n22863;
wire n22864;
wire n22865;
wire n22866;
wire n22867;
wire n22868;
wire n22869;
wire n2287;
wire n22870;
wire n22871;
wire n22872;
wire n22873;
wire n22874;
wire n22875;
wire n22876;
wire n22877;
wire n22878;
wire n22879;
wire n22880;
wire n22881;
wire n22882;
wire n22883;
wire n22884;
wire n22885;
wire n22886;
wire n22887;
wire n22888;
wire n22889;
wire n22890;
wire n22891;
wire n22892;
wire n22893;
wire n22894;
wire n22895;
wire n22896;
wire n22897;
wire n22898;
wire n22899;
wire n22900;
wire n22901;
wire n22902;
wire n22903;
wire n22904;
wire n22905;
wire n22906;
wire n22907;
wire n22908;
wire n22909;
wire n22910;
wire n22911;
wire n22912;
wire n22913;
wire n22914;
wire n22915;
wire n22916;
wire n22917;
wire n22918;
wire n22919;
wire n2292;
wire n22920;
wire n22921;
wire n22922;
wire n22923;
wire n22924;
wire n22925;
wire n22926;
wire n22927;
wire n22928;
wire n22929;
wire n22930;
wire n22931;
wire n22932;
wire n22933;
wire n22934;
wire n22935;
wire n22936;
wire n22937;
wire n22938;
wire n22939;
wire n22940;
wire n22941;
wire n22942;
wire n22943;
wire n22944;
wire n22945;
wire n22946;
wire n22947;
wire n22948;
wire n22949;
wire n22950;
wire n22951;
wire n22952;
wire n22953;
wire n22954;
wire n22955;
wire n22956;
wire n22957;
wire n22958;
wire n22959;
wire n22960;
wire n22961;
wire n22962;
wire n22963;
wire n22964;
wire n22965;
wire n22966;
wire n22967;
wire n22968;
wire n22969;
wire n2297;
wire n22970;
wire n22971;
wire n22972;
wire n22973;
wire n22974;
wire n22975;
wire n22976;
wire n22977;
wire n22978;
wire n22979;
wire n22980;
wire n22981;
wire n22982;
wire n22983;
wire n22984;
wire n22985;
wire n22986;
wire n22987;
wire n22988;
wire n22989;
wire n22990;
wire n22991;
wire n22992;
wire n22993;
wire n22994;
wire n22995;
wire n22996;
wire n22997;
wire n22998;
wire n22999;
wire n23000;
wire n23001;
wire n23002;
wire n23003;
wire n23004;
wire n23005;
wire n23006;
wire n23007;
wire n23008;
wire n23009;
wire n23010;
wire n23011;
wire n23012;
wire n23013;
wire n23014;
wire n23015;
wire n23016;
wire n23017;
wire n23018;
wire n23019;
wire n2302;
wire n23020;
wire n23021;
wire n23022;
wire n23023;
wire n23024;
wire n23025;
wire n23026;
wire n23027;
wire n23028;
wire n23029;
wire n23030;
wire n23031;
wire n23032;
wire n23033;
wire n23034;
wire n23035;
wire n23036;
wire n23037;
wire n23038;
wire n23039;
wire n23040;
wire n23041;
wire n23042;
wire n23043;
wire n23044;
wire n23045;
wire n23046;
wire n23047;
wire n23048;
wire n23049;
wire n23050;
wire n23051;
wire n23052;
wire n23053;
wire n23054;
wire n23055;
wire n23056;
wire n23057;
wire n23058;
wire n23059;
wire n23060;
wire n23061;
wire n23062;
wire n23063;
wire n23064;
wire n23065;
wire n23066;
wire n23067;
wire n23068;
wire n23069;
wire n2307;
wire n23070;
wire n23071;
wire n23072;
wire n23073;
wire n23074;
wire n23075;
wire n23076;
wire n23077;
wire n23078;
wire n23079;
wire n23080;
wire n23081;
wire n23082;
wire n23083;
wire n23084;
wire n23085;
wire n23086;
wire n23087;
wire n23088;
wire n23089;
wire n23090;
wire n23091;
wire n23092;
wire n23093;
wire n23094;
wire n23095;
wire n23096;
wire n23097;
wire n23098;
wire n23099;
wire n23100;
wire n23101;
wire n23102;
wire n23103;
wire n23104;
wire n23105;
wire n23106;
wire n23107;
wire n23108;
wire n23109;
wire n23110;
wire n23111;
wire n23112;
wire n23113;
wire n23114;
wire n23115;
wire n23116;
wire n23117;
wire n23118;
wire n23119;
wire n2312;
wire n23120;
wire n23121;
wire n23122;
wire n23123;
wire n23124;
wire n23125;
wire n23126;
wire n23127;
wire n23128;
wire n23129;
wire n23130;
wire n23131;
wire n23132;
wire n23133;
wire n23134;
wire n23135;
wire n23136;
wire n23137;
wire n23138;
wire n23139;
wire n23140;
wire n23141;
wire n23142;
wire n23143;
wire n23144;
wire n23145;
wire n23146;
wire n23147;
wire n23148;
wire n23149;
wire n23150;
wire n23151;
wire n23152;
wire n23153;
wire n23154;
wire n23155;
wire n23156;
wire n23157;
wire n23158;
wire n23159;
wire n23160;
wire n23161;
wire n23162;
wire n23163;
wire n23164;
wire n23165;
wire n23166;
wire n23167;
wire n23168;
wire n23169;
wire n2317;
wire n23170;
wire n23171;
wire n23172;
wire n23173;
wire n23174;
wire n23175;
wire n23176;
wire n23177;
wire n23178;
wire n23179;
wire n23180;
wire n23181;
wire n23182;
wire n23183;
wire n23184;
wire n23185;
wire n23186;
wire n23187;
wire n23188;
wire n23189;
wire n23190;
wire n23191;
wire n23192;
wire n23193;
wire n23194;
wire n23195;
wire n23196;
wire n23197;
wire n23198;
wire n23199;
wire n23200;
wire n23201;
wire n23202;
wire n23203;
wire n23204;
wire n23205;
wire n23206;
wire n23207;
wire n23208;
wire n23209;
wire n23210;
wire n23211;
wire n23212;
wire n23213;
wire n23214;
wire n23215;
wire n23216;
wire n23217;
wire n23218;
wire n23219;
wire n2322;
wire n23220;
wire n23221;
wire n23222;
wire n23223;
wire n23224;
wire n23225;
wire n23226;
wire n23227;
wire n23228;
wire n23229;
wire n23230;
wire n23231;
wire n23232;
wire n23233;
wire n23234;
wire n23235;
wire n23236;
wire n23237;
wire n23238;
wire n23239;
wire n23240;
wire n23241;
wire n23242;
wire n23243;
wire n23244;
wire n23245;
wire n23246;
wire n23247;
wire n23248;
wire n23249;
wire n23250;
wire n23251;
wire n23252;
wire n23253;
wire n23254;
wire n23255;
wire n23256;
wire n23257;
wire n23258;
wire n23259;
wire n23260;
wire n23261;
wire n23262;
wire n23263;
wire n23264;
wire n23265;
wire n23266;
wire n23267;
wire n23268;
wire n23269;
wire n2327;
wire n23270;
wire n23271;
wire n23272;
wire n23273;
wire n23274;
wire n23275;
wire n23276;
wire n23277;
wire n23278;
wire n23279;
wire n23280;
wire n23281;
wire n23282;
wire n23283;
wire n23284;
wire n23285;
wire n23286;
wire n23287;
wire n23288;
wire n23289;
wire n23290;
wire n23291;
wire n23292;
wire n23293;
wire n23294;
wire n23295;
wire n23296;
wire n23297;
wire n23298;
wire n23299;
wire n233;
wire n23300;
wire n23301;
wire n23302;
wire n23303;
wire n23304;
wire n23305;
wire n23306;
wire n23307;
wire n23308;
wire n23309;
wire n23310;
wire n23311;
wire n23312;
wire n23313;
wire n23314;
wire n23315;
wire n23316;
wire n23317;
wire n23318;
wire n23319;
wire n2332;
wire n23320;
wire n23321;
wire n23322;
wire n23323;
wire n23324;
wire n23325;
wire n23326;
wire n23327;
wire n23328;
wire n23329;
wire n23330;
wire n23331;
wire n23332;
wire n23333;
wire n23334;
wire n23335;
wire n23336;
wire n23337;
wire n23338;
wire n23339;
wire n23340;
wire n23341;
wire n23342;
wire n23343;
wire n23344;
wire n23345;
wire n23346;
wire n23347;
wire n23348;
wire n23349;
wire n23350;
wire n23351;
wire n23352;
wire n23353;
wire n23354;
wire n23355;
wire n23356;
wire n23357;
wire n23359;
wire n23360;
wire n23361;
wire n23362;
wire n23363;
wire n23364;
wire n23365;
wire n23366;
wire n23367;
wire n23368;
wire n23369;
wire n2337;
wire n23370;
wire n23371;
wire n23372;
wire n23373;
wire n23374;
wire n23375;
wire n23376;
wire n23377;
wire n23378;
wire n23379;
wire n23380;
wire n23381;
wire n23382;
wire n23383;
wire n23384;
wire n23385;
wire n23386;
wire n23387;
wire n23388;
wire n23389;
wire n23390;
wire n23391;
wire n23392;
wire n23393;
wire n23394;
wire n23395;
wire n23396;
wire n23397;
wire n23398;
wire n23399;
wire n23400;
wire n23401;
wire n23402;
wire n23403;
wire n23404;
wire n23405;
wire n23406;
wire n23407;
wire n23408;
wire n23409;
wire n23410;
wire n23411;
wire n23412;
wire n23413;
wire n23414;
wire n23415;
wire n23416;
wire n23417;
wire n23418;
wire n23419;
wire n2342;
wire n23420;
wire n23421;
wire n23422;
wire n23423;
wire n23424;
wire n23425;
wire n23426;
wire n23427;
wire n23428;
wire n23429;
wire n23430;
wire n23431;
wire n23432;
wire n23433;
wire n23434;
wire n23435;
wire n23436;
wire n23437;
wire n23438;
wire n23439;
wire n23440;
wire n23441;
wire n23442;
wire n23443;
wire n23444;
wire n23445;
wire n23446;
wire n23447;
wire n23448;
wire n23449;
wire n23450;
wire n23451;
wire n23452;
wire n23453;
wire n23454;
wire n23455;
wire n23456;
wire n23457;
wire n23458;
wire n23459;
wire n23460;
wire n23461;
wire n23462;
wire n23463;
wire n23464;
wire n23465;
wire n23466;
wire n23467;
wire n23468;
wire n23469;
wire n2347;
wire n23470;
wire n23471;
wire n23472;
wire n23473;
wire n23474;
wire n23475;
wire n23476;
wire n23477;
wire n23478;
wire n23479;
wire n23480;
wire n23481;
wire n23482;
wire n23483;
wire n23484;
wire n23485;
wire n23486;
wire n23487;
wire n23488;
wire n23489;
wire n23490;
wire n23491;
wire n23492;
wire n23493;
wire n23494;
wire n23495;
wire n23496;
wire n23497;
wire n23498;
wire n23499;
wire n23500;
wire n23501;
wire n23502;
wire n23503;
wire n23504;
wire n23505;
wire n23506;
wire n23507;
wire n23508;
wire n23509;
wire n23510;
wire n23511;
wire n23512;
wire n23513;
wire n23514;
wire n23515;
wire n23516;
wire n23517;
wire n23518;
wire n23519;
wire n2352;
wire n23520;
wire n23521;
wire n23522;
wire n23523;
wire n23524;
wire n23525;
wire n23526;
wire n23527;
wire n23528;
wire n23529;
wire n23530;
wire n23531;
wire n23532;
wire n23533;
wire n23534;
wire n23535;
wire n23536;
wire n23537;
wire n23538;
wire n23539;
wire n23540;
wire n23541;
wire n23542;
wire n23543;
wire n23544;
wire n23545;
wire n23546;
wire n23547;
wire n23548;
wire n23549;
wire n23550;
wire n23551;
wire n23552;
wire n23553;
wire n23554;
wire n23555;
wire n23556;
wire n23557;
wire n23558;
wire n23559;
wire n23560;
wire n23561;
wire n23562;
wire n23563;
wire n23564;
wire n23565;
wire n23566;
wire n23567;
wire n23568;
wire n23569;
wire n2357;
wire n23570;
wire n23571;
wire n23572;
wire n23573;
wire n23574;
wire n23575;
wire n23576;
wire n23577;
wire n23578;
wire n23579;
wire n23580;
wire n23581;
wire n23582;
wire n23583;
wire n23584;
wire n23585;
wire n23586;
wire n23587;
wire n23588;
wire n23589;
wire n23590;
wire n23591;
wire n23592;
wire n23593;
wire n23594;
wire n23595;
wire n23596;
wire n23597;
wire n23598;
wire n23599;
wire n23600;
wire n23601;
wire n23602;
wire n23603;
wire n23604;
wire n23605;
wire n23606;
wire n23607;
wire n23608;
wire n23609;
wire n23610;
wire n23611;
wire n23612;
wire n23613;
wire n23614;
wire n23615;
wire n23616;
wire n23617;
wire n23618;
wire n23619;
wire n2362;
wire n23620;
wire n23621;
wire n23622;
wire n23623;
wire n23624;
wire n23625;
wire n23626;
wire n23627;
wire n23628;
wire n23629;
wire n23630;
wire n23631;
wire n23632;
wire n23633;
wire n23634;
wire n23635;
wire n23636;
wire n23637;
wire n23638;
wire n23639;
wire n23640;
wire n23641;
wire n23642;
wire n23643;
wire n23644;
wire n23645;
wire n23646;
wire n23647;
wire n23648;
wire n23649;
wire n23650;
wire n23651;
wire n23652;
wire n23653;
wire n23654;
wire n23655;
wire n23656;
wire n23657;
wire n23658;
wire n23659;
wire n23660;
wire n23661;
wire n23662;
wire n23663;
wire n23664;
wire n23665;
wire n23666;
wire n23667;
wire n23668;
wire n23669;
wire n2367;
wire n23670;
wire n23671;
wire n23672;
wire n23673;
wire n23674;
wire n23675;
wire n23676;
wire n23677;
wire n23678;
wire n23679;
wire n23680;
wire n23681;
wire n23682;
wire n23683;
wire n23684;
wire n23685;
wire n23686;
wire n23687;
wire n23688;
wire n23689;
wire n23690;
wire n23691;
wire n23692;
wire n23693;
wire n23694;
wire n23695;
wire n23696;
wire n23697;
wire n23698;
wire n23699;
wire n23700;
wire n23701;
wire n23702;
wire n23703;
wire n23704;
wire n23705;
wire n23706;
wire n23707;
wire n23708;
wire n23709;
wire n23710;
wire n23711;
wire n23712;
wire n23713;
wire n23714;
wire n23715;
wire n23716;
wire n23717;
wire n23718;
wire n23719;
wire n2372;
wire n23720;
wire n23721;
wire n23722;
wire n23723;
wire n23724;
wire n23725;
wire n23726;
wire n23727;
wire n23728;
wire n23729;
wire n23730;
wire n23731;
wire n23732;
wire n23733;
wire n23734;
wire n23735;
wire n23736;
wire n23737;
wire n23738;
wire n23739;
wire n23740;
wire n23741;
wire n23742;
wire n23743;
wire n23744;
wire n23745;
wire n23746;
wire n23747;
wire n23748;
wire n23749;
wire n23750;
wire n23751;
wire n23752;
wire n23753;
wire n23754;
wire n23755;
wire n23756;
wire n23757;
wire n23758;
wire n23759;
wire n23760;
wire n23761;
wire n23762;
wire n23763;
wire n23764;
wire n23765;
wire n23766;
wire n23767;
wire n23768;
wire n23769;
wire n2377;
wire n23770;
wire n23771;
wire n23772;
wire n23773;
wire n23774;
wire n23775;
wire n23776;
wire n23777;
wire n23778;
wire n23779;
wire n23780;
wire n23781;
wire n23782;
wire n23783;
wire n23784;
wire n23785;
wire n23786;
wire n23787;
wire n23788;
wire n23789;
wire n23790;
wire n23791;
wire n23792;
wire n23793;
wire n23794;
wire n23795;
wire n23796;
wire n23797;
wire n23798;
wire n23799;
wire n238;
wire n23800;
wire n23801;
wire n23802;
wire n23803;
wire n23804;
wire n23805;
wire n23806;
wire n23807;
wire n23808;
wire n23809;
wire n23810;
wire n23811;
wire n23812;
wire n23813;
wire n23814;
wire n23815;
wire n23816;
wire n23817;
wire n23818;
wire n23819;
wire n2382;
wire n23820;
wire n23821;
wire n23822;
wire n23823;
wire n23824;
wire n23825;
wire n23826;
wire n23827;
wire n23828;
wire n23829;
wire n23830;
wire n23831;
wire n23832;
wire n23833;
wire n23834;
wire n23835;
wire n23836;
wire n23837;
wire n23838;
wire n23839;
wire n23840;
wire n23841;
wire n23842;
wire n23843;
wire n23844;
wire n23845;
wire n23846;
wire n23847;
wire n23848;
wire n23849;
wire n23850;
wire n23851;
wire n23852;
wire n23853;
wire n23854;
wire n23855;
wire n23856;
wire n23857;
wire n23858;
wire n23859;
wire n23860;
wire n23861;
wire n23862;
wire n23863;
wire n23864;
wire n23865;
wire n23866;
wire n23867;
wire n23868;
wire n23869;
wire n2387;
wire n23870;
wire n23871;
wire n23872;
wire n23873;
wire n23874;
wire n23875;
wire n23876;
wire n23877;
wire n23878;
wire n23879;
wire n23880;
wire n23881;
wire n23882;
wire n23883;
wire n23884;
wire n23885;
wire n23886;
wire n23887;
wire n23888;
wire n23889;
wire n23890;
wire n23891;
wire n23892;
wire n23893;
wire n23894;
wire n23895;
wire n23896;
wire n23897;
wire n23898;
wire n23899;
wire n23900;
wire n23901;
wire n23902;
wire n23903;
wire n23904;
wire n23905;
wire n23906;
wire n23907;
wire n23908;
wire n23909;
wire n23910;
wire n23911;
wire n23912;
wire n23913;
wire n23914;
wire n23915;
wire n23916;
wire n23917;
wire n23918;
wire n23919;
wire n2392;
wire n23920;
wire n23921;
wire n23922;
wire n23923;
wire n23924;
wire n23925;
wire n23926;
wire n23927;
wire n23928;
wire n23929;
wire n23930;
wire n23931;
wire n23932;
wire n23933;
wire n23934;
wire n23935;
wire n23936;
wire n23937;
wire n23938;
wire n23939;
wire n23940;
wire n23941;
wire n23942;
wire n23943;
wire n23944;
wire n23945;
wire n23946;
wire n23947;
wire n23948;
wire n23949;
wire n23950;
wire n23951;
wire n23952;
wire n23953;
wire n23954;
wire n23955;
wire n23956;
wire n23957;
wire n23958;
wire n23959;
wire n23960;
wire n23961;
wire n23962;
wire n23963;
wire n23964;
wire n23965;
wire n23966;
wire n23967;
wire n23968;
wire n23969;
wire n2397;
wire n23970;
wire n23971;
wire n23972;
wire n23973;
wire n23974;
wire n23975;
wire n23976;
wire n23977;
wire n23978;
wire n23979;
wire n23980;
wire n23981;
wire n23982;
wire n23983;
wire n23984;
wire n23985;
wire n23986;
wire n23987;
wire n23988;
wire n23989;
wire n23990;
wire n23991;
wire n23992;
wire n23993;
wire n23994;
wire n23995;
wire n23996;
wire n23997;
wire n23998;
wire n23999;
wire n24000;
wire n24001;
wire n24002;
wire n24003;
wire n24004;
wire n24005;
wire n24006;
wire n24007;
wire n24008;
wire n24009;
wire n24010;
wire n24011;
wire n24012;
wire n24013;
wire n24014;
wire n24015;
wire n24016;
wire n24017;
wire n24018;
wire n24019;
wire n2402;
wire n24020;
wire n24021;
wire n24022;
wire n24023;
wire n24024;
wire n24025;
wire n24026;
wire n24027;
wire n24028;
wire n24029;
wire n24030;
wire n24031;
wire n24032;
wire n24033;
wire n24034;
wire n24035;
wire n24036;
wire n24037;
wire n24038;
wire n24039;
wire n24040;
wire n24041;
wire n24042;
wire n24043;
wire n24044;
wire n24045;
wire n24046;
wire n24047;
wire n24048;
wire n24049;
wire n24050;
wire n24051;
wire n24052;
wire n24053;
wire n24054;
wire n24055;
wire n24056;
wire n24057;
wire n24058;
wire n24059;
wire n24060;
wire n24061;
wire n24062;
wire n24063;
wire n24064;
wire n24065;
wire n24066;
wire n24067;
wire n24068;
wire n24069;
wire n2407;
wire n24070;
wire n24071;
wire n24072;
wire n24073;
wire n24074;
wire n24075;
wire n24076;
wire n24077;
wire n24078;
wire n24079;
wire n24080;
wire n24081;
wire n24082;
wire n24083;
wire n24084;
wire n24085;
wire n24086;
wire n24087;
wire n24088;
wire n24089;
wire n24090;
wire n24091;
wire n24092;
wire n24093;
wire n24094;
wire n24095;
wire n24096;
wire n24097;
wire n24098;
wire n24099;
wire n24100;
wire n24101;
wire n24102;
wire n24103;
wire n24104;
wire n24105;
wire n24106;
wire n24107;
wire n24108;
wire n24109;
wire n24110;
wire n24111;
wire n24112;
wire n24113;
wire n24114;
wire n24115;
wire n24116;
wire n24117;
wire n24118;
wire n24119;
wire n2412;
wire n24120;
wire n24121;
wire n24122;
wire n24123;
wire n24124;
wire n24125;
wire n24126;
wire n24127;
wire n24128;
wire n24129;
wire n24130;
wire n24131;
wire n24132;
wire n24133;
wire n24134;
wire n24135;
wire n24136;
wire n24137;
wire n24138;
wire n24139;
wire n24140;
wire n24141;
wire n24142;
wire n24143;
wire n24144;
wire n24145;
wire n24146;
wire n24147;
wire n24148;
wire n24149;
wire n24150;
wire n24151;
wire n24152;
wire n24153;
wire n24154;
wire n24155;
wire n24156;
wire n24157;
wire n24158;
wire n24159;
wire n24160;
wire n24161;
wire n24162;
wire n24163;
wire n24164;
wire n24165;
wire n24166;
wire n24167;
wire n24168;
wire n24169;
wire n2417;
wire n24170;
wire n24171;
wire n24172;
wire n24173;
wire n24174;
wire n24175;
wire n24176;
wire n24177;
wire n24178;
wire n24179;
wire n24180;
wire n24181;
wire n24182;
wire n24183;
wire n24184;
wire n24185;
wire n24186;
wire n24187;
wire n24188;
wire n24189;
wire n24190;
wire n24191;
wire n24192;
wire n24193;
wire n24194;
wire n24195;
wire n24196;
wire n24197;
wire n24198;
wire n24199;
wire n24200;
wire n24201;
wire n24202;
wire n24203;
wire n24204;
wire n24205;
wire n24206;
wire n24207;
wire n24208;
wire n24209;
wire n24210;
wire n24211;
wire n24212;
wire n24213;
wire n24214;
wire n24215;
wire n24216;
wire n24217;
wire n24218;
wire n24219;
wire n2422;
wire n24220;
wire n24221;
wire n24222;
wire n24223;
wire n24224;
wire n24225;
wire n24226;
wire n24227;
wire n24228;
wire n24229;
wire n24230;
wire n24231;
wire n24232;
wire n24233;
wire n24234;
wire n24235;
wire n24236;
wire n24237;
wire n24238;
wire n24239;
wire n24240;
wire n24241;
wire n24242;
wire n24243;
wire n24244;
wire n24245;
wire n24246;
wire n24247;
wire n24248;
wire n24249;
wire n24250;
wire n24251;
wire n24252;
wire n24253;
wire n24254;
wire n24255;
wire n24256;
wire n24257;
wire n24258;
wire n24259;
wire n24260;
wire n24261;
wire n24262;
wire n24263;
wire n24264;
wire n24265;
wire n24266;
wire n24267;
wire n24268;
wire n24269;
wire n2427;
wire n24270;
wire n24271;
wire n24272;
wire n24273;
wire n24274;
wire n24275;
wire n24276;
wire n24277;
wire n24278;
wire n24279;
wire n24280;
wire n24281;
wire n24282;
wire n24283;
wire n24284;
wire n24285;
wire n24286;
wire n24287;
wire n24288;
wire n24289;
wire n24290;
wire n24291;
wire n24292;
wire n24293;
wire n24294;
wire n24295;
wire n24296;
wire n24297;
wire n24298;
wire n24299;
wire n243;
wire n24300;
wire n24301;
wire n24302;
wire n24303;
wire n24304;
wire n24305;
wire n24306;
wire n24307;
wire n24308;
wire n24309;
wire n24310;
wire n24311;
wire n24312;
wire n24313;
wire n24314;
wire n24315;
wire n24316;
wire n24317;
wire n24318;
wire n24319;
wire n2432;
wire n24320;
wire n24321;
wire n24322;
wire n24323;
wire n24324;
wire n24325;
wire n24326;
wire n24327;
wire n24328;
wire n24329;
wire n24330;
wire n24331;
wire n24332;
wire n24333;
wire n24334;
wire n24335;
wire n24336;
wire n24337;
wire n24338;
wire n24339;
wire n24340;
wire n24341;
wire n24342;
wire n24343;
wire n24344;
wire n24345;
wire n24346;
wire n24347;
wire n24348;
wire n24349;
wire n24350;
wire n24351;
wire n24352;
wire n24353;
wire n24354;
wire n24355;
wire n24356;
wire n24357;
wire n24358;
wire n24359;
wire n24360;
wire n24361;
wire n24362;
wire n24363;
wire n24364;
wire n24365;
wire n24366;
wire n24367;
wire n24368;
wire n24369;
wire n2437;
wire n24370;
wire n24371;
wire n24372;
wire n24373;
wire n24374;
wire n24375;
wire n24376;
wire n24377;
wire n24378;
wire n24379;
wire n24380;
wire n24381;
wire n24382;
wire n24383;
wire n24384;
wire n24385;
wire n24386;
wire n24387;
wire n24388;
wire n24389;
wire n24390;
wire n24391;
wire n24392;
wire n24393;
wire n24394;
wire n24395;
wire n24396;
wire n24397;
wire n24398;
wire n24399;
wire n24400;
wire n24401;
wire n24402;
wire n24403;
wire n24404;
wire n24405;
wire n24406;
wire n24407;
wire n24408;
wire n24409;
wire n24410;
wire n24411;
wire n24412;
wire n24413;
wire n24414;
wire n24415;
wire n24416;
wire n24417;
wire n24418;
wire n24419;
wire n2442;
wire n24420;
wire n24421;
wire n24422;
wire n24423;
wire n24424;
wire n24425;
wire n24426;
wire n24427;
wire n24428;
wire n24429;
wire n24430;
wire n24431;
wire n24432;
wire n24433;
wire n24434;
wire n24435;
wire n24436;
wire n24437;
wire n24438;
wire n24439;
wire n24440;
wire n24441;
wire n24442;
wire n24443;
wire n24444;
wire n24445;
wire n24446;
wire n24447;
wire n24448;
wire n24449;
wire n24450;
wire n24451;
wire n24452;
wire n24453;
wire n24454;
wire n24455;
wire n24456;
wire n24457;
wire n24458;
wire n24459;
wire n24460;
wire n24461;
wire n24462;
wire n24463;
wire n24464;
wire n24465;
wire n24466;
wire n24467;
wire n24468;
wire n24469;
wire n2447;
wire n24470;
wire n24471;
wire n24472;
wire n24473;
wire n24474;
wire n24475;
wire n24476;
wire n24477;
wire n24478;
wire n24479;
wire n24480;
wire n24481;
wire n24482;
wire n24483;
wire n24484;
wire n24485;
wire n24486;
wire n24487;
wire n24488;
wire n24489;
wire n24490;
wire n24491;
wire n24492;
wire n24493;
wire n24494;
wire n24495;
wire n24496;
wire n24497;
wire n24498;
wire n24499;
wire n24500;
wire n24501;
wire n24502;
wire n24503;
wire n24504;
wire n24505;
wire n24506;
wire n24507;
wire n24508;
wire n24509;
wire n2451;
wire n24510;
wire n24511;
wire n24512;
wire n24513;
wire n24514;
wire n24515;
wire n24516;
wire n24517;
wire n24518;
wire n24519;
wire n24520;
wire n24521;
wire n24522;
wire n24523;
wire n24524;
wire n24525;
wire n24526;
wire n24527;
wire n24528;
wire n24529;
wire n24530;
wire n24531;
wire n24532;
wire n24533;
wire n24534;
wire n24535;
wire n24536;
wire n24537;
wire n24538;
wire n24539;
wire n24540;
wire n24541;
wire n24542;
wire n24543;
wire n24544;
wire n24545;
wire n24546;
wire n24547;
wire n24548;
wire n24549;
wire n24550;
wire n24551;
wire n24552;
wire n24553;
wire n24554;
wire n24555;
wire n24556;
wire n24557;
wire n24558;
wire n24559;
wire n2456;
wire n24560;
wire n24561;
wire n24562;
wire n24563;
wire n24564;
wire n24565;
wire n24566;
wire n24567;
wire n24568;
wire n24569;
wire n24570;
wire n24571;
wire n24572;
wire n24573;
wire n24574;
wire n24575;
wire n24576;
wire n24577;
wire n24578;
wire n24579;
wire n24580;
wire n24581;
wire n24582;
wire n24583;
wire n24584;
wire n24585;
wire n24586;
wire n24587;
wire n24588;
wire n24589;
wire n24590;
wire n24591;
wire n24592;
wire n24593;
wire n24594;
wire n24595;
wire n24596;
wire n24597;
wire n24598;
wire n24599;
wire n24600;
wire n24601;
wire n24602;
wire n24603;
wire n24604;
wire n24605;
wire n24606;
wire n24607;
wire n24608;
wire n24609;
wire n2461;
wire n24610;
wire n24611;
wire n24612;
wire n24613;
wire n24614;
wire n24615;
wire n24616;
wire n24617;
wire n24618;
wire n24619;
wire n24620;
wire n24621;
wire n24622;
wire n24623;
wire n24624;
wire n24625;
wire n24626;
wire n24627;
wire n24628;
wire n24629;
wire n24630;
wire n24631;
wire n24632;
wire n24633;
wire n24634;
wire n24635;
wire n24636;
wire n24637;
wire n24638;
wire n24639;
wire n24640;
wire n24641;
wire n24642;
wire n24643;
wire n24644;
wire n24645;
wire n24646;
wire n24647;
wire n24648;
wire n24649;
wire n24650;
wire n24651;
wire n24652;
wire n24653;
wire n24654;
wire n24655;
wire n24656;
wire n24657;
wire n24659;
wire n2466;
wire n24660;
wire n24661;
wire n24662;
wire n24663;
wire n24664;
wire n24665;
wire n24666;
wire n24667;
wire n24668;
wire n24669;
wire n24670;
wire n24671;
wire n24672;
wire n24673;
wire n24674;
wire n24675;
wire n24676;
wire n24677;
wire n24678;
wire n24679;
wire n24680;
wire n24681;
wire n24682;
wire n24683;
wire n24684;
wire n24685;
wire n24686;
wire n24687;
wire n24688;
wire n24689;
wire n24690;
wire n24691;
wire n24692;
wire n24693;
wire n24694;
wire n24695;
wire n24696;
wire n24697;
wire n24698;
wire n24699;
wire n24700;
wire n24701;
wire n24702;
wire n24703;
wire n24704;
wire n24705;
wire n24706;
wire n24707;
wire n24708;
wire n24709;
wire n2471;
wire n24710;
wire n24711;
wire n24712;
wire n24713;
wire n24714;
wire n24715;
wire n24716;
wire n24717;
wire n24718;
wire n24719;
wire n24720;
wire n24721;
wire n24722;
wire n24723;
wire n24724;
wire n24725;
wire n24726;
wire n24727;
wire n24728;
wire n24729;
wire n24730;
wire n24731;
wire n24732;
wire n24733;
wire n24734;
wire n24735;
wire n24736;
wire n24737;
wire n24738;
wire n24739;
wire n24740;
wire n24741;
wire n24742;
wire n24743;
wire n24744;
wire n24745;
wire n24746;
wire n24747;
wire n24748;
wire n24749;
wire n24750;
wire n24751;
wire n24752;
wire n24753;
wire n24754;
wire n24755;
wire n24756;
wire n24757;
wire n24758;
wire n24759;
wire n2476;
wire n24760;
wire n24761;
wire n24762;
wire n24763;
wire n24764;
wire n24765;
wire n24766;
wire n24767;
wire n24768;
wire n24769;
wire n24770;
wire n24771;
wire n24772;
wire n24773;
wire n24774;
wire n24775;
wire n24776;
wire n24777;
wire n24778;
wire n24779;
wire n24780;
wire n24781;
wire n24782;
wire n24783;
wire n24784;
wire n24785;
wire n24786;
wire n24787;
wire n24788;
wire n24789;
wire n24790;
wire n24791;
wire n24792;
wire n24793;
wire n24794;
wire n24795;
wire n24796;
wire n24797;
wire n24798;
wire n24799;
wire n248;
wire n24800;
wire n24801;
wire n24802;
wire n24803;
wire n24804;
wire n24805;
wire n24806;
wire n24807;
wire n24808;
wire n24809;
wire n2481;
wire n24810;
wire n24811;
wire n24812;
wire n24813;
wire n24814;
wire n24815;
wire n24816;
wire n24817;
wire n24818;
wire n24819;
wire n24820;
wire n24821;
wire n24822;
wire n24823;
wire n24824;
wire n24825;
wire n24826;
wire n24827;
wire n24828;
wire n24829;
wire n24830;
wire n24831;
wire n24832;
wire n24833;
wire n24834;
wire n24835;
wire n24836;
wire n24837;
wire n24838;
wire n24839;
wire n24840;
wire n24841;
wire n24842;
wire n24843;
wire n24844;
wire n24845;
wire n24846;
wire n24847;
wire n24848;
wire n24849;
wire n24850;
wire n24851;
wire n24852;
wire n24853;
wire n24854;
wire n24855;
wire n24856;
wire n24857;
wire n24858;
wire n24859;
wire n2486;
wire n24860;
wire n24861;
wire n24862;
wire n24863;
wire n24864;
wire n24865;
wire n24866;
wire n24867;
wire n24868;
wire n24869;
wire n24870;
wire n24871;
wire n24872;
wire n24873;
wire n24874;
wire n24875;
wire n24876;
wire n24877;
wire n24878;
wire n24879;
wire n24880;
wire n24881;
wire n24882;
wire n24883;
wire n24884;
wire n24885;
wire n24886;
wire n24887;
wire n24888;
wire n24889;
wire n24890;
wire n24891;
wire n24892;
wire n24893;
wire n24894;
wire n24895;
wire n24896;
wire n24897;
wire n24898;
wire n24899;
wire n24900;
wire n24901;
wire n24902;
wire n24903;
wire n24904;
wire n24905;
wire n24906;
wire n24907;
wire n24908;
wire n24909;
wire n2491;
wire n24910;
wire n24911;
wire n24912;
wire n24913;
wire n24914;
wire n24915;
wire n24916;
wire n24917;
wire n24918;
wire n24919;
wire n24920;
wire n24921;
wire n24922;
wire n24923;
wire n24924;
wire n24925;
wire n24926;
wire n24927;
wire n24928;
wire n24929;
wire n24930;
wire n24931;
wire n24932;
wire n24933;
wire n24934;
wire n24935;
wire n24936;
wire n24937;
wire n24938;
wire n24939;
wire n24940;
wire n24941;
wire n24942;
wire n24943;
wire n24944;
wire n24945;
wire n24946;
wire n24947;
wire n24948;
wire n24949;
wire n24950;
wire n24951;
wire n24952;
wire n24953;
wire n24954;
wire n24955;
wire n24956;
wire n24957;
wire n24958;
wire n24959;
wire n2496;
wire n24960;
wire n24961;
wire n24962;
wire n24963;
wire n24964;
wire n24965;
wire n24966;
wire n24967;
wire n24968;
wire n24969;
wire n24970;
wire n24971;
wire n24972;
wire n24973;
wire n24974;
wire n24975;
wire n24976;
wire n24977;
wire n24978;
wire n24979;
wire n24980;
wire n24981;
wire n24982;
wire n24983;
wire n24984;
wire n24985;
wire n24986;
wire n24987;
wire n24988;
wire n24989;
wire n24990;
wire n24991;
wire n24992;
wire n24993;
wire n24994;
wire n24995;
wire n24996;
wire n24997;
wire n24998;
wire n24999;
wire n25000;
wire n25001;
wire n25002;
wire n25003;
wire n25004;
wire n25005;
wire n25006;
wire n25007;
wire n25008;
wire n25009;
wire n2501;
wire n25010;
wire n25011;
wire n25012;
wire n25013;
wire n25014;
wire n25015;
wire n25016;
wire n25017;
wire n25018;
wire n25019;
wire n25020;
wire n25021;
wire n25022;
wire n25023;
wire n25024;
wire n25025;
wire n25026;
wire n25027;
wire n25028;
wire n25029;
wire n25030;
wire n25031;
wire n25032;
wire n25033;
wire n25034;
wire n25035;
wire n25036;
wire n25037;
wire n25038;
wire n25039;
wire n25040;
wire n25041;
wire n25042;
wire n25043;
wire n25044;
wire n25045;
wire n25046;
wire n25047;
wire n25048;
wire n25049;
wire n25050;
wire n25051;
wire n25052;
wire n25053;
wire n25054;
wire n25055;
wire n25056;
wire n25057;
wire n25058;
wire n25059;
wire n2506;
wire n25060;
wire n25061;
wire n25062;
wire n25063;
wire n25064;
wire n25065;
wire n25066;
wire n25067;
wire n25068;
wire n25069;
wire n25070;
wire n25071;
wire n25072;
wire n25073;
wire n25074;
wire n25075;
wire n25076;
wire n25077;
wire n25078;
wire n25079;
wire n25080;
wire n25081;
wire n25082;
wire n25083;
wire n25084;
wire n25085;
wire n25086;
wire n25087;
wire n25088;
wire n25089;
wire n25090;
wire n25091;
wire n25092;
wire n25093;
wire n25094;
wire n25095;
wire n25096;
wire n25097;
wire n25098;
wire n25099;
wire n25100;
wire n25101;
wire n25102;
wire n25103;
wire n25104;
wire n25105;
wire n25106;
wire n25107;
wire n25108;
wire n25109;
wire n2511;
wire n25110;
wire n25111;
wire n25112;
wire n25113;
wire n25114;
wire n25115;
wire n25116;
wire n25117;
wire n25118;
wire n25119;
wire n25120;
wire n25121;
wire n25122;
wire n25123;
wire n25124;
wire n25125;
wire n25126;
wire n25127;
wire n25128;
wire n25129;
wire n25130;
wire n25131;
wire n25132;
wire n25133;
wire n25134;
wire n25135;
wire n25136;
wire n25137;
wire n25138;
wire n25139;
wire n25140;
wire n25141;
wire n25142;
wire n25143;
wire n25144;
wire n25145;
wire n25146;
wire n25147;
wire n25148;
wire n25149;
wire n25150;
wire n25151;
wire n25152;
wire n25153;
wire n25154;
wire n25155;
wire n25156;
wire n25157;
wire n25158;
wire n25159;
wire n2516;
wire n25160;
wire n25161;
wire n25162;
wire n25163;
wire n25164;
wire n25165;
wire n25166;
wire n25167;
wire n25168;
wire n25169;
wire n25170;
wire n25171;
wire n25172;
wire n25173;
wire n25174;
wire n25175;
wire n25176;
wire n25177;
wire n25178;
wire n25179;
wire n25180;
wire n25181;
wire n25182;
wire n25183;
wire n25184;
wire n25185;
wire n25186;
wire n25187;
wire n25188;
wire n25189;
wire n25190;
wire n25191;
wire n25192;
wire n25193;
wire n25194;
wire n25195;
wire n25196;
wire n25197;
wire n25198;
wire n25199;
wire n25200;
wire n25201;
wire n25202;
wire n25203;
wire n25204;
wire n25205;
wire n25206;
wire n25207;
wire n25208;
wire n25209;
wire n2521;
wire n25210;
wire n25211;
wire n25212;
wire n25213;
wire n25214;
wire n25215;
wire n25216;
wire n25217;
wire n25218;
wire n25219;
wire n25220;
wire n25221;
wire n25222;
wire n25223;
wire n25224;
wire n25225;
wire n25226;
wire n25227;
wire n25228;
wire n25229;
wire n25230;
wire n25231;
wire n25232;
wire n25233;
wire n25234;
wire n25235;
wire n25236;
wire n25237;
wire n25238;
wire n25239;
wire n25240;
wire n25241;
wire n25242;
wire n25243;
wire n25244;
wire n25245;
wire n25246;
wire n25247;
wire n25248;
wire n25249;
wire n2525;
wire n25250;
wire n25251;
wire n25252;
wire n25253;
wire n25254;
wire n25255;
wire n25256;
wire n25257;
wire n25258;
wire n25259;
wire n25260;
wire n25261;
wire n25262;
wire n25263;
wire n25264;
wire n25265;
wire n25266;
wire n25267;
wire n25268;
wire n25269;
wire n25270;
wire n25271;
wire n25272;
wire n25273;
wire n25274;
wire n25275;
wire n25276;
wire n25277;
wire n25278;
wire n25279;
wire n25280;
wire n25281;
wire n25282;
wire n25283;
wire n25284;
wire n25285;
wire n25286;
wire n25287;
wire n25288;
wire n25289;
wire n25290;
wire n25291;
wire n25292;
wire n25293;
wire n25294;
wire n25295;
wire n25296;
wire n25297;
wire n25298;
wire n25299;
wire n253;
wire n2530;
wire n25300;
wire n25301;
wire n25302;
wire n25303;
wire n25304;
wire n25305;
wire n25306;
wire n25307;
wire n25308;
wire n25309;
wire n25310;
wire n25311;
wire n25312;
wire n25313;
wire n25314;
wire n25315;
wire n25316;
wire n25317;
wire n25318;
wire n25319;
wire n25320;
wire n25321;
wire n25322;
wire n25323;
wire n25324;
wire n25325;
wire n25326;
wire n25327;
wire n25328;
wire n25329;
wire n25330;
wire n25331;
wire n25332;
wire n25333;
wire n25334;
wire n25335;
wire n25336;
wire n25337;
wire n25338;
wire n25339;
wire n25340;
wire n25341;
wire n25342;
wire n25343;
wire n25344;
wire n25345;
wire n25346;
wire n25347;
wire n25348;
wire n25349;
wire n2535;
wire n25350;
wire n25351;
wire n25352;
wire n25353;
wire n25354;
wire n25355;
wire n25356;
wire n25357;
wire n25358;
wire n25359;
wire n25360;
wire n25361;
wire n25362;
wire n25363;
wire n25364;
wire n25365;
wire n25366;
wire n25367;
wire n25368;
wire n25369;
wire n25370;
wire n25371;
wire n25372;
wire n25373;
wire n25374;
wire n25375;
wire n25376;
wire n25377;
wire n25378;
wire n25379;
wire n25380;
wire n25381;
wire n25382;
wire n25383;
wire n25384;
wire n25385;
wire n25386;
wire n25387;
wire n25388;
wire n25389;
wire n25390;
wire n25391;
wire n25392;
wire n25393;
wire n25394;
wire n25395;
wire n25396;
wire n25397;
wire n25398;
wire n25399;
wire n2540;
wire n25400;
wire n25401;
wire n25402;
wire n25403;
wire n25404;
wire n25405;
wire n25406;
wire n25407;
wire n25408;
wire n25409;
wire n25410;
wire n25411;
wire n25412;
wire n25413;
wire n25414;
wire n25415;
wire n25416;
wire n25417;
wire n25418;
wire n25419;
wire n25420;
wire n25421;
wire n25422;
wire n25423;
wire n25424;
wire n25425;
wire n25426;
wire n25427;
wire n25428;
wire n25429;
wire n25430;
wire n25431;
wire n25432;
wire n25433;
wire n25434;
wire n25435;
wire n25436;
wire n25437;
wire n25438;
wire n25439;
wire n25440;
wire n25441;
wire n25442;
wire n25443;
wire n25444;
wire n25445;
wire n25446;
wire n25447;
wire n25448;
wire n25449;
wire n2545;
wire n25450;
wire n25451;
wire n25452;
wire n25453;
wire n25454;
wire n25455;
wire n25456;
wire n25457;
wire n25458;
wire n25459;
wire n25460;
wire n25461;
wire n25462;
wire n25463;
wire n25464;
wire n25465;
wire n25466;
wire n25467;
wire n25468;
wire n25469;
wire n25470;
wire n25471;
wire n25472;
wire n25473;
wire n25474;
wire n25475;
wire n25476;
wire n25477;
wire n25478;
wire n25479;
wire n25480;
wire n25481;
wire n25482;
wire n25483;
wire n25484;
wire n25485;
wire n25486;
wire n25487;
wire n25488;
wire n25489;
wire n25490;
wire n25491;
wire n25492;
wire n25493;
wire n25494;
wire n25495;
wire n25496;
wire n25497;
wire n25498;
wire n25499;
wire n2550;
wire n25500;
wire n25501;
wire n25502;
wire n25503;
wire n25504;
wire n25505;
wire n25506;
wire n25507;
wire n25508;
wire n25509;
wire n25510;
wire n25511;
wire n25512;
wire n25513;
wire n25514;
wire n25515;
wire n25516;
wire n25517;
wire n25518;
wire n25519;
wire n25520;
wire n25521;
wire n25522;
wire n25523;
wire n25524;
wire n25525;
wire n25526;
wire n25527;
wire n25528;
wire n25529;
wire n25530;
wire n25531;
wire n25532;
wire n25533;
wire n25534;
wire n25535;
wire n25536;
wire n25537;
wire n25538;
wire n25539;
wire n25540;
wire n25541;
wire n25542;
wire n25543;
wire n25544;
wire n25545;
wire n25546;
wire n25547;
wire n25548;
wire n25549;
wire n2555;
wire n25550;
wire n25551;
wire n25552;
wire n25553;
wire n25554;
wire n25555;
wire n25556;
wire n25557;
wire n25558;
wire n25559;
wire n25560;
wire n25561;
wire n25562;
wire n25563;
wire n25564;
wire n25565;
wire n25566;
wire n25567;
wire n25568;
wire n25569;
wire n25570;
wire n25571;
wire n25572;
wire n25573;
wire n25574;
wire n25575;
wire n25576;
wire n25577;
wire n25578;
wire n25579;
wire n25580;
wire n25582;
wire n25583;
wire n25584;
wire n25585;
wire n25586;
wire n25587;
wire n25588;
wire n25589;
wire n25590;
wire n25591;
wire n25592;
wire n25593;
wire n25594;
wire n25595;
wire n25596;
wire n25597;
wire n25598;
wire n25599;
wire n2560;
wire n25600;
wire n25601;
wire n25602;
wire n25603;
wire n25604;
wire n25605;
wire n25606;
wire n25607;
wire n25608;
wire n25609;
wire n25610;
wire n25611;
wire n25612;
wire n25613;
wire n25614;
wire n25615;
wire n25616;
wire n25617;
wire n25618;
wire n25619;
wire n25620;
wire n25621;
wire n25622;
wire n25623;
wire n25624;
wire n25626;
wire n25627;
wire n25629;
wire n25630;
wire n25631;
wire n25632;
wire n25633;
wire n25634;
wire n25635;
wire n25636;
wire n25637;
wire n25639;
wire n25640;
wire n25641;
wire n25642;
wire n25643;
wire n25644;
wire n25645;
wire n25646;
wire n25647;
wire n25649;
wire n2565;
wire n25651;
wire n25652;
wire n25653;
wire n25654;
wire n25655;
wire n25656;
wire n25657;
wire n25658;
wire n25659;
wire n25660;
wire n25661;
wire n25662;
wire n25663;
wire n25664;
wire n25665;
wire n25666;
wire n25667;
wire n25668;
wire n25670;
wire n25671;
wire n25672;
wire n25673;
wire n25674;
wire n25675;
wire n25676;
wire n25677;
wire n25678;
wire n25679;
wire n25680;
wire n25681;
wire n25682;
wire n25683;
wire n25684;
wire n25685;
wire n25686;
wire n25687;
wire n25688;
wire n25689;
wire n25690;
wire n25691;
wire n25692;
wire n25693;
wire n25694;
wire n25695;
wire n25696;
wire n25697;
wire n25698;
wire n25699;
wire n2570;
wire n25700;
wire n25701;
wire n25702;
wire n25703;
wire n25704;
wire n25705;
wire n25706;
wire n25707;
wire n25708;
wire n25709;
wire n25710;
wire n25711;
wire n25712;
wire n25713;
wire n25714;
wire n25715;
wire n25716;
wire n25717;
wire n25718;
wire n25719;
wire n25720;
wire n25721;
wire n25722;
wire n25723;
wire n25724;
wire n25725;
wire n25726;
wire n25727;
wire n25728;
wire n25729;
wire n25730;
wire n25731;
wire n25732;
wire n25733;
wire n25734;
wire n25735;
wire n25736;
wire n25737;
wire n25738;
wire n25739;
wire n25740;
wire n25741;
wire n25742;
wire n25743;
wire n25744;
wire n25745;
wire n25746;
wire n25747;
wire n25748;
wire n25749;
wire n2575;
wire n25750;
wire n25751;
wire n25752;
wire n25753;
wire n25754;
wire n25755;
wire n25756;
wire n25757;
wire n25758;
wire n25759;
wire n25760;
wire n25761;
wire n25762;
wire n25763;
wire n25764;
wire n25765;
wire n25766;
wire n25767;
wire n25768;
wire n25769;
wire n25770;
wire n25771;
wire n25772;
wire n25773;
wire n25774;
wire n25775;
wire n25776;
wire n25777;
wire n25778;
wire n25779;
wire n25780;
wire n25781;
wire n25782;
wire n25783;
wire n25784;
wire n25785;
wire n25786;
wire n25787;
wire n25788;
wire n25789;
wire n2579;
wire n25790;
wire n25791;
wire n25792;
wire n25793;
wire n25794;
wire n25795;
wire n25796;
wire n25797;
wire n25798;
wire n25799;
wire n258;
wire n25800;
wire n25801;
wire n25802;
wire n25803;
wire n25804;
wire n25805;
wire n25806;
wire n25807;
wire n25808;
wire n25809;
wire n25810;
wire n25811;
wire n25812;
wire n25813;
wire n25814;
wire n25815;
wire n25816;
wire n25817;
wire n25818;
wire n25819;
wire n25820;
wire n25821;
wire n25822;
wire n25823;
wire n25824;
wire n25825;
wire n25826;
wire n25827;
wire n25828;
wire n25829;
wire n25830;
wire n25831;
wire n25832;
wire n25833;
wire n25834;
wire n25835;
wire n25836;
wire n25837;
wire n25838;
wire n25839;
wire n2584;
wire n25840;
wire n25841;
wire n25842;
wire n25843;
wire n25844;
wire n25845;
wire n25846;
wire n25847;
wire n25848;
wire n25849;
wire n25850;
wire n25851;
wire n25852;
wire n25853;
wire n25854;
wire n25855;
wire n25856;
wire n25857;
wire n25858;
wire n25859;
wire n25860;
wire n25861;
wire n25862;
wire n25863;
wire n25864;
wire n25865;
wire n25866;
wire n25867;
wire n25868;
wire n25869;
wire n25870;
wire n25871;
wire n25872;
wire n25873;
wire n25874;
wire n25875;
wire n25876;
wire n25877;
wire n25878;
wire n25879;
wire n25880;
wire n25881;
wire n25882;
wire n25883;
wire n25884;
wire n25885;
wire n25886;
wire n25887;
wire n25888;
wire n25889;
wire n2589;
wire n25890;
wire n25891;
wire n25892;
wire n25893;
wire n25894;
wire n25895;
wire n25896;
wire n25897;
wire n25898;
wire n25899;
wire n25900;
wire n25901;
wire n25902;
wire n25903;
wire n25904;
wire n25905;
wire n25906;
wire n25907;
wire n25908;
wire n25909;
wire n25910;
wire n25911;
wire n25912;
wire n25913;
wire n25914;
wire n25915;
wire n25916;
wire n25917;
wire n25918;
wire n25919;
wire n25920;
wire n25921;
wire n25922;
wire n25923;
wire n25924;
wire n25925;
wire n25926;
wire n25927;
wire n25929;
wire n25931;
wire n25932;
wire n25933;
wire n25934;
wire n25935;
wire n25937;
wire n25938;
wire n2594;
wire n25940;
wire n25941;
wire n25942;
wire n25943;
wire n25944;
wire n25945;
wire n25946;
wire n25947;
wire n25948;
wire n25949;
wire n25950;
wire n25951;
wire n25952;
wire n25953;
wire n25954;
wire n25955;
wire n25956;
wire n25957;
wire n25958;
wire n25959;
wire n25960;
wire n25961;
wire n25962;
wire n25963;
wire n25964;
wire n25965;
wire n25966;
wire n25967;
wire n25968;
wire n25969;
wire n25970;
wire n25971;
wire n25972;
wire n25973;
wire n25974;
wire n25975;
wire n25976;
wire n25977;
wire n25978;
wire n25979;
wire n25980;
wire n25981;
wire n25982;
wire n25983;
wire n25984;
wire n25985;
wire n25986;
wire n25987;
wire n25988;
wire n25989;
wire n2599;
wire n25990;
wire n25991;
wire n25992;
wire n25993;
wire n25994;
wire n25995;
wire n25996;
wire n25997;
wire n25998;
wire n25999;
wire n26000;
wire n26001;
wire n26002;
wire n26003;
wire n26004;
wire n26005;
wire n26006;
wire n26007;
wire n26008;
wire n26009;
wire n26010;
wire n26011;
wire n26012;
wire n26013;
wire n26014;
wire n26015;
wire n26016;
wire n26017;
wire n26018;
wire n26019;
wire n26020;
wire n26021;
wire n26022;
wire n26023;
wire n26024;
wire n26025;
wire n26026;
wire n26027;
wire n26028;
wire n26029;
wire n26030;
wire n26031;
wire n26032;
wire n26033;
wire n26034;
wire n26035;
wire n26036;
wire n26037;
wire n26038;
wire n26039;
wire n2604;
wire n26040;
wire n26041;
wire n26042;
wire n26043;
wire n26044;
wire n26045;
wire n26046;
wire n26047;
wire n26048;
wire n26049;
wire n26050;
wire n26051;
wire n26052;
wire n26053;
wire n26054;
wire n26055;
wire n26056;
wire n26057;
wire n26058;
wire n26059;
wire n26060;
wire n26061;
wire n26062;
wire n26063;
wire n26064;
wire n26065;
wire n26066;
wire n26067;
wire n26068;
wire n26069;
wire n26070;
wire n26071;
wire n26072;
wire n26073;
wire n26074;
wire n26075;
wire n26076;
wire n26077;
wire n26078;
wire n26079;
wire n26080;
wire n26081;
wire n26082;
wire n26083;
wire n26084;
wire n26085;
wire n26086;
wire n26087;
wire n26088;
wire n26089;
wire n2609;
wire n26090;
wire n26091;
wire n26092;
wire n26093;
wire n26094;
wire n26095;
wire n26096;
wire n26097;
wire n26098;
wire n26099;
wire n26100;
wire n26101;
wire n26102;
wire n26103;
wire n26104;
wire n26105;
wire n26106;
wire n26107;
wire n26108;
wire n26109;
wire n26110;
wire n26111;
wire n26112;
wire n26113;
wire n26114;
wire n26115;
wire n26116;
wire n26117;
wire n26118;
wire n26119;
wire n26120;
wire n26121;
wire n26122;
wire n26123;
wire n26124;
wire n26125;
wire n26126;
wire n26127;
wire n26128;
wire n26129;
wire n26130;
wire n26131;
wire n26132;
wire n26133;
wire n26134;
wire n26135;
wire n26136;
wire n26137;
wire n26138;
wire n26139;
wire n2614;
wire n26140;
wire n26141;
wire n26142;
wire n26143;
wire n26144;
wire n26145;
wire n26146;
wire n26147;
wire n26148;
wire n26149;
wire n26150;
wire n26151;
wire n26152;
wire n26153;
wire n26154;
wire n26155;
wire n26156;
wire n26157;
wire n26158;
wire n26159;
wire n26160;
wire n26161;
wire n26162;
wire n26163;
wire n26164;
wire n26165;
wire n26166;
wire n26167;
wire n26168;
wire n26169;
wire n26170;
wire n26171;
wire n26172;
wire n26173;
wire n26174;
wire n26175;
wire n26176;
wire n26177;
wire n26178;
wire n26179;
wire n2618;
wire n26180;
wire n26181;
wire n26182;
wire n26183;
wire n26184;
wire n26185;
wire n26186;
wire n26187;
wire n26188;
wire n26189;
wire n26190;
wire n26191;
wire n26192;
wire n26193;
wire n26194;
wire n26195;
wire n26196;
wire n26197;
wire n26198;
wire n26199;
wire n26200;
wire n26201;
wire n26202;
wire n26203;
wire n26204;
wire n26205;
wire n26206;
wire n26207;
wire n26208;
wire n26209;
wire n26210;
wire n26211;
wire n26212;
wire n26213;
wire n26214;
wire n26215;
wire n26216;
wire n26217;
wire n26218;
wire n26219;
wire n26220;
wire n26221;
wire n26222;
wire n26223;
wire n26224;
wire n26225;
wire n26226;
wire n26227;
wire n26228;
wire n26229;
wire n2623;
wire n26230;
wire n26231;
wire n26232;
wire n26233;
wire n26234;
wire n26235;
wire n26236;
wire n26237;
wire n26238;
wire n26239;
wire n26240;
wire n26241;
wire n26242;
wire n26243;
wire n26244;
wire n26245;
wire n26246;
wire n26247;
wire n26248;
wire n26249;
wire n26250;
wire n26251;
wire n26252;
wire n26253;
wire n26254;
wire n26255;
wire n26256;
wire n26257;
wire n26258;
wire n26259;
wire n26260;
wire n26261;
wire n26262;
wire n26263;
wire n26264;
wire n26265;
wire n26266;
wire n26267;
wire n26268;
wire n26269;
wire n26270;
wire n26271;
wire n26272;
wire n26273;
wire n26274;
wire n26275;
wire n26276;
wire n26277;
wire n26278;
wire n26279;
wire n2628;
wire n26280;
wire n26281;
wire n26282;
wire n26283;
wire n26284;
wire n26285;
wire n26286;
wire n26287;
wire n26288;
wire n26289;
wire n26290;
wire n26291;
wire n26292;
wire n26293;
wire n26294;
wire n26295;
wire n26296;
wire n26297;
wire n26298;
wire n26299;
wire n263;
wire n26300;
wire n26301;
wire n26302;
wire n26303;
wire n26304;
wire n26305;
wire n26306;
wire n26307;
wire n26308;
wire n26309;
wire n26310;
wire n26311;
wire n26312;
wire n26313;
wire n26314;
wire n26315;
wire n26316;
wire n26317;
wire n26318;
wire n26319;
wire n26320;
wire n26321;
wire n26322;
wire n26323;
wire n26324;
wire n26325;
wire n26326;
wire n26327;
wire n26328;
wire n26329;
wire n2633;
wire n26330;
wire n26331;
wire n26332;
wire n26333;
wire n26334;
wire n26335;
wire n26336;
wire n26337;
wire n26338;
wire n26339;
wire n26340;
wire n26341;
wire n26342;
wire n26343;
wire n26344;
wire n26345;
wire n26346;
wire n26347;
wire n26348;
wire n26349;
wire n26350;
wire n26351;
wire n26352;
wire n26353;
wire n26354;
wire n26355;
wire n26356;
wire n26357;
wire n26358;
wire n26359;
wire n26360;
wire n26361;
wire n26362;
wire n26363;
wire n26364;
wire n26365;
wire n26366;
wire n26367;
wire n26368;
wire n26369;
wire n2637;
wire n26370;
wire n26371;
wire n26372;
wire n26373;
wire n26374;
wire n26375;
wire n26376;
wire n26377;
wire n26378;
wire n26379;
wire n26380;
wire n26381;
wire n26382;
wire n26383;
wire n26384;
wire n26385;
wire n26386;
wire n26387;
wire n26388;
wire n26389;
wire n26390;
wire n26391;
wire n26392;
wire n26393;
wire n26394;
wire n26395;
wire n26396;
wire n26397;
wire n26398;
wire n26399;
wire n26400;
wire n26401;
wire n26402;
wire n26403;
wire n26404;
wire n26405;
wire n26406;
wire n26407;
wire n26408;
wire n26409;
wire n26410;
wire n26411;
wire n26412;
wire n26413;
wire n26414;
wire n26415;
wire n26416;
wire n26417;
wire n26418;
wire n26419;
wire n2642;
wire n26420;
wire n26421;
wire n26422;
wire n26423;
wire n26424;
wire n26425;
wire n26426;
wire n26427;
wire n26428;
wire n26429;
wire n26430;
wire n26431;
wire n26432;
wire n26433;
wire n26434;
wire n26435;
wire n26436;
wire n26437;
wire n26438;
wire n26439;
wire n26440;
wire n26441;
wire n26442;
wire n26443;
wire n26444;
wire n26445;
wire n26446;
wire n26447;
wire n26448;
wire n26449;
wire n26450;
wire n26451;
wire n26452;
wire n26453;
wire n26454;
wire n26455;
wire n26456;
wire n26457;
wire n26458;
wire n26459;
wire n26460;
wire n26461;
wire n26462;
wire n26463;
wire n26464;
wire n26465;
wire n26466;
wire n26467;
wire n26468;
wire n26469;
wire n2647;
wire n26470;
wire n26471;
wire n26472;
wire n26473;
wire n26474;
wire n26475;
wire n26476;
wire n26477;
wire n26478;
wire n26479;
wire n26480;
wire n26481;
wire n26482;
wire n26483;
wire n26484;
wire n26485;
wire n26486;
wire n26487;
wire n26488;
wire n26489;
wire n26490;
wire n26491;
wire n26492;
wire n26493;
wire n26494;
wire n26495;
wire n26496;
wire n26497;
wire n26498;
wire n26499;
wire n26500;
wire n26501;
wire n26502;
wire n26503;
wire n26504;
wire n26505;
wire n26506;
wire n26507;
wire n26508;
wire n26509;
wire n26510;
wire n26511;
wire n26512;
wire n26513;
wire n26514;
wire n26515;
wire n26516;
wire n26517;
wire n26518;
wire n26519;
wire n2652;
wire n26520;
wire n26521;
wire n26522;
wire n26523;
wire n26524;
wire n26525;
wire n26526;
wire n26527;
wire n26528;
wire n26529;
wire n26530;
wire n26531;
wire n26532;
wire n26533;
wire n26534;
wire n26535;
wire n26536;
wire n26537;
wire n26538;
wire n26539;
wire n26540;
wire n26541;
wire n26542;
wire n26543;
wire n26544;
wire n26545;
wire n26546;
wire n26547;
wire n26548;
wire n26549;
wire n26550;
wire n26551;
wire n26552;
wire n26553;
wire n26554;
wire n26555;
wire n26556;
wire n26557;
wire n26558;
wire n26559;
wire n26560;
wire n26561;
wire n26562;
wire n26563;
wire n26564;
wire n26565;
wire n26566;
wire n26567;
wire n26568;
wire n26569;
wire n2657;
wire n26570;
wire n26571;
wire n26572;
wire n26573;
wire n26574;
wire n26575;
wire n26576;
wire n26577;
wire n26578;
wire n26579;
wire n26580;
wire n26581;
wire n26582;
wire n26583;
wire n26584;
wire n26585;
wire n26586;
wire n26587;
wire n26588;
wire n26589;
wire n26590;
wire n26591;
wire n26592;
wire n26593;
wire n26594;
wire n26595;
wire n26596;
wire n26597;
wire n26598;
wire n26599;
wire n26600;
wire n26601;
wire n26602;
wire n26603;
wire n26604;
wire n26605;
wire n26606;
wire n26607;
wire n26608;
wire n26609;
wire n26610;
wire n26611;
wire n26612;
wire n26613;
wire n26614;
wire n26615;
wire n26616;
wire n26617;
wire n26618;
wire n26619;
wire n2662;
wire n26620;
wire n26621;
wire n26622;
wire n26623;
wire n26624;
wire n26625;
wire n26626;
wire n26627;
wire n26628;
wire n26629;
wire n26630;
wire n26631;
wire n26632;
wire n26633;
wire n26634;
wire n26635;
wire n26636;
wire n26637;
wire n26638;
wire n26639;
wire n26640;
wire n26641;
wire n26642;
wire n26643;
wire n26644;
wire n26645;
wire n26646;
wire n26647;
wire n26648;
wire n26649;
wire n26650;
wire n26651;
wire n26652;
wire n26653;
wire n26654;
wire n26655;
wire n26656;
wire n26657;
wire n26658;
wire n26659;
wire n26660;
wire n26661;
wire n26662;
wire n26663;
wire n26664;
wire n26665;
wire n26666;
wire n26667;
wire n26668;
wire n26669;
wire n2667;
wire n26670;
wire n26671;
wire n26672;
wire n26673;
wire n26674;
wire n26675;
wire n26676;
wire n26677;
wire n26678;
wire n26679;
wire n26680;
wire n26681;
wire n26682;
wire n26683;
wire n26684;
wire n26685;
wire n26686;
wire n26687;
wire n26688;
wire n26689;
wire n26690;
wire n26691;
wire n26692;
wire n26693;
wire n26694;
wire n26695;
wire n26696;
wire n26697;
wire n26698;
wire n26699;
wire n26700;
wire n26701;
wire n26702;
wire n26703;
wire n26704;
wire n26705;
wire n26706;
wire n26707;
wire n26708;
wire n26709;
wire n26710;
wire n26711;
wire n26712;
wire n26713;
wire n26714;
wire n26715;
wire n26716;
wire n26717;
wire n26718;
wire n26719;
wire n2672;
wire n26720;
wire n26721;
wire n26722;
wire n26723;
wire n26724;
wire n26725;
wire n26726;
wire n26727;
wire n26728;
wire n26729;
wire n26730;
wire n26731;
wire n26732;
wire n26733;
wire n26734;
wire n26735;
wire n26736;
wire n26737;
wire n26738;
wire n26739;
wire n26740;
wire n26741;
wire n26742;
wire n26743;
wire n26744;
wire n26745;
wire n26746;
wire n26747;
wire n26748;
wire n26749;
wire n26750;
wire n26751;
wire n26752;
wire n26753;
wire n26754;
wire n26755;
wire n26756;
wire n26757;
wire n26758;
wire n26759;
wire n26760;
wire n26761;
wire n26762;
wire n26763;
wire n26764;
wire n26765;
wire n26766;
wire n26767;
wire n26768;
wire n26769;
wire n2677;
wire n26770;
wire n26771;
wire n26772;
wire n26773;
wire n26774;
wire n26775;
wire n26776;
wire n26777;
wire n26778;
wire n26779;
wire n26780;
wire n26781;
wire n26782;
wire n26783;
wire n26784;
wire n26785;
wire n26786;
wire n26787;
wire n26788;
wire n26789;
wire n26790;
wire n26791;
wire n26792;
wire n26793;
wire n26794;
wire n26795;
wire n26796;
wire n26797;
wire n26798;
wire n26799;
wire n268;
wire n26800;
wire n26801;
wire n26802;
wire n26803;
wire n26804;
wire n26805;
wire n26806;
wire n26807;
wire n26808;
wire n26809;
wire n26810;
wire n26811;
wire n26812;
wire n26813;
wire n26814;
wire n26815;
wire n26816;
wire n26817;
wire n26818;
wire n26819;
wire n2682;
wire n26820;
wire n26821;
wire n26822;
wire n26823;
wire n26824;
wire n26825;
wire n26826;
wire n26827;
wire n26828;
wire n26829;
wire n26830;
wire n26831;
wire n26832;
wire n26833;
wire n26834;
wire n26835;
wire n26836;
wire n26837;
wire n26838;
wire n26839;
wire n26840;
wire n26841;
wire n26842;
wire n26843;
wire n26844;
wire n26845;
wire n26846;
wire n26847;
wire n26848;
wire n26849;
wire n26850;
wire n26851;
wire n26852;
wire n26853;
wire n26854;
wire n26855;
wire n26856;
wire n26857;
wire n26858;
wire n26859;
wire n26860;
wire n26861;
wire n26862;
wire n26863;
wire n26864;
wire n26865;
wire n26866;
wire n26867;
wire n26868;
wire n26869;
wire n2687;
wire n26870;
wire n26871;
wire n26872;
wire n26873;
wire n26874;
wire n26875;
wire n26876;
wire n26877;
wire n26878;
wire n26879;
wire n26880;
wire n26881;
wire n26882;
wire n26883;
wire n26884;
wire n26885;
wire n26886;
wire n26887;
wire n26888;
wire n26889;
wire n26890;
wire n26891;
wire n26892;
wire n26893;
wire n26894;
wire n26895;
wire n26896;
wire n26897;
wire n26898;
wire n26899;
wire n26900;
wire n26901;
wire n26902;
wire n26903;
wire n26904;
wire n26905;
wire n26906;
wire n26907;
wire n26908;
wire n26909;
wire n26910;
wire n26911;
wire n26912;
wire n26913;
wire n26914;
wire n26915;
wire n26916;
wire n26917;
wire n26918;
wire n26919;
wire n2692;
wire n26920;
wire n26921;
wire n26922;
wire n26923;
wire n26924;
wire n26925;
wire n26926;
wire n26927;
wire n26928;
wire n26929;
wire n26930;
wire n26931;
wire n26932;
wire n26933;
wire n26934;
wire n26935;
wire n26936;
wire n26937;
wire n26938;
wire n26939;
wire n26940;
wire n26941;
wire n26942;
wire n26943;
wire n26944;
wire n26945;
wire n26946;
wire n26947;
wire n26948;
wire n26949;
wire n26950;
wire n26951;
wire n26952;
wire n26953;
wire n26954;
wire n26955;
wire n26956;
wire n26957;
wire n26958;
wire n26959;
wire n26960;
wire n26961;
wire n26962;
wire n26963;
wire n26964;
wire n26965;
wire n26966;
wire n26967;
wire n26968;
wire n26969;
wire n2697;
wire n26970;
wire n26971;
wire n26972;
wire n26973;
wire n26974;
wire n26975;
wire n26976;
wire n26977;
wire n26978;
wire n26979;
wire n26980;
wire n26981;
wire n26982;
wire n26983;
wire n26984;
wire n26985;
wire n26986;
wire n26987;
wire n26988;
wire n26989;
wire n26990;
wire n26991;
wire n26992;
wire n26993;
wire n26994;
wire n26995;
wire n26996;
wire n26997;
wire n26998;
wire n26999;
wire n27000;
wire n27001;
wire n27002;
wire n27003;
wire n27004;
wire n27005;
wire n27006;
wire n27007;
wire n27008;
wire n27009;
wire n27010;
wire n27011;
wire n27012;
wire n27013;
wire n27014;
wire n27015;
wire n27016;
wire n27017;
wire n27018;
wire n27019;
wire n2702;
wire n27020;
wire n27021;
wire n27022;
wire n27023;
wire n27024;
wire n27025;
wire n27026;
wire n27027;
wire n27028;
wire n27029;
wire n27030;
wire n27031;
wire n27032;
wire n27033;
wire n27034;
wire n27035;
wire n27036;
wire n27037;
wire n27038;
wire n27039;
wire n27040;
wire n27041;
wire n27042;
wire n27043;
wire n27044;
wire n27045;
wire n27046;
wire n27047;
wire n27048;
wire n27049;
wire n27050;
wire n27051;
wire n27052;
wire n27053;
wire n27054;
wire n27055;
wire n27056;
wire n27057;
wire n27058;
wire n27059;
wire n27060;
wire n27061;
wire n27062;
wire n27063;
wire n27064;
wire n27065;
wire n27066;
wire n27067;
wire n27068;
wire n27069;
wire n2707;
wire n27070;
wire n27071;
wire n27072;
wire n27073;
wire n27074;
wire n27075;
wire n27076;
wire n27077;
wire n27078;
wire n27079;
wire n27080;
wire n27081;
wire n27082;
wire n27083;
wire n27084;
wire n27085;
wire n27086;
wire n27087;
wire n27088;
wire n27089;
wire n27090;
wire n27091;
wire n27092;
wire n27093;
wire n27094;
wire n27095;
wire n27096;
wire n27097;
wire n27098;
wire n27099;
wire n27100;
wire n27101;
wire n27102;
wire n27103;
wire n27104;
wire n27105;
wire n27106;
wire n27107;
wire n27108;
wire n27109;
wire n27110;
wire n27111;
wire n27112;
wire n27113;
wire n27114;
wire n27115;
wire n27116;
wire n27117;
wire n27118;
wire n27119;
wire n2712;
wire n27120;
wire n27121;
wire n27122;
wire n27123;
wire n27124;
wire n27125;
wire n27126;
wire n27127;
wire n27128;
wire n27129;
wire n27130;
wire n27131;
wire n27132;
wire n27133;
wire n27134;
wire n27135;
wire n27136;
wire n27137;
wire n27138;
wire n27139;
wire n27140;
wire n27141;
wire n27142;
wire n27143;
wire n27144;
wire n27145;
wire n27146;
wire n27147;
wire n27148;
wire n27149;
wire n27150;
wire n27151;
wire n27152;
wire n27153;
wire n27154;
wire n27155;
wire n27156;
wire n27157;
wire n27158;
wire n27159;
wire n27160;
wire n27161;
wire n27162;
wire n27163;
wire n27164;
wire n27165;
wire n27166;
wire n27167;
wire n27168;
wire n27169;
wire n2717;
wire n27170;
wire n27171;
wire n27172;
wire n27173;
wire n27174;
wire n27175;
wire n27176;
wire n27177;
wire n27178;
wire n27179;
wire n27180;
wire n27181;
wire n27182;
wire n27183;
wire n27184;
wire n27185;
wire n27186;
wire n27187;
wire n27188;
wire n27189;
wire n27190;
wire n27191;
wire n27192;
wire n27193;
wire n27194;
wire n27195;
wire n27196;
wire n27197;
wire n27198;
wire n27199;
wire n27200;
wire n27201;
wire n27202;
wire n27203;
wire n27204;
wire n27205;
wire n27206;
wire n27207;
wire n27208;
wire n27209;
wire n27210;
wire n27211;
wire n27212;
wire n27213;
wire n27214;
wire n27215;
wire n27216;
wire n27217;
wire n27218;
wire n27219;
wire n2722;
wire n27220;
wire n27221;
wire n27222;
wire n27223;
wire n27224;
wire n27225;
wire n27226;
wire n27227;
wire n27228;
wire n27229;
wire n27230;
wire n27231;
wire n27232;
wire n27233;
wire n27234;
wire n27235;
wire n27236;
wire n27237;
wire n27238;
wire n27239;
wire n27240;
wire n27241;
wire n27242;
wire n27243;
wire n27244;
wire n27245;
wire n27246;
wire n27247;
wire n27248;
wire n27249;
wire n27250;
wire n27251;
wire n27252;
wire n27253;
wire n27254;
wire n27255;
wire n27256;
wire n27257;
wire n27259;
wire n27260;
wire n27261;
wire n27262;
wire n27263;
wire n27264;
wire n27265;
wire n27266;
wire n27267;
wire n27268;
wire n27269;
wire n2727;
wire n27270;
wire n27271;
wire n27272;
wire n27273;
wire n27274;
wire n27275;
wire n27276;
wire n27277;
wire n27278;
wire n27279;
wire n27280;
wire n27281;
wire n27282;
wire n27283;
wire n27284;
wire n27285;
wire n27286;
wire n27287;
wire n27288;
wire n27289;
wire n27290;
wire n27291;
wire n27292;
wire n27293;
wire n27294;
wire n27295;
wire n27296;
wire n27297;
wire n27298;
wire n27299;
wire n273;
wire n27300;
wire n27301;
wire n27302;
wire n27303;
wire n27304;
wire n27305;
wire n27306;
wire n27307;
wire n27308;
wire n27309;
wire n2731;
wire n27310;
wire n27311;
wire n27312;
wire n27313;
wire n27314;
wire n27315;
wire n27316;
wire n27317;
wire n27318;
wire n27319;
wire n27320;
wire n27321;
wire n27322;
wire n27323;
wire n27324;
wire n27325;
wire n27326;
wire n27327;
wire n27328;
wire n27329;
wire n27330;
wire n27331;
wire n27332;
wire n27333;
wire n27334;
wire n27335;
wire n27336;
wire n27337;
wire n27338;
wire n27339;
wire n27340;
wire n27341;
wire n27342;
wire n27343;
wire n27344;
wire n27345;
wire n27346;
wire n27347;
wire n27348;
wire n27349;
wire n27350;
wire n27351;
wire n27352;
wire n27353;
wire n27354;
wire n27355;
wire n27356;
wire n27357;
wire n27358;
wire n27359;
wire n2736;
wire n27360;
wire n27361;
wire n27362;
wire n27363;
wire n27364;
wire n27365;
wire n27366;
wire n27367;
wire n27368;
wire n27369;
wire n27370;
wire n27371;
wire n27372;
wire n27373;
wire n27374;
wire n27375;
wire n27376;
wire n27377;
wire n27378;
wire n27379;
wire n27380;
wire n27381;
wire n27382;
wire n27383;
wire n27384;
wire n27385;
wire n27386;
wire n27387;
wire n27388;
wire n27389;
wire n27390;
wire n27391;
wire n27392;
wire n27393;
wire n27394;
wire n27395;
wire n27396;
wire n27397;
wire n27398;
wire n27399;
wire n27400;
wire n27401;
wire n27402;
wire n27403;
wire n27404;
wire n27405;
wire n27406;
wire n27407;
wire n27408;
wire n27409;
wire n2741;
wire n27410;
wire n27411;
wire n27412;
wire n27413;
wire n27414;
wire n27415;
wire n27416;
wire n27417;
wire n27418;
wire n27419;
wire n27420;
wire n27421;
wire n27422;
wire n27423;
wire n27424;
wire n27425;
wire n27426;
wire n27427;
wire n27428;
wire n27429;
wire n27430;
wire n27431;
wire n27432;
wire n27433;
wire n27434;
wire n27435;
wire n27436;
wire n27437;
wire n27438;
wire n27439;
wire n27440;
wire n27441;
wire n27442;
wire n27443;
wire n27444;
wire n27445;
wire n27446;
wire n27447;
wire n27448;
wire n27449;
wire n27450;
wire n27451;
wire n27452;
wire n27453;
wire n27454;
wire n27455;
wire n27456;
wire n27457;
wire n27458;
wire n27459;
wire n2746;
wire n27460;
wire n27461;
wire n27462;
wire n27463;
wire n27464;
wire n27465;
wire n27466;
wire n27467;
wire n27468;
wire n27469;
wire n27470;
wire n27471;
wire n27472;
wire n27473;
wire n27474;
wire n27475;
wire n27476;
wire n27477;
wire n27478;
wire n27479;
wire n27480;
wire n27481;
wire n27482;
wire n27483;
wire n27484;
wire n27485;
wire n27486;
wire n27487;
wire n27488;
wire n27489;
wire n27490;
wire n27491;
wire n27492;
wire n27493;
wire n27494;
wire n27495;
wire n27496;
wire n27497;
wire n27498;
wire n27499;
wire n27500;
wire n27501;
wire n27502;
wire n27503;
wire n27504;
wire n27505;
wire n27506;
wire n27507;
wire n27508;
wire n27509;
wire n2751;
wire n27510;
wire n27511;
wire n27512;
wire n27513;
wire n27514;
wire n27515;
wire n27516;
wire n27517;
wire n27518;
wire n27519;
wire n27520;
wire n27521;
wire n27522;
wire n27523;
wire n27524;
wire n27525;
wire n27526;
wire n27527;
wire n27528;
wire n27529;
wire n27530;
wire n27531;
wire n27532;
wire n27533;
wire n27534;
wire n27535;
wire n27536;
wire n27537;
wire n27538;
wire n27539;
wire n27540;
wire n27541;
wire n27542;
wire n27543;
wire n27544;
wire n27545;
wire n27546;
wire n27547;
wire n27548;
wire n27549;
wire n27550;
wire n27551;
wire n27552;
wire n27553;
wire n27554;
wire n27555;
wire n27556;
wire n27557;
wire n27558;
wire n27559;
wire n2756;
wire n27560;
wire n27561;
wire n27562;
wire n27563;
wire n27564;
wire n27565;
wire n27566;
wire n27567;
wire n27568;
wire n27569;
wire n27570;
wire n27571;
wire n27572;
wire n27573;
wire n27574;
wire n27575;
wire n27576;
wire n27577;
wire n27578;
wire n27579;
wire n27580;
wire n27581;
wire n27582;
wire n27583;
wire n27584;
wire n27585;
wire n27586;
wire n27587;
wire n27588;
wire n27589;
wire n27590;
wire n27591;
wire n27592;
wire n27593;
wire n27594;
wire n27595;
wire n27596;
wire n27597;
wire n27598;
wire n27599;
wire n27600;
wire n27601;
wire n27602;
wire n27603;
wire n27604;
wire n27605;
wire n27606;
wire n27607;
wire n27608;
wire n27609;
wire n2761;
wire n27610;
wire n27611;
wire n27612;
wire n27613;
wire n27614;
wire n27615;
wire n27616;
wire n27617;
wire n27618;
wire n27619;
wire n27620;
wire n27621;
wire n27622;
wire n27623;
wire n27624;
wire n27625;
wire n27626;
wire n27627;
wire n27628;
wire n27629;
wire n27630;
wire n27631;
wire n27632;
wire n27633;
wire n27634;
wire n27635;
wire n27636;
wire n27637;
wire n27638;
wire n27639;
wire n27640;
wire n27641;
wire n27642;
wire n27643;
wire n27644;
wire n27645;
wire n27646;
wire n27647;
wire n27648;
wire n27649;
wire n27650;
wire n27651;
wire n27652;
wire n27653;
wire n27654;
wire n27655;
wire n27656;
wire n27657;
wire n27658;
wire n27659;
wire n2766;
wire n27660;
wire n27661;
wire n27662;
wire n27663;
wire n27664;
wire n27665;
wire n27666;
wire n27667;
wire n27668;
wire n27669;
wire n27670;
wire n27671;
wire n27672;
wire n27673;
wire n27674;
wire n27675;
wire n27676;
wire n27677;
wire n27678;
wire n27679;
wire n27681;
wire n27682;
wire n27683;
wire n27684;
wire n27685;
wire n27686;
wire n27687;
wire n27688;
wire n27689;
wire n27690;
wire n27691;
wire n27692;
wire n27693;
wire n27694;
wire n27695;
wire n27696;
wire n27697;
wire n27698;
wire n27699;
wire n27700;
wire n27701;
wire n27702;
wire n27703;
wire n27704;
wire n27705;
wire n27706;
wire n27707;
wire n27708;
wire n27709;
wire n2771;
wire n27710;
wire n27711;
wire n27712;
wire n27713;
wire n27714;
wire n27715;
wire n27716;
wire n27717;
wire n27718;
wire n27719;
wire n27720;
wire n27721;
wire n27722;
wire n27723;
wire n27724;
wire n27725;
wire n27726;
wire n27727;
wire n27728;
wire n27729;
wire n27730;
wire n27731;
wire n27732;
wire n27733;
wire n27734;
wire n27735;
wire n27736;
wire n27737;
wire n27738;
wire n27739;
wire n27740;
wire n27741;
wire n27742;
wire n27743;
wire n27744;
wire n27745;
wire n27746;
wire n27747;
wire n27748;
wire n27749;
wire n27750;
wire n27751;
wire n27752;
wire n27753;
wire n27754;
wire n27755;
wire n27756;
wire n27757;
wire n27758;
wire n27759;
wire n2776;
wire n27760;
wire n27761;
wire n27762;
wire n27763;
wire n27764;
wire n27765;
wire n27766;
wire n27767;
wire n27768;
wire n27769;
wire n27770;
wire n27771;
wire n27772;
wire n27773;
wire n27774;
wire n27775;
wire n27776;
wire n27777;
wire n27778;
wire n27779;
wire n27780;
wire n27781;
wire n27782;
wire n27783;
wire n27784;
wire n27785;
wire n27786;
wire n27787;
wire n27788;
wire n27789;
wire n27790;
wire n27791;
wire n27792;
wire n27793;
wire n27794;
wire n27795;
wire n27796;
wire n27797;
wire n27798;
wire n27799;
wire n278;
wire n27800;
wire n27801;
wire n27802;
wire n27803;
wire n27804;
wire n27805;
wire n27806;
wire n27807;
wire n27808;
wire n27809;
wire n2781;
wire n27810;
wire n27811;
wire n27812;
wire n27813;
wire n27814;
wire n27815;
wire n27816;
wire n27817;
wire n27818;
wire n27819;
wire n27820;
wire n27821;
wire n27822;
wire n27823;
wire n27824;
wire n27825;
wire n27826;
wire n27827;
wire n27828;
wire n27829;
wire n27830;
wire n27831;
wire n27832;
wire n27833;
wire n27834;
wire n27835;
wire n27836;
wire n27837;
wire n27838;
wire n27839;
wire n27840;
wire n27841;
wire n27842;
wire n27843;
wire n27844;
wire n27845;
wire n27846;
wire n27847;
wire n27848;
wire n27849;
wire n27850;
wire n27851;
wire n27852;
wire n27853;
wire n27854;
wire n27855;
wire n27856;
wire n27857;
wire n27858;
wire n27859;
wire n2786;
wire n27860;
wire n27861;
wire n27862;
wire n27863;
wire n27864;
wire n27865;
wire n27866;
wire n27867;
wire n27868;
wire n27869;
wire n27870;
wire n27871;
wire n27872;
wire n27873;
wire n27874;
wire n27875;
wire n27876;
wire n27877;
wire n27878;
wire n27879;
wire n27880;
wire n27881;
wire n27882;
wire n27883;
wire n27884;
wire n27885;
wire n27886;
wire n27887;
wire n27888;
wire n27889;
wire n27890;
wire n27891;
wire n27892;
wire n27893;
wire n27894;
wire n27895;
wire n27896;
wire n27897;
wire n27898;
wire n27899;
wire n27900;
wire n27901;
wire n27902;
wire n27903;
wire n27904;
wire n27905;
wire n27906;
wire n27907;
wire n27908;
wire n27909;
wire n2791;
wire n27910;
wire n27911;
wire n27912;
wire n27913;
wire n27914;
wire n27915;
wire n27916;
wire n27917;
wire n27918;
wire n27919;
wire n27920;
wire n27921;
wire n27922;
wire n27923;
wire n27924;
wire n27925;
wire n27926;
wire n27927;
wire n27928;
wire n27929;
wire n27930;
wire n27931;
wire n27932;
wire n27933;
wire n27934;
wire n27935;
wire n27936;
wire n27937;
wire n27938;
wire n27939;
wire n27940;
wire n27941;
wire n27942;
wire n27943;
wire n27944;
wire n27945;
wire n27946;
wire n27947;
wire n27948;
wire n27949;
wire n27950;
wire n27951;
wire n27952;
wire n27953;
wire n27954;
wire n27955;
wire n27956;
wire n27957;
wire n27958;
wire n27959;
wire n2796;
wire n27960;
wire n27961;
wire n27962;
wire n27963;
wire n27964;
wire n27965;
wire n27966;
wire n27967;
wire n27968;
wire n27969;
wire n27970;
wire n27971;
wire n27972;
wire n27973;
wire n27974;
wire n27975;
wire n27976;
wire n27977;
wire n27978;
wire n27979;
wire n27980;
wire n27981;
wire n27982;
wire n27983;
wire n27984;
wire n27985;
wire n27986;
wire n27987;
wire n27988;
wire n27989;
wire n27990;
wire n27991;
wire n27992;
wire n27993;
wire n27994;
wire n27995;
wire n27996;
wire n27997;
wire n27998;
wire n27999;
wire n28000;
wire n28001;
wire n28002;
wire n28003;
wire n28004;
wire n28005;
wire n28006;
wire n28007;
wire n28008;
wire n28009;
wire n2801;
wire n28010;
wire n28011;
wire n28012;
wire n28013;
wire n28014;
wire n28015;
wire n28016;
wire n28017;
wire n28018;
wire n28019;
wire n28020;
wire n28021;
wire n28022;
wire n28023;
wire n28024;
wire n28025;
wire n28026;
wire n28027;
wire n28028;
wire n28029;
wire n28030;
wire n28031;
wire n28032;
wire n28033;
wire n28034;
wire n28035;
wire n28036;
wire n28037;
wire n28038;
wire n28039;
wire n28040;
wire n28041;
wire n28042;
wire n28043;
wire n28044;
wire n28045;
wire n28046;
wire n28047;
wire n28048;
wire n28049;
wire n28050;
wire n28051;
wire n28052;
wire n28053;
wire n28054;
wire n28055;
wire n28056;
wire n28057;
wire n28058;
wire n28059;
wire n2806;
wire n28060;
wire n28061;
wire n28062;
wire n28063;
wire n28064;
wire n28065;
wire n28066;
wire n28067;
wire n28068;
wire n28069;
wire n28070;
wire n28071;
wire n28072;
wire n28073;
wire n28074;
wire n28075;
wire n28076;
wire n28077;
wire n28078;
wire n28079;
wire n28080;
wire n28081;
wire n28082;
wire n28083;
wire n28084;
wire n28085;
wire n28086;
wire n28087;
wire n28088;
wire n28089;
wire n28090;
wire n28091;
wire n28092;
wire n28093;
wire n28094;
wire n28095;
wire n28096;
wire n28097;
wire n28098;
wire n28099;
wire n28100;
wire n28101;
wire n28102;
wire n28103;
wire n28104;
wire n28105;
wire n28106;
wire n28107;
wire n28108;
wire n28109;
wire n2811;
wire n28110;
wire n28111;
wire n28112;
wire n28113;
wire n28114;
wire n28115;
wire n28116;
wire n28117;
wire n28118;
wire n28119;
wire n28120;
wire n28121;
wire n28122;
wire n28123;
wire n28124;
wire n28125;
wire n28126;
wire n28127;
wire n28128;
wire n28129;
wire n28130;
wire n28131;
wire n28132;
wire n28133;
wire n28134;
wire n28135;
wire n28136;
wire n28137;
wire n28138;
wire n28139;
wire n28140;
wire n28141;
wire n28142;
wire n28143;
wire n28144;
wire n28145;
wire n28146;
wire n28147;
wire n28148;
wire n28149;
wire n28150;
wire n28151;
wire n28152;
wire n28153;
wire n28154;
wire n28155;
wire n28156;
wire n28157;
wire n28158;
wire n28159;
wire n2816;
wire n28160;
wire n28161;
wire n28162;
wire n28163;
wire n28164;
wire n28165;
wire n28166;
wire n28167;
wire n28168;
wire n28169;
wire n28170;
wire n28171;
wire n28172;
wire n28173;
wire n28174;
wire n28175;
wire n28176;
wire n28177;
wire n28178;
wire n28179;
wire n28180;
wire n28181;
wire n28182;
wire n28183;
wire n28184;
wire n28185;
wire n28186;
wire n28187;
wire n28188;
wire n28189;
wire n28190;
wire n28191;
wire n28192;
wire n28193;
wire n28194;
wire n28195;
wire n28196;
wire n28197;
wire n28198;
wire n28199;
wire n28200;
wire n28201;
wire n28202;
wire n28203;
wire n28204;
wire n28205;
wire n28206;
wire n28207;
wire n28208;
wire n28209;
wire n2821;
wire n28210;
wire n28211;
wire n28212;
wire n28213;
wire n28214;
wire n28215;
wire n28216;
wire n28217;
wire n28218;
wire n28219;
wire n28220;
wire n28221;
wire n28222;
wire n28223;
wire n28224;
wire n28225;
wire n28226;
wire n28227;
wire n28228;
wire n28229;
wire n28230;
wire n28231;
wire n28232;
wire n28233;
wire n28234;
wire n28235;
wire n28236;
wire n28237;
wire n28238;
wire n28239;
wire n28240;
wire n28241;
wire n28242;
wire n28243;
wire n28244;
wire n28245;
wire n28246;
wire n28247;
wire n28248;
wire n28249;
wire n28250;
wire n28251;
wire n28252;
wire n28253;
wire n28254;
wire n28255;
wire n28256;
wire n28257;
wire n28258;
wire n28259;
wire n2826;
wire n28260;
wire n28261;
wire n28262;
wire n28263;
wire n28264;
wire n28265;
wire n28266;
wire n28267;
wire n28268;
wire n28269;
wire n28270;
wire n28271;
wire n28272;
wire n28273;
wire n28274;
wire n28275;
wire n28276;
wire n28277;
wire n28278;
wire n28279;
wire n28280;
wire n28281;
wire n28282;
wire n28283;
wire n28284;
wire n28285;
wire n28286;
wire n28287;
wire n28288;
wire n28289;
wire n28290;
wire n28291;
wire n28292;
wire n28293;
wire n28294;
wire n28295;
wire n28296;
wire n28297;
wire n28298;
wire n28299;
wire n283;
wire n28300;
wire n28301;
wire n28302;
wire n28303;
wire n28304;
wire n28305;
wire n28306;
wire n28307;
wire n28308;
wire n28309;
wire n2831;
wire n28310;
wire n28311;
wire n28312;
wire n28313;
wire n28314;
wire n28315;
wire n28316;
wire n28317;
wire n28318;
wire n28319;
wire n28320;
wire n28321;
wire n28322;
wire n28323;
wire n28324;
wire n28325;
wire n28326;
wire n28327;
wire n28328;
wire n28329;
wire n28330;
wire n28331;
wire n28332;
wire n28333;
wire n28334;
wire n28335;
wire n28336;
wire n28337;
wire n28338;
wire n28339;
wire n28340;
wire n28341;
wire n28342;
wire n28343;
wire n28344;
wire n28345;
wire n28346;
wire n28347;
wire n28348;
wire n28349;
wire n28350;
wire n28351;
wire n28352;
wire n28353;
wire n28354;
wire n28355;
wire n28356;
wire n28357;
wire n28358;
wire n28359;
wire n2836;
wire n28360;
wire n28361;
wire n28362;
wire n28363;
wire n28364;
wire n28365;
wire n28366;
wire n28367;
wire n28368;
wire n28369;
wire n28370;
wire n28371;
wire n28372;
wire n28373;
wire n28374;
wire n28375;
wire n28376;
wire n28377;
wire n28378;
wire n28379;
wire n28380;
wire n28381;
wire n28382;
wire n28383;
wire n28384;
wire n28385;
wire n28386;
wire n28387;
wire n28388;
wire n28389;
wire n28390;
wire n28391;
wire n28392;
wire n28393;
wire n28394;
wire n28395;
wire n28396;
wire n28397;
wire n28398;
wire n28399;
wire n28400;
wire n28401;
wire n28402;
wire n28403;
wire n28404;
wire n28405;
wire n28406;
wire n28407;
wire n28408;
wire n28409;
wire n2841;
wire n28410;
wire n28411;
wire n28412;
wire n28413;
wire n28414;
wire n28415;
wire n28416;
wire n28417;
wire n28418;
wire n28419;
wire n28420;
wire n28421;
wire n28422;
wire n28423;
wire n28424;
wire n28425;
wire n28426;
wire n28427;
wire n28428;
wire n28429;
wire n28430;
wire n28431;
wire n28432;
wire n28433;
wire n28434;
wire n28435;
wire n28436;
wire n28437;
wire n28438;
wire n28439;
wire n28440;
wire n28441;
wire n28442;
wire n28443;
wire n28444;
wire n28445;
wire n28446;
wire n28447;
wire n28448;
wire n28449;
wire n28450;
wire n28451;
wire n28452;
wire n28453;
wire n28454;
wire n28455;
wire n28456;
wire n28457;
wire n28458;
wire n28459;
wire n2846;
wire n28460;
wire n28461;
wire n28462;
wire n28463;
wire n28464;
wire n28465;
wire n28466;
wire n28467;
wire n28468;
wire n28469;
wire n28470;
wire n28471;
wire n28472;
wire n28473;
wire n28474;
wire n28475;
wire n28476;
wire n28477;
wire n28478;
wire n28479;
wire n28480;
wire n28481;
wire n28482;
wire n28483;
wire n28484;
wire n28485;
wire n28486;
wire n28487;
wire n28488;
wire n28489;
wire n28490;
wire n28491;
wire n28492;
wire n28493;
wire n28494;
wire n28495;
wire n28496;
wire n28497;
wire n28498;
wire n28499;
wire n28500;
wire n28501;
wire n28502;
wire n28503;
wire n28504;
wire n28505;
wire n28506;
wire n28507;
wire n28508;
wire n28509;
wire n2851;
wire n28510;
wire n28511;
wire n28512;
wire n28513;
wire n28514;
wire n28515;
wire n28516;
wire n28517;
wire n28518;
wire n28519;
wire n28520;
wire n28521;
wire n28522;
wire n28523;
wire n28524;
wire n28525;
wire n28526;
wire n28527;
wire n28528;
wire n28529;
wire n28530;
wire n28531;
wire n28532;
wire n28533;
wire n28534;
wire n28535;
wire n28536;
wire n28537;
wire n28538;
wire n28539;
wire n28540;
wire n28541;
wire n28542;
wire n28543;
wire n28544;
wire n28545;
wire n28546;
wire n28547;
wire n28548;
wire n28549;
wire n28550;
wire n28551;
wire n28552;
wire n28553;
wire n28554;
wire n28555;
wire n28556;
wire n28557;
wire n28558;
wire n28559;
wire n2856;
wire n28560;
wire n28561;
wire n28562;
wire n28563;
wire n28564;
wire n28565;
wire n28566;
wire n28567;
wire n28568;
wire n28569;
wire n28570;
wire n28571;
wire n28572;
wire n28573;
wire n28574;
wire n28575;
wire n28576;
wire n28577;
wire n28578;
wire n28579;
wire n28580;
wire n28581;
wire n28582;
wire n28583;
wire n28584;
wire n28585;
wire n28586;
wire n28587;
wire n28588;
wire n28589;
wire n28590;
wire n28591;
wire n28592;
wire n28593;
wire n28594;
wire n28595;
wire n28596;
wire n28597;
wire n28598;
wire n28599;
wire n28600;
wire n28601;
wire n28602;
wire n28603;
wire n28604;
wire n28605;
wire n28606;
wire n28607;
wire n28608;
wire n28609;
wire n2861;
wire n28610;
wire n28611;
wire n28612;
wire n28613;
wire n28614;
wire n28615;
wire n28616;
wire n28617;
wire n28618;
wire n28619;
wire n28620;
wire n28621;
wire n28622;
wire n28623;
wire n28624;
wire n28625;
wire n28626;
wire n28627;
wire n28628;
wire n28629;
wire n28630;
wire n28631;
wire n28632;
wire n28633;
wire n28634;
wire n28635;
wire n28636;
wire n28637;
wire n28638;
wire n28639;
wire n28640;
wire n28641;
wire n28642;
wire n28643;
wire n28644;
wire n28645;
wire n28646;
wire n28647;
wire n28648;
wire n28649;
wire n28650;
wire n28651;
wire n28652;
wire n28653;
wire n28654;
wire n28655;
wire n28656;
wire n28657;
wire n28658;
wire n28659;
wire n2866;
wire n28660;
wire n28661;
wire n28662;
wire n28663;
wire n28664;
wire n28665;
wire n28666;
wire n28667;
wire n28668;
wire n28669;
wire n28670;
wire n28671;
wire n28672;
wire n28673;
wire n28674;
wire n28675;
wire n28676;
wire n28677;
wire n28678;
wire n28679;
wire n28680;
wire n28681;
wire n28682;
wire n28683;
wire n28684;
wire n28685;
wire n28686;
wire n28687;
wire n28688;
wire n28689;
wire n28690;
wire n28691;
wire n28692;
wire n28693;
wire n28694;
wire n28695;
wire n28696;
wire n28697;
wire n28698;
wire n28699;
wire n28700;
wire n28701;
wire n28702;
wire n28703;
wire n28704;
wire n28705;
wire n28706;
wire n28707;
wire n28708;
wire n28709;
wire n2871;
wire n28710;
wire n28711;
wire n28712;
wire n28713;
wire n28714;
wire n28715;
wire n28716;
wire n28717;
wire n28718;
wire n28719;
wire n28720;
wire n28721;
wire n28722;
wire n28723;
wire n28724;
wire n28725;
wire n28726;
wire n28727;
wire n28728;
wire n28729;
wire n28730;
wire n28731;
wire n28732;
wire n28733;
wire n28734;
wire n28735;
wire n28736;
wire n28737;
wire n28738;
wire n28739;
wire n28740;
wire n28741;
wire n28742;
wire n28743;
wire n28744;
wire n28745;
wire n28746;
wire n28747;
wire n28748;
wire n28749;
wire n28750;
wire n28751;
wire n28752;
wire n28753;
wire n28754;
wire n28755;
wire n28756;
wire n28757;
wire n28758;
wire n28759;
wire n2876;
wire n28760;
wire n28761;
wire n28762;
wire n28763;
wire n28764;
wire n28765;
wire n28766;
wire n28767;
wire n28768;
wire n28769;
wire n28770;
wire n28771;
wire n28772;
wire n28773;
wire n28774;
wire n28775;
wire n28776;
wire n28777;
wire n28778;
wire n28779;
wire n28780;
wire n28781;
wire n28782;
wire n28783;
wire n28784;
wire n28785;
wire n28786;
wire n28787;
wire n28788;
wire n28789;
wire n28790;
wire n28791;
wire n28792;
wire n28793;
wire n28794;
wire n28795;
wire n28796;
wire n28797;
wire n28798;
wire n28799;
wire n288;
wire n28800;
wire n28801;
wire n28802;
wire n28803;
wire n28804;
wire n28805;
wire n28806;
wire n28807;
wire n28808;
wire n28809;
wire n2881;
wire n28810;
wire n28811;
wire n28812;
wire n28813;
wire n28814;
wire n28815;
wire n28816;
wire n28817;
wire n28818;
wire n28819;
wire n28820;
wire n28821;
wire n28822;
wire n28823;
wire n28824;
wire n28825;
wire n28826;
wire n28827;
wire n28828;
wire n28829;
wire n28830;
wire n28831;
wire n28832;
wire n28833;
wire n28834;
wire n28835;
wire n28836;
wire n28837;
wire n28838;
wire n28839;
wire n28840;
wire n28841;
wire n28842;
wire n28843;
wire n28844;
wire n28845;
wire n28846;
wire n28847;
wire n28848;
wire n28849;
wire n28850;
wire n28851;
wire n28852;
wire n28853;
wire n28854;
wire n28855;
wire n28856;
wire n28857;
wire n28858;
wire n28859;
wire n2886;
wire n28860;
wire n28861;
wire n28862;
wire n28863;
wire n28864;
wire n28865;
wire n28866;
wire n28867;
wire n28868;
wire n28869;
wire n28870;
wire n28871;
wire n28872;
wire n28873;
wire n28874;
wire n28875;
wire n28876;
wire n28877;
wire n28878;
wire n28879;
wire n28880;
wire n28881;
wire n28882;
wire n28883;
wire n28884;
wire n28885;
wire n28886;
wire n28887;
wire n28888;
wire n28889;
wire n28890;
wire n28891;
wire n28892;
wire n28893;
wire n28894;
wire n28895;
wire n28896;
wire n28897;
wire n28898;
wire n28899;
wire n28900;
wire n28901;
wire n28902;
wire n28903;
wire n28904;
wire n28905;
wire n28906;
wire n28907;
wire n28908;
wire n28909;
wire n2891;
wire n28910;
wire n28911;
wire n28912;
wire n28913;
wire n28914;
wire n28915;
wire n28916;
wire n28917;
wire n28918;
wire n28919;
wire n28920;
wire n28921;
wire n28922;
wire n28923;
wire n28924;
wire n28925;
wire n28926;
wire n28927;
wire n28928;
wire n28929;
wire n28930;
wire n28931;
wire n28932;
wire n28933;
wire n28934;
wire n28935;
wire n28936;
wire n28937;
wire n28938;
wire n28939;
wire n28940;
wire n28941;
wire n28942;
wire n28943;
wire n28944;
wire n28945;
wire n28946;
wire n28947;
wire n28948;
wire n28949;
wire n28950;
wire n28951;
wire n28952;
wire n28953;
wire n28954;
wire n28955;
wire n28956;
wire n28957;
wire n28958;
wire n28959;
wire n2896;
wire n28960;
wire n28961;
wire n28962;
wire n28963;
wire n28964;
wire n28965;
wire n28966;
wire n28967;
wire n28968;
wire n28969;
wire n28970;
wire n28971;
wire n28972;
wire n28973;
wire n28974;
wire n28975;
wire n28976;
wire n28977;
wire n28978;
wire n28979;
wire n28980;
wire n28981;
wire n28982;
wire n28983;
wire n28984;
wire n28985;
wire n28986;
wire n28987;
wire n28988;
wire n28989;
wire n28990;
wire n28991;
wire n28992;
wire n28993;
wire n28994;
wire n28995;
wire n28996;
wire n28997;
wire n28998;
wire n28999;
wire n29000;
wire n29001;
wire n29002;
wire n29003;
wire n29004;
wire n29005;
wire n29006;
wire n29007;
wire n29008;
wire n29009;
wire n2901;
wire n29010;
wire n29011;
wire n29012;
wire n29013;
wire n29014;
wire n29015;
wire n29016;
wire n29017;
wire n29018;
wire n29019;
wire n29020;
wire n29021;
wire n29022;
wire n29023;
wire n29024;
wire n29025;
wire n29026;
wire n29027;
wire n29028;
wire n29029;
wire n29030;
wire n29031;
wire n29032;
wire n29033;
wire n29034;
wire n29035;
wire n29036;
wire n29037;
wire n29038;
wire n29039;
wire n29040;
wire n29041;
wire n29042;
wire n29043;
wire n29044;
wire n29045;
wire n29046;
wire n29047;
wire n29048;
wire n29049;
wire n29050;
wire n29051;
wire n29052;
wire n29053;
wire n29054;
wire n29055;
wire n29056;
wire n29057;
wire n29058;
wire n29059;
wire n2906;
wire n29060;
wire n29061;
wire n29062;
wire n29063;
wire n29064;
wire n29065;
wire n29066;
wire n29067;
wire n29068;
wire n29069;
wire n29070;
wire n29071;
wire n29072;
wire n29073;
wire n29074;
wire n29075;
wire n29076;
wire n29077;
wire n29078;
wire n29079;
wire n29080;
wire n29081;
wire n29082;
wire n29083;
wire n29084;
wire n29085;
wire n29086;
wire n29087;
wire n29088;
wire n29089;
wire n29090;
wire n29091;
wire n29092;
wire n29093;
wire n29094;
wire n29095;
wire n29096;
wire n29097;
wire n29098;
wire n29099;
wire n29100;
wire n29101;
wire n29102;
wire n29103;
wire n29104;
wire n29105;
wire n29106;
wire n29107;
wire n29108;
wire n29109;
wire n2911;
wire n29110;
wire n29111;
wire n29112;
wire n29113;
wire n29114;
wire n29115;
wire n29116;
wire n29117;
wire n29118;
wire n29119;
wire n29120;
wire n29121;
wire n29122;
wire n29123;
wire n29124;
wire n29125;
wire n29126;
wire n29127;
wire n29128;
wire n29129;
wire n29130;
wire n29131;
wire n29132;
wire n29133;
wire n29134;
wire n29135;
wire n29136;
wire n29137;
wire n29138;
wire n29139;
wire n29140;
wire n29141;
wire n29142;
wire n29143;
wire n29144;
wire n29145;
wire n29146;
wire n29147;
wire n29148;
wire n29149;
wire n29150;
wire n29151;
wire n29152;
wire n29153;
wire n29154;
wire n29155;
wire n29156;
wire n29157;
wire n29158;
wire n29159;
wire n2916;
wire n29160;
wire n29161;
wire n29162;
wire n29163;
wire n29164;
wire n29165;
wire n29166;
wire n29167;
wire n29168;
wire n29169;
wire n29170;
wire n29171;
wire n29172;
wire n29173;
wire n29174;
wire n29175;
wire n29176;
wire n29177;
wire n29178;
wire n29179;
wire n29180;
wire n29181;
wire n29182;
wire n29183;
wire n29184;
wire n29185;
wire n29186;
wire n29187;
wire n29188;
wire n29189;
wire n29190;
wire n29191;
wire n29192;
wire n29193;
wire n29194;
wire n29195;
wire n29196;
wire n29197;
wire n29198;
wire n29199;
wire n29200;
wire n29201;
wire n29202;
wire n29203;
wire n29204;
wire n29205;
wire n29206;
wire n29207;
wire n29208;
wire n29209;
wire n2921;
wire n29210;
wire n29211;
wire n29212;
wire n29213;
wire n29214;
wire n29215;
wire n29216;
wire n29217;
wire n29218;
wire n29219;
wire n29220;
wire n29221;
wire n29222;
wire n29223;
wire n29224;
wire n29225;
wire n29226;
wire n29227;
wire n29228;
wire n29229;
wire n29230;
wire n29231;
wire n29232;
wire n29233;
wire n29234;
wire n29235;
wire n29236;
wire n29237;
wire n29238;
wire n29239;
wire n29240;
wire n29241;
wire n29242;
wire n29243;
wire n29244;
wire n29245;
wire n29246;
wire n29247;
wire n29248;
wire n29249;
wire n29250;
wire n29251;
wire n29252;
wire n29253;
wire n29254;
wire n29255;
wire n29256;
wire n29257;
wire n29258;
wire n29259;
wire n2926;
wire n29260;
wire n29261;
wire n29262;
wire n29263;
wire n29264;
wire n29265;
wire n29266;
wire n29267;
wire n29268;
wire n29269;
wire n29270;
wire n29271;
wire n29272;
wire n29273;
wire n29274;
wire n29275;
wire n29276;
wire n29277;
wire n29278;
wire n29279;
wire n29280;
wire n29281;
wire n29282;
wire n29283;
wire n29284;
wire n29285;
wire n29286;
wire n29287;
wire n29288;
wire n29289;
wire n29290;
wire n29291;
wire n29292;
wire n29293;
wire n29294;
wire n29295;
wire n29296;
wire n29297;
wire n29298;
wire n29299;
wire n293;
wire n29300;
wire n29301;
wire n29302;
wire n29303;
wire n29304;
wire n29305;
wire n29306;
wire n29307;
wire n29308;
wire n29309;
wire n2931;
wire n29310;
wire n29311;
wire n29312;
wire n29313;
wire n29314;
wire n29315;
wire n29316;
wire n29317;
wire n29318;
wire n29319;
wire n29320;
wire n29321;
wire n29322;
wire n29323;
wire n29324;
wire n29325;
wire n29326;
wire n29327;
wire n29328;
wire n29329;
wire n29330;
wire n29331;
wire n29332;
wire n29333;
wire n29334;
wire n29335;
wire n29336;
wire n29337;
wire n29338;
wire n29339;
wire n29340;
wire n29341;
wire n29342;
wire n29343;
wire n29344;
wire n29345;
wire n29346;
wire n29347;
wire n29348;
wire n29349;
wire n29350;
wire n29351;
wire n29352;
wire n29353;
wire n29354;
wire n29355;
wire n29356;
wire n29357;
wire n29358;
wire n29359;
wire n2936;
wire n29360;
wire n29361;
wire n29362;
wire n29363;
wire n29364;
wire n29365;
wire n29366;
wire n29367;
wire n29368;
wire n29369;
wire n29370;
wire n29371;
wire n29372;
wire n29373;
wire n29374;
wire n29375;
wire n29376;
wire n29377;
wire n29378;
wire n29379;
wire n29380;
wire n29381;
wire n29382;
wire n29383;
wire n29384;
wire n29385;
wire n29386;
wire n29387;
wire n29388;
wire n29389;
wire n29390;
wire n29391;
wire n29392;
wire n29393;
wire n29394;
wire n29395;
wire n29396;
wire n29397;
wire n29398;
wire n29399;
wire n29400;
wire n29401;
wire n29402;
wire n29403;
wire n29404;
wire n29405;
wire n29406;
wire n29407;
wire n29408;
wire n29409;
wire n2941;
wire n29410;
wire n29411;
wire n29412;
wire n29413;
wire n29414;
wire n29415;
wire n29416;
wire n29417;
wire n29418;
wire n29419;
wire n29420;
wire n29421;
wire n29422;
wire n29423;
wire n29424;
wire n29425;
wire n29426;
wire n29427;
wire n29428;
wire n29429;
wire n29430;
wire n29431;
wire n29432;
wire n29433;
wire n29434;
wire n29435;
wire n29436;
wire n29437;
wire n29438;
wire n29439;
wire n29440;
wire n29441;
wire n29442;
wire n29443;
wire n29444;
wire n29445;
wire n29446;
wire n29447;
wire n29448;
wire n29449;
wire n29450;
wire n29451;
wire n29452;
wire n29453;
wire n29454;
wire n29455;
wire n29456;
wire n29457;
wire n29458;
wire n29459;
wire n2946;
wire n29460;
wire n29461;
wire n29462;
wire n29463;
wire n29464;
wire n29465;
wire n29466;
wire n29467;
wire n29468;
wire n29469;
wire n29470;
wire n29471;
wire n29472;
wire n29473;
wire n29474;
wire n29475;
wire n29476;
wire n29477;
wire n29478;
wire n29479;
wire n29480;
wire n29481;
wire n29482;
wire n29483;
wire n29484;
wire n29485;
wire n29486;
wire n29487;
wire n29488;
wire n29489;
wire n29490;
wire n29491;
wire n29492;
wire n29493;
wire n29494;
wire n29495;
wire n29496;
wire n29497;
wire n29498;
wire n29499;
wire n29500;
wire n29501;
wire n29502;
wire n29503;
wire n29504;
wire n29505;
wire n29506;
wire n29507;
wire n29508;
wire n29509;
wire n2951;
wire n29510;
wire n29511;
wire n29512;
wire n29513;
wire n29514;
wire n29515;
wire n29516;
wire n29517;
wire n29518;
wire n29519;
wire n29520;
wire n29521;
wire n29522;
wire n29523;
wire n29524;
wire n29525;
wire n29526;
wire n29527;
wire n29528;
wire n29529;
wire n29530;
wire n29531;
wire n29532;
wire n29533;
wire n29534;
wire n29535;
wire n29536;
wire n29537;
wire n29538;
wire n29539;
wire n29540;
wire n29541;
wire n29542;
wire n29543;
wire n29544;
wire n29545;
wire n29546;
wire n29547;
wire n29548;
wire n29549;
wire n29550;
wire n29551;
wire n29552;
wire n29553;
wire n29554;
wire n29555;
wire n29556;
wire n29557;
wire n29558;
wire n29559;
wire n2956;
wire n29560;
wire n29561;
wire n29562;
wire n29563;
wire n29564;
wire n29565;
wire n29566;
wire n29567;
wire n29568;
wire n29569;
wire n29570;
wire n29571;
wire n29572;
wire n29573;
wire n29574;
wire n29575;
wire n29576;
wire n29577;
wire n29578;
wire n29579;
wire n29580;
wire n29581;
wire n29582;
wire n29583;
wire n29584;
wire n29585;
wire n29586;
wire n29587;
wire n29588;
wire n29589;
wire n29590;
wire n29591;
wire n29592;
wire n29593;
wire n29594;
wire n29595;
wire n29596;
wire n29597;
wire n29598;
wire n29599;
wire n29600;
wire n29601;
wire n29602;
wire n29603;
wire n29604;
wire n29605;
wire n29606;
wire n29607;
wire n29608;
wire n29609;
wire n2961;
wire n29610;
wire n29611;
wire n29612;
wire n29613;
wire n29614;
wire n29615;
wire n29616;
wire n29617;
wire n29618;
wire n29619;
wire n29620;
wire n29621;
wire n29622;
wire n29623;
wire n29624;
wire n29625;
wire n29626;
wire n29627;
wire n29628;
wire n29629;
wire n29630;
wire n29631;
wire n29632;
wire n29633;
wire n29634;
wire n29635;
wire n29636;
wire n29637;
wire n29638;
wire n29639;
wire n29640;
wire n29641;
wire n29642;
wire n29643;
wire n29644;
wire n29645;
wire n29646;
wire n29647;
wire n29648;
wire n29649;
wire n29650;
wire n29651;
wire n29652;
wire n29653;
wire n29654;
wire n29655;
wire n29656;
wire n29657;
wire n29658;
wire n29659;
wire n2966;
wire n29660;
wire n29661;
wire n29662;
wire n29663;
wire n29664;
wire n29665;
wire n29666;
wire n29667;
wire n29668;
wire n29669;
wire n29670;
wire n29671;
wire n29672;
wire n29673;
wire n29674;
wire n29675;
wire n29676;
wire n29677;
wire n29678;
wire n29679;
wire n29680;
wire n29681;
wire n29682;
wire n29683;
wire n29684;
wire n29685;
wire n29686;
wire n29687;
wire n29688;
wire n29689;
wire n29690;
wire n29691;
wire n29692;
wire n29693;
wire n29694;
wire n29695;
wire n29696;
wire n29697;
wire n29698;
wire n29699;
wire n29700;
wire n29701;
wire n29702;
wire n29703;
wire n29704;
wire n29705;
wire n29706;
wire n29707;
wire n29708;
wire n29709;
wire n2971;
wire n29710;
wire n29711;
wire n29712;
wire n29713;
wire n29714;
wire n29715;
wire n29716;
wire n29717;
wire n29718;
wire n29719;
wire n29720;
wire n29721;
wire n29722;
wire n29723;
wire n29724;
wire n29725;
wire n29727;
wire n29728;
wire n29730;
wire n29731;
wire n29732;
wire n29733;
wire n29734;
wire n29735;
wire n29736;
wire n29738;
wire n29739;
wire n29740;
wire n29741;
wire n29742;
wire n29743;
wire n29744;
wire n29745;
wire n29746;
wire n29747;
wire n29748;
wire n29749;
wire n29750;
wire n29751;
wire n29752;
wire n29753;
wire n29754;
wire n29755;
wire n29756;
wire n29757;
wire n29758;
wire n29759;
wire n2976;
wire n29760;
wire n29761;
wire n29762;
wire n29763;
wire n29764;
wire n29765;
wire n29766;
wire n29767;
wire n29768;
wire n29769;
wire n29770;
wire n29771;
wire n29772;
wire n29773;
wire n29774;
wire n29775;
wire n29776;
wire n29777;
wire n29778;
wire n29779;
wire n29780;
wire n29781;
wire n29782;
wire n29783;
wire n29784;
wire n29785;
wire n29786;
wire n29787;
wire n29788;
wire n29789;
wire n29790;
wire n29791;
wire n29792;
wire n29793;
wire n29794;
wire n29795;
wire n29796;
wire n29797;
wire n29798;
wire n29799;
wire n298;
wire n29800;
wire n29801;
wire n29802;
wire n29803;
wire n29804;
wire n29805;
wire n29806;
wire n29807;
wire n29808;
wire n29809;
wire n2981;
wire n29810;
wire n29811;
wire n29812;
wire n29813;
wire n29814;
wire n29815;
wire n29816;
wire n29817;
wire n29818;
wire n29819;
wire n29820;
wire n29821;
wire n29822;
wire n29823;
wire n29824;
wire n29825;
wire n29826;
wire n29827;
wire n29828;
wire n29829;
wire n29830;
wire n29831;
wire n29832;
wire n29833;
wire n29834;
wire n29836;
wire n29837;
wire n29838;
wire n29839;
wire n29841;
wire n29842;
wire n29843;
wire n29844;
wire n29845;
wire n29847;
wire n29849;
wire n29850;
wire n29851;
wire n29852;
wire n29853;
wire n29854;
wire n29855;
wire n29856;
wire n29857;
wire n29858;
wire n29859;
wire n2986;
wire n29860;
wire n29861;
wire n29862;
wire n29863;
wire n29864;
wire n29865;
wire n29866;
wire n29867;
wire n29868;
wire n29869;
wire n29870;
wire n29871;
wire n29872;
wire n29873;
wire n29874;
wire n29875;
wire n29876;
wire n29877;
wire n29878;
wire n29880;
wire n29881;
wire n29882;
wire n29883;
wire n29884;
wire n29886;
wire n29887;
wire n29888;
wire n29889;
wire n29890;
wire n29891;
wire n29892;
wire n29893;
wire n29894;
wire n29895;
wire n29896;
wire n29897;
wire n29898;
wire n29899;
wire n29900;
wire n29901;
wire n29902;
wire n29903;
wire n29904;
wire n29905;
wire n29906;
wire n29907;
wire n29908;
wire n29909;
wire n2991;
wire n29910;
wire n29911;
wire n29912;
wire n29913;
wire n29914;
wire n29915;
wire n29916;
wire n29917;
wire n29918;
wire n29919;
wire n29920;
wire n29921;
wire n29922;
wire n29923;
wire n29924;
wire n29925;
wire n29926;
wire n29927;
wire n29928;
wire n29929;
wire n29930;
wire n29931;
wire n29932;
wire n29933;
wire n29934;
wire n29935;
wire n29936;
wire n29937;
wire n29938;
wire n29939;
wire n29940;
wire n29941;
wire n29942;
wire n29943;
wire n29944;
wire n29945;
wire n29946;
wire n29947;
wire n29948;
wire n29949;
wire n29950;
wire n29951;
wire n29952;
wire n29953;
wire n29954;
wire n29955;
wire n29956;
wire n29957;
wire n29958;
wire n29959;
wire n2996;
wire n29960;
wire n29961;
wire n29962;
wire n29963;
wire n29964;
wire n29965;
wire n29966;
wire n29967;
wire n29968;
wire n29969;
wire n29970;
wire n29971;
wire n29972;
wire n29973;
wire n29974;
wire n29975;
wire n29976;
wire n29977;
wire n29978;
wire n29979;
wire n29980;
wire n29981;
wire n29982;
wire n29983;
wire n29984;
wire n29985;
wire n29986;
wire n29987;
wire n29988;
wire n29989;
wire n29990;
wire n29991;
wire n29992;
wire n29993;
wire n29994;
wire n29995;
wire n29996;
wire n29997;
wire n29998;
wire n29999;
wire n30000;
wire n30001;
wire n30002;
wire n30003;
wire n30004;
wire n30005;
wire n30006;
wire n30007;
wire n30008;
wire n30009;
wire n3001;
wire n30010;
wire n30011;
wire n30012;
wire n30013;
wire n30014;
wire n30015;
wire n30016;
wire n30017;
wire n30018;
wire n30019;
wire n30020;
wire n30021;
wire n30022;
wire n30023;
wire n30024;
wire n30025;
wire n30026;
wire n30027;
wire n30028;
wire n30029;
wire n30030;
wire n30031;
wire n30032;
wire n30033;
wire n30034;
wire n30035;
wire n30036;
wire n30037;
wire n30038;
wire n30039;
wire n30040;
wire n30041;
wire n30042;
wire n30043;
wire n30044;
wire n30045;
wire n30046;
wire n30047;
wire n30048;
wire n30049;
wire n3005;
wire n30050;
wire n30051;
wire n30052;
wire n30053;
wire n30054;
wire n30055;
wire n30056;
wire n30057;
wire n30058;
wire n30059;
wire n30060;
wire n30061;
wire n30062;
wire n30063;
wire n30064;
wire n30065;
wire n30066;
wire n30067;
wire n30068;
wire n30069;
wire n30070;
wire n30071;
wire n30072;
wire n30073;
wire n30074;
wire n30075;
wire n30076;
wire n30077;
wire n30078;
wire n30079;
wire n30080;
wire n30081;
wire n30082;
wire n30083;
wire n30084;
wire n30085;
wire n30086;
wire n30087;
wire n30088;
wire n30089;
wire n30090;
wire n30091;
wire n30092;
wire n30093;
wire n30094;
wire n30095;
wire n30096;
wire n30097;
wire n30098;
wire n30099;
wire n3010;
wire n30100;
wire n30101;
wire n30102;
wire n30103;
wire n30104;
wire n30105;
wire n30106;
wire n30107;
wire n30108;
wire n30109;
wire n30110;
wire n30111;
wire n30112;
wire n30113;
wire n30114;
wire n30115;
wire n30116;
wire n30117;
wire n30118;
wire n30119;
wire n30120;
wire n30121;
wire n30122;
wire n30123;
wire n30124;
wire n30125;
wire n30126;
wire n30127;
wire n30128;
wire n30129;
wire n30130;
wire n30131;
wire n30132;
wire n30133;
wire n30134;
wire n30135;
wire n30136;
wire n30138;
wire n30140;
wire n30141;
wire n30142;
wire n30143;
wire n30144;
wire n30146;
wire n30147;
wire n30148;
wire n30149;
wire n3015;
wire n30150;
wire n30151;
wire n30152;
wire n30153;
wire n30154;
wire n30155;
wire n30156;
wire n30157;
wire n30158;
wire n30159;
wire n30160;
wire n30161;
wire n30162;
wire n30163;
wire n30164;
wire n30165;
wire n30166;
wire n30167;
wire n30168;
wire n30169;
wire n30170;
wire n30171;
wire n30172;
wire n30173;
wire n30174;
wire n30175;
wire n30176;
wire n30177;
wire n30178;
wire n30179;
wire n30180;
wire n30181;
wire n30182;
wire n30183;
wire n30184;
wire n30185;
wire n30186;
wire n30187;
wire n30188;
wire n30189;
wire n30190;
wire n30191;
wire n30192;
wire n30193;
wire n30194;
wire n30195;
wire n30196;
wire n30197;
wire n30198;
wire n30199;
wire n3020;
wire n30200;
wire n30201;
wire n30202;
wire n30203;
wire n30204;
wire n30205;
wire n30206;
wire n30207;
wire n30208;
wire n30209;
wire n30210;
wire n30211;
wire n30212;
wire n30213;
wire n30214;
wire n30215;
wire n30216;
wire n30217;
wire n30218;
wire n30219;
wire n30220;
wire n30221;
wire n30222;
wire n30223;
wire n30224;
wire n30225;
wire n30226;
wire n30227;
wire n30228;
wire n30229;
wire n30230;
wire n30231;
wire n30232;
wire n30233;
wire n30234;
wire n30235;
wire n30236;
wire n30237;
wire n30238;
wire n30239;
wire n30240;
wire n30241;
wire n30242;
wire n30243;
wire n30244;
wire n30245;
wire n30246;
wire n30247;
wire n30248;
wire n30249;
wire n3025;
wire n30250;
wire n30251;
wire n30252;
wire n30253;
wire n30254;
wire n30255;
wire n30256;
wire n30257;
wire n30258;
wire n30259;
wire n30260;
wire n30261;
wire n30262;
wire n30263;
wire n30264;
wire n30265;
wire n30266;
wire n30267;
wire n30268;
wire n30269;
wire n30270;
wire n30271;
wire n30272;
wire n30273;
wire n30274;
wire n30275;
wire n30276;
wire n30277;
wire n30278;
wire n30279;
wire n30280;
wire n30281;
wire n30282;
wire n30283;
wire n30284;
wire n30285;
wire n30286;
wire n30287;
wire n30288;
wire n30289;
wire n30290;
wire n30291;
wire n30292;
wire n30293;
wire n30294;
wire n30295;
wire n30296;
wire n30297;
wire n30298;
wire n30299;
wire n303;
wire n3030;
wire n30300;
wire n30301;
wire n30302;
wire n30303;
wire n30304;
wire n30305;
wire n30306;
wire n30307;
wire n30308;
wire n30309;
wire n30310;
wire n30311;
wire n30312;
wire n30313;
wire n30314;
wire n30315;
wire n30316;
wire n30317;
wire n30318;
wire n30319;
wire n30320;
wire n30321;
wire n30322;
wire n30323;
wire n30324;
wire n30325;
wire n30326;
wire n30327;
wire n30328;
wire n30329;
wire n30330;
wire n30331;
wire n30332;
wire n30333;
wire n30334;
wire n30335;
wire n30336;
wire n30337;
wire n30338;
wire n30339;
wire n30340;
wire n30341;
wire n30342;
wire n30343;
wire n30344;
wire n30345;
wire n30346;
wire n30347;
wire n30348;
wire n30349;
wire n3035;
wire n30350;
wire n30351;
wire n30352;
wire n30353;
wire n30354;
wire n30355;
wire n30356;
wire n30357;
wire n30358;
wire n30359;
wire n30360;
wire n30361;
wire n30362;
wire n30363;
wire n30364;
wire n30365;
wire n30366;
wire n30367;
wire n30368;
wire n30369;
wire n30370;
wire n30371;
wire n30372;
wire n30373;
wire n30374;
wire n30375;
wire n30376;
wire n30377;
wire n30378;
wire n30379;
wire n30380;
wire n30381;
wire n30382;
wire n30383;
wire n30384;
wire n30385;
wire n30386;
wire n30387;
wire n30388;
wire n30389;
wire n30390;
wire n30391;
wire n30392;
wire n30393;
wire n30394;
wire n30395;
wire n30396;
wire n30397;
wire n30398;
wire n30399;
wire n3040;
wire n30400;
wire n30401;
wire n30402;
wire n30403;
wire n30404;
wire n30405;
wire n30406;
wire n30407;
wire n30408;
wire n30409;
wire n30410;
wire n30411;
wire n30412;
wire n30413;
wire n30414;
wire n30415;
wire n30416;
wire n30417;
wire n30418;
wire n30419;
wire n30420;
wire n30421;
wire n30422;
wire n30423;
wire n30424;
wire n30425;
wire n30426;
wire n30427;
wire n30428;
wire n30429;
wire n30430;
wire n30431;
wire n30432;
wire n30433;
wire n30434;
wire n30435;
wire n30436;
wire n30437;
wire n30438;
wire n30439;
wire n30440;
wire n30441;
wire n30442;
wire n30443;
wire n30444;
wire n30445;
wire n30446;
wire n30447;
wire n30448;
wire n30449;
wire n3045;
wire n30450;
wire n30451;
wire n30452;
wire n30453;
wire n30454;
wire n30455;
wire n30456;
wire n30457;
wire n30458;
wire n30459;
wire n30460;
wire n30461;
wire n30462;
wire n30463;
wire n30464;
wire n30465;
wire n30466;
wire n30467;
wire n30468;
wire n30469;
wire n30470;
wire n30471;
wire n30472;
wire n30473;
wire n30474;
wire n30475;
wire n30476;
wire n30477;
wire n30478;
wire n30479;
wire n30480;
wire n30481;
wire n30482;
wire n30483;
wire n30484;
wire n30485;
wire n30486;
wire n30487;
wire n30488;
wire n30489;
wire n30490;
wire n30491;
wire n30492;
wire n30493;
wire n30494;
wire n30495;
wire n30496;
wire n30497;
wire n30498;
wire n30499;
wire n3050;
wire n30500;
wire n30501;
wire n30502;
wire n30503;
wire n30504;
wire n30505;
wire n30506;
wire n30507;
wire n30508;
wire n30509;
wire n30510;
wire n30511;
wire n30512;
wire n30513;
wire n30514;
wire n30515;
wire n30516;
wire n30517;
wire n30518;
wire n30519;
wire n30520;
wire n30521;
wire n30522;
wire n30523;
wire n30524;
wire n30525;
wire n30526;
wire n30527;
wire n30528;
wire n30529;
wire n30530;
wire n30531;
wire n30532;
wire n30533;
wire n30534;
wire n30535;
wire n30536;
wire n30537;
wire n30538;
wire n30539;
wire n30540;
wire n30541;
wire n30542;
wire n30543;
wire n30544;
wire n30545;
wire n30546;
wire n30547;
wire n30548;
wire n30549;
wire n3055;
wire n30550;
wire n30551;
wire n30552;
wire n30553;
wire n30554;
wire n30555;
wire n30556;
wire n30557;
wire n30558;
wire n30559;
wire n30560;
wire n30561;
wire n30562;
wire n30563;
wire n30564;
wire n30565;
wire n30566;
wire n30567;
wire n30568;
wire n30569;
wire n30570;
wire n30571;
wire n30572;
wire n30573;
wire n30574;
wire n30575;
wire n30576;
wire n30577;
wire n30578;
wire n30579;
wire n30580;
wire n30581;
wire n30582;
wire n30583;
wire n30584;
wire n30585;
wire n30586;
wire n30587;
wire n30588;
wire n30589;
wire n30590;
wire n30591;
wire n30592;
wire n30593;
wire n30594;
wire n30595;
wire n30596;
wire n30597;
wire n30598;
wire n30599;
wire n3060;
wire n30600;
wire n30601;
wire n30602;
wire n30603;
wire n30604;
wire n30605;
wire n30606;
wire n30607;
wire n30608;
wire n30609;
wire n30610;
wire n30611;
wire n30612;
wire n30613;
wire n30614;
wire n30615;
wire n30616;
wire n30617;
wire n30618;
wire n30619;
wire n30620;
wire n30621;
wire n30622;
wire n30623;
wire n30624;
wire n30625;
wire n30626;
wire n30627;
wire n30628;
wire n30629;
wire n30630;
wire n30631;
wire n30632;
wire n30633;
wire n30634;
wire n30635;
wire n30636;
wire n30637;
wire n30638;
wire n30639;
wire n30640;
wire n30641;
wire n30642;
wire n30643;
wire n30644;
wire n30645;
wire n30646;
wire n30647;
wire n30648;
wire n30649;
wire n3065;
wire n30650;
wire n30651;
wire n30652;
wire n30653;
wire n30654;
wire n30655;
wire n30656;
wire n30657;
wire n30658;
wire n30659;
wire n30660;
wire n30661;
wire n30662;
wire n30663;
wire n30664;
wire n30665;
wire n30666;
wire n30667;
wire n30668;
wire n30669;
wire n30670;
wire n30671;
wire n30672;
wire n30673;
wire n30674;
wire n30675;
wire n30676;
wire n30677;
wire n30678;
wire n30679;
wire n30680;
wire n30681;
wire n30682;
wire n30683;
wire n30684;
wire n30685;
wire n30686;
wire n30687;
wire n30688;
wire n30689;
wire n30690;
wire n30691;
wire n30692;
wire n30693;
wire n30694;
wire n30695;
wire n30696;
wire n30697;
wire n30698;
wire n30699;
wire n3070;
wire n30700;
wire n30701;
wire n30702;
wire n30703;
wire n30704;
wire n30705;
wire n30706;
wire n30707;
wire n30708;
wire n30709;
wire n30710;
wire n30711;
wire n30712;
wire n30713;
wire n30714;
wire n30715;
wire n30716;
wire n30717;
wire n30718;
wire n30719;
wire n30720;
wire n30721;
wire n30722;
wire n30723;
wire n30724;
wire n30725;
wire n30726;
wire n30727;
wire n30728;
wire n30729;
wire n30730;
wire n30731;
wire n30732;
wire n30733;
wire n30734;
wire n30735;
wire n30736;
wire n30737;
wire n30738;
wire n30739;
wire n30740;
wire n30741;
wire n30742;
wire n30743;
wire n30744;
wire n30745;
wire n30746;
wire n30747;
wire n30748;
wire n30749;
wire n3075;
wire n30750;
wire n30751;
wire n30752;
wire n30753;
wire n30754;
wire n30755;
wire n30756;
wire n30757;
wire n30758;
wire n30759;
wire n30760;
wire n30761;
wire n30762;
wire n30763;
wire n30764;
wire n30765;
wire n30766;
wire n30767;
wire n30768;
wire n30769;
wire n30770;
wire n30771;
wire n30772;
wire n30773;
wire n30774;
wire n30775;
wire n30776;
wire n30777;
wire n30778;
wire n30779;
wire n30780;
wire n30781;
wire n30782;
wire n30783;
wire n30784;
wire n30785;
wire n30786;
wire n30787;
wire n30788;
wire n30789;
wire n30790;
wire n30791;
wire n30792;
wire n30793;
wire n30794;
wire n30795;
wire n30796;
wire n30797;
wire n30798;
wire n30799;
wire n308;
wire n3080;
wire n30800;
wire n30801;
wire n30802;
wire n30803;
wire n30804;
wire n30805;
wire n30806;
wire n30807;
wire n30808;
wire n30809;
wire n30810;
wire n30811;
wire n30812;
wire n30813;
wire n30814;
wire n30815;
wire n30816;
wire n30817;
wire n30818;
wire n30819;
wire n30820;
wire n30821;
wire n30822;
wire n30823;
wire n30824;
wire n30825;
wire n30826;
wire n30827;
wire n30828;
wire n30829;
wire n30830;
wire n30831;
wire n30832;
wire n30833;
wire n30834;
wire n30835;
wire n30836;
wire n30837;
wire n30838;
wire n30839;
wire n30840;
wire n30841;
wire n30842;
wire n30843;
wire n30844;
wire n30845;
wire n30846;
wire n30847;
wire n30848;
wire n30849;
wire n3085;
wire n30850;
wire n30851;
wire n30852;
wire n30853;
wire n30854;
wire n30855;
wire n30856;
wire n30857;
wire n30858;
wire n30859;
wire n30860;
wire n30861;
wire n30862;
wire n30863;
wire n30864;
wire n30865;
wire n30866;
wire n30867;
wire n30868;
wire n30869;
wire n30870;
wire n30871;
wire n30872;
wire n30873;
wire n30874;
wire n30875;
wire n30876;
wire n30877;
wire n30878;
wire n30879;
wire n30880;
wire n30881;
wire n30882;
wire n30883;
wire n30884;
wire n30885;
wire n30886;
wire n30887;
wire n30888;
wire n30889;
wire n30890;
wire n30891;
wire n30892;
wire n30893;
wire n30894;
wire n30895;
wire n30896;
wire n30897;
wire n30898;
wire n30899;
wire n3090;
wire n30900;
wire n30901;
wire n30902;
wire n30903;
wire n30904;
wire n30905;
wire n30906;
wire n30907;
wire n30908;
wire n30909;
wire n30910;
wire n30911;
wire n30912;
wire n30913;
wire n30914;
wire n30915;
wire n30916;
wire n30917;
wire n30918;
wire n30919;
wire n30920;
wire n30921;
wire n30922;
wire n30923;
wire n30924;
wire n30925;
wire n30926;
wire n30927;
wire n30928;
wire n30929;
wire n30930;
wire n30931;
wire n30932;
wire n30933;
wire n30934;
wire n30935;
wire n30936;
wire n30937;
wire n30938;
wire n30939;
wire n30940;
wire n30941;
wire n30942;
wire n30943;
wire n30944;
wire n30945;
wire n30946;
wire n30947;
wire n30948;
wire n30949;
wire n3095;
wire n30950;
wire n30951;
wire n30952;
wire n30953;
wire n30954;
wire n30955;
wire n30956;
wire n30957;
wire n30958;
wire n30959;
wire n30960;
wire n30961;
wire n30962;
wire n30963;
wire n30964;
wire n30965;
wire n30966;
wire n30967;
wire n30968;
wire n30969;
wire n30970;
wire n30971;
wire n30972;
wire n30973;
wire n30974;
wire n30975;
wire n30976;
wire n30977;
wire n30978;
wire n30979;
wire n30980;
wire n30981;
wire n30982;
wire n30983;
wire n30984;
wire n30985;
wire n30986;
wire n30987;
wire n30988;
wire n30989;
wire n30990;
wire n30991;
wire n30992;
wire n30993;
wire n30994;
wire n30995;
wire n30996;
wire n30997;
wire n30998;
wire n30999;
wire n3100;
wire n31000;
wire n31001;
wire n31002;
wire n31003;
wire n31004;
wire n31005;
wire n31006;
wire n31007;
wire n31008;
wire n31009;
wire n31010;
wire n31011;
wire n31012;
wire n31013;
wire n31014;
wire n31015;
wire n31016;
wire n31017;
wire n31018;
wire n31019;
wire n31020;
wire n31021;
wire n31022;
wire n31023;
wire n31024;
wire n31025;
wire n31026;
wire n31027;
wire n31028;
wire n31029;
wire n31030;
wire n31031;
wire n31032;
wire n31033;
wire n31034;
wire n31035;
wire n31036;
wire n31037;
wire n31038;
wire n31039;
wire n31040;
wire n31041;
wire n31042;
wire n31043;
wire n31044;
wire n31045;
wire n31046;
wire n31047;
wire n31048;
wire n31049;
wire n3105;
wire n31050;
wire n31051;
wire n31052;
wire n31053;
wire n31054;
wire n31055;
wire n31056;
wire n31057;
wire n31058;
wire n31059;
wire n31060;
wire n31061;
wire n31062;
wire n31063;
wire n31064;
wire n31065;
wire n31066;
wire n31067;
wire n31068;
wire n31069;
wire n31070;
wire n31071;
wire n31072;
wire n31073;
wire n31074;
wire n31075;
wire n31076;
wire n31077;
wire n31078;
wire n31079;
wire n31080;
wire n31081;
wire n31082;
wire n31083;
wire n31084;
wire n31085;
wire n31086;
wire n31087;
wire n31088;
wire n31089;
wire n31090;
wire n31091;
wire n31092;
wire n31093;
wire n31094;
wire n31095;
wire n31096;
wire n31097;
wire n31098;
wire n31099;
wire n3110;
wire n31100;
wire n31101;
wire n31102;
wire n31103;
wire n31104;
wire n31105;
wire n31106;
wire n31107;
wire n31108;
wire n31109;
wire n31110;
wire n31111;
wire n31112;
wire n31113;
wire n31114;
wire n31115;
wire n31116;
wire n31117;
wire n31118;
wire n31119;
wire n31120;
wire n31121;
wire n31122;
wire n31123;
wire n31124;
wire n31125;
wire n31126;
wire n31127;
wire n31128;
wire n31129;
wire n31130;
wire n31131;
wire n31132;
wire n31133;
wire n31134;
wire n31135;
wire n31136;
wire n31137;
wire n31138;
wire n31139;
wire n31140;
wire n31141;
wire n31142;
wire n31143;
wire n31144;
wire n31145;
wire n31146;
wire n31147;
wire n31148;
wire n31149;
wire n3115;
wire n31150;
wire n31151;
wire n31152;
wire n31153;
wire n31154;
wire n31155;
wire n31156;
wire n31157;
wire n31158;
wire n31159;
wire n31160;
wire n31161;
wire n31162;
wire n31163;
wire n31164;
wire n31165;
wire n31166;
wire n31167;
wire n31168;
wire n31169;
wire n31170;
wire n31171;
wire n31172;
wire n31173;
wire n31174;
wire n31175;
wire n31176;
wire n31177;
wire n31178;
wire n31179;
wire n31180;
wire n31181;
wire n31182;
wire n31183;
wire n31184;
wire n31185;
wire n31186;
wire n31187;
wire n31188;
wire n31189;
wire n31190;
wire n31191;
wire n31192;
wire n31193;
wire n31194;
wire n31195;
wire n31196;
wire n31197;
wire n31198;
wire n31199;
wire n3120;
wire n31200;
wire n31201;
wire n31202;
wire n31203;
wire n31204;
wire n31205;
wire n31206;
wire n31207;
wire n31208;
wire n31209;
wire n31210;
wire n31211;
wire n31212;
wire n31213;
wire n31214;
wire n31215;
wire n31216;
wire n31217;
wire n31218;
wire n31219;
wire n31220;
wire n31221;
wire n31222;
wire n31223;
wire n31224;
wire n31225;
wire n31226;
wire n31227;
wire n31228;
wire n31229;
wire n31230;
wire n31231;
wire n31232;
wire n31233;
wire n31234;
wire n31235;
wire n31236;
wire n31237;
wire n31238;
wire n31239;
wire n31240;
wire n31241;
wire n31242;
wire n31243;
wire n31244;
wire n31245;
wire n31246;
wire n31247;
wire n31248;
wire n31249;
wire n3125;
wire n31250;
wire n31251;
wire n31252;
wire n31253;
wire n31254;
wire n31255;
wire n31256;
wire n31257;
wire n31258;
wire n31259;
wire n31260;
wire n31261;
wire n31262;
wire n31263;
wire n31264;
wire n31265;
wire n31266;
wire n31267;
wire n31268;
wire n31269;
wire n31270;
wire n31271;
wire n31272;
wire n31273;
wire n31274;
wire n31275;
wire n31276;
wire n31277;
wire n31278;
wire n31279;
wire n31280;
wire n31281;
wire n31282;
wire n31283;
wire n31284;
wire n31285;
wire n31286;
wire n31287;
wire n31288;
wire n31289;
wire n31290;
wire n31291;
wire n31292;
wire n31293;
wire n31294;
wire n31295;
wire n31296;
wire n31297;
wire n31298;
wire n31299;
wire n313;
wire n3130;
wire n31300;
wire n31301;
wire n31302;
wire n31303;
wire n31304;
wire n31305;
wire n31306;
wire n31307;
wire n31308;
wire n31309;
wire n31310;
wire n31311;
wire n31312;
wire n31313;
wire n31314;
wire n31315;
wire n31316;
wire n31317;
wire n31318;
wire n31319;
wire n31320;
wire n31321;
wire n31322;
wire n31323;
wire n31324;
wire n31325;
wire n31326;
wire n31327;
wire n31328;
wire n31329;
wire n31330;
wire n31331;
wire n31332;
wire n31333;
wire n31334;
wire n31335;
wire n31336;
wire n31337;
wire n31338;
wire n31339;
wire n31340;
wire n31341;
wire n31342;
wire n31343;
wire n31344;
wire n31345;
wire n31346;
wire n31347;
wire n31348;
wire n31349;
wire n3135;
wire n31350;
wire n31351;
wire n31352;
wire n31353;
wire n31354;
wire n31355;
wire n31356;
wire n31357;
wire n31358;
wire n31359;
wire n31360;
wire n31361;
wire n31362;
wire n31363;
wire n31364;
wire n31365;
wire n31366;
wire n31367;
wire n31368;
wire n31369;
wire n31370;
wire n31371;
wire n31372;
wire n31373;
wire n31374;
wire n31375;
wire n31376;
wire n31377;
wire n31378;
wire n31379;
wire n31380;
wire n31381;
wire n31382;
wire n31383;
wire n31384;
wire n31385;
wire n31386;
wire n31387;
wire n31388;
wire n31389;
wire n31390;
wire n31391;
wire n31392;
wire n31393;
wire n31394;
wire n31395;
wire n31396;
wire n31397;
wire n31398;
wire n31399;
wire n3140;
wire n31400;
wire n31401;
wire n31402;
wire n31403;
wire n31404;
wire n31405;
wire n31406;
wire n31407;
wire n31408;
wire n31409;
wire n31410;
wire n31411;
wire n31412;
wire n31413;
wire n31414;
wire n31415;
wire n31416;
wire n31417;
wire n31418;
wire n31419;
wire n31420;
wire n31421;
wire n31422;
wire n31423;
wire n31424;
wire n31425;
wire n31426;
wire n31427;
wire n31428;
wire n31429;
wire n31430;
wire n31431;
wire n31432;
wire n31433;
wire n31434;
wire n31435;
wire n31436;
wire n31437;
wire n31438;
wire n31439;
wire n31440;
wire n31441;
wire n31442;
wire n31443;
wire n31444;
wire n31445;
wire n31446;
wire n31447;
wire n31448;
wire n31449;
wire n3145;
wire n31450;
wire n31451;
wire n31452;
wire n31453;
wire n31454;
wire n31455;
wire n31456;
wire n31457;
wire n31458;
wire n31459;
wire n31460;
wire n31461;
wire n31462;
wire n31463;
wire n31464;
wire n31465;
wire n31466;
wire n31467;
wire n31468;
wire n31469;
wire n31470;
wire n31471;
wire n31472;
wire n31473;
wire n31474;
wire n31475;
wire n31476;
wire n31477;
wire n31478;
wire n31479;
wire n31480;
wire n31481;
wire n31482;
wire n31483;
wire n31484;
wire n31485;
wire n31486;
wire n31487;
wire n31488;
wire n31489;
wire n31490;
wire n31491;
wire n31492;
wire n31493;
wire n31494;
wire n31495;
wire n31496;
wire n31497;
wire n31498;
wire n31499;
wire n3150;
wire n31500;
wire n31501;
wire n31502;
wire n31503;
wire n31504;
wire n31505;
wire n31506;
wire n31507;
wire n31508;
wire n31509;
wire n31510;
wire n31511;
wire n31512;
wire n31513;
wire n31514;
wire n31515;
wire n31516;
wire n31517;
wire n31518;
wire n31519;
wire n31520;
wire n31521;
wire n31522;
wire n31523;
wire n31524;
wire n31525;
wire n31526;
wire n31527;
wire n31528;
wire n31529;
wire n31530;
wire n31531;
wire n31532;
wire n31533;
wire n31534;
wire n31535;
wire n31536;
wire n31537;
wire n31538;
wire n31539;
wire n31540;
wire n31541;
wire n31542;
wire n31543;
wire n31544;
wire n31545;
wire n31546;
wire n31547;
wire n31548;
wire n31549;
wire n3155;
wire n31550;
wire n31551;
wire n31552;
wire n31553;
wire n31554;
wire n31555;
wire n31556;
wire n31557;
wire n31558;
wire n31559;
wire n31560;
wire n31561;
wire n31562;
wire n31563;
wire n31564;
wire n31565;
wire n31566;
wire n31567;
wire n31568;
wire n31569;
wire n31570;
wire n31571;
wire n31572;
wire n31573;
wire n31574;
wire n31575;
wire n31576;
wire n31577;
wire n31578;
wire n31579;
wire n31580;
wire n31581;
wire n31582;
wire n31583;
wire n31584;
wire n31585;
wire n31586;
wire n31587;
wire n31588;
wire n31589;
wire n31590;
wire n31591;
wire n31592;
wire n31593;
wire n31594;
wire n31595;
wire n31596;
wire n31597;
wire n31598;
wire n31599;
wire n3160;
wire n31600;
wire n31601;
wire n31602;
wire n31603;
wire n31604;
wire n31605;
wire n31606;
wire n31607;
wire n31608;
wire n31609;
wire n31610;
wire n31611;
wire n31612;
wire n31613;
wire n31614;
wire n31615;
wire n31616;
wire n31617;
wire n31618;
wire n31619;
wire n31620;
wire n31621;
wire n31622;
wire n31623;
wire n31624;
wire n31625;
wire n31626;
wire n31627;
wire n31628;
wire n31629;
wire n31630;
wire n31631;
wire n31632;
wire n31633;
wire n31634;
wire n31635;
wire n31636;
wire n31637;
wire n31638;
wire n31639;
wire n31640;
wire n31641;
wire n31642;
wire n31643;
wire n31644;
wire n31645;
wire n31646;
wire n31647;
wire n31648;
wire n31649;
wire n3165;
wire n31650;
wire n31651;
wire n31652;
wire n31653;
wire n31654;
wire n31655;
wire n31656;
wire n31657;
wire n31658;
wire n31659;
wire n31660;
wire n31661;
wire n31662;
wire n31663;
wire n31664;
wire n31665;
wire n31666;
wire n31667;
wire n31668;
wire n31669;
wire n31670;
wire n31671;
wire n31672;
wire n31673;
wire n31674;
wire n31675;
wire n31676;
wire n31677;
wire n31678;
wire n31679;
wire n31680;
wire n31681;
wire n31682;
wire n31683;
wire n31684;
wire n31685;
wire n31686;
wire n31687;
wire n31688;
wire n31689;
wire n31690;
wire n31691;
wire n31692;
wire n31693;
wire n31694;
wire n31695;
wire n31696;
wire n31697;
wire n31698;
wire n31699;
wire n3170;
wire n31700;
wire n31701;
wire n31702;
wire n31703;
wire n31704;
wire n31705;
wire n31706;
wire n31707;
wire n31708;
wire n31709;
wire n31710;
wire n31711;
wire n31712;
wire n31713;
wire n31714;
wire n31715;
wire n31716;
wire n31717;
wire n31718;
wire n31719;
wire n31720;
wire n31721;
wire n31722;
wire n31723;
wire n31724;
wire n31725;
wire n31726;
wire n31727;
wire n31728;
wire n31729;
wire n31730;
wire n31731;
wire n31732;
wire n31733;
wire n31734;
wire n31735;
wire n31736;
wire n31737;
wire n31738;
wire n31739;
wire n31740;
wire n31741;
wire n31742;
wire n31743;
wire n31744;
wire n31745;
wire n31746;
wire n31747;
wire n31748;
wire n31749;
wire n3175;
wire n31750;
wire n31751;
wire n31752;
wire n31753;
wire n31754;
wire n31755;
wire n31756;
wire n31757;
wire n31758;
wire n31759;
wire n31760;
wire n31761;
wire n31762;
wire n31763;
wire n31764;
wire n31765;
wire n31766;
wire n31767;
wire n31768;
wire n31769;
wire n31770;
wire n31771;
wire n31772;
wire n31773;
wire n31774;
wire n31775;
wire n31776;
wire n31777;
wire n31778;
wire n31779;
wire n31780;
wire n31781;
wire n31782;
wire n31783;
wire n31784;
wire n31785;
wire n31786;
wire n31787;
wire n31788;
wire n31789;
wire n31790;
wire n31791;
wire n31792;
wire n31793;
wire n31794;
wire n31795;
wire n31796;
wire n31797;
wire n31798;
wire n31799;
wire n318;
wire n3180;
wire n31800;
wire n31801;
wire n31802;
wire n31803;
wire n31804;
wire n31805;
wire n31806;
wire n31807;
wire n31808;
wire n31809;
wire n31810;
wire n31811;
wire n31812;
wire n31813;
wire n31814;
wire n31815;
wire n31816;
wire n31817;
wire n31818;
wire n31819;
wire n31820;
wire n31821;
wire n31822;
wire n31823;
wire n31824;
wire n31825;
wire n31826;
wire n31827;
wire n31828;
wire n31829;
wire n31830;
wire n31831;
wire n31832;
wire n31833;
wire n31834;
wire n31835;
wire n31836;
wire n31837;
wire n31838;
wire n31839;
wire n31840;
wire n31841;
wire n31842;
wire n31843;
wire n31844;
wire n31845;
wire n31846;
wire n31847;
wire n31848;
wire n31849;
wire n3185;
wire n31850;
wire n31851;
wire n31852;
wire n31853;
wire n31854;
wire n31855;
wire n31856;
wire n31857;
wire n31858;
wire n31859;
wire n31860;
wire n31861;
wire n31862;
wire n31863;
wire n31864;
wire n31865;
wire n31866;
wire n31867;
wire n31868;
wire n31869;
wire n31870;
wire n31871;
wire n31872;
wire n31873;
wire n31874;
wire n31875;
wire n31876;
wire n31877;
wire n31878;
wire n31879;
wire n31880;
wire n31881;
wire n31882;
wire n31883;
wire n31884;
wire n31885;
wire n31886;
wire n31887;
wire n31888;
wire n31889;
wire n31890;
wire n31891;
wire n31892;
wire n31893;
wire n31894;
wire n31895;
wire n31896;
wire n31897;
wire n31898;
wire n31899;
wire n3190;
wire n31900;
wire n31901;
wire n31902;
wire n31903;
wire n31904;
wire n31905;
wire n31906;
wire n31907;
wire n31908;
wire n31909;
wire n31910;
wire n31911;
wire n31912;
wire n31913;
wire n31914;
wire n31915;
wire n31916;
wire n31917;
wire n31918;
wire n31919;
wire n31920;
wire n31921;
wire n31922;
wire n31923;
wire n31924;
wire n31925;
wire n31926;
wire n31927;
wire n31928;
wire n31929;
wire n31930;
wire n31931;
wire n31932;
wire n31933;
wire n31934;
wire n31935;
wire n31936;
wire n31937;
wire n31938;
wire n31939;
wire n3194;
wire n31940;
wire n31941;
wire n31942;
wire n31943;
wire n31944;
wire n31945;
wire n31946;
wire n31947;
wire n31948;
wire n31949;
wire n31950;
wire n31951;
wire n31952;
wire n31953;
wire n31954;
wire n31955;
wire n31956;
wire n31957;
wire n31958;
wire n31959;
wire n31960;
wire n31961;
wire n31962;
wire n31963;
wire n31964;
wire n31965;
wire n31966;
wire n31967;
wire n31968;
wire n31969;
wire n31970;
wire n31971;
wire n31972;
wire n31973;
wire n31974;
wire n31975;
wire n31976;
wire n31977;
wire n31978;
wire n31979;
wire n31980;
wire n31981;
wire n31982;
wire n31983;
wire n31984;
wire n31985;
wire n31986;
wire n31987;
wire n31988;
wire n31989;
wire n3199;
wire n31990;
wire n31991;
wire n31992;
wire n31993;
wire n31994;
wire n31995;
wire n31996;
wire n31997;
wire n31998;
wire n31999;
wire n32000;
wire n32001;
wire n32002;
wire n32003;
wire n32004;
wire n32005;
wire n32006;
wire n32007;
wire n32008;
wire n32009;
wire n32010;
wire n32011;
wire n32012;
wire n32013;
wire n32014;
wire n32015;
wire n32016;
wire n32017;
wire n32018;
wire n32019;
wire n32020;
wire n32021;
wire n32022;
wire n32023;
wire n32024;
wire n32025;
wire n32026;
wire n32027;
wire n32028;
wire n32029;
wire n32030;
wire n32031;
wire n32032;
wire n32033;
wire n32034;
wire n32035;
wire n32036;
wire n32037;
wire n32038;
wire n32039;
wire n3204;
wire n32040;
wire n32041;
wire n32042;
wire n32043;
wire n32044;
wire n32045;
wire n32046;
wire n32047;
wire n32048;
wire n32049;
wire n32050;
wire n32051;
wire n32052;
wire n32053;
wire n32054;
wire n32055;
wire n32056;
wire n32057;
wire n32058;
wire n32059;
wire n32060;
wire n32061;
wire n32062;
wire n32063;
wire n32064;
wire n32065;
wire n32066;
wire n32067;
wire n32068;
wire n32069;
wire n32070;
wire n32071;
wire n32072;
wire n32073;
wire n32074;
wire n32075;
wire n32076;
wire n32077;
wire n32078;
wire n32079;
wire n32080;
wire n32081;
wire n32082;
wire n32083;
wire n32084;
wire n32085;
wire n32086;
wire n32087;
wire n32088;
wire n32089;
wire n3209;
wire n32090;
wire n32091;
wire n32092;
wire n32093;
wire n32094;
wire n32095;
wire n32096;
wire n32097;
wire n32098;
wire n32099;
wire n32100;
wire n32101;
wire n32102;
wire n32103;
wire n32104;
wire n32105;
wire n32106;
wire n32107;
wire n32108;
wire n32109;
wire n32110;
wire n32111;
wire n32112;
wire n32113;
wire n32114;
wire n32115;
wire n32116;
wire n32117;
wire n32118;
wire n32119;
wire n32120;
wire n32121;
wire n32122;
wire n32123;
wire n32124;
wire n32125;
wire n32126;
wire n32127;
wire n32128;
wire n32129;
wire n32130;
wire n32131;
wire n32132;
wire n32133;
wire n32134;
wire n32135;
wire n32136;
wire n32137;
wire n32138;
wire n32139;
wire n3214;
wire n32140;
wire n32141;
wire n32142;
wire n32143;
wire n32144;
wire n32145;
wire n32146;
wire n32147;
wire n32148;
wire n32149;
wire n32150;
wire n32151;
wire n32152;
wire n32153;
wire n32154;
wire n32155;
wire n32156;
wire n32157;
wire n32158;
wire n32159;
wire n32160;
wire n32161;
wire n32162;
wire n32163;
wire n32164;
wire n32165;
wire n32166;
wire n32167;
wire n32168;
wire n32169;
wire n32170;
wire n32171;
wire n32172;
wire n32173;
wire n32174;
wire n32175;
wire n32176;
wire n32177;
wire n32178;
wire n32179;
wire n32180;
wire n32181;
wire n32182;
wire n32183;
wire n32184;
wire n32185;
wire n32186;
wire n32187;
wire n32188;
wire n32189;
wire n3219;
wire n32190;
wire n32191;
wire n32192;
wire n32193;
wire n32194;
wire n32195;
wire n32196;
wire n32197;
wire n32198;
wire n32199;
wire n32200;
wire n32201;
wire n32202;
wire n32203;
wire n32204;
wire n32205;
wire n32206;
wire n32207;
wire n32208;
wire n32209;
wire n32210;
wire n32211;
wire n32212;
wire n32213;
wire n32214;
wire n32215;
wire n32216;
wire n32217;
wire n32218;
wire n32219;
wire n32220;
wire n32221;
wire n32222;
wire n32223;
wire n32224;
wire n32225;
wire n32226;
wire n32227;
wire n32228;
wire n32229;
wire n32230;
wire n32231;
wire n32232;
wire n32233;
wire n32234;
wire n32235;
wire n32236;
wire n32237;
wire n32238;
wire n32239;
wire n3224;
wire n32240;
wire n32241;
wire n32242;
wire n32243;
wire n32244;
wire n32245;
wire n32246;
wire n32247;
wire n32248;
wire n32249;
wire n32250;
wire n32251;
wire n32252;
wire n32253;
wire n32254;
wire n32255;
wire n32256;
wire n32257;
wire n32258;
wire n32259;
wire n32260;
wire n32261;
wire n32262;
wire n32263;
wire n32264;
wire n32265;
wire n32266;
wire n32267;
wire n32268;
wire n32269;
wire n32270;
wire n32271;
wire n32272;
wire n32273;
wire n32274;
wire n32275;
wire n32276;
wire n32277;
wire n32278;
wire n32279;
wire n3228;
wire n32280;
wire n32281;
wire n32282;
wire n32283;
wire n32284;
wire n32285;
wire n32286;
wire n32287;
wire n32288;
wire n32289;
wire n32290;
wire n32291;
wire n32292;
wire n32293;
wire n32294;
wire n32295;
wire n32296;
wire n32297;
wire n32298;
wire n32299;
wire n323;
wire n32300;
wire n32301;
wire n32302;
wire n32303;
wire n32304;
wire n32305;
wire n32306;
wire n32307;
wire n32308;
wire n32309;
wire n32310;
wire n32311;
wire n32312;
wire n32313;
wire n32314;
wire n32315;
wire n32316;
wire n32317;
wire n32318;
wire n32319;
wire n32320;
wire n32321;
wire n32322;
wire n32323;
wire n32324;
wire n32325;
wire n32326;
wire n32327;
wire n32328;
wire n32329;
wire n3233;
wire n32330;
wire n32331;
wire n32332;
wire n32333;
wire n32334;
wire n32335;
wire n32336;
wire n32337;
wire n32338;
wire n32339;
wire n32340;
wire n32341;
wire n32342;
wire n32343;
wire n32344;
wire n32345;
wire n32346;
wire n32347;
wire n32348;
wire n32349;
wire n32350;
wire n32351;
wire n32352;
wire n32353;
wire n32354;
wire n32355;
wire n32356;
wire n32357;
wire n32358;
wire n32359;
wire n32360;
wire n32361;
wire n32362;
wire n32363;
wire n32364;
wire n32365;
wire n32366;
wire n32367;
wire n32368;
wire n32369;
wire n32370;
wire n32371;
wire n32372;
wire n32373;
wire n32374;
wire n32375;
wire n32376;
wire n32377;
wire n32378;
wire n32379;
wire n3238;
wire n32380;
wire n32381;
wire n32382;
wire n32383;
wire n32384;
wire n32385;
wire n32386;
wire n32387;
wire n32388;
wire n32389;
wire n32390;
wire n32391;
wire n32392;
wire n32393;
wire n32394;
wire n32395;
wire n32396;
wire n32397;
wire n32398;
wire n32399;
wire n32400;
wire n32401;
wire n32402;
wire n32403;
wire n32404;
wire n32405;
wire n32406;
wire n32407;
wire n32408;
wire n32409;
wire n32410;
wire n32411;
wire n32412;
wire n32413;
wire n32414;
wire n32415;
wire n32416;
wire n32417;
wire n32418;
wire n32419;
wire n32420;
wire n32421;
wire n32422;
wire n32423;
wire n32424;
wire n32425;
wire n32426;
wire n32427;
wire n32428;
wire n32429;
wire n3243;
wire n32430;
wire n32431;
wire n32432;
wire n32433;
wire n32434;
wire n32435;
wire n32436;
wire n32437;
wire n32438;
wire n32439;
wire n32440;
wire n32441;
wire n32442;
wire n32443;
wire n32444;
wire n32445;
wire n32446;
wire n32447;
wire n32448;
wire n32449;
wire n32450;
wire n32451;
wire n32452;
wire n32453;
wire n32454;
wire n32455;
wire n32456;
wire n32457;
wire n32458;
wire n32459;
wire n32460;
wire n32461;
wire n32462;
wire n32463;
wire n32464;
wire n32465;
wire n32466;
wire n32467;
wire n32468;
wire n32469;
wire n32470;
wire n32471;
wire n32472;
wire n32473;
wire n32474;
wire n32475;
wire n32476;
wire n32477;
wire n32478;
wire n32479;
wire n3248;
wire n32480;
wire n32481;
wire n32482;
wire n32483;
wire n32484;
wire n32485;
wire n32486;
wire n32487;
wire n32488;
wire n32489;
wire n32490;
wire n32491;
wire n32492;
wire n32493;
wire n32494;
wire n32495;
wire n32496;
wire n32497;
wire n32499;
wire n32500;
wire n32501;
wire n32502;
wire n32503;
wire n32504;
wire n32505;
wire n32506;
wire n32507;
wire n32509;
wire n32510;
wire n32511;
wire n32512;
wire n32513;
wire n32514;
wire n32515;
wire n32516;
wire n32517;
wire n32518;
wire n32519;
wire n3252;
wire n32520;
wire n32521;
wire n32522;
wire n32523;
wire n32524;
wire n32525;
wire n32526;
wire n32527;
wire n32528;
wire n32529;
wire n32530;
wire n32531;
wire n32532;
wire n32533;
wire n32534;
wire n32535;
wire n32536;
wire n32537;
wire n32538;
wire n32539;
wire n32540;
wire n32541;
wire n32542;
wire n32543;
wire n32544;
wire n32545;
wire n32546;
wire n32547;
wire n32548;
wire n32549;
wire n32550;
wire n32551;
wire n32552;
wire n32553;
wire n32554;
wire n32555;
wire n32556;
wire n32557;
wire n32558;
wire n32559;
wire n32560;
wire n32561;
wire n32562;
wire n32563;
wire n32564;
wire n32565;
wire n32566;
wire n32567;
wire n32568;
wire n32569;
wire n3257;
wire n32570;
wire n32571;
wire n32572;
wire n32573;
wire n32574;
wire n32575;
wire n32576;
wire n32577;
wire n32578;
wire n32579;
wire n32580;
wire n32581;
wire n32582;
wire n32583;
wire n32584;
wire n32585;
wire n32586;
wire n32587;
wire n32588;
wire n32589;
wire n32590;
wire n32591;
wire n32592;
wire n32593;
wire n32594;
wire n32595;
wire n32596;
wire n32597;
wire n32598;
wire n32599;
wire n32600;
wire n32601;
wire n32602;
wire n32603;
wire n32604;
wire n32605;
wire n32606;
wire n32607;
wire n32608;
wire n32609;
wire n32610;
wire n32611;
wire n32612;
wire n32613;
wire n32614;
wire n32615;
wire n32616;
wire n32617;
wire n32618;
wire n32619;
wire n3262;
wire n32620;
wire n32621;
wire n32622;
wire n32623;
wire n32624;
wire n32625;
wire n32626;
wire n32627;
wire n32628;
wire n32629;
wire n32630;
wire n32631;
wire n32632;
wire n32633;
wire n32634;
wire n32635;
wire n32636;
wire n32637;
wire n32638;
wire n32639;
wire n32640;
wire n32641;
wire n32642;
wire n32643;
wire n32644;
wire n32645;
wire n32646;
wire n32647;
wire n32648;
wire n32649;
wire n32650;
wire n32651;
wire n32652;
wire n32653;
wire n32654;
wire n32655;
wire n32656;
wire n32657;
wire n32658;
wire n32659;
wire n32660;
wire n32661;
wire n32662;
wire n32663;
wire n32664;
wire n32665;
wire n32666;
wire n32667;
wire n32668;
wire n32669;
wire n3267;
wire n32670;
wire n32671;
wire n32672;
wire n32673;
wire n32674;
wire n32675;
wire n32676;
wire n32677;
wire n32678;
wire n32679;
wire n32680;
wire n32681;
wire n32682;
wire n32683;
wire n32684;
wire n32685;
wire n32686;
wire n32687;
wire n32688;
wire n32689;
wire n32690;
wire n32691;
wire n32692;
wire n32693;
wire n32694;
wire n32695;
wire n32696;
wire n32697;
wire n32698;
wire n32699;
wire n32700;
wire n32701;
wire n32702;
wire n32703;
wire n32704;
wire n32705;
wire n32706;
wire n32707;
wire n32708;
wire n32709;
wire n32710;
wire n32711;
wire n32712;
wire n32713;
wire n32714;
wire n32715;
wire n32716;
wire n32717;
wire n32718;
wire n32719;
wire n3272;
wire n32720;
wire n32721;
wire n32722;
wire n32723;
wire n32724;
wire n32725;
wire n32726;
wire n32727;
wire n32728;
wire n32729;
wire n32730;
wire n32732;
wire n32733;
wire n32734;
wire n32735;
wire n32736;
wire n32737;
wire n32738;
wire n32739;
wire n32740;
wire n32741;
wire n32742;
wire n32743;
wire n32744;
wire n32745;
wire n32746;
wire n32747;
wire n32748;
wire n32749;
wire n32750;
wire n32751;
wire n32752;
wire n32753;
wire n32754;
wire n32755;
wire n32756;
wire n32757;
wire n32758;
wire n32759;
wire n32760;
wire n32761;
wire n32762;
wire n32763;
wire n32764;
wire n32765;
wire n32766;
wire n32767;
wire n32768;
wire n32769;
wire n3277;
wire n32770;
wire n32771;
wire n32772;
wire n32773;
wire n32774;
wire n32775;
wire n32776;
wire n32777;
wire n32778;
wire n32779;
wire n32780;
wire n32781;
wire n32782;
wire n32783;
wire n32784;
wire n32785;
wire n32786;
wire n32787;
wire n32788;
wire n32789;
wire n32790;
wire n32791;
wire n32792;
wire n32793;
wire n32794;
wire n32795;
wire n32796;
wire n32797;
wire n32798;
wire n32799;
wire n328;
wire n32800;
wire n32801;
wire n32802;
wire n32803;
wire n32804;
wire n32805;
wire n32806;
wire n32807;
wire n32808;
wire n32809;
wire n32810;
wire n32811;
wire n32812;
wire n32813;
wire n32814;
wire n32815;
wire n32816;
wire n32817;
wire n32818;
wire n32819;
wire n3282;
wire n32820;
wire n32821;
wire n32822;
wire n32823;
wire n32824;
wire n32825;
wire n32826;
wire n32827;
wire n32828;
wire n32829;
wire n32830;
wire n32831;
wire n32832;
wire n32833;
wire n32834;
wire n32835;
wire n32836;
wire n32837;
wire n32838;
wire n32839;
wire n32840;
wire n32841;
wire n32842;
wire n32843;
wire n32844;
wire n32845;
wire n32846;
wire n32847;
wire n32848;
wire n32849;
wire n32850;
wire n32851;
wire n32852;
wire n32853;
wire n32854;
wire n32855;
wire n32856;
wire n32857;
wire n32858;
wire n32859;
wire n32860;
wire n32861;
wire n32862;
wire n32863;
wire n32864;
wire n32865;
wire n32866;
wire n32867;
wire n32868;
wire n32869;
wire n3287;
wire n32870;
wire n32871;
wire n32872;
wire n32873;
wire n32874;
wire n32875;
wire n32876;
wire n32877;
wire n32878;
wire n32879;
wire n32880;
wire n32881;
wire n32882;
wire n32883;
wire n32884;
wire n32885;
wire n32886;
wire n32887;
wire n32888;
wire n32889;
wire n32890;
wire n32891;
wire n32892;
wire n32893;
wire n32894;
wire n32895;
wire n32896;
wire n32897;
wire n32898;
wire n32899;
wire n32900;
wire n32901;
wire n32902;
wire n32903;
wire n32904;
wire n32905;
wire n32906;
wire n32907;
wire n32908;
wire n32909;
wire n32910;
wire n32911;
wire n32912;
wire n32913;
wire n32914;
wire n32915;
wire n32916;
wire n32917;
wire n32918;
wire n32919;
wire n3292;
wire n32920;
wire n32921;
wire n32922;
wire n32923;
wire n32924;
wire n32925;
wire n32926;
wire n32927;
wire n32928;
wire n32929;
wire n32930;
wire n32931;
wire n32932;
wire n32933;
wire n32934;
wire n32935;
wire n32936;
wire n32937;
wire n32938;
wire n32939;
wire n32940;
wire n32941;
wire n32942;
wire n32943;
wire n32944;
wire n32945;
wire n32946;
wire n32947;
wire n32948;
wire n32949;
wire n32950;
wire n32951;
wire n32952;
wire n32953;
wire n32954;
wire n32955;
wire n32956;
wire n32957;
wire n32958;
wire n32959;
wire n32960;
wire n32961;
wire n32962;
wire n32963;
wire n32964;
wire n32965;
wire n32966;
wire n32967;
wire n32968;
wire n32969;
wire n3297;
wire n32970;
wire n32971;
wire n32972;
wire n32973;
wire n32974;
wire n32975;
wire n32976;
wire n32977;
wire n32978;
wire n32979;
wire n32980;
wire n32981;
wire n32982;
wire n32983;
wire n32984;
wire n32985;
wire n32986;
wire n32987;
wire n32988;
wire n32989;
wire n32990;
wire n32991;
wire n32992;
wire n32993;
wire n32994;
wire n32995;
wire n32996;
wire n32997;
wire n32998;
wire n32999;
wire n33000;
wire n33001;
wire n33002;
wire n33003;
wire n33004;
wire n33005;
wire n33006;
wire n33007;
wire n33008;
wire n33009;
wire n33010;
wire n33011;
wire n33012;
wire n33013;
wire n33014;
wire n33015;
wire n33016;
wire n33017;
wire n33018;
wire n33019;
wire n3302;
wire n33020;
wire n33021;
wire n33022;
wire n33023;
wire n33024;
wire n33025;
wire n33026;
wire n33027;
wire n33028;
wire n33029;
wire n33030;
wire n33031;
wire n33032;
wire n33033;
wire n33034;
wire n33035;
wire n33036;
wire n33037;
wire n33038;
wire n33039;
wire n33040;
wire n33041;
wire n33042;
wire n33043;
wire n33044;
wire n33045;
wire n33046;
wire n33047;
wire n33048;
wire n33049;
wire n33050;
wire n33051;
wire n33052;
wire n33053;
wire n33054;
wire n33055;
wire n33056;
wire n33057;
wire n33058;
wire n33059;
wire n33060;
wire n33061;
wire n33062;
wire n33063;
wire n33064;
wire n33065;
wire n33066;
wire n33067;
wire n33068;
wire n33069;
wire n3307;
wire n33070;
wire n33071;
wire n33072;
wire n33073;
wire n33074;
wire n33075;
wire n33076;
wire n33077;
wire n33078;
wire n33079;
wire n33080;
wire n33081;
wire n33082;
wire n33083;
wire n33084;
wire n33085;
wire n33086;
wire n33087;
wire n33088;
wire n33089;
wire n33090;
wire n33091;
wire n33092;
wire n33093;
wire n33094;
wire n33095;
wire n33096;
wire n33097;
wire n33098;
wire n33099;
wire n33100;
wire n33101;
wire n33102;
wire n33103;
wire n33104;
wire n33105;
wire n33106;
wire n33107;
wire n33108;
wire n33109;
wire n33110;
wire n33111;
wire n33112;
wire n33113;
wire n33114;
wire n33115;
wire n33116;
wire n33117;
wire n33118;
wire n33119;
wire n3312;
wire n33120;
wire n33121;
wire n33122;
wire n33123;
wire n33124;
wire n33125;
wire n33126;
wire n33127;
wire n33128;
wire n33129;
wire n33130;
wire n33131;
wire n33132;
wire n33133;
wire n33134;
wire n33135;
wire n33136;
wire n33137;
wire n33138;
wire n33139;
wire n33140;
wire n33141;
wire n33142;
wire n33143;
wire n33144;
wire n33145;
wire n33146;
wire n33147;
wire n33148;
wire n33149;
wire n33150;
wire n33151;
wire n33152;
wire n33153;
wire n33154;
wire n33155;
wire n33156;
wire n33157;
wire n33158;
wire n33159;
wire n33160;
wire n33161;
wire n33162;
wire n33163;
wire n33164;
wire n33165;
wire n33166;
wire n33167;
wire n33168;
wire n33169;
wire n3317;
wire n33170;
wire n33171;
wire n33172;
wire n33173;
wire n33174;
wire n33175;
wire n33176;
wire n33177;
wire n33178;
wire n33179;
wire n33180;
wire n33181;
wire n33182;
wire n33183;
wire n33184;
wire n33185;
wire n33186;
wire n33187;
wire n33188;
wire n33189;
wire n33190;
wire n33191;
wire n33192;
wire n33193;
wire n33194;
wire n33195;
wire n33196;
wire n33197;
wire n33198;
wire n33199;
wire n33200;
wire n33201;
wire n33202;
wire n33203;
wire n33204;
wire n33205;
wire n33206;
wire n33207;
wire n33208;
wire n33209;
wire n33210;
wire n33211;
wire n33212;
wire n33213;
wire n33214;
wire n33215;
wire n33216;
wire n33217;
wire n33218;
wire n33219;
wire n3322;
wire n33220;
wire n33221;
wire n33222;
wire n33223;
wire n33224;
wire n33225;
wire n33226;
wire n33227;
wire n33228;
wire n33229;
wire n33230;
wire n33231;
wire n33232;
wire n33233;
wire n33234;
wire n33235;
wire n33236;
wire n33237;
wire n33238;
wire n33239;
wire n33240;
wire n33241;
wire n33242;
wire n33243;
wire n33244;
wire n33245;
wire n33246;
wire n33247;
wire n33248;
wire n33249;
wire n33250;
wire n33251;
wire n33252;
wire n33253;
wire n33254;
wire n33255;
wire n33256;
wire n33257;
wire n33258;
wire n33259;
wire n33260;
wire n33261;
wire n33262;
wire n33263;
wire n33264;
wire n33265;
wire n33266;
wire n33267;
wire n33268;
wire n33269;
wire n3327;
wire n33270;
wire n33271;
wire n33272;
wire n33273;
wire n33274;
wire n33275;
wire n33276;
wire n33277;
wire n33278;
wire n33279;
wire n33280;
wire n33281;
wire n33282;
wire n33283;
wire n33284;
wire n33285;
wire n33286;
wire n33287;
wire n33288;
wire n33289;
wire n33290;
wire n33291;
wire n33292;
wire n33293;
wire n33294;
wire n33295;
wire n33296;
wire n33297;
wire n33298;
wire n33299;
wire n333;
wire n33300;
wire n33301;
wire n33302;
wire n33303;
wire n33304;
wire n33305;
wire n33306;
wire n33307;
wire n33308;
wire n33309;
wire n33310;
wire n33311;
wire n33312;
wire n33313;
wire n33314;
wire n33315;
wire n33316;
wire n33317;
wire n33318;
wire n33319;
wire n3332;
wire n33320;
wire n33321;
wire n33322;
wire n33323;
wire n33324;
wire n33325;
wire n33326;
wire n33327;
wire n33328;
wire n33329;
wire n33330;
wire n33331;
wire n33332;
wire n33333;
wire n33334;
wire n33335;
wire n33336;
wire n33337;
wire n33338;
wire n33339;
wire n33340;
wire n33341;
wire n33342;
wire n33343;
wire n33344;
wire n33345;
wire n33346;
wire n33347;
wire n33348;
wire n33349;
wire n33350;
wire n33351;
wire n33352;
wire n33353;
wire n33354;
wire n33355;
wire n33356;
wire n33357;
wire n33358;
wire n33359;
wire n33360;
wire n33361;
wire n33362;
wire n33363;
wire n33364;
wire n33365;
wire n33366;
wire n33367;
wire n33368;
wire n33369;
wire n3337;
wire n33370;
wire n33371;
wire n33372;
wire n33373;
wire n33374;
wire n33375;
wire n33376;
wire n33377;
wire n33378;
wire n33379;
wire n33380;
wire n33381;
wire n33382;
wire n33383;
wire n33384;
wire n33385;
wire n33386;
wire n33387;
wire n33388;
wire n33389;
wire n33390;
wire n33391;
wire n33392;
wire n33393;
wire n33394;
wire n33395;
wire n33396;
wire n33397;
wire n33398;
wire n33399;
wire n33400;
wire n33401;
wire n33402;
wire n33403;
wire n33404;
wire n33405;
wire n33406;
wire n33407;
wire n33408;
wire n33409;
wire n33410;
wire n33411;
wire n33412;
wire n33413;
wire n33414;
wire n33415;
wire n33416;
wire n33417;
wire n33418;
wire n33419;
wire n3342;
wire n33420;
wire n33421;
wire n33422;
wire n33423;
wire n33424;
wire n33425;
wire n33426;
wire n33427;
wire n33428;
wire n33429;
wire n33430;
wire n33431;
wire n33432;
wire n33433;
wire n33434;
wire n33435;
wire n33436;
wire n33437;
wire n33438;
wire n33439;
wire n33440;
wire n33441;
wire n33442;
wire n33443;
wire n33444;
wire n33445;
wire n33446;
wire n33447;
wire n33448;
wire n33449;
wire n33450;
wire n33451;
wire n33452;
wire n33453;
wire n33454;
wire n33455;
wire n33456;
wire n33457;
wire n33458;
wire n33459;
wire n33460;
wire n33461;
wire n33462;
wire n33463;
wire n33464;
wire n33465;
wire n33466;
wire n33467;
wire n33468;
wire n33469;
wire n3347;
wire n33470;
wire n33471;
wire n33472;
wire n33473;
wire n33474;
wire n33475;
wire n33476;
wire n33477;
wire n33478;
wire n33479;
wire n33480;
wire n33481;
wire n33482;
wire n33483;
wire n33484;
wire n33485;
wire n33486;
wire n33487;
wire n33488;
wire n33489;
wire n33490;
wire n33491;
wire n33492;
wire n33493;
wire n33494;
wire n33495;
wire n33496;
wire n33497;
wire n33498;
wire n33499;
wire n33500;
wire n33501;
wire n33502;
wire n33503;
wire n33504;
wire n33505;
wire n33506;
wire n33507;
wire n33508;
wire n33509;
wire n33510;
wire n33511;
wire n33512;
wire n33513;
wire n33514;
wire n33515;
wire n33516;
wire n33517;
wire n33518;
wire n33519;
wire n3352;
wire n33520;
wire n33521;
wire n33522;
wire n33523;
wire n33524;
wire n33525;
wire n33526;
wire n33527;
wire n33528;
wire n33529;
wire n33530;
wire n33531;
wire n33532;
wire n33533;
wire n33534;
wire n33535;
wire n33536;
wire n33537;
wire n33538;
wire n33539;
wire n33540;
wire n33541;
wire n33542;
wire n33543;
wire n33544;
wire n33545;
wire n33546;
wire n33547;
wire n33548;
wire n33549;
wire n33550;
wire n33551;
wire n33552;
wire n33553;
wire n33554;
wire n33555;
wire n33556;
wire n33557;
wire n33558;
wire n33559;
wire n33560;
wire n33561;
wire n33562;
wire n33563;
wire n33564;
wire n33565;
wire n33566;
wire n33567;
wire n33568;
wire n33569;
wire n3357;
wire n33570;
wire n33571;
wire n33572;
wire n33573;
wire n33574;
wire n33575;
wire n33576;
wire n33577;
wire n33578;
wire n33579;
wire n33580;
wire n33581;
wire n33582;
wire n33583;
wire n33584;
wire n33585;
wire n33586;
wire n33587;
wire n33588;
wire n33589;
wire n33590;
wire n33591;
wire n33592;
wire n33593;
wire n33594;
wire n33595;
wire n33596;
wire n33597;
wire n33598;
wire n33599;
wire n33600;
wire n33601;
wire n33602;
wire n33603;
wire n33604;
wire n33605;
wire n33606;
wire n33607;
wire n33608;
wire n33609;
wire n33610;
wire n33611;
wire n33612;
wire n33613;
wire n33614;
wire n33615;
wire n33616;
wire n33617;
wire n33618;
wire n33619;
wire n3362;
wire n33620;
wire n33621;
wire n33622;
wire n33623;
wire n33624;
wire n33625;
wire n33626;
wire n33627;
wire n33628;
wire n33629;
wire n33630;
wire n33631;
wire n33632;
wire n33633;
wire n33634;
wire n33635;
wire n33636;
wire n33637;
wire n33638;
wire n33639;
wire n33640;
wire n33641;
wire n33642;
wire n33643;
wire n33644;
wire n33645;
wire n33646;
wire n33647;
wire n33648;
wire n33649;
wire n33650;
wire n33651;
wire n33652;
wire n33653;
wire n33654;
wire n33655;
wire n33656;
wire n33657;
wire n33658;
wire n33659;
wire n33660;
wire n33661;
wire n33662;
wire n33663;
wire n33664;
wire n33665;
wire n33666;
wire n33667;
wire n33668;
wire n33669;
wire n3367;
wire n33670;
wire n33671;
wire n33672;
wire n33673;
wire n33674;
wire n33675;
wire n33676;
wire n33677;
wire n33678;
wire n33679;
wire n33680;
wire n33681;
wire n33682;
wire n33683;
wire n33684;
wire n33685;
wire n33686;
wire n33687;
wire n33688;
wire n33689;
wire n33690;
wire n33691;
wire n33692;
wire n33693;
wire n33694;
wire n33695;
wire n33696;
wire n33697;
wire n33698;
wire n33699;
wire n33700;
wire n33701;
wire n33702;
wire n33703;
wire n33704;
wire n33705;
wire n33706;
wire n33707;
wire n33708;
wire n33709;
wire n33710;
wire n33711;
wire n33712;
wire n33713;
wire n33714;
wire n33715;
wire n33716;
wire n33717;
wire n33718;
wire n33719;
wire n3372;
wire n33720;
wire n33721;
wire n33722;
wire n33723;
wire n33724;
wire n33725;
wire n33726;
wire n33727;
wire n33728;
wire n33729;
wire n33730;
wire n33731;
wire n33732;
wire n33733;
wire n33734;
wire n33735;
wire n33736;
wire n33737;
wire n33738;
wire n33739;
wire n33740;
wire n33741;
wire n33742;
wire n33743;
wire n33744;
wire n33745;
wire n33746;
wire n33747;
wire n33748;
wire n33749;
wire n33750;
wire n33751;
wire n33752;
wire n33753;
wire n33754;
wire n33755;
wire n33756;
wire n33757;
wire n33758;
wire n33759;
wire n33760;
wire n33761;
wire n33762;
wire n33763;
wire n33764;
wire n33765;
wire n33766;
wire n33767;
wire n33768;
wire n33769;
wire n3377;
wire n33770;
wire n33771;
wire n33772;
wire n33773;
wire n33774;
wire n33775;
wire n33776;
wire n33777;
wire n33778;
wire n33779;
wire n33780;
wire n33781;
wire n33782;
wire n33783;
wire n33784;
wire n33785;
wire n33786;
wire n33787;
wire n33788;
wire n33789;
wire n33790;
wire n33791;
wire n33792;
wire n33793;
wire n33794;
wire n33795;
wire n33796;
wire n33797;
wire n33798;
wire n33799;
wire n338;
wire n33800;
wire n33801;
wire n33802;
wire n33803;
wire n33804;
wire n33805;
wire n33806;
wire n33807;
wire n33808;
wire n33809;
wire n33810;
wire n33811;
wire n33812;
wire n33813;
wire n33814;
wire n33815;
wire n33816;
wire n33817;
wire n33818;
wire n33819;
wire n3382;
wire n33820;
wire n33821;
wire n33822;
wire n33823;
wire n33824;
wire n33825;
wire n33826;
wire n33827;
wire n33828;
wire n33829;
wire n33830;
wire n33831;
wire n33832;
wire n33833;
wire n33834;
wire n33835;
wire n33836;
wire n33837;
wire n33838;
wire n33839;
wire n33840;
wire n33841;
wire n33842;
wire n33843;
wire n33844;
wire n33845;
wire n33846;
wire n33847;
wire n33848;
wire n33849;
wire n33850;
wire n33851;
wire n33852;
wire n33853;
wire n33854;
wire n33855;
wire n33856;
wire n33857;
wire n33858;
wire n33859;
wire n33860;
wire n33861;
wire n33862;
wire n33863;
wire n33864;
wire n33865;
wire n33866;
wire n33867;
wire n33868;
wire n33869;
wire n3387;
wire n33870;
wire n33871;
wire n33872;
wire n33873;
wire n33874;
wire n33875;
wire n33876;
wire n33877;
wire n33878;
wire n33879;
wire n33880;
wire n33881;
wire n33882;
wire n33883;
wire n33884;
wire n33885;
wire n33886;
wire n33887;
wire n33888;
wire n33889;
wire n33890;
wire n33891;
wire n33892;
wire n33893;
wire n33894;
wire n33895;
wire n33896;
wire n33897;
wire n33898;
wire n33899;
wire n33900;
wire n33901;
wire n33902;
wire n33903;
wire n33904;
wire n33905;
wire n33906;
wire n33907;
wire n33908;
wire n33909;
wire n33910;
wire n33911;
wire n33912;
wire n33913;
wire n33914;
wire n33915;
wire n33916;
wire n33917;
wire n33918;
wire n33919;
wire n3392;
wire n33920;
wire n33921;
wire n33922;
wire n33923;
wire n33924;
wire n33925;
wire n33926;
wire n33927;
wire n33928;
wire n33929;
wire n33930;
wire n33931;
wire n33932;
wire n33933;
wire n33934;
wire n33935;
wire n33936;
wire n33937;
wire n33938;
wire n33939;
wire n33940;
wire n33941;
wire n33942;
wire n33943;
wire n33944;
wire n33945;
wire n33946;
wire n33947;
wire n33948;
wire n33949;
wire n33950;
wire n33951;
wire n33952;
wire n33953;
wire n33954;
wire n33955;
wire n33956;
wire n33957;
wire n33958;
wire n33959;
wire n33960;
wire n33961;
wire n33962;
wire n33963;
wire n33964;
wire n33965;
wire n33966;
wire n33967;
wire n33968;
wire n33969;
wire n3397;
wire n33970;
wire n33971;
wire n33972;
wire n33973;
wire n33974;
wire n33975;
wire n33976;
wire n33977;
wire n33978;
wire n33979;
wire n33980;
wire n33981;
wire n33982;
wire n33983;
wire n33984;
wire n33985;
wire n33986;
wire n33987;
wire n33988;
wire n33989;
wire n33990;
wire n33991;
wire n33992;
wire n33993;
wire n33994;
wire n33995;
wire n33996;
wire n33997;
wire n33998;
wire n33999;
wire n34000;
wire n34001;
wire n34002;
wire n34003;
wire n34004;
wire n34005;
wire n34006;
wire n34007;
wire n34008;
wire n34009;
wire n34010;
wire n34011;
wire n34012;
wire n34013;
wire n34014;
wire n34015;
wire n34016;
wire n34017;
wire n34018;
wire n34019;
wire n3402;
wire n34020;
wire n34021;
wire n34022;
wire n34023;
wire n34024;
wire n34025;
wire n34026;
wire n34027;
wire n34028;
wire n34029;
wire n34030;
wire n34031;
wire n34032;
wire n34033;
wire n34034;
wire n34035;
wire n34036;
wire n34037;
wire n34038;
wire n34039;
wire n34040;
wire n34041;
wire n34042;
wire n34043;
wire n34044;
wire n34045;
wire n34046;
wire n34047;
wire n34048;
wire n34049;
wire n34050;
wire n34051;
wire n34052;
wire n34053;
wire n34054;
wire n34055;
wire n34056;
wire n34057;
wire n34058;
wire n34059;
wire n34060;
wire n34061;
wire n34062;
wire n34063;
wire n34064;
wire n34065;
wire n34066;
wire n34067;
wire n34068;
wire n34069;
wire n3407;
wire n34070;
wire n34071;
wire n34072;
wire n34073;
wire n34074;
wire n34075;
wire n34076;
wire n34077;
wire n34078;
wire n34079;
wire n34080;
wire n34081;
wire n34082;
wire n34083;
wire n34084;
wire n34085;
wire n34086;
wire n34087;
wire n34088;
wire n34089;
wire n34090;
wire n34091;
wire n34092;
wire n34093;
wire n34094;
wire n34095;
wire n34096;
wire n34097;
wire n34098;
wire n34099;
wire n34100;
wire n34101;
wire n34102;
wire n34103;
wire n34104;
wire n34105;
wire n34106;
wire n34107;
wire n34108;
wire n34109;
wire n3411;
wire n34110;
wire n34111;
wire n34112;
wire n34113;
wire n34114;
wire n34115;
wire n34116;
wire n34117;
wire n34118;
wire n34119;
wire n34120;
wire n34121;
wire n34122;
wire n34123;
wire n34124;
wire n34125;
wire n34126;
wire n34127;
wire n34128;
wire n34129;
wire n34130;
wire n34131;
wire n34132;
wire n34133;
wire n34134;
wire n34135;
wire n34136;
wire n34137;
wire n34138;
wire n34139;
wire n34140;
wire n34141;
wire n34142;
wire n34143;
wire n34144;
wire n34145;
wire n34146;
wire n34147;
wire n34148;
wire n34149;
wire n34150;
wire n34151;
wire n34152;
wire n34153;
wire n34154;
wire n34155;
wire n34156;
wire n34157;
wire n34158;
wire n34159;
wire n3416;
wire n34160;
wire n34161;
wire n34162;
wire n34163;
wire n34164;
wire n34165;
wire n34166;
wire n34167;
wire n34168;
wire n34169;
wire n34170;
wire n34171;
wire n34172;
wire n34173;
wire n34174;
wire n34175;
wire n34176;
wire n34177;
wire n34178;
wire n34179;
wire n34180;
wire n34181;
wire n34182;
wire n34183;
wire n34184;
wire n34185;
wire n34186;
wire n34187;
wire n34188;
wire n34189;
wire n34190;
wire n34191;
wire n34192;
wire n34193;
wire n34194;
wire n34195;
wire n34196;
wire n34197;
wire n34198;
wire n34199;
wire n34200;
wire n34201;
wire n34202;
wire n34203;
wire n34204;
wire n34205;
wire n34206;
wire n34207;
wire n34208;
wire n34209;
wire n3421;
wire n34210;
wire n34211;
wire n34212;
wire n34213;
wire n34214;
wire n34215;
wire n34216;
wire n34217;
wire n34218;
wire n34219;
wire n34220;
wire n34221;
wire n34222;
wire n34223;
wire n34224;
wire n34225;
wire n34226;
wire n34227;
wire n34228;
wire n34229;
wire n34230;
wire n34231;
wire n34232;
wire n34233;
wire n34234;
wire n34235;
wire n34236;
wire n34237;
wire n34238;
wire n34239;
wire n34240;
wire n34241;
wire n34242;
wire n34243;
wire n34244;
wire n34245;
wire n34246;
wire n34247;
wire n34248;
wire n34249;
wire n34250;
wire n34251;
wire n34252;
wire n34253;
wire n34254;
wire n34255;
wire n34256;
wire n34257;
wire n34258;
wire n34259;
wire n3426;
wire n34260;
wire n34261;
wire n34262;
wire n34263;
wire n34264;
wire n34265;
wire n34266;
wire n34267;
wire n34268;
wire n34269;
wire n34270;
wire n34271;
wire n34272;
wire n34273;
wire n34274;
wire n34275;
wire n34276;
wire n34277;
wire n34278;
wire n34279;
wire n34280;
wire n34281;
wire n34282;
wire n34283;
wire n34284;
wire n34285;
wire n34286;
wire n34287;
wire n34288;
wire n34289;
wire n34290;
wire n34291;
wire n34292;
wire n34293;
wire n34294;
wire n34295;
wire n34296;
wire n34297;
wire n34298;
wire n34299;
wire n343;
wire n34300;
wire n34301;
wire n34302;
wire n34303;
wire n34304;
wire n34305;
wire n34306;
wire n34307;
wire n34308;
wire n34309;
wire n3431;
wire n34310;
wire n34311;
wire n34312;
wire n34313;
wire n34314;
wire n34315;
wire n34316;
wire n34317;
wire n34318;
wire n34319;
wire n34320;
wire n34321;
wire n34322;
wire n34323;
wire n34324;
wire n34325;
wire n34326;
wire n34327;
wire n34328;
wire n34329;
wire n34330;
wire n34331;
wire n34332;
wire n34333;
wire n34334;
wire n34335;
wire n34336;
wire n34337;
wire n34338;
wire n34339;
wire n34340;
wire n34341;
wire n34342;
wire n34343;
wire n34344;
wire n34345;
wire n34346;
wire n34347;
wire n34348;
wire n34349;
wire n34350;
wire n34351;
wire n34352;
wire n34353;
wire n34354;
wire n34355;
wire n34356;
wire n34357;
wire n34358;
wire n34359;
wire n3436;
wire n34360;
wire n34361;
wire n34362;
wire n34363;
wire n34364;
wire n34365;
wire n34366;
wire n34367;
wire n34368;
wire n34369;
wire n34370;
wire n34371;
wire n34372;
wire n34373;
wire n34374;
wire n34375;
wire n34376;
wire n34377;
wire n34378;
wire n34379;
wire n34380;
wire n34381;
wire n34382;
wire n34383;
wire n34384;
wire n34385;
wire n34386;
wire n34387;
wire n34388;
wire n34389;
wire n34390;
wire n34391;
wire n34392;
wire n34393;
wire n34394;
wire n34395;
wire n34396;
wire n34397;
wire n34398;
wire n34399;
wire n34401;
wire n34402;
wire n34403;
wire n34404;
wire n34405;
wire n34406;
wire n34407;
wire n3441;
wire n34411;
wire n34412;
wire n34413;
wire n34414;
wire n34415;
wire n34416;
wire n34417;
wire n34418;
wire n34420;
wire n34421;
wire n34422;
wire n34423;
wire n34424;
wire n34425;
wire n34426;
wire n34427;
wire n34428;
wire n34429;
wire n34430;
wire n34431;
wire n34432;
wire n34433;
wire n34434;
wire n34435;
wire n34436;
wire n34437;
wire n34438;
wire n34439;
wire n34440;
wire n34441;
wire n34442;
wire n34443;
wire n34444;
wire n34445;
wire n34446;
wire n34447;
wire n34448;
wire n34449;
wire n34450;
wire n34451;
wire n34452;
wire n34453;
wire n34454;
wire n34455;
wire n34456;
wire n34457;
wire n34458;
wire n34459;
wire n3446;
wire n34460;
wire n34461;
wire n34462;
wire n34463;
wire n34464;
wire n34465;
wire n34466;
wire n34467;
wire n34468;
wire n34469;
wire n34470;
wire n34471;
wire n34472;
wire n34473;
wire n34474;
wire n34475;
wire n34476;
wire n34477;
wire n34478;
wire n34479;
wire n34480;
wire n34481;
wire n34482;
wire n34483;
wire n34484;
wire n34485;
wire n34486;
wire n34487;
wire n34488;
wire n34489;
wire n34490;
wire n34491;
wire n34492;
wire n34493;
wire n34494;
wire n34495;
wire n34496;
wire n34497;
wire n34498;
wire n34499;
wire n34500;
wire n34501;
wire n34502;
wire n34503;
wire n34504;
wire n34505;
wire n34506;
wire n34507;
wire n34508;
wire n34509;
wire n3451;
wire n34510;
wire n34511;
wire n34512;
wire n34513;
wire n34514;
wire n34515;
wire n34516;
wire n34517;
wire n34518;
wire n34519;
wire n34520;
wire n34521;
wire n34522;
wire n34523;
wire n34524;
wire n34525;
wire n34526;
wire n34527;
wire n34528;
wire n34529;
wire n34530;
wire n34531;
wire n34532;
wire n34533;
wire n34534;
wire n34535;
wire n34536;
wire n34537;
wire n34538;
wire n34539;
wire n34540;
wire n34541;
wire n34542;
wire n34543;
wire n34544;
wire n34545;
wire n34546;
wire n34547;
wire n34548;
wire n34549;
wire n34550;
wire n34551;
wire n34552;
wire n34553;
wire n34554;
wire n34555;
wire n34556;
wire n34558;
wire n34559;
wire n3456;
wire n34560;
wire n34561;
wire n34562;
wire n34563;
wire n34564;
wire n34565;
wire n34566;
wire n34567;
wire n34568;
wire n34569;
wire n34570;
wire n34571;
wire n34572;
wire n34573;
wire n34574;
wire n34575;
wire n34576;
wire n34577;
wire n34578;
wire n34579;
wire n34580;
wire n34581;
wire n34582;
wire n34583;
wire n34584;
wire n34585;
wire n34586;
wire n34587;
wire n34588;
wire n34589;
wire n34590;
wire n34591;
wire n34592;
wire n34593;
wire n34594;
wire n34595;
wire n34596;
wire n34597;
wire n34598;
wire n34599;
wire n34600;
wire n34601;
wire n34602;
wire n34603;
wire n34604;
wire n34605;
wire n34606;
wire n34607;
wire n34608;
wire n34609;
wire n3461;
wire n34610;
wire n34611;
wire n34612;
wire n34613;
wire n34614;
wire n34615;
wire n34616;
wire n34617;
wire n34618;
wire n34619;
wire n34620;
wire n34621;
wire n34622;
wire n34623;
wire n34624;
wire n34625;
wire n34626;
wire n34627;
wire n34628;
wire n34629;
wire n34630;
wire n34631;
wire n34632;
wire n34633;
wire n34634;
wire n34635;
wire n34636;
wire n34637;
wire n34638;
wire n34639;
wire n34640;
wire n34641;
wire n34642;
wire n34643;
wire n34644;
wire n34645;
wire n34646;
wire n34647;
wire n34648;
wire n34649;
wire n34650;
wire n34651;
wire n34652;
wire n34653;
wire n34654;
wire n34655;
wire n34656;
wire n34657;
wire n34658;
wire n34659;
wire n3466;
wire n34660;
wire n34661;
wire n34662;
wire n34663;
wire n34664;
wire n34665;
wire n34666;
wire n34667;
wire n34668;
wire n34669;
wire n34670;
wire n34671;
wire n34672;
wire n34673;
wire n34674;
wire n34675;
wire n34676;
wire n34677;
wire n34678;
wire n34679;
wire n34680;
wire n34681;
wire n34682;
wire n34683;
wire n34684;
wire n34685;
wire n34686;
wire n34687;
wire n34688;
wire n34689;
wire n34690;
wire n34691;
wire n34692;
wire n34693;
wire n34694;
wire n34695;
wire n34696;
wire n34697;
wire n34698;
wire n34699;
wire n34700;
wire n34701;
wire n34702;
wire n34703;
wire n34704;
wire n34705;
wire n34706;
wire n34707;
wire n34708;
wire n34709;
wire n3471;
wire n34710;
wire n34711;
wire n34712;
wire n34713;
wire n34714;
wire n34715;
wire n34716;
wire n34717;
wire n34718;
wire n34719;
wire n34720;
wire n34721;
wire n34722;
wire n34723;
wire n34724;
wire n34725;
wire n34726;
wire n34727;
wire n34728;
wire n34729;
wire n34730;
wire n34731;
wire n34732;
wire n34733;
wire n34734;
wire n34735;
wire n34736;
wire n34737;
wire n34738;
wire n34739;
wire n34740;
wire n34741;
wire n34742;
wire n34743;
wire n34744;
wire n34745;
wire n34746;
wire n34747;
wire n34748;
wire n34749;
wire n34750;
wire n34751;
wire n34752;
wire n34753;
wire n34754;
wire n34755;
wire n34756;
wire n34757;
wire n34758;
wire n34759;
wire n3476;
wire n34760;
wire n34761;
wire n34762;
wire n34763;
wire n34764;
wire n34765;
wire n34766;
wire n34767;
wire n34768;
wire n34769;
wire n34770;
wire n34771;
wire n34772;
wire n34773;
wire n34774;
wire n34775;
wire n34776;
wire n34777;
wire n34778;
wire n34779;
wire n34780;
wire n34781;
wire n34782;
wire n34783;
wire n34784;
wire n34785;
wire n34786;
wire n34787;
wire n34788;
wire n34789;
wire n34790;
wire n34791;
wire n34792;
wire n34793;
wire n34794;
wire n34795;
wire n34796;
wire n34797;
wire n34798;
wire n34799;
wire n348;
wire n34800;
wire n34801;
wire n34802;
wire n34803;
wire n34804;
wire n34805;
wire n34806;
wire n34807;
wire n34808;
wire n34809;
wire n3481;
wire n34810;
wire n34811;
wire n34812;
wire n34813;
wire n34814;
wire n34815;
wire n34816;
wire n34817;
wire n34818;
wire n34819;
wire n34820;
wire n34821;
wire n34822;
wire n34823;
wire n34824;
wire n34825;
wire n34826;
wire n34827;
wire n34828;
wire n34829;
wire n34830;
wire n34831;
wire n34832;
wire n34833;
wire n34834;
wire n34835;
wire n34836;
wire n34837;
wire n34838;
wire n34839;
wire n34840;
wire n34841;
wire n34842;
wire n34843;
wire n34844;
wire n34845;
wire n34846;
wire n34847;
wire n34848;
wire n34849;
wire n34850;
wire n34851;
wire n34852;
wire n34853;
wire n34854;
wire n34855;
wire n34856;
wire n34857;
wire n34858;
wire n34859;
wire n3486;
wire n34860;
wire n34861;
wire n34862;
wire n34863;
wire n34864;
wire n34865;
wire n34866;
wire n34867;
wire n34868;
wire n34869;
wire n34870;
wire n34871;
wire n34872;
wire n34873;
wire n34874;
wire n34875;
wire n34876;
wire n34877;
wire n34878;
wire n34879;
wire n34880;
wire n34881;
wire n34882;
wire n34883;
wire n34884;
wire n34885;
wire n34886;
wire n34887;
wire n34888;
wire n34889;
wire n34890;
wire n34891;
wire n34892;
wire n34893;
wire n34894;
wire n34895;
wire n34896;
wire n34897;
wire n34898;
wire n34899;
wire n34900;
wire n34901;
wire n34902;
wire n34903;
wire n34904;
wire n34905;
wire n34906;
wire n34907;
wire n34908;
wire n34909;
wire n3491;
wire n34910;
wire n34911;
wire n34912;
wire n34913;
wire n34914;
wire n34915;
wire n34916;
wire n34917;
wire n34918;
wire n34919;
wire n34920;
wire n34921;
wire n34922;
wire n34923;
wire n34924;
wire n34925;
wire n34926;
wire n34927;
wire n34928;
wire n34929;
wire n34930;
wire n34931;
wire n34932;
wire n34933;
wire n34934;
wire n34935;
wire n34937;
wire n34938;
wire n34939;
wire n34940;
wire n34941;
wire n34942;
wire n34943;
wire n34944;
wire n34945;
wire n34946;
wire n34947;
wire n34948;
wire n34949;
wire n34950;
wire n34951;
wire n34952;
wire n34953;
wire n34954;
wire n34955;
wire n34956;
wire n34957;
wire n34958;
wire n34959;
wire n3496;
wire n34960;
wire n34961;
wire n34962;
wire n34963;
wire n34964;
wire n34965;
wire n34966;
wire n34967;
wire n34968;
wire n34969;
wire n34970;
wire n34971;
wire n34972;
wire n34973;
wire n34974;
wire n34975;
wire n34976;
wire n34977;
wire n34978;
wire n34979;
wire n34980;
wire n34981;
wire n34982;
wire n34983;
wire n34984;
wire n34985;
wire n34986;
wire n34987;
wire n34988;
wire n34989;
wire n34990;
wire n34991;
wire n34992;
wire n34993;
wire n34994;
wire n34995;
wire n34996;
wire n34997;
wire n34998;
wire n34999;
wire n35000;
wire n35001;
wire n35002;
wire n35003;
wire n35004;
wire n35005;
wire n35006;
wire n35007;
wire n35008;
wire n35009;
wire n3501;
wire n35010;
wire n35011;
wire n35012;
wire n35013;
wire n35014;
wire n35015;
wire n35016;
wire n35017;
wire n35018;
wire n35019;
wire n35020;
wire n35021;
wire n35022;
wire n35023;
wire n35024;
wire n35025;
wire n35026;
wire n35027;
wire n35028;
wire n35029;
wire n35030;
wire n35031;
wire n35032;
wire n35033;
wire n35034;
wire n35035;
wire n35036;
wire n35037;
wire n35038;
wire n35039;
wire n35040;
wire n35041;
wire n35042;
wire n35043;
wire n35044;
wire n35045;
wire n35046;
wire n35047;
wire n35048;
wire n35049;
wire n35050;
wire n35051;
wire n35052;
wire n35053;
wire n35054;
wire n35055;
wire n35056;
wire n35057;
wire n35058;
wire n35059;
wire n3506;
wire n35060;
wire n35061;
wire n35062;
wire n35063;
wire n35064;
wire n35065;
wire n35066;
wire n35067;
wire n35068;
wire n35069;
wire n35070;
wire n35071;
wire n35072;
wire n35073;
wire n35074;
wire n35075;
wire n35076;
wire n35077;
wire n35078;
wire n35079;
wire n35080;
wire n35081;
wire n35082;
wire n35083;
wire n35084;
wire n35085;
wire n35086;
wire n35087;
wire n35088;
wire n35089;
wire n35090;
wire n35091;
wire n35092;
wire n35093;
wire n35094;
wire n35095;
wire n35096;
wire n35097;
wire n35098;
wire n35099;
wire n35100;
wire n35101;
wire n35102;
wire n35103;
wire n35104;
wire n35105;
wire n35106;
wire n35107;
wire n35108;
wire n35109;
wire n3511;
wire n35110;
wire n35111;
wire n35112;
wire n35113;
wire n35114;
wire n35115;
wire n35116;
wire n35117;
wire n35118;
wire n35119;
wire n35120;
wire n35121;
wire n35122;
wire n35123;
wire n35124;
wire n35125;
wire n35126;
wire n35127;
wire n35128;
wire n35129;
wire n35130;
wire n35131;
wire n35132;
wire n35133;
wire n35134;
wire n35135;
wire n35136;
wire n35137;
wire n35138;
wire n35139;
wire n35140;
wire n35141;
wire n35142;
wire n35143;
wire n35144;
wire n35145;
wire n35146;
wire n35147;
wire n35148;
wire n35149;
wire n35150;
wire n35151;
wire n35152;
wire n35153;
wire n35154;
wire n35155;
wire n35156;
wire n35157;
wire n35158;
wire n35159;
wire n3516;
wire n35160;
wire n35161;
wire n35162;
wire n35163;
wire n35164;
wire n35165;
wire n35166;
wire n35167;
wire n35168;
wire n35169;
wire n35170;
wire n35171;
wire n35172;
wire n35173;
wire n35174;
wire n35175;
wire n35176;
wire n35177;
wire n35178;
wire n35179;
wire n35180;
wire n35181;
wire n35182;
wire n35183;
wire n35184;
wire n35185;
wire n35186;
wire n35187;
wire n35188;
wire n35189;
wire n35190;
wire n35191;
wire n35192;
wire n35193;
wire n35194;
wire n35195;
wire n35196;
wire n35197;
wire n35198;
wire n35199;
wire n35200;
wire n35201;
wire n35202;
wire n35203;
wire n35204;
wire n35205;
wire n35206;
wire n35207;
wire n35208;
wire n35209;
wire n3521;
wire n35210;
wire n35211;
wire n35212;
wire n35213;
wire n35214;
wire n35215;
wire n35216;
wire n35217;
wire n35218;
wire n35219;
wire n35220;
wire n35221;
wire n35222;
wire n35223;
wire n35224;
wire n35225;
wire n35226;
wire n35227;
wire n35228;
wire n35229;
wire n35230;
wire n35231;
wire n35232;
wire n35233;
wire n35234;
wire n35235;
wire n35236;
wire n35237;
wire n35238;
wire n35239;
wire n35240;
wire n35241;
wire n35242;
wire n35243;
wire n35244;
wire n35245;
wire n35246;
wire n35247;
wire n35248;
wire n35249;
wire n35250;
wire n35251;
wire n35252;
wire n35253;
wire n35254;
wire n35255;
wire n35256;
wire n35258;
wire n35259;
wire n3526;
wire n35260;
wire n35261;
wire n35262;
wire n35263;
wire n35264;
wire n35265;
wire n35266;
wire n35267;
wire n35268;
wire n35269;
wire n35270;
wire n35271;
wire n35272;
wire n35273;
wire n35274;
wire n35275;
wire n35276;
wire n35277;
wire n35278;
wire n35279;
wire n35280;
wire n35281;
wire n35282;
wire n35283;
wire n35284;
wire n35285;
wire n35286;
wire n35287;
wire n35288;
wire n35289;
wire n35290;
wire n35291;
wire n35292;
wire n35293;
wire n35294;
wire n35295;
wire n35296;
wire n35297;
wire n35298;
wire n35299;
wire n353;
wire n35300;
wire n35301;
wire n35302;
wire n35303;
wire n35304;
wire n35305;
wire n35306;
wire n35307;
wire n35308;
wire n35309;
wire n3531;
wire n35310;
wire n35311;
wire n35312;
wire n35313;
wire n35314;
wire n35315;
wire n35316;
wire n35317;
wire n35318;
wire n35319;
wire n35320;
wire n35321;
wire n35322;
wire n35323;
wire n35324;
wire n35325;
wire n35326;
wire n35327;
wire n35328;
wire n35329;
wire n35330;
wire n35331;
wire n35332;
wire n35333;
wire n35334;
wire n35335;
wire n35336;
wire n35337;
wire n35338;
wire n35339;
wire n35340;
wire n35341;
wire n35342;
wire n35343;
wire n35344;
wire n35345;
wire n35346;
wire n35347;
wire n35348;
wire n35349;
wire n3535;
wire n35350;
wire n35351;
wire n35352;
wire n35353;
wire n35354;
wire n35355;
wire n35356;
wire n35357;
wire n35358;
wire n35359;
wire n35360;
wire n35361;
wire n35362;
wire n35363;
wire n35364;
wire n35365;
wire n35366;
wire n35367;
wire n35368;
wire n35369;
wire n35370;
wire n35371;
wire n35372;
wire n35373;
wire n35374;
wire n35375;
wire n35376;
wire n35377;
wire n35378;
wire n35379;
wire n35380;
wire n35381;
wire n35382;
wire n35383;
wire n35384;
wire n35385;
wire n35386;
wire n35387;
wire n35388;
wire n35389;
wire n35390;
wire n35391;
wire n35392;
wire n35393;
wire n35394;
wire n35395;
wire n35396;
wire n35397;
wire n35398;
wire n35399;
wire n3540;
wire n35400;
wire n35401;
wire n35402;
wire n35403;
wire n35404;
wire n35405;
wire n35406;
wire n35407;
wire n35408;
wire n35409;
wire n35410;
wire n35411;
wire n35412;
wire n35413;
wire n35414;
wire n35415;
wire n35416;
wire n35417;
wire n35418;
wire n35419;
wire n35420;
wire n35421;
wire n35422;
wire n35423;
wire n35424;
wire n35425;
wire n35426;
wire n35427;
wire n35428;
wire n35429;
wire n35430;
wire n35431;
wire n35432;
wire n35433;
wire n35434;
wire n35435;
wire n35436;
wire n35437;
wire n35438;
wire n35439;
wire n35440;
wire n35441;
wire n35442;
wire n35443;
wire n35444;
wire n35445;
wire n35446;
wire n35447;
wire n35448;
wire n35449;
wire n3545;
wire n35450;
wire n35451;
wire n35452;
wire n35453;
wire n35454;
wire n35455;
wire n35456;
wire n35457;
wire n35458;
wire n35459;
wire n35460;
wire n35461;
wire n35462;
wire n35463;
wire n35464;
wire n35465;
wire n35466;
wire n35467;
wire n35468;
wire n35469;
wire n35470;
wire n35471;
wire n35472;
wire n35473;
wire n35474;
wire n35475;
wire n35476;
wire n35477;
wire n35478;
wire n35479;
wire n35480;
wire n35481;
wire n35482;
wire n35483;
wire n35484;
wire n35485;
wire n35486;
wire n35487;
wire n35488;
wire n35489;
wire n35490;
wire n35491;
wire n35492;
wire n35493;
wire n35494;
wire n35495;
wire n35496;
wire n35497;
wire n35498;
wire n35499;
wire n3550;
wire n35500;
wire n35501;
wire n35502;
wire n35503;
wire n35504;
wire n35505;
wire n35506;
wire n35507;
wire n35508;
wire n35509;
wire n35510;
wire n35511;
wire n35512;
wire n35513;
wire n35514;
wire n35515;
wire n35516;
wire n35517;
wire n35518;
wire n35519;
wire n35520;
wire n35521;
wire n35522;
wire n35523;
wire n35524;
wire n35525;
wire n35526;
wire n35527;
wire n35528;
wire n35529;
wire n35530;
wire n35531;
wire n35532;
wire n35533;
wire n35534;
wire n35535;
wire n35536;
wire n35537;
wire n35538;
wire n35539;
wire n35540;
wire n35541;
wire n35542;
wire n35543;
wire n35544;
wire n35545;
wire n35546;
wire n35547;
wire n35548;
wire n35549;
wire n3555;
wire n35550;
wire n35551;
wire n35552;
wire n35553;
wire n35554;
wire n35555;
wire n35556;
wire n35557;
wire n35558;
wire n35559;
wire n35560;
wire n35561;
wire n35562;
wire n35564;
wire n35565;
wire n35566;
wire n35567;
wire n35569;
wire n35570;
wire n35571;
wire n35572;
wire n35573;
wire n35575;
wire n35576;
wire n35577;
wire n35578;
wire n35579;
wire n35580;
wire n35581;
wire n35582;
wire n35583;
wire n35585;
wire n35586;
wire n35588;
wire n35589;
wire n35590;
wire n35591;
wire n35592;
wire n35593;
wire n35595;
wire n35596;
wire n35597;
wire n35598;
wire n35599;
wire n3560;
wire n35600;
wire n35601;
wire n35602;
wire n35603;
wire n35604;
wire n35605;
wire n35606;
wire n35607;
wire n35608;
wire n35609;
wire n35610;
wire n35611;
wire n35612;
wire n35613;
wire n35614;
wire n35615;
wire n35616;
wire n35617;
wire n35618;
wire n35619;
wire n35620;
wire n35621;
wire n35622;
wire n35623;
wire n35624;
wire n35625;
wire n35626;
wire n35627;
wire n35628;
wire n35629;
wire n35630;
wire n35631;
wire n35632;
wire n35633;
wire n35634;
wire n35635;
wire n35636;
wire n35637;
wire n35638;
wire n35639;
wire n35640;
wire n35641;
wire n35642;
wire n35643;
wire n35644;
wire n35645;
wire n35646;
wire n35647;
wire n35648;
wire n35649;
wire n3565;
wire n35650;
wire n35651;
wire n35652;
wire n35653;
wire n35654;
wire n35655;
wire n35656;
wire n35657;
wire n35658;
wire n35659;
wire n35660;
wire n35661;
wire n35662;
wire n35663;
wire n35664;
wire n35665;
wire n35666;
wire n35667;
wire n35668;
wire n35669;
wire n35670;
wire n35671;
wire n35672;
wire n35673;
wire n35674;
wire n35675;
wire n35676;
wire n35677;
wire n35678;
wire n35679;
wire n35680;
wire n35681;
wire n35682;
wire n35683;
wire n35684;
wire n35685;
wire n35686;
wire n35687;
wire n35688;
wire n35689;
wire n35690;
wire n35691;
wire n35692;
wire n35693;
wire n35694;
wire n35695;
wire n35696;
wire n35697;
wire n35698;
wire n35699;
wire n3570;
wire n35700;
wire n35701;
wire n35702;
wire n35703;
wire n35704;
wire n35705;
wire n35706;
wire n35707;
wire n35708;
wire n35709;
wire n35710;
wire n35711;
wire n35712;
wire n35713;
wire n35714;
wire n35715;
wire n35716;
wire n35717;
wire n35718;
wire n35719;
wire n35720;
wire n35721;
wire n35722;
wire n35723;
wire n35724;
wire n35725;
wire n35726;
wire n35727;
wire n35728;
wire n35729;
wire n35730;
wire n35731;
wire n35732;
wire n35733;
wire n35734;
wire n35735;
wire n35736;
wire n35737;
wire n35738;
wire n35739;
wire n35740;
wire n35741;
wire n35742;
wire n35743;
wire n35744;
wire n35745;
wire n35746;
wire n35747;
wire n35748;
wire n35749;
wire n3575;
wire n35750;
wire n35751;
wire n35752;
wire n35753;
wire n35754;
wire n35755;
wire n35756;
wire n35757;
wire n35758;
wire n35759;
wire n35760;
wire n35761;
wire n35762;
wire n35763;
wire n35764;
wire n35765;
wire n35766;
wire n35767;
wire n35768;
wire n35769;
wire n35770;
wire n35771;
wire n35772;
wire n35773;
wire n35774;
wire n35775;
wire n35776;
wire n35777;
wire n35778;
wire n35779;
wire n35780;
wire n35781;
wire n35782;
wire n35783;
wire n35784;
wire n35785;
wire n35786;
wire n35787;
wire n35788;
wire n35789;
wire n35790;
wire n35791;
wire n35792;
wire n35793;
wire n35794;
wire n35795;
wire n35796;
wire n35797;
wire n35798;
wire n35799;
wire n358;
wire n3580;
wire n35800;
wire n35801;
wire n35802;
wire n35803;
wire n35804;
wire n35805;
wire n35806;
wire n35807;
wire n35808;
wire n35809;
wire n35810;
wire n35811;
wire n35812;
wire n35813;
wire n35814;
wire n35815;
wire n35816;
wire n35817;
wire n35818;
wire n35819;
wire n35820;
wire n35821;
wire n35822;
wire n35823;
wire n35824;
wire n35825;
wire n35826;
wire n35827;
wire n35828;
wire n35829;
wire n35830;
wire n35831;
wire n35832;
wire n35833;
wire n35834;
wire n35835;
wire n35836;
wire n35837;
wire n35838;
wire n35839;
wire n35840;
wire n35841;
wire n35842;
wire n35843;
wire n35844;
wire n35845;
wire n35846;
wire n35847;
wire n35848;
wire n35849;
wire n3585;
wire n35850;
wire n35851;
wire n35852;
wire n35853;
wire n35854;
wire n35855;
wire n35856;
wire n35857;
wire n35858;
wire n35859;
wire n35860;
wire n35861;
wire n35862;
wire n35863;
wire n35864;
wire n35865;
wire n35866;
wire n35867;
wire n35868;
wire n35869;
wire n35870;
wire n35871;
wire n35872;
wire n35873;
wire n35874;
wire n35875;
wire n35876;
wire n35877;
wire n35878;
wire n35879;
wire n35880;
wire n35881;
wire n35882;
wire n35883;
wire n35884;
wire n35885;
wire n35886;
wire n35887;
wire n35888;
wire n35889;
wire n35890;
wire n35891;
wire n35892;
wire n35893;
wire n35894;
wire n35895;
wire n35896;
wire n35897;
wire n35898;
wire n35899;
wire n3590;
wire n35900;
wire n35901;
wire n35902;
wire n35903;
wire n35904;
wire n35905;
wire n35906;
wire n35907;
wire n35908;
wire n35909;
wire n35910;
wire n35911;
wire n35912;
wire n35913;
wire n35914;
wire n35915;
wire n35916;
wire n35917;
wire n35918;
wire n35919;
wire n35920;
wire n35921;
wire n35922;
wire n35923;
wire n35924;
wire n35925;
wire n35926;
wire n35927;
wire n35928;
wire n35929;
wire n35930;
wire n35931;
wire n35932;
wire n35933;
wire n35934;
wire n35935;
wire n35936;
wire n35937;
wire n35938;
wire n35939;
wire n35940;
wire n35941;
wire n35942;
wire n35943;
wire n35944;
wire n35945;
wire n35946;
wire n35947;
wire n35948;
wire n35949;
wire n3595;
wire n35950;
wire n35951;
wire n35952;
wire n35953;
wire n35954;
wire n35955;
wire n35956;
wire n35957;
wire n35958;
wire n35959;
wire n35960;
wire n35961;
wire n35962;
wire n35963;
wire n35964;
wire n35965;
wire n35966;
wire n35967;
wire n35968;
wire n35969;
wire n35970;
wire n35971;
wire n35972;
wire n35973;
wire n35974;
wire n35975;
wire n35976;
wire n35977;
wire n35978;
wire n35979;
wire n35980;
wire n35982;
wire n35983;
wire n35984;
wire n35985;
wire n35986;
wire n35987;
wire n35988;
wire n35989;
wire n35990;
wire n35991;
wire n35992;
wire n35993;
wire n35994;
wire n35995;
wire n35996;
wire n35997;
wire n35998;
wire n35999;
wire n3600;
wire n36000;
wire n36001;
wire n36002;
wire n36003;
wire n36004;
wire n36005;
wire n36006;
wire n36007;
wire n36008;
wire n36009;
wire n36010;
wire n36011;
wire n36012;
wire n36013;
wire n36014;
wire n36015;
wire n36016;
wire n36017;
wire n36018;
wire n36019;
wire n36020;
wire n36021;
wire n36022;
wire n36023;
wire n36024;
wire n36025;
wire n36026;
wire n36027;
wire n36028;
wire n36029;
wire n36030;
wire n36031;
wire n36032;
wire n36033;
wire n36034;
wire n36035;
wire n36036;
wire n36037;
wire n36038;
wire n36039;
wire n3604;
wire n36040;
wire n36041;
wire n36042;
wire n36043;
wire n36044;
wire n36045;
wire n36046;
wire n36047;
wire n36048;
wire n36049;
wire n36050;
wire n36051;
wire n36052;
wire n36053;
wire n36054;
wire n36055;
wire n36056;
wire n36057;
wire n36058;
wire n36059;
wire n36060;
wire n36061;
wire n36062;
wire n36063;
wire n36064;
wire n36065;
wire n36066;
wire n36067;
wire n36068;
wire n36069;
wire n36070;
wire n36071;
wire n36072;
wire n36073;
wire n36074;
wire n36075;
wire n36076;
wire n36077;
wire n36078;
wire n36079;
wire n36080;
wire n36081;
wire n36082;
wire n36083;
wire n36084;
wire n36085;
wire n36086;
wire n36087;
wire n36088;
wire n36089;
wire n3609;
wire n36090;
wire n36091;
wire n36092;
wire n36093;
wire n36094;
wire n36095;
wire n36096;
wire n36097;
wire n36098;
wire n36099;
wire n36100;
wire n36101;
wire n36102;
wire n36103;
wire n36104;
wire n36105;
wire n36106;
wire n36107;
wire n36108;
wire n36109;
wire n36110;
wire n36111;
wire n36112;
wire n36113;
wire n36114;
wire n36115;
wire n36116;
wire n36117;
wire n36118;
wire n36119;
wire n36120;
wire n36121;
wire n36122;
wire n36123;
wire n36124;
wire n36125;
wire n36126;
wire n36127;
wire n36128;
wire n36129;
wire n36130;
wire n36131;
wire n36132;
wire n36133;
wire n36134;
wire n36135;
wire n36136;
wire n36137;
wire n36138;
wire n36139;
wire n3614;
wire n36140;
wire n36141;
wire n36142;
wire n36143;
wire n36144;
wire n36145;
wire n36146;
wire n36147;
wire n36148;
wire n36149;
wire n36150;
wire n36151;
wire n36152;
wire n36153;
wire n36154;
wire n36155;
wire n36156;
wire n36157;
wire n36158;
wire n36159;
wire n36160;
wire n36161;
wire n36162;
wire n36163;
wire n36164;
wire n36165;
wire n36166;
wire n36167;
wire n36168;
wire n36169;
wire n36170;
wire n36171;
wire n36172;
wire n36173;
wire n36174;
wire n36175;
wire n36176;
wire n36177;
wire n36178;
wire n36179;
wire n36180;
wire n36181;
wire n36182;
wire n36183;
wire n36184;
wire n36185;
wire n36186;
wire n36187;
wire n36188;
wire n36189;
wire n3619;
wire n36190;
wire n36191;
wire n36192;
wire n36193;
wire n36194;
wire n36195;
wire n36196;
wire n36197;
wire n36198;
wire n36199;
wire n36200;
wire n36201;
wire n36202;
wire n36203;
wire n36204;
wire n36205;
wire n36206;
wire n36207;
wire n36208;
wire n36209;
wire n36210;
wire n36211;
wire n36212;
wire n36213;
wire n36214;
wire n36215;
wire n36216;
wire n36217;
wire n36218;
wire n36219;
wire n36220;
wire n36222;
wire n36223;
wire n36224;
wire n36225;
wire n36226;
wire n36227;
wire n36228;
wire n36229;
wire n3623;
wire n36230;
wire n36231;
wire n36232;
wire n36233;
wire n36234;
wire n36235;
wire n36236;
wire n36237;
wire n36238;
wire n36239;
wire n36240;
wire n36241;
wire n36242;
wire n36243;
wire n36244;
wire n36245;
wire n36246;
wire n36247;
wire n36248;
wire n36249;
wire n36250;
wire n36251;
wire n36252;
wire n36253;
wire n36254;
wire n36255;
wire n36256;
wire n36257;
wire n36258;
wire n36259;
wire n36260;
wire n36261;
wire n36262;
wire n36263;
wire n36264;
wire n36265;
wire n36266;
wire n36267;
wire n36268;
wire n36269;
wire n36270;
wire n36271;
wire n36272;
wire n36273;
wire n36274;
wire n36275;
wire n36276;
wire n36277;
wire n36278;
wire n36279;
wire n3628;
wire n36280;
wire n36281;
wire n36282;
wire n36283;
wire n36284;
wire n36285;
wire n36286;
wire n36287;
wire n36288;
wire n36289;
wire n36290;
wire n36291;
wire n36292;
wire n36293;
wire n36294;
wire n36295;
wire n36296;
wire n36297;
wire n36298;
wire n36299;
wire n363;
wire n36300;
wire n36301;
wire n36302;
wire n36303;
wire n36304;
wire n36305;
wire n36306;
wire n36307;
wire n36308;
wire n36309;
wire n36310;
wire n36311;
wire n36312;
wire n36313;
wire n36314;
wire n36315;
wire n36316;
wire n36317;
wire n36318;
wire n36319;
wire n36320;
wire n36321;
wire n36322;
wire n36323;
wire n36324;
wire n36325;
wire n36326;
wire n36327;
wire n36328;
wire n36329;
wire n3633;
wire n36330;
wire n36331;
wire n36332;
wire n36333;
wire n36334;
wire n36335;
wire n36336;
wire n36337;
wire n36338;
wire n36339;
wire n36340;
wire n36341;
wire n36342;
wire n36343;
wire n36344;
wire n36345;
wire n36346;
wire n36347;
wire n36348;
wire n36349;
wire n36350;
wire n36351;
wire n36352;
wire n36353;
wire n36354;
wire n36355;
wire n36356;
wire n36357;
wire n36358;
wire n36359;
wire n36360;
wire n36361;
wire n36362;
wire n36363;
wire n36364;
wire n36365;
wire n36366;
wire n36367;
wire n36368;
wire n36369;
wire n36370;
wire n36371;
wire n36372;
wire n36373;
wire n36374;
wire n36375;
wire n36376;
wire n36377;
wire n36378;
wire n36379;
wire n3638;
wire n36380;
wire n36381;
wire n36382;
wire n36383;
wire n36384;
wire n36385;
wire n36386;
wire n36387;
wire n36388;
wire n36389;
wire n36390;
wire n36391;
wire n36392;
wire n36393;
wire n36394;
wire n36395;
wire n36396;
wire n36398;
wire n36399;
wire n36401;
wire n36402;
wire n36403;
wire n36404;
wire n36406;
wire n36407;
wire n36408;
wire n36409;
wire n36410;
wire n36411;
wire n36412;
wire n36413;
wire n36414;
wire n36415;
wire n36416;
wire n36417;
wire n36418;
wire n36419;
wire n36420;
wire n36421;
wire n36422;
wire n36423;
wire n36424;
wire n36425;
wire n36426;
wire n36427;
wire n36428;
wire n36429;
wire n3643;
wire n36430;
wire n36431;
wire n36432;
wire n36433;
wire n36434;
wire n36435;
wire n36436;
wire n36437;
wire n36438;
wire n36439;
wire n36440;
wire n36441;
wire n36442;
wire n36443;
wire n36444;
wire n36445;
wire n36446;
wire n36447;
wire n36448;
wire n36449;
wire n36450;
wire n36451;
wire n36452;
wire n36453;
wire n36454;
wire n36455;
wire n36456;
wire n36457;
wire n36458;
wire n36459;
wire n36460;
wire n36461;
wire n36462;
wire n36463;
wire n36464;
wire n36465;
wire n36466;
wire n36467;
wire n36468;
wire n36469;
wire n36470;
wire n36471;
wire n36472;
wire n36473;
wire n36474;
wire n36475;
wire n36476;
wire n36477;
wire n36478;
wire n36479;
wire n3648;
wire n36480;
wire n36481;
wire n36482;
wire n36483;
wire n36484;
wire n36485;
wire n36486;
wire n36487;
wire n36488;
wire n36489;
wire n36490;
wire n36491;
wire n36492;
wire n36493;
wire n36494;
wire n36495;
wire n36496;
wire n36497;
wire n36498;
wire n36499;
wire n36500;
wire n36501;
wire n36502;
wire n36503;
wire n36504;
wire n36505;
wire n36506;
wire n36507;
wire n36508;
wire n36509;
wire n36510;
wire n36511;
wire n36512;
wire n36513;
wire n36515;
wire n36516;
wire n36517;
wire n36518;
wire n36519;
wire n36520;
wire n36521;
wire n36522;
wire n36523;
wire n36524;
wire n36525;
wire n36526;
wire n36528;
wire n36529;
wire n3653;
wire n36530;
wire n36531;
wire n36532;
wire n36533;
wire n36534;
wire n36535;
wire n36536;
wire n36537;
wire n36538;
wire n36539;
wire n36540;
wire n36541;
wire n36543;
wire n36544;
wire n36545;
wire n36546;
wire n36547;
wire n36548;
wire n36549;
wire n36550;
wire n36551;
wire n36552;
wire n36553;
wire n36554;
wire n36555;
wire n36556;
wire n36557;
wire n36558;
wire n36559;
wire n36560;
wire n36561;
wire n36562;
wire n36563;
wire n36564;
wire n36565;
wire n36566;
wire n36567;
wire n36568;
wire n36569;
wire n36570;
wire n36571;
wire n36572;
wire n36573;
wire n36574;
wire n36575;
wire n36576;
wire n36577;
wire n36578;
wire n36579;
wire n3658;
wire n36580;
wire n36581;
wire n36582;
wire n36583;
wire n36584;
wire n36585;
wire n36586;
wire n36587;
wire n36588;
wire n36589;
wire n36590;
wire n36591;
wire n36592;
wire n36593;
wire n36594;
wire n36595;
wire n36596;
wire n36597;
wire n36598;
wire n36599;
wire n36600;
wire n36601;
wire n36602;
wire n36603;
wire n36604;
wire n36605;
wire n36606;
wire n36607;
wire n36608;
wire n36609;
wire n36610;
wire n36611;
wire n36612;
wire n36613;
wire n36614;
wire n36615;
wire n36616;
wire n36617;
wire n36618;
wire n36620;
wire n36621;
wire n36622;
wire n36623;
wire n36624;
wire n36625;
wire n36626;
wire n36627;
wire n36628;
wire n36629;
wire n3663;
wire n36630;
wire n36631;
wire n36632;
wire n36633;
wire n36634;
wire n36635;
wire n36636;
wire n36637;
wire n36638;
wire n36639;
wire n36640;
wire n36641;
wire n36642;
wire n36643;
wire n36644;
wire n36645;
wire n36646;
wire n36647;
wire n36648;
wire n36649;
wire n36650;
wire n36651;
wire n36652;
wire n36653;
wire n36654;
wire n36655;
wire n36656;
wire n36657;
wire n36658;
wire n36659;
wire n36660;
wire n36661;
wire n36662;
wire n36663;
wire n36664;
wire n36665;
wire n36666;
wire n36667;
wire n36668;
wire n36669;
wire n36670;
wire n36671;
wire n36672;
wire n36673;
wire n36675;
wire n36677;
wire n36678;
wire n36679;
wire n3668;
wire n36680;
wire n36681;
wire n36682;
wire n36683;
wire n36685;
wire n36687;
wire n36688;
wire n36689;
wire n36690;
wire n36691;
wire n36692;
wire n36693;
wire n36694;
wire n36695;
wire n36696;
wire n36697;
wire n36698;
wire n36699;
wire n36700;
wire n36701;
wire n36702;
wire n36703;
wire n36704;
wire n36705;
wire n36706;
wire n36707;
wire n36708;
wire n36709;
wire n36710;
wire n36711;
wire n36712;
wire n36713;
wire n36714;
wire n36715;
wire n36716;
wire n36717;
wire n36718;
wire n36719;
wire n36720;
wire n36721;
wire n36722;
wire n36723;
wire n36724;
wire n36725;
wire n36726;
wire n36727;
wire n36728;
wire n36729;
wire n3673;
wire n36730;
wire n36731;
wire n36732;
wire n36733;
wire n36734;
wire n36735;
wire n36736;
wire n36737;
wire n36738;
wire n36739;
wire n36740;
wire n36741;
wire n36742;
wire n36743;
wire n36744;
wire n36745;
wire n36746;
wire n36747;
wire n36748;
wire n36749;
wire n36750;
wire n36751;
wire n36752;
wire n36753;
wire n36754;
wire n36755;
wire n36756;
wire n36757;
wire n36758;
wire n36759;
wire n36760;
wire n36761;
wire n36762;
wire n36763;
wire n36764;
wire n36765;
wire n36766;
wire n36767;
wire n36768;
wire n36769;
wire n36770;
wire n36771;
wire n36772;
wire n36773;
wire n36774;
wire n36775;
wire n36776;
wire n36777;
wire n36778;
wire n36779;
wire n3678;
wire n36780;
wire n36781;
wire n36782;
wire n36783;
wire n36784;
wire n36785;
wire n36786;
wire n36787;
wire n36788;
wire n36789;
wire n36790;
wire n36791;
wire n36792;
wire n36793;
wire n36794;
wire n36795;
wire n36796;
wire n36797;
wire n36798;
wire n36799;
wire n368;
wire n36800;
wire n36801;
wire n36803;
wire n36804;
wire n36805;
wire n36806;
wire n36807;
wire n36808;
wire n36809;
wire n36810;
wire n36811;
wire n36812;
wire n36813;
wire n36814;
wire n36815;
wire n36816;
wire n36817;
wire n36818;
wire n36819;
wire n36820;
wire n36821;
wire n36822;
wire n36823;
wire n36824;
wire n36825;
wire n36826;
wire n36827;
wire n36828;
wire n36829;
wire n3683;
wire n36830;
wire n36831;
wire n36832;
wire n36833;
wire n36834;
wire n36835;
wire n36836;
wire n36837;
wire n36838;
wire n36839;
wire n36840;
wire n36841;
wire n36842;
wire n36843;
wire n36844;
wire n36845;
wire n36846;
wire n36847;
wire n36848;
wire n36849;
wire n36850;
wire n36851;
wire n36852;
wire n36853;
wire n36854;
wire n36855;
wire n36856;
wire n36857;
wire n36858;
wire n36859;
wire n36860;
wire n36861;
wire n36862;
wire n36863;
wire n36864;
wire n36865;
wire n36866;
wire n36867;
wire n36868;
wire n36869;
wire n36870;
wire n36871;
wire n36872;
wire n36873;
wire n36874;
wire n36875;
wire n36876;
wire n36877;
wire n36878;
wire n36879;
wire n3688;
wire n36880;
wire n36881;
wire n36882;
wire n36883;
wire n36884;
wire n36885;
wire n36886;
wire n36887;
wire n36888;
wire n36889;
wire n36890;
wire n36891;
wire n36892;
wire n36893;
wire n36895;
wire n36896;
wire n36897;
wire n36898;
wire n36899;
wire n36900;
wire n36901;
wire n36902;
wire n36903;
wire n36904;
wire n36905;
wire n36906;
wire n36907;
wire n36908;
wire n36909;
wire n36910;
wire n36911;
wire n36912;
wire n36913;
wire n36914;
wire n36915;
wire n36916;
wire n36917;
wire n36918;
wire n36919;
wire n36920;
wire n36921;
wire n36922;
wire n36923;
wire n36924;
wire n36925;
wire n36926;
wire n36927;
wire n36928;
wire n36929;
wire n3693;
wire n36930;
wire n36931;
wire n36932;
wire n36933;
wire n36934;
wire n36935;
wire n36936;
wire n36937;
wire n36938;
wire n36939;
wire n36940;
wire n36941;
wire n36942;
wire n36943;
wire n36944;
wire n36945;
wire n36946;
wire n36947;
wire n36948;
wire n36949;
wire n36950;
wire n36951;
wire n36952;
wire n36953;
wire n36954;
wire n36955;
wire n36956;
wire n36957;
wire n36958;
wire n36959;
wire n36960;
wire n36961;
wire n36962;
wire n36963;
wire n36964;
wire n36965;
wire n36966;
wire n36967;
wire n36968;
wire n36969;
wire n36970;
wire n36971;
wire n36972;
wire n36973;
wire n36974;
wire n36975;
wire n36976;
wire n36977;
wire n36978;
wire n36979;
wire n3698;
wire n36980;
wire n36981;
wire n36982;
wire n36983;
wire n36984;
wire n36985;
wire n36986;
wire n36987;
wire n36988;
wire n36989;
wire n36990;
wire n36991;
wire n36992;
wire n36993;
wire n36994;
wire n36995;
wire n36996;
wire n36997;
wire n36998;
wire n36999;
wire n37000;
wire n37001;
wire n37002;
wire n37003;
wire n37004;
wire n37005;
wire n37006;
wire n37007;
wire n37008;
wire n37009;
wire n37010;
wire n37011;
wire n37012;
wire n37013;
wire n37014;
wire n37015;
wire n37016;
wire n37017;
wire n37018;
wire n37019;
wire n37020;
wire n37021;
wire n37022;
wire n37023;
wire n37024;
wire n37025;
wire n37026;
wire n37027;
wire n37028;
wire n37029;
wire n3703;
wire n37030;
wire n37031;
wire n37032;
wire n37033;
wire n37034;
wire n37035;
wire n37036;
wire n37037;
wire n37038;
wire n37039;
wire n37040;
wire n37041;
wire n37042;
wire n37043;
wire n37044;
wire n37045;
wire n37046;
wire n37047;
wire n37048;
wire n37049;
wire n37050;
wire n37051;
wire n37052;
wire n37053;
wire n37054;
wire n37055;
wire n37056;
wire n37057;
wire n37058;
wire n37059;
wire n37060;
wire n37061;
wire n37062;
wire n37063;
wire n37064;
wire n37065;
wire n37066;
wire n37067;
wire n37068;
wire n37069;
wire n3707;
wire n37070;
wire n37071;
wire n37072;
wire n37073;
wire n37074;
wire n37075;
wire n37076;
wire n37077;
wire n37078;
wire n37079;
wire n37080;
wire n37081;
wire n37082;
wire n37083;
wire n37084;
wire n37085;
wire n37086;
wire n37087;
wire n37088;
wire n37089;
wire n37090;
wire n37091;
wire n37092;
wire n37093;
wire n37094;
wire n37095;
wire n37096;
wire n37097;
wire n37098;
wire n37099;
wire n37100;
wire n37101;
wire n37102;
wire n37103;
wire n37104;
wire n37105;
wire n37106;
wire n37107;
wire n37108;
wire n37109;
wire n37110;
wire n37111;
wire n37112;
wire n37113;
wire n37114;
wire n37115;
wire n37116;
wire n37117;
wire n37118;
wire n37119;
wire n3712;
wire n37120;
wire n37121;
wire n37122;
wire n37123;
wire n37124;
wire n37125;
wire n37126;
wire n37127;
wire n37128;
wire n37129;
wire n37131;
wire n37132;
wire n37133;
wire n37134;
wire n37135;
wire n37136;
wire n37137;
wire n37138;
wire n37139;
wire n37140;
wire n37141;
wire n37142;
wire n37143;
wire n37144;
wire n37145;
wire n37146;
wire n37147;
wire n37149;
wire n37150;
wire n37151;
wire n37152;
wire n37153;
wire n37154;
wire n37155;
wire n37156;
wire n37157;
wire n37158;
wire n37159;
wire n37160;
wire n37161;
wire n37162;
wire n37163;
wire n37164;
wire n37165;
wire n37166;
wire n37167;
wire n37168;
wire n37169;
wire n3717;
wire n37170;
wire n37171;
wire n37172;
wire n37173;
wire n37174;
wire n37175;
wire n37176;
wire n37177;
wire n37178;
wire n37179;
wire n37180;
wire n37181;
wire n37182;
wire n37183;
wire n37184;
wire n37185;
wire n37186;
wire n37187;
wire n37188;
wire n37189;
wire n37190;
wire n37191;
wire n37192;
wire n37193;
wire n37194;
wire n37195;
wire n37196;
wire n37197;
wire n37198;
wire n37199;
wire n37200;
wire n37201;
wire n37202;
wire n37203;
wire n37204;
wire n37205;
wire n37206;
wire n37207;
wire n37208;
wire n37209;
wire n37210;
wire n37211;
wire n37212;
wire n37213;
wire n37214;
wire n37215;
wire n37216;
wire n37217;
wire n37218;
wire n37219;
wire n3722;
wire n37220;
wire n37221;
wire n37222;
wire n37223;
wire n37224;
wire n37225;
wire n37226;
wire n37227;
wire n37228;
wire n37229;
wire n37230;
wire n37231;
wire n37232;
wire n37233;
wire n37234;
wire n37235;
wire n37236;
wire n37237;
wire n37238;
wire n37239;
wire n37240;
wire n37241;
wire n37242;
wire n37243;
wire n37244;
wire n37245;
wire n37246;
wire n37247;
wire n37248;
wire n37249;
wire n37250;
wire n37251;
wire n37252;
wire n37253;
wire n37254;
wire n37255;
wire n37256;
wire n37257;
wire n37258;
wire n37259;
wire n37260;
wire n37261;
wire n37262;
wire n37263;
wire n37264;
wire n37265;
wire n37266;
wire n37267;
wire n37268;
wire n37269;
wire n3727;
wire n37270;
wire n37271;
wire n37272;
wire n37273;
wire n37274;
wire n37275;
wire n37276;
wire n37277;
wire n37278;
wire n37279;
wire n37280;
wire n37281;
wire n37282;
wire n37283;
wire n37284;
wire n37285;
wire n37286;
wire n37287;
wire n37288;
wire n37289;
wire n37290;
wire n37291;
wire n37292;
wire n37293;
wire n37294;
wire n37295;
wire n37296;
wire n37297;
wire n37298;
wire n37299;
wire n373;
wire n37300;
wire n37301;
wire n37302;
wire n37303;
wire n37304;
wire n37305;
wire n37306;
wire n37307;
wire n37308;
wire n37309;
wire n37310;
wire n37312;
wire n37313;
wire n37314;
wire n37315;
wire n37316;
wire n37317;
wire n37318;
wire n37319;
wire n3732;
wire n37320;
wire n37321;
wire n37322;
wire n37323;
wire n37324;
wire n37325;
wire n37326;
wire n37327;
wire n37328;
wire n37329;
wire n37330;
wire n37331;
wire n37332;
wire n37333;
wire n37334;
wire n37335;
wire n37336;
wire n37337;
wire n37338;
wire n37339;
wire n37340;
wire n37341;
wire n37342;
wire n37343;
wire n37344;
wire n37345;
wire n37346;
wire n37347;
wire n37348;
wire n37349;
wire n37350;
wire n37351;
wire n37352;
wire n37353;
wire n37354;
wire n37355;
wire n37356;
wire n37357;
wire n37358;
wire n37359;
wire n37360;
wire n37361;
wire n37362;
wire n37363;
wire n37364;
wire n37365;
wire n37366;
wire n37367;
wire n37369;
wire n3737;
wire n37370;
wire n37371;
wire n37372;
wire n37373;
wire n37375;
wire n37376;
wire n37377;
wire n37378;
wire n37379;
wire n37380;
wire n37382;
wire n37383;
wire n37384;
wire n37385;
wire n37386;
wire n37387;
wire n37388;
wire n37389;
wire n37390;
wire n37391;
wire n37393;
wire n37394;
wire n37395;
wire n37396;
wire n37398;
wire n37399;
wire n37400;
wire n37402;
wire n37403;
wire n37404;
wire n37405;
wire n37406;
wire n37407;
wire n37408;
wire n37409;
wire n37410;
wire n37411;
wire n37412;
wire n37413;
wire n37414;
wire n37415;
wire n37416;
wire n37417;
wire n37418;
wire n37419;
wire n3742;
wire n37420;
wire n37421;
wire n37423;
wire n37425;
wire n37426;
wire n37427;
wire n37428;
wire n37429;
wire n37430;
wire n37431;
wire n37432;
wire n37433;
wire n37434;
wire n37435;
wire n37436;
wire n37437;
wire n37438;
wire n37439;
wire n37440;
wire n37441;
wire n37442;
wire n37443;
wire n37444;
wire n37445;
wire n37447;
wire n37448;
wire n37449;
wire n37450;
wire n37451;
wire n37452;
wire n37453;
wire n37454;
wire n37455;
wire n37456;
wire n37457;
wire n37458;
wire n37459;
wire n37460;
wire n37461;
wire n37462;
wire n37463;
wire n37464;
wire n37465;
wire n37466;
wire n37467;
wire n37468;
wire n37469;
wire n3747;
wire n37470;
wire n37471;
wire n37472;
wire n37473;
wire n37474;
wire n37475;
wire n37476;
wire n37477;
wire n37478;
wire n37479;
wire n37480;
wire n37481;
wire n37482;
wire n37483;
wire n37484;
wire n37485;
wire n37486;
wire n37487;
wire n37488;
wire n37489;
wire n37490;
wire n37491;
wire n37492;
wire n37493;
wire n37494;
wire n37495;
wire n37496;
wire n37497;
wire n37498;
wire n37499;
wire n37500;
wire n37501;
wire n37502;
wire n37503;
wire n37504;
wire n37505;
wire n37506;
wire n37507;
wire n37508;
wire n37509;
wire n37510;
wire n37511;
wire n37512;
wire n37513;
wire n37514;
wire n37515;
wire n37516;
wire n37517;
wire n37518;
wire n37519;
wire n3752;
wire n37520;
wire n37521;
wire n37522;
wire n37523;
wire n37524;
wire n37525;
wire n37526;
wire n37527;
wire n37528;
wire n37529;
wire n37530;
wire n37531;
wire n37532;
wire n37533;
wire n37534;
wire n37535;
wire n37536;
wire n37537;
wire n37538;
wire n37539;
wire n37540;
wire n37541;
wire n37542;
wire n37543;
wire n37544;
wire n37545;
wire n37546;
wire n37547;
wire n37548;
wire n37549;
wire n37550;
wire n37551;
wire n37552;
wire n37553;
wire n37554;
wire n37555;
wire n37556;
wire n37557;
wire n37558;
wire n37559;
wire n37560;
wire n37561;
wire n37562;
wire n37563;
wire n37564;
wire n37565;
wire n37566;
wire n37567;
wire n37568;
wire n37569;
wire n3757;
wire n37570;
wire n37571;
wire n37572;
wire n37573;
wire n37574;
wire n37575;
wire n37576;
wire n37577;
wire n37578;
wire n37579;
wire n37580;
wire n37581;
wire n37582;
wire n37583;
wire n37584;
wire n37585;
wire n37586;
wire n37587;
wire n37588;
wire n37589;
wire n37590;
wire n37591;
wire n37592;
wire n37593;
wire n37594;
wire n37595;
wire n37596;
wire n37597;
wire n37598;
wire n37599;
wire n37600;
wire n37601;
wire n37602;
wire n37603;
wire n37604;
wire n37605;
wire n37606;
wire n37607;
wire n37608;
wire n37609;
wire n37610;
wire n37611;
wire n37612;
wire n37613;
wire n37614;
wire n37615;
wire n37616;
wire n37617;
wire n37618;
wire n37619;
wire n3762;
wire n37620;
wire n37621;
wire n37622;
wire n37623;
wire n37624;
wire n37625;
wire n37626;
wire n37627;
wire n37628;
wire n37629;
wire n37630;
wire n37631;
wire n37632;
wire n37633;
wire n37634;
wire n37635;
wire n37636;
wire n37637;
wire n37638;
wire n37639;
wire n37640;
wire n37641;
wire n37642;
wire n37643;
wire n37644;
wire n37645;
wire n37646;
wire n37647;
wire n37648;
wire n37649;
wire n37650;
wire n37651;
wire n37652;
wire n37653;
wire n37654;
wire n37655;
wire n37656;
wire n37657;
wire n37658;
wire n37659;
wire n37660;
wire n37661;
wire n37662;
wire n37663;
wire n37664;
wire n37665;
wire n37666;
wire n37667;
wire n37669;
wire n3767;
wire n37670;
wire n37671;
wire n37672;
wire n37673;
wire n37674;
wire n37675;
wire n37676;
wire n37677;
wire n37678;
wire n37679;
wire n37680;
wire n37681;
wire n37682;
wire n37683;
wire n37684;
wire n37685;
wire n37686;
wire n37687;
wire n37688;
wire n37689;
wire n37690;
wire n37691;
wire n37692;
wire n37693;
wire n37694;
wire n37695;
wire n37696;
wire n37697;
wire n37698;
wire n37699;
wire n37700;
wire n37701;
wire n37702;
wire n37703;
wire n37704;
wire n37705;
wire n37706;
wire n37707;
wire n37708;
wire n37709;
wire n37710;
wire n37711;
wire n37712;
wire n37713;
wire n37714;
wire n37715;
wire n37716;
wire n37717;
wire n37718;
wire n37719;
wire n3772;
wire n37720;
wire n37721;
wire n37722;
wire n37723;
wire n37724;
wire n37725;
wire n37726;
wire n37727;
wire n37728;
wire n37729;
wire n37730;
wire n37731;
wire n37732;
wire n37733;
wire n37734;
wire n37735;
wire n37736;
wire n37737;
wire n37738;
wire n37739;
wire n37740;
wire n37741;
wire n37742;
wire n37743;
wire n37744;
wire n37745;
wire n37746;
wire n37747;
wire n37748;
wire n37749;
wire n37750;
wire n37751;
wire n37752;
wire n37753;
wire n37754;
wire n37755;
wire n37756;
wire n37757;
wire n37758;
wire n37759;
wire n37760;
wire n37761;
wire n37762;
wire n37763;
wire n37764;
wire n37765;
wire n37766;
wire n37767;
wire n37768;
wire n37769;
wire n3777;
wire n37770;
wire n37771;
wire n37772;
wire n37773;
wire n37774;
wire n37775;
wire n37776;
wire n37777;
wire n37778;
wire n37779;
wire n37780;
wire n37781;
wire n37782;
wire n37783;
wire n37784;
wire n37785;
wire n37786;
wire n37787;
wire n37788;
wire n37789;
wire n37790;
wire n37791;
wire n37792;
wire n37793;
wire n37794;
wire n37795;
wire n37797;
wire n37798;
wire n37799;
wire n378;
wire n37800;
wire n37801;
wire n37802;
wire n37803;
wire n37804;
wire n37805;
wire n37806;
wire n37807;
wire n37808;
wire n37809;
wire n37810;
wire n37812;
wire n37813;
wire n37814;
wire n37815;
wire n37816;
wire n37817;
wire n37818;
wire n37819;
wire n3782;
wire n37820;
wire n37821;
wire n37822;
wire n37823;
wire n37824;
wire n37825;
wire n37826;
wire n37827;
wire n37828;
wire n37829;
wire n37830;
wire n37831;
wire n37832;
wire n37833;
wire n37834;
wire n37835;
wire n37836;
wire n37837;
wire n37838;
wire n37839;
wire n37840;
wire n37841;
wire n37842;
wire n37843;
wire n37844;
wire n37845;
wire n37846;
wire n37847;
wire n37848;
wire n37849;
wire n37850;
wire n37851;
wire n37852;
wire n37853;
wire n37854;
wire n37855;
wire n37856;
wire n37857;
wire n37858;
wire n37859;
wire n37860;
wire n37861;
wire n37862;
wire n37863;
wire n37864;
wire n37865;
wire n37866;
wire n37867;
wire n37868;
wire n37869;
wire n3787;
wire n37870;
wire n37871;
wire n37872;
wire n37873;
wire n37874;
wire n37875;
wire n37876;
wire n37877;
wire n37878;
wire n37879;
wire n37880;
wire n37881;
wire n37882;
wire n37883;
wire n37884;
wire n37885;
wire n37886;
wire n37887;
wire n37888;
wire n37889;
wire n3789;
wire n37890;
wire n37891;
wire n37892;
wire n37893;
wire n37894;
wire n37895;
wire n37896;
wire n37897;
wire n37898;
wire n37899;
wire n3790;
wire n37900;
wire n37901;
wire n37902;
wire n37903;
wire n37904;
wire n37905;
wire n37906;
wire n37907;
wire n37908;
wire n37909;
wire n3791;
wire n37910;
wire n37911;
wire n37912;
wire n37913;
wire n37914;
wire n37915;
wire n37916;
wire n37917;
wire n37918;
wire n37919;
wire n3792;
wire n37920;
wire n37921;
wire n37922;
wire n37923;
wire n37924;
wire n37925;
wire n37926;
wire n37927;
wire n37928;
wire n37929;
wire n3792_1;
wire n3793;
wire n37930;
wire n37931;
wire n37932;
wire n37933;
wire n37934;
wire n37935;
wire n37936;
wire n37937;
wire n37938;
wire n37939;
wire n3794;
wire n37940;
wire n37941;
wire n37942;
wire n37943;
wire n37944;
wire n37945;
wire n37946;
wire n37947;
wire n37948;
wire n37949;
wire n3795;
wire n37950;
wire n37951;
wire n37952;
wire n37953;
wire n37954;
wire n37955;
wire n37956;
wire n37957;
wire n37958;
wire n37959;
wire n3796;
wire n37960;
wire n37961;
wire n37962;
wire n37963;
wire n37964;
wire n37965;
wire n37966;
wire n37967;
wire n37968;
wire n37969;
wire n3797;
wire n37970;
wire n37971;
wire n37972;
wire n37973;
wire n37974;
wire n37975;
wire n37976;
wire n37977;
wire n37978;
wire n37979;
wire n3797_1;
wire n3798;
wire n37980;
wire n37981;
wire n37982;
wire n37983;
wire n37984;
wire n37985;
wire n37986;
wire n37987;
wire n37988;
wire n37989;
wire n3799;
wire n37990;
wire n37991;
wire n37992;
wire n37993;
wire n37994;
wire n37995;
wire n37996;
wire n37997;
wire n37998;
wire n37999;
wire n3800;
wire n38000;
wire n38001;
wire n38002;
wire n38003;
wire n38004;
wire n38005;
wire n38006;
wire n38007;
wire n38008;
wire n38009;
wire n3801;
wire n38010;
wire n38011;
wire n38012;
wire n38013;
wire n38014;
wire n38015;
wire n38016;
wire n38017;
wire n38018;
wire n38019;
wire n3802;
wire n38020;
wire n38021;
wire n38022;
wire n38023;
wire n38024;
wire n38025;
wire n38026;
wire n38027;
wire n38028;
wire n38029;
wire n3802_1;
wire n3803;
wire n38030;
wire n38031;
wire n38032;
wire n38033;
wire n38034;
wire n38035;
wire n38036;
wire n38037;
wire n38038;
wire n38039;
wire n3804;
wire n38040;
wire n38041;
wire n38042;
wire n38043;
wire n38044;
wire n38045;
wire n38046;
wire n38047;
wire n38048;
wire n38049;
wire n3805;
wire n38050;
wire n38051;
wire n38052;
wire n38054;
wire n38056;
wire n38057;
wire n38058;
wire n38059;
wire n3806;
wire n38060;
wire n38061;
wire n38062;
wire n38063;
wire n38064;
wire n38065;
wire n38066;
wire n38067;
wire n38068;
wire n38069;
wire n3806_1;
wire n3807;
wire n38070;
wire n38071;
wire n38072;
wire n38073;
wire n38074;
wire n38076;
wire n38077;
wire n38078;
wire n38079;
wire n3808;
wire n38080;
wire n38081;
wire n38082;
wire n38083;
wire n38085;
wire n38086;
wire n38087;
wire n38088;
wire n38089;
wire n3809;
wire n38090;
wire n38091;
wire n38092;
wire n38093;
wire n38094;
wire n38095;
wire n38096;
wire n38097;
wire n38098;
wire n38099;
wire n3810;
wire n38100;
wire n38101;
wire n38102;
wire n38103;
wire n38104;
wire n38105;
wire n38106;
wire n38107;
wire n38108;
wire n38109;
wire n3811;
wire n38110;
wire n38111;
wire n38112;
wire n38113;
wire n38114;
wire n38115;
wire n38116;
wire n38117;
wire n38118;
wire n38119;
wire n3811_1;
wire n3812;
wire n38120;
wire n38121;
wire n38122;
wire n38123;
wire n38124;
wire n38125;
wire n38126;
wire n38127;
wire n38128;
wire n38129;
wire n3813;
wire n38130;
wire n38131;
wire n38132;
wire n38133;
wire n38134;
wire n38135;
wire n38136;
wire n38137;
wire n38138;
wire n38139;
wire n3814;
wire n38140;
wire n38141;
wire n38142;
wire n38143;
wire n38144;
wire n38145;
wire n38146;
wire n38147;
wire n38148;
wire n38149;
wire n3815;
wire n38150;
wire n38151;
wire n38152;
wire n38153;
wire n38154;
wire n38155;
wire n38156;
wire n38157;
wire n38158;
wire n38159;
wire n3816;
wire n38160;
wire n38161;
wire n38162;
wire n38163;
wire n38164;
wire n38166;
wire n38167;
wire n38168;
wire n38169;
wire n3816_1;
wire n3817;
wire n38170;
wire n38171;
wire n38172;
wire n38173;
wire n38175;
wire n38176;
wire n38177;
wire n38178;
wire n38179;
wire n3818;
wire n38180;
wire n38181;
wire n38182;
wire n38183;
wire n38185;
wire n38186;
wire n38187;
wire n38188;
wire n38189;
wire n3819;
wire n38190;
wire n38191;
wire n38193;
wire n38194;
wire n38195;
wire n38196;
wire n38197;
wire n38198;
wire n38199;
wire n3820;
wire n38200;
wire n38201;
wire n38202;
wire n38203;
wire n38204;
wire n38205;
wire n38206;
wire n38207;
wire n38208;
wire n38209;
wire n3821;
wire n38211;
wire n38212;
wire n38213;
wire n38214;
wire n38215;
wire n38216;
wire n38217;
wire n38218;
wire n38219;
wire n3821_1;
wire n3822;
wire n38220;
wire n38221;
wire n38222;
wire n38223;
wire n38224;
wire n38225;
wire n38226;
wire n38227;
wire n38228;
wire n38229;
wire n3823;
wire n38230;
wire n38231;
wire n38232;
wire n38233;
wire n38234;
wire n38235;
wire n38236;
wire n38237;
wire n38238;
wire n38239;
wire n3824;
wire n38240;
wire n38241;
wire n38242;
wire n38243;
wire n38244;
wire n38245;
wire n38246;
wire n38247;
wire n38248;
wire n38249;
wire n3825;
wire n38250;
wire n38251;
wire n38252;
wire n38253;
wire n38254;
wire n38255;
wire n38256;
wire n38257;
wire n38258;
wire n38259;
wire n3826;
wire n38260;
wire n38261;
wire n38262;
wire n38263;
wire n38264;
wire n38265;
wire n38266;
wire n38267;
wire n38268;
wire n38269;
wire n3826_1;
wire n3827;
wire n38270;
wire n38271;
wire n38272;
wire n38273;
wire n38274;
wire n38275;
wire n38276;
wire n38277;
wire n38278;
wire n38279;
wire n3828;
wire n38280;
wire n38281;
wire n38282;
wire n38283;
wire n38284;
wire n38285;
wire n38286;
wire n38287;
wire n38288;
wire n38289;
wire n3829;
wire n38290;
wire n38291;
wire n38292;
wire n38293;
wire n38294;
wire n38295;
wire n38296;
wire n38297;
wire n38298;
wire n38299;
wire n383;
wire n3830;
wire n38300;
wire n38301;
wire n38302;
wire n38303;
wire n38304;
wire n38305;
wire n38306;
wire n38307;
wire n38308;
wire n38309;
wire n3831;
wire n38310;
wire n38311;
wire n38312;
wire n38313;
wire n38314;
wire n38315;
wire n38316;
wire n38317;
wire n38318;
wire n38319;
wire n3831_1;
wire n3832;
wire n38320;
wire n38321;
wire n38322;
wire n38323;
wire n38324;
wire n38325;
wire n38326;
wire n38327;
wire n38328;
wire n38329;
wire n3833;
wire n38330;
wire n38331;
wire n38332;
wire n38333;
wire n38334;
wire n38335;
wire n38336;
wire n38337;
wire n38338;
wire n38339;
wire n3834;
wire n38340;
wire n38341;
wire n38342;
wire n38343;
wire n38344;
wire n38345;
wire n38346;
wire n38347;
wire n38348;
wire n38349;
wire n3835;
wire n38350;
wire n38351;
wire n38352;
wire n38353;
wire n38354;
wire n38355;
wire n38356;
wire n38357;
wire n38358;
wire n38359;
wire n3836;
wire n38360;
wire n38361;
wire n38362;
wire n38363;
wire n38364;
wire n38365;
wire n38366;
wire n38367;
wire n38368;
wire n38369;
wire n3836_1;
wire n3837;
wire n38370;
wire n38371;
wire n38372;
wire n38373;
wire n38374;
wire n38375;
wire n38376;
wire n38377;
wire n38378;
wire n38379;
wire n3838;
wire n38380;
wire n38381;
wire n38382;
wire n38383;
wire n38384;
wire n38385;
wire n38386;
wire n38387;
wire n38388;
wire n38389;
wire n3839;
wire n38390;
wire n38391;
wire n38392;
wire n38393;
wire n38394;
wire n38395;
wire n38396;
wire n38397;
wire n38398;
wire n38399;
wire n3840;
wire n38400;
wire n38401;
wire n38402;
wire n38403;
wire n38404;
wire n38405;
wire n38406;
wire n38407;
wire n38408;
wire n38409;
wire n3841;
wire n38410;
wire n38411;
wire n38412;
wire n38413;
wire n38414;
wire n38415;
wire n38416;
wire n38417;
wire n38418;
wire n38419;
wire n3841_1;
wire n3842;
wire n38420;
wire n38421;
wire n38422;
wire n38423;
wire n38424;
wire n38425;
wire n38426;
wire n38427;
wire n38428;
wire n38429;
wire n3843;
wire n38430;
wire n38431;
wire n38432;
wire n38433;
wire n38434;
wire n38435;
wire n38436;
wire n38437;
wire n38438;
wire n38439;
wire n3844;
wire n38440;
wire n38441;
wire n38442;
wire n38443;
wire n38444;
wire n38445;
wire n38446;
wire n38447;
wire n38448;
wire n38449;
wire n3845;
wire n38450;
wire n38451;
wire n38452;
wire n38453;
wire n38454;
wire n38455;
wire n38456;
wire n38457;
wire n38458;
wire n38459;
wire n3846;
wire n38460;
wire n38461;
wire n38462;
wire n38463;
wire n38464;
wire n38465;
wire n38466;
wire n38467;
wire n38468;
wire n38469;
wire n3846_1;
wire n3847;
wire n38470;
wire n38471;
wire n38472;
wire n38473;
wire n38474;
wire n38475;
wire n38476;
wire n38477;
wire n38478;
wire n38479;
wire n3848;
wire n38480;
wire n38481;
wire n38482;
wire n38483;
wire n38484;
wire n38485;
wire n38486;
wire n38487;
wire n38488;
wire n38489;
wire n3849;
wire n38490;
wire n38491;
wire n38492;
wire n38493;
wire n38494;
wire n38495;
wire n38496;
wire n38497;
wire n38498;
wire n38499;
wire n3850;
wire n38500;
wire n38501;
wire n38502;
wire n38503;
wire n38504;
wire n38505;
wire n38506;
wire n38507;
wire n38508;
wire n38509;
wire n3850_1;
wire n3851;
wire n38510;
wire n38511;
wire n38512;
wire n38513;
wire n38514;
wire n38515;
wire n38516;
wire n38517;
wire n38518;
wire n38519;
wire n3852;
wire n38520;
wire n38521;
wire n38522;
wire n38523;
wire n38524;
wire n38525;
wire n38526;
wire n38527;
wire n38528;
wire n38529;
wire n3853;
wire n38530;
wire n38531;
wire n38532;
wire n38533;
wire n38534;
wire n38535;
wire n38536;
wire n38537;
wire n38538;
wire n38539;
wire n3854;
wire n38540;
wire n38541;
wire n38542;
wire n38543;
wire n38544;
wire n38545;
wire n38547;
wire n38548;
wire n38549;
wire n3855;
wire n38550;
wire n38551;
wire n38552;
wire n38553;
wire n38554;
wire n38555;
wire n38556;
wire n38557;
wire n38558;
wire n38559;
wire n3855_1;
wire n3856;
wire n38560;
wire n38561;
wire n38562;
wire n38563;
wire n38564;
wire n38566;
wire n38567;
wire n38569;
wire n3857;
wire n38570;
wire n38571;
wire n38572;
wire n38573;
wire n38574;
wire n38575;
wire n38578;
wire n38579;
wire n3858;
wire n38580;
wire n38581;
wire n38582;
wire n38583;
wire n38584;
wire n38585;
wire n38586;
wire n38587;
wire n38589;
wire n3859;
wire n38591;
wire n38592;
wire n38593;
wire n38594;
wire n38595;
wire n38596;
wire n38597;
wire n38598;
wire n38599;
wire n3860;
wire n38600;
wire n38601;
wire n38602;
wire n38603;
wire n38604;
wire n38605;
wire n38606;
wire n38607;
wire n38608;
wire n38609;
wire n3860_1;
wire n3861;
wire n38610;
wire n38611;
wire n38612;
wire n38613;
wire n38614;
wire n38615;
wire n38616;
wire n38617;
wire n38618;
wire n38619;
wire n3862;
wire n38620;
wire n38621;
wire n38622;
wire n38623;
wire n38624;
wire n38625;
wire n38626;
wire n38627;
wire n38628;
wire n38629;
wire n3863;
wire n38630;
wire n38631;
wire n38632;
wire n38633;
wire n38635;
wire n38636;
wire n38637;
wire n38638;
wire n38639;
wire n3864;
wire n38640;
wire n38641;
wire n38642;
wire n38643;
wire n38644;
wire n38645;
wire n38647;
wire n38648;
wire n38649;
wire n3865;
wire n38650;
wire n38651;
wire n38653;
wire n38654;
wire n38655;
wire n38656;
wire n38657;
wire n38658;
wire n38659;
wire n3865_1;
wire n3866;
wire n38660;
wire n38662;
wire n38663;
wire n38664;
wire n38665;
wire n38666;
wire n38667;
wire n38668;
wire n38669;
wire n3867;
wire n38670;
wire n38671;
wire n38672;
wire n38674;
wire n38675;
wire n38676;
wire n38677;
wire n38678;
wire n38679;
wire n3868;
wire n38680;
wire n38681;
wire n38682;
wire n38683;
wire n38684;
wire n38685;
wire n38686;
wire n38687;
wire n38688;
wire n38689;
wire n3869;
wire n38690;
wire n38691;
wire n38692;
wire n38693;
wire n38694;
wire n38695;
wire n38696;
wire n38697;
wire n38698;
wire n38699;
wire n3870;
wire n38700;
wire n38701;
wire n38702;
wire n38703;
wire n38704;
wire n38705;
wire n38706;
wire n38707;
wire n38708;
wire n38709;
wire n3870_1;
wire n3871;
wire n38710;
wire n38711;
wire n38712;
wire n38713;
wire n38714;
wire n38715;
wire n38716;
wire n38717;
wire n38718;
wire n38719;
wire n3872;
wire n38720;
wire n38721;
wire n38722;
wire n38723;
wire n38724;
wire n38725;
wire n38726;
wire n38727;
wire n38728;
wire n38729;
wire n3873;
wire n38730;
wire n38731;
wire n38732;
wire n38733;
wire n38734;
wire n38735;
wire n38736;
wire n38737;
wire n38738;
wire n38739;
wire n3874;
wire n38740;
wire n38741;
wire n38742;
wire n38743;
wire n38744;
wire n38745;
wire n38746;
wire n38747;
wire n38748;
wire n38749;
wire n3875;
wire n38750;
wire n38751;
wire n38752;
wire n38753;
wire n38754;
wire n38756;
wire n38757;
wire n38758;
wire n38759;
wire n3875_1;
wire n3876;
wire n38760;
wire n38761;
wire n38762;
wire n38763;
wire n38764;
wire n38765;
wire n38766;
wire n38767;
wire n38768;
wire n38769;
wire n3877;
wire n38770;
wire n38771;
wire n38772;
wire n38773;
wire n38774;
wire n38775;
wire n38776;
wire n38777;
wire n38778;
wire n38779;
wire n3878;
wire n38780;
wire n38781;
wire n38782;
wire n38783;
wire n38784;
wire n38785;
wire n38786;
wire n38787;
wire n38788;
wire n38789;
wire n3879;
wire n38790;
wire n38791;
wire n38792;
wire n38793;
wire n38794;
wire n38795;
wire n38796;
wire n38797;
wire n38798;
wire n38799;
wire n388;
wire n3880;
wire n38800;
wire n38801;
wire n38802;
wire n38803;
wire n38804;
wire n38805;
wire n38806;
wire n38807;
wire n38808;
wire n38809;
wire n3880_1;
wire n3881;
wire n38810;
wire n38811;
wire n38812;
wire n38813;
wire n38814;
wire n38815;
wire n38816;
wire n38817;
wire n38818;
wire n38819;
wire n3882;
wire n38820;
wire n38821;
wire n38822;
wire n38823;
wire n38824;
wire n38825;
wire n38826;
wire n38827;
wire n38828;
wire n38829;
wire n3883;
wire n38830;
wire n38831;
wire n38832;
wire n38833;
wire n38834;
wire n38835;
wire n38836;
wire n38837;
wire n38838;
wire n38839;
wire n3884;
wire n38840;
wire n38841;
wire n38842;
wire n38843;
wire n38844;
wire n38845;
wire n38846;
wire n38847;
wire n38848;
wire n38849;
wire n3885;
wire n38850;
wire n38851;
wire n38852;
wire n38853;
wire n38854;
wire n38855;
wire n38856;
wire n38858;
wire n3885_1;
wire n3886;
wire n38860;
wire n38861;
wire n38862;
wire n38863;
wire n38864;
wire n38865;
wire n38866;
wire n38868;
wire n38869;
wire n3887;
wire n38870;
wire n38871;
wire n38873;
wire n38874;
wire n38875;
wire n38876;
wire n38877;
wire n38879;
wire n3888;
wire n38880;
wire n38881;
wire n38882;
wire n38883;
wire n38884;
wire n38885;
wire n38886;
wire n38887;
wire n38888;
wire n38889;
wire n3889;
wire n38890;
wire n38891;
wire n38892;
wire n38893;
wire n38894;
wire n38895;
wire n38896;
wire n38897;
wire n38898;
wire n38899;
wire n3890;
wire n38900;
wire n38901;
wire n38902;
wire n38903;
wire n38904;
wire n38905;
wire n38906;
wire n38907;
wire n38908;
wire n38909;
wire n3890_1;
wire n3891;
wire n38910;
wire n38911;
wire n38912;
wire n38913;
wire n38914;
wire n38915;
wire n38916;
wire n38917;
wire n38918;
wire n38919;
wire n3892;
wire n38920;
wire n38921;
wire n38922;
wire n38923;
wire n38924;
wire n38925;
wire n38926;
wire n38927;
wire n38928;
wire n38929;
wire n3893;
wire n38930;
wire n38931;
wire n38932;
wire n38933;
wire n38934;
wire n38935;
wire n38936;
wire n38937;
wire n38938;
wire n38939;
wire n3894;
wire n38940;
wire n38941;
wire n38942;
wire n38943;
wire n38944;
wire n38945;
wire n38946;
wire n38947;
wire n38948;
wire n38949;
wire n3895;
wire n38950;
wire n38951;
wire n38952;
wire n38953;
wire n38954;
wire n38955;
wire n38956;
wire n38957;
wire n38958;
wire n38959;
wire n3895_1;
wire n3896;
wire n38960;
wire n38961;
wire n38962;
wire n38965;
wire n38967;
wire n38969;
wire n3897;
wire n38970;
wire n38972;
wire n38973;
wire n38974;
wire n38975;
wire n38976;
wire n38977;
wire n38979;
wire n3898;
wire n38980;
wire n38981;
wire n38982;
wire n38983;
wire n38984;
wire n38985;
wire n38986;
wire n38987;
wire n38988;
wire n3899;
wire n38990;
wire n38991;
wire n38992;
wire n38993;
wire n38995;
wire n38997;
wire n38998;
wire n38999;
wire n3900;
wire n39000;
wire n39001;
wire n39002;
wire n39003;
wire n39004;
wire n39005;
wire n39007;
wire n39008;
wire n39009;
wire n3900_1;
wire n3901;
wire n39010;
wire n39011;
wire n39012;
wire n39013;
wire n39014;
wire n39016;
wire n39017;
wire n39018;
wire n39019;
wire n3902;
wire n39020;
wire n39021;
wire n39022;
wire n39023;
wire n39024;
wire n39026;
wire n39028;
wire n39029;
wire n3903;
wire n39030;
wire n39031;
wire n39032;
wire n39033;
wire n39034;
wire n39035;
wire n39036;
wire n39037;
wire n39039;
wire n3904;
wire n39040;
wire n39042;
wire n39043;
wire n39044;
wire n39045;
wire n39046;
wire n39047;
wire n39048;
wire n39049;
wire n3905;
wire n39050;
wire n39052;
wire n39053;
wire n39054;
wire n39055;
wire n39056;
wire n39057;
wire n39058;
wire n39059;
wire n3905_1;
wire n3906;
wire n39060;
wire n39061;
wire n39062;
wire n39063;
wire n39064;
wire n39065;
wire n39066;
wire n39067;
wire n39068;
wire n39069;
wire n3907;
wire n39070;
wire n39071;
wire n39072;
wire n39073;
wire n39074;
wire n39075;
wire n39076;
wire n39077;
wire n39078;
wire n39079;
wire n3908;
wire n39080;
wire n39081;
wire n39082;
wire n39083;
wire n39084;
wire n39085;
wire n39086;
wire n39087;
wire n39088;
wire n39089;
wire n3909;
wire n39090;
wire n39091;
wire n39092;
wire n39093;
wire n39094;
wire n39095;
wire n39096;
wire n39097;
wire n39098;
wire n39099;
wire n3910;
wire n39100;
wire n39101;
wire n39102;
wire n39103;
wire n39104;
wire n39105;
wire n39106;
wire n39107;
wire n39108;
wire n39109;
wire n3910_1;
wire n3911;
wire n39110;
wire n39111;
wire n39112;
wire n39113;
wire n39114;
wire n39115;
wire n39116;
wire n39117;
wire n39118;
wire n39119;
wire n3912;
wire n39120;
wire n39121;
wire n39122;
wire n39123;
wire n39124;
wire n39125;
wire n39126;
wire n39127;
wire n39128;
wire n39129;
wire n3913;
wire n39130;
wire n39131;
wire n39132;
wire n39133;
wire n39134;
wire n39135;
wire n39136;
wire n39137;
wire n39138;
wire n39139;
wire n3914;
wire n39140;
wire n39141;
wire n39142;
wire n39143;
wire n39144;
wire n39145;
wire n39146;
wire n39147;
wire n39148;
wire n39149;
wire n3915;
wire n39150;
wire n39151;
wire n39152;
wire n39153;
wire n39154;
wire n39155;
wire n39156;
wire n39157;
wire n39158;
wire n39159;
wire n3915_1;
wire n3916;
wire n39160;
wire n39161;
wire n39162;
wire n39163;
wire n39164;
wire n39165;
wire n39166;
wire n39167;
wire n39168;
wire n39169;
wire n3917;
wire n39170;
wire n39171;
wire n39172;
wire n39173;
wire n39174;
wire n39175;
wire n39177;
wire n39178;
wire n39179;
wire n3918;
wire n39180;
wire n39181;
wire n39182;
wire n39183;
wire n39184;
wire n39185;
wire n39186;
wire n39187;
wire n39189;
wire n3919;
wire n39190;
wire n39191;
wire n39192;
wire n39193;
wire n39194;
wire n39195;
wire n39196;
wire n39197;
wire n39198;
wire n39199;
wire n3920;
wire n39200;
wire n39201;
wire n39202;
wire n39203;
wire n39204;
wire n39205;
wire n39207;
wire n39208;
wire n39209;
wire n3920_1;
wire n3921;
wire n39210;
wire n39211;
wire n39212;
wire n39213;
wire n39214;
wire n39215;
wire n39216;
wire n39217;
wire n39218;
wire n3922;
wire n39220;
wire n39221;
wire n39222;
wire n39223;
wire n39224;
wire n39225;
wire n39226;
wire n39227;
wire n39228;
wire n39229;
wire n3923;
wire n39230;
wire n39231;
wire n39232;
wire n39233;
wire n39234;
wire n39235;
wire n39236;
wire n39237;
wire n39238;
wire n39239;
wire n3924;
wire n39240;
wire n39241;
wire n39242;
wire n39243;
wire n39244;
wire n39245;
wire n39246;
wire n39247;
wire n39248;
wire n39249;
wire n3925;
wire n39250;
wire n39251;
wire n39252;
wire n39253;
wire n39254;
wire n39255;
wire n39256;
wire n39257;
wire n39258;
wire n39259;
wire n3925_1;
wire n3926;
wire n39260;
wire n39261;
wire n39262;
wire n39263;
wire n39264;
wire n39265;
wire n39266;
wire n39267;
wire n39268;
wire n39269;
wire n3927;
wire n39270;
wire n39271;
wire n39272;
wire n39273;
wire n39274;
wire n39275;
wire n39276;
wire n39277;
wire n39278;
wire n39279;
wire n3928;
wire n39280;
wire n39281;
wire n39282;
wire n39283;
wire n39284;
wire n39285;
wire n39286;
wire n39287;
wire n39288;
wire n39289;
wire n3929;
wire n39290;
wire n39291;
wire n39292;
wire n39293;
wire n39294;
wire n39295;
wire n39296;
wire n39297;
wire n39298;
wire n39299;
wire n393;
wire n3930;
wire n39300;
wire n39301;
wire n39302;
wire n39303;
wire n39304;
wire n39305;
wire n39306;
wire n39307;
wire n39308;
wire n39309;
wire n3930_1;
wire n3931;
wire n39310;
wire n39311;
wire n39312;
wire n39313;
wire n39314;
wire n39315;
wire n39316;
wire n39317;
wire n39318;
wire n39319;
wire n3932;
wire n39320;
wire n39321;
wire n39322;
wire n39323;
wire n39324;
wire n39325;
wire n39326;
wire n39327;
wire n39328;
wire n39329;
wire n3933;
wire n39330;
wire n39331;
wire n39332;
wire n39333;
wire n39334;
wire n39335;
wire n39336;
wire n39337;
wire n39338;
wire n39339;
wire n3934;
wire n39340;
wire n39341;
wire n39342;
wire n39343;
wire n39344;
wire n39345;
wire n39346;
wire n39347;
wire n39348;
wire n39349;
wire n3935;
wire n39350;
wire n39351;
wire n39352;
wire n39353;
wire n39354;
wire n39355;
wire n39356;
wire n39357;
wire n39358;
wire n39359;
wire n3935_1;
wire n3936;
wire n39360;
wire n39361;
wire n39362;
wire n39363;
wire n39364;
wire n39365;
wire n39366;
wire n39367;
wire n39368;
wire n39369;
wire n3937;
wire n39370;
wire n39371;
wire n39372;
wire n39373;
wire n39374;
wire n39375;
wire n39376;
wire n39377;
wire n39378;
wire n39379;
wire n3938;
wire n39380;
wire n39381;
wire n39382;
wire n39383;
wire n39384;
wire n39385;
wire n39386;
wire n39387;
wire n39388;
wire n39389;
wire n3939;
wire n39390;
wire n39391;
wire n39392;
wire n39393;
wire n39394;
wire n39395;
wire n39396;
wire n39397;
wire n39398;
wire n39399;
wire n3940;
wire n39400;
wire n39401;
wire n39402;
wire n39403;
wire n39404;
wire n39405;
wire n39406;
wire n39407;
wire n39408;
wire n39409;
wire n3940_1;
wire n3941;
wire n39410;
wire n39411;
wire n39412;
wire n39413;
wire n39414;
wire n39415;
wire n39416;
wire n39417;
wire n39418;
wire n39419;
wire n3942;
wire n39420;
wire n39421;
wire n39422;
wire n39423;
wire n39424;
wire n39425;
wire n39426;
wire n39427;
wire n39428;
wire n39429;
wire n3943;
wire n39430;
wire n39431;
wire n39432;
wire n39433;
wire n39434;
wire n39435;
wire n39436;
wire n39437;
wire n39438;
wire n39439;
wire n3944;
wire n39440;
wire n39441;
wire n39442;
wire n39443;
wire n39444;
wire n39445;
wire n39446;
wire n39447;
wire n39448;
wire n39449;
wire n3945;
wire n39450;
wire n39451;
wire n39452;
wire n39453;
wire n39454;
wire n39455;
wire n39456;
wire n39457;
wire n39458;
wire n39459;
wire n3945_1;
wire n3946;
wire n39460;
wire n39461;
wire n39462;
wire n39463;
wire n39464;
wire n39465;
wire n39466;
wire n39467;
wire n39468;
wire n39469;
wire n3947;
wire n39470;
wire n39471;
wire n39472;
wire n39473;
wire n39474;
wire n39475;
wire n39476;
wire n39477;
wire n39478;
wire n39479;
wire n3948;
wire n39480;
wire n39481;
wire n39482;
wire n39483;
wire n39484;
wire n39485;
wire n39487;
wire n39488;
wire n39489;
wire n3949;
wire n39490;
wire n39491;
wire n39493;
wire n39494;
wire n39495;
wire n39496;
wire n39497;
wire n39498;
wire n39499;
wire n3950;
wire n39500;
wire n39501;
wire n39502;
wire n39503;
wire n39504;
wire n39505;
wire n39506;
wire n39507;
wire n39508;
wire n39509;
wire n3950_1;
wire n3951;
wire n39510;
wire n39511;
wire n39512;
wire n39513;
wire n39514;
wire n39515;
wire n39516;
wire n39517;
wire n39518;
wire n3952;
wire n39520;
wire n39521;
wire n39522;
wire n39523;
wire n39524;
wire n39525;
wire n39526;
wire n39527;
wire n39528;
wire n39529;
wire n3953;
wire n39530;
wire n39532;
wire n39534;
wire n39535;
wire n39536;
wire n39537;
wire n39538;
wire n39539;
wire n3954;
wire n39540;
wire n39542;
wire n39543;
wire n39545;
wire n39546;
wire n39547;
wire n39548;
wire n39549;
wire n3955;
wire n39550;
wire n39551;
wire n39552;
wire n39553;
wire n39554;
wire n39555;
wire n39556;
wire n39557;
wire n39558;
wire n39559;
wire n3955_1;
wire n3956;
wire n39560;
wire n39561;
wire n39562;
wire n39563;
wire n39564;
wire n39565;
wire n39566;
wire n39567;
wire n39568;
wire n39569;
wire n3957;
wire n39570;
wire n39571;
wire n39572;
wire n39573;
wire n39574;
wire n39575;
wire n39576;
wire n39577;
wire n39578;
wire n39579;
wire n3958;
wire n39580;
wire n39581;
wire n39582;
wire n39583;
wire n39584;
wire n39585;
wire n39586;
wire n39587;
wire n39588;
wire n39589;
wire n3959;
wire n39590;
wire n39591;
wire n39592;
wire n39593;
wire n39594;
wire n39595;
wire n39596;
wire n39597;
wire n39598;
wire n39599;
wire n3960;
wire n39600;
wire n39601;
wire n39602;
wire n39603;
wire n39604;
wire n39605;
wire n39606;
wire n39607;
wire n39608;
wire n39609;
wire n3960_1;
wire n3961;
wire n39610;
wire n39611;
wire n39612;
wire n39613;
wire n39614;
wire n39615;
wire n39616;
wire n39617;
wire n39618;
wire n39619;
wire n3962;
wire n39621;
wire n39622;
wire n39623;
wire n39624;
wire n39625;
wire n39626;
wire n39627;
wire n39628;
wire n39629;
wire n3963;
wire n39630;
wire n39631;
wire n39632;
wire n39633;
wire n39634;
wire n39636;
wire n39639;
wire n3964;
wire n39640;
wire n39642;
wire n39643;
wire n39644;
wire n39645;
wire n39646;
wire n39647;
wire n39648;
wire n39649;
wire n3965;
wire n39650;
wire n39651;
wire n39652;
wire n39653;
wire n39654;
wire n39655;
wire n39656;
wire n39658;
wire n39659;
wire n3965_1;
wire n3966;
wire n39660;
wire n39661;
wire n39662;
wire n39663;
wire n39664;
wire n39665;
wire n39666;
wire n39667;
wire n39668;
wire n39669;
wire n3967;
wire n39670;
wire n39671;
wire n39672;
wire n39673;
wire n39674;
wire n39675;
wire n39676;
wire n39677;
wire n39678;
wire n39679;
wire n3968;
wire n39680;
wire n39681;
wire n39682;
wire n39683;
wire n39684;
wire n39685;
wire n39686;
wire n39687;
wire n39688;
wire n39689;
wire n3969;
wire n39690;
wire n39691;
wire n39692;
wire n39693;
wire n39694;
wire n39695;
wire n39696;
wire n39697;
wire n39698;
wire n39699;
wire n3970;
wire n39700;
wire n39701;
wire n39702;
wire n39703;
wire n39704;
wire n39705;
wire n39706;
wire n39707;
wire n39708;
wire n39709;
wire n3970_1;
wire n3971;
wire n39710;
wire n39711;
wire n39712;
wire n39713;
wire n39714;
wire n39716;
wire n39717;
wire n39718;
wire n3972;
wire n39720;
wire n39721;
wire n39722;
wire n39723;
wire n39724;
wire n39725;
wire n39727;
wire n39728;
wire n39729;
wire n3973;
wire n39730;
wire n39731;
wire n39733;
wire n39734;
wire n39735;
wire n39737;
wire n39738;
wire n39739;
wire n3974;
wire n39740;
wire n39742;
wire n39743;
wire n39744;
wire n39745;
wire n39746;
wire n39747;
wire n39748;
wire n39749;
wire n3975;
wire n39750;
wire n39751;
wire n39752;
wire n39754;
wire n39755;
wire n39756;
wire n39757;
wire n39758;
wire n3975_1;
wire n3976;
wire n39760;
wire n39762;
wire n39763;
wire n39764;
wire n39765;
wire n39766;
wire n39768;
wire n3977;
wire n39770;
wire n39771;
wire n39772;
wire n39773;
wire n39774;
wire n39775;
wire n39776;
wire n39777;
wire n39779;
wire n3978;
wire n39780;
wire n39782;
wire n39783;
wire n39784;
wire n39785;
wire n39786;
wire n39787;
wire n39788;
wire n39789;
wire n3979;
wire n39790;
wire n39791;
wire n39792;
wire n39794;
wire n39795;
wire n39796;
wire n39797;
wire n39798;
wire n398;
wire n3980;
wire n39800;
wire n39801;
wire n39802;
wire n39803;
wire n39804;
wire n39805;
wire n39806;
wire n39807;
wire n39808;
wire n39809;
wire n3980_1;
wire n3981;
wire n39810;
wire n39811;
wire n39813;
wire n39814;
wire n39815;
wire n39816;
wire n39817;
wire n39818;
wire n39819;
wire n3982;
wire n39820;
wire n39821;
wire n39822;
wire n39823;
wire n39825;
wire n39826;
wire n39827;
wire n39828;
wire n3983;
wire n39830;
wire n39831;
wire n39832;
wire n39833;
wire n39834;
wire n39835;
wire n39836;
wire n39837;
wire n39839;
wire n3984;
wire n39840;
wire n39841;
wire n39842;
wire n39843;
wire n39844;
wire n39845;
wire n39846;
wire n39847;
wire n39848;
wire n39849;
wire n3985;
wire n39850;
wire n39851;
wire n39852;
wire n39853;
wire n39854;
wire n39855;
wire n39856;
wire n39857;
wire n39858;
wire n39859;
wire n3985_1;
wire n3986;
wire n39860;
wire n39861;
wire n39862;
wire n39863;
wire n39864;
wire n39865;
wire n39866;
wire n39867;
wire n39868;
wire n39869;
wire n3987;
wire n39870;
wire n39871;
wire n39872;
wire n39873;
wire n39874;
wire n39875;
wire n39876;
wire n39877;
wire n39878;
wire n39879;
wire n3988;
wire n39880;
wire n39881;
wire n39882;
wire n39883;
wire n39884;
wire n39885;
wire n39886;
wire n39887;
wire n39888;
wire n39889;
wire n3989;
wire n39890;
wire n39891;
wire n39892;
wire n39893;
wire n39894;
wire n39895;
wire n39896;
wire n39897;
wire n39898;
wire n39899;
wire n3990;
wire n39900;
wire n39901;
wire n39902;
wire n39903;
wire n39904;
wire n39905;
wire n39906;
wire n39907;
wire n39908;
wire n39909;
wire n3990_1;
wire n3991;
wire n39910;
wire n39911;
wire n39912;
wire n39913;
wire n39914;
wire n39915;
wire n39916;
wire n39917;
wire n39918;
wire n39919;
wire n3992;
wire n39920;
wire n39921;
wire n39922;
wire n39923;
wire n39924;
wire n39925;
wire n39926;
wire n39927;
wire n39928;
wire n39929;
wire n3993;
wire n39930;
wire n39931;
wire n39932;
wire n39933;
wire n39934;
wire n39935;
wire n39936;
wire n39937;
wire n39938;
wire n39939;
wire n3994;
wire n39940;
wire n39941;
wire n39942;
wire n39943;
wire n39944;
wire n39945;
wire n39946;
wire n39947;
wire n39948;
wire n39949;
wire n3994_1;
wire n3995;
wire n39950;
wire n39951;
wire n39952;
wire n39953;
wire n39954;
wire n39955;
wire n39956;
wire n39957;
wire n39958;
wire n39959;
wire n3996;
wire n39960;
wire n39961;
wire n39962;
wire n39963;
wire n39964;
wire n39965;
wire n39966;
wire n39967;
wire n39968;
wire n39969;
wire n3997;
wire n39970;
wire n39971;
wire n39972;
wire n39973;
wire n39974;
wire n39975;
wire n39976;
wire n39977;
wire n39978;
wire n39979;
wire n3998;
wire n39980;
wire n39981;
wire n39982;
wire n39983;
wire n39984;
wire n39985;
wire n39986;
wire n39987;
wire n39988;
wire n39989;
wire n3999;
wire n39990;
wire n39991;
wire n39992;
wire n39993;
wire n39994;
wire n39995;
wire n39996;
wire n39997;
wire n39998;
wire n39999;
wire n3999_1;
wire n4000;
wire n40000;
wire n40001;
wire n40002;
wire n40003;
wire n40004;
wire n40005;
wire n40006;
wire n40007;
wire n40008;
wire n40009;
wire n4001;
wire n40010;
wire n40011;
wire n40012;
wire n40013;
wire n40014;
wire n40015;
wire n40016;
wire n40017;
wire n40018;
wire n40019;
wire n4002;
wire n40020;
wire n40021;
wire n40022;
wire n40023;
wire n40024;
wire n40025;
wire n40026;
wire n40027;
wire n40028;
wire n40029;
wire n4003;
wire n40030;
wire n40031;
wire n40032;
wire n40033;
wire n40034;
wire n40035;
wire n40036;
wire n40037;
wire n40038;
wire n40039;
wire n4004;
wire n40040;
wire n40041;
wire n40042;
wire n40043;
wire n40044;
wire n40045;
wire n40046;
wire n40047;
wire n40048;
wire n40049;
wire n4004_1;
wire n4005;
wire n40050;
wire n40052;
wire n40053;
wire n40054;
wire n40055;
wire n40056;
wire n40057;
wire n40058;
wire n40059;
wire n4006;
wire n40060;
wire n40061;
wire n40062;
wire n40063;
wire n40064;
wire n40065;
wire n40067;
wire n40068;
wire n40069;
wire n4007;
wire n40070;
wire n40072;
wire n40073;
wire n40074;
wire n40075;
wire n40076;
wire n40077;
wire n40078;
wire n40079;
wire n4008;
wire n40080;
wire n40081;
wire n40082;
wire n40083;
wire n40085;
wire n40086;
wire n40087;
wire n40088;
wire n40089;
wire n4009;
wire n40090;
wire n40091;
wire n40092;
wire n40093;
wire n40094;
wire n40095;
wire n40096;
wire n40097;
wire n40098;
wire n40099;
wire n4009_1;
wire n4010;
wire n40100;
wire n40101;
wire n40102;
wire n40103;
wire n40104;
wire n40105;
wire n40106;
wire n40107;
wire n40108;
wire n40109;
wire n4011;
wire n40110;
wire n40111;
wire n40112;
wire n40113;
wire n40114;
wire n40115;
wire n40116;
wire n40117;
wire n40118;
wire n40119;
wire n4012;
wire n40120;
wire n40121;
wire n40122;
wire n40123;
wire n40124;
wire n40125;
wire n40126;
wire n40127;
wire n40128;
wire n40129;
wire n4013;
wire n40130;
wire n40131;
wire n40132;
wire n40133;
wire n40134;
wire n40135;
wire n40136;
wire n40137;
wire n40138;
wire n40139;
wire n4014;
wire n40140;
wire n40141;
wire n40142;
wire n40143;
wire n40144;
wire n40145;
wire n40146;
wire n40147;
wire n40148;
wire n40149;
wire n4014_1;
wire n4015;
wire n40150;
wire n40151;
wire n40152;
wire n40153;
wire n40154;
wire n40155;
wire n40156;
wire n40157;
wire n40158;
wire n40159;
wire n4016;
wire n40160;
wire n40161;
wire n40162;
wire n40163;
wire n40164;
wire n40165;
wire n40166;
wire n40167;
wire n40168;
wire n40169;
wire n4017;
wire n40170;
wire n40171;
wire n40172;
wire n40173;
wire n40174;
wire n40175;
wire n40176;
wire n40177;
wire n40178;
wire n40179;
wire n4018;
wire n40180;
wire n40181;
wire n40182;
wire n40183;
wire n40184;
wire n40185;
wire n40186;
wire n40187;
wire n40188;
wire n40189;
wire n4019;
wire n40190;
wire n40191;
wire n40192;
wire n40193;
wire n40194;
wire n40195;
wire n40196;
wire n40197;
wire n40198;
wire n40199;
wire n4019_1;
wire n4020;
wire n40200;
wire n40202;
wire n40203;
wire n40204;
wire n40205;
wire n40206;
wire n40207;
wire n40208;
wire n40209;
wire n4021;
wire n40210;
wire n40211;
wire n40213;
wire n40214;
wire n40215;
wire n40216;
wire n40217;
wire n40218;
wire n4022;
wire n40220;
wire n40222;
wire n40223;
wire n40226;
wire n40227;
wire n40228;
wire n40229;
wire n4023;
wire n40230;
wire n40232;
wire n40233;
wire n40234;
wire n40235;
wire n40237;
wire n40238;
wire n40239;
wire n4024;
wire n40240;
wire n40241;
wire n40242;
wire n40244;
wire n40246;
wire n40247;
wire n40248;
wire n40249;
wire n4024_1;
wire n4025;
wire n40250;
wire n40251;
wire n40252;
wire n40253;
wire n40254;
wire n40255;
wire n40256;
wire n40257;
wire n40258;
wire n40259;
wire n4026;
wire n40260;
wire n40261;
wire n40262;
wire n40263;
wire n40264;
wire n40265;
wire n40266;
wire n40267;
wire n40268;
wire n40269;
wire n4027;
wire n40270;
wire n40271;
wire n40272;
wire n40273;
wire n40274;
wire n40275;
wire n40276;
wire n40277;
wire n40278;
wire n40279;
wire n4028;
wire n40280;
wire n40281;
wire n40282;
wire n40283;
wire n40284;
wire n40285;
wire n40286;
wire n40287;
wire n40288;
wire n40289;
wire n4028_1;
wire n4029;
wire n40290;
wire n40291;
wire n40292;
wire n40293;
wire n40294;
wire n40295;
wire n40296;
wire n40297;
wire n40298;
wire n40299;
wire n403;
wire n4030;
wire n40300;
wire n40301;
wire n40302;
wire n40303;
wire n40304;
wire n40305;
wire n40306;
wire n40307;
wire n40308;
wire n40309;
wire n4031;
wire n40310;
wire n40311;
wire n40312;
wire n40313;
wire n40314;
wire n40315;
wire n40316;
wire n40317;
wire n40318;
wire n4032;
wire n40321;
wire n40322;
wire n40323;
wire n40324;
wire n40325;
wire n40326;
wire n40327;
wire n40328;
wire n40329;
wire n4033;
wire n40331;
wire n40332;
wire n40333;
wire n40334;
wire n40335;
wire n40336;
wire n40338;
wire n40339;
wire n4033_1;
wire n4034;
wire n40341;
wire n40342;
wire n40343;
wire n40344;
wire n40345;
wire n40346;
wire n40348;
wire n40349;
wire n4035;
wire n40350;
wire n40351;
wire n40352;
wire n40354;
wire n40355;
wire n40356;
wire n40357;
wire n40358;
wire n40359;
wire n4036;
wire n40360;
wire n40361;
wire n40362;
wire n40363;
wire n40365;
wire n40367;
wire n40368;
wire n40369;
wire n4037;
wire n40370;
wire n40372;
wire n40373;
wire n40375;
wire n40376;
wire n40377;
wire n40378;
wire n40379;
wire n4038;
wire n40380;
wire n40381;
wire n40382;
wire n40383;
wire n40385;
wire n40386;
wire n40387;
wire n40388;
wire n40389;
wire n4038_1;
wire n4039;
wire n40390;
wire n40391;
wire n40392;
wire n40393;
wire n40394;
wire n40396;
wire n40397;
wire n40398;
wire n40399;
wire n4040;
wire n40400;
wire n40401;
wire n40402;
wire n40403;
wire n40405;
wire n40406;
wire n40407;
wire n40408;
wire n40409;
wire n4041;
wire n40410;
wire n40412;
wire n40413;
wire n40414;
wire n40415;
wire n40416;
wire n40418;
wire n40419;
wire n4042;
wire n40420;
wire n40421;
wire n40422;
wire n40423;
wire n40425;
wire n40426;
wire n40427;
wire n40428;
wire n4043;
wire n40430;
wire n40431;
wire n40432;
wire n40433;
wire n40434;
wire n40435;
wire n40436;
wire n40437;
wire n40439;
wire n4043_1;
wire n4044;
wire n40440;
wire n40441;
wire n40442;
wire n40443;
wire n40444;
wire n40446;
wire n40447;
wire n40448;
wire n40449;
wire n4045;
wire n40450;
wire n40451;
wire n40452;
wire n40453;
wire n40454;
wire n40456;
wire n40457;
wire n40458;
wire n40459;
wire n4046;
wire n40461;
wire n40462;
wire n40463;
wire n40464;
wire n40465;
wire n40467;
wire n40469;
wire n4047;
wire n40470;
wire n40471;
wire n40472;
wire n40473;
wire n40474;
wire n40476;
wire n40477;
wire n40478;
wire n40479;
wire n4048;
wire n40481;
wire n40482;
wire n40483;
wire n40484;
wire n40486;
wire n40487;
wire n40488;
wire n40489;
wire n4048_1;
wire n4049;
wire n40490;
wire n40491;
wire n40493;
wire n40494;
wire n40496;
wire n40497;
wire n40499;
wire n4050;
wire n40500;
wire n40502;
wire n40503;
wire n40504;
wire n40505;
wire n40506;
wire n40507;
wire n40508;
wire n40509;
wire n4051;
wire n40510;
wire n40511;
wire n40512;
wire n40513;
wire n40514;
wire n40516;
wire n40517;
wire n40518;
wire n40519;
wire n4052;
wire n40520;
wire n40522;
wire n40523;
wire n40524;
wire n40525;
wire n40527;
wire n40528;
wire n40529;
wire n4053;
wire n40530;
wire n40531;
wire n40532;
wire n40533;
wire n40534;
wire n40535;
wire n40536;
wire n40537;
wire n40539;
wire n4053_1;
wire n4054;
wire n40540;
wire n40541;
wire n40542;
wire n40543;
wire n40545;
wire n40546;
wire n40547;
wire n40548;
wire n40549;
wire n4055;
wire n40550;
wire n40551;
wire n40553;
wire n40554;
wire n40556;
wire n40557;
wire n40559;
wire n4056;
wire n40561;
wire n40563;
wire n40564;
wire n40565;
wire n40566;
wire n40567;
wire n40568;
wire n40569;
wire n4057;
wire n40570;
wire n40571;
wire n40572;
wire n40573;
wire n40574;
wire n40575;
wire n40576;
wire n40577;
wire n40578;
wire n40579;
wire n4058;
wire n40580;
wire n40581;
wire n40582;
wire n40583;
wire n40584;
wire n40585;
wire n40586;
wire n40587;
wire n40588;
wire n40589;
wire n4058_1;
wire n4059;
wire n40590;
wire n40591;
wire n40592;
wire n40593;
wire n40594;
wire n40595;
wire n40596;
wire n40597;
wire n40599;
wire n4060;
wire n40600;
wire n40601;
wire n40602;
wire n40603;
wire n40604;
wire n40606;
wire n40608;
wire n40609;
wire n4061;
wire n40610;
wire n40611;
wire n40612;
wire n40613;
wire n40615;
wire n40616;
wire n40618;
wire n40619;
wire n4062;
wire n40620;
wire n40621;
wire n40622;
wire n40623;
wire n40624;
wire n40625;
wire n40626;
wire n40627;
wire n40628;
wire n40629;
wire n4063;
wire n40630;
wire n40631;
wire n40632;
wire n40633;
wire n40634;
wire n40635;
wire n40636;
wire n40637;
wire n40638;
wire n40639;
wire n4063_1;
wire n4064;
wire n40640;
wire n40641;
wire n40642;
wire n40643;
wire n40644;
wire n40645;
wire n40646;
wire n40647;
wire n40648;
wire n40649;
wire n4065;
wire n40650;
wire n40651;
wire n40652;
wire n40653;
wire n40654;
wire n40655;
wire n40656;
wire n40657;
wire n40658;
wire n40659;
wire n4066;
wire n40660;
wire n40661;
wire n40662;
wire n40663;
wire n40664;
wire n40665;
wire n40666;
wire n40667;
wire n40668;
wire n40669;
wire n4067;
wire n40670;
wire n40671;
wire n40672;
wire n40673;
wire n40674;
wire n40675;
wire n40676;
wire n40677;
wire n40678;
wire n40679;
wire n4068;
wire n40680;
wire n40681;
wire n40682;
wire n40683;
wire n40684;
wire n40685;
wire n40686;
wire n40687;
wire n40688;
wire n40689;
wire n4068_1;
wire n4069;
wire n40690;
wire n40691;
wire n40692;
wire n40693;
wire n40694;
wire n40695;
wire n40696;
wire n40697;
wire n40698;
wire n40699;
wire n4070;
wire n40700;
wire n40701;
wire n40702;
wire n40703;
wire n40704;
wire n40705;
wire n40706;
wire n40707;
wire n40708;
wire n40709;
wire n4071;
wire n40710;
wire n40711;
wire n40712;
wire n40713;
wire n40714;
wire n40715;
wire n40716;
wire n40717;
wire n40718;
wire n40719;
wire n4072;
wire n40720;
wire n40721;
wire n40722;
wire n40723;
wire n40724;
wire n40725;
wire n40726;
wire n40727;
wire n40728;
wire n40729;
wire n4073;
wire n40730;
wire n40731;
wire n40732;
wire n40733;
wire n40734;
wire n40735;
wire n40736;
wire n40737;
wire n40738;
wire n40739;
wire n4073_1;
wire n4074;
wire n40740;
wire n40741;
wire n40742;
wire n40743;
wire n40744;
wire n40745;
wire n40746;
wire n40747;
wire n40748;
wire n40749;
wire n4075;
wire n40750;
wire n40751;
wire n40752;
wire n40753;
wire n40754;
wire n40755;
wire n40756;
wire n40757;
wire n40758;
wire n40759;
wire n4076;
wire n40760;
wire n40761;
wire n40762;
wire n40763;
wire n40764;
wire n40765;
wire n40766;
wire n40767;
wire n40768;
wire n40769;
wire n4077;
wire n40770;
wire n40771;
wire n40772;
wire n40773;
wire n40774;
wire n40775;
wire n40776;
wire n40777;
wire n40778;
wire n40779;
wire n4078;
wire n40780;
wire n40781;
wire n40782;
wire n40783;
wire n40784;
wire n40785;
wire n40786;
wire n40787;
wire n40788;
wire n40789;
wire n4078_1;
wire n4079;
wire n40790;
wire n40791;
wire n40792;
wire n40793;
wire n40794;
wire n40795;
wire n40796;
wire n40797;
wire n40798;
wire n40799;
wire n408;
wire n4080;
wire n40800;
wire n40801;
wire n40802;
wire n40803;
wire n40804;
wire n40805;
wire n40806;
wire n40807;
wire n40808;
wire n40809;
wire n4081;
wire n40810;
wire n40811;
wire n40812;
wire n40813;
wire n40814;
wire n40815;
wire n40816;
wire n40817;
wire n40818;
wire n40819;
wire n4082;
wire n40820;
wire n40821;
wire n40822;
wire n40823;
wire n40824;
wire n40825;
wire n40826;
wire n40827;
wire n40828;
wire n40829;
wire n4083;
wire n40830;
wire n40831;
wire n40832;
wire n40833;
wire n40834;
wire n40835;
wire n40836;
wire n40837;
wire n40838;
wire n40839;
wire n4083_1;
wire n4084;
wire n40840;
wire n40841;
wire n40842;
wire n40843;
wire n40844;
wire n40845;
wire n40846;
wire n40847;
wire n40848;
wire n40849;
wire n4085;
wire n40850;
wire n40851;
wire n40852;
wire n40853;
wire n40854;
wire n40855;
wire n40856;
wire n40857;
wire n40858;
wire n40859;
wire n4086;
wire n40860;
wire n40861;
wire n40862;
wire n40863;
wire n40864;
wire n40865;
wire n40866;
wire n40867;
wire n40868;
wire n40869;
wire n4087;
wire n40870;
wire n40871;
wire n40872;
wire n40873;
wire n40874;
wire n40875;
wire n40876;
wire n40877;
wire n40878;
wire n40879;
wire n4088;
wire n40880;
wire n40881;
wire n40882;
wire n40883;
wire n40884;
wire n40885;
wire n40886;
wire n40887;
wire n40888;
wire n40889;
wire n4088_1;
wire n4089;
wire n40890;
wire n40891;
wire n40892;
wire n40893;
wire n40894;
wire n40895;
wire n40896;
wire n40897;
wire n40898;
wire n40899;
wire n4090;
wire n40900;
wire n40901;
wire n40902;
wire n40903;
wire n40904;
wire n40905;
wire n40906;
wire n40907;
wire n40908;
wire n40909;
wire n4091;
wire n40910;
wire n40911;
wire n40912;
wire n40913;
wire n40914;
wire n40915;
wire n40916;
wire n40917;
wire n40918;
wire n40919;
wire n4092;
wire n40920;
wire n40921;
wire n40922;
wire n40923;
wire n40924;
wire n40925;
wire n40926;
wire n40927;
wire n40928;
wire n40929;
wire n4093;
wire n40930;
wire n40931;
wire n40932;
wire n40933;
wire n40934;
wire n40935;
wire n40936;
wire n40937;
wire n40938;
wire n40939;
wire n4093_1;
wire n4094;
wire n40940;
wire n40941;
wire n40942;
wire n40943;
wire n40944;
wire n40945;
wire n40946;
wire n40947;
wire n40948;
wire n40949;
wire n4095;
wire n40950;
wire n40951;
wire n40952;
wire n40954;
wire n40956;
wire n40957;
wire n40958;
wire n40959;
wire n4096;
wire n40960;
wire n40961;
wire n40962;
wire n40963;
wire n40964;
wire n40965;
wire n40967;
wire n40968;
wire n40969;
wire n4097;
wire n40971;
wire n40972;
wire n40973;
wire n40974;
wire n40975;
wire n40976;
wire n40978;
wire n4098;
wire n40980;
wire n40981;
wire n40982;
wire n40983;
wire n40984;
wire n40986;
wire n40987;
wire n40988;
wire n40989;
wire n4098_1;
wire n4099;
wire n40990;
wire n40991;
wire n40992;
wire n40993;
wire n40994;
wire n40995;
wire n40996;
wire n40997;
wire n40999;
wire n4100;
wire n41000;
wire n41002;
wire n41003;
wire n41005;
wire n41006;
wire n41007;
wire n41008;
wire n41009;
wire n4101;
wire n41010;
wire n41011;
wire n41012;
wire n41013;
wire n41014;
wire n41015;
wire n41016;
wire n41017;
wire n41018;
wire n41019;
wire n4102;
wire n41020;
wire n41021;
wire n41022;
wire n41023;
wire n41024;
wire n41025;
wire n41026;
wire n41027;
wire n41028;
wire n41029;
wire n4103;
wire n41030;
wire n41031;
wire n41032;
wire n41033;
wire n41034;
wire n41035;
wire n41036;
wire n41037;
wire n41038;
wire n41039;
wire n4103_1;
wire n4104;
wire n41040;
wire n41042;
wire n41043;
wire n41044;
wire n41045;
wire n41046;
wire n41047;
wire n41048;
wire n41049;
wire n4105;
wire n41050;
wire n41051;
wire n41052;
wire n41053;
wire n41055;
wire n41056;
wire n41057;
wire n41058;
wire n4106;
wire n41060;
wire n41061;
wire n41062;
wire n41063;
wire n41064;
wire n41065;
wire n41066;
wire n41067;
wire n41068;
wire n41069;
wire n4107;
wire n41071;
wire n41073;
wire n41074;
wire n41075;
wire n41076;
wire n41077;
wire n41078;
wire n41079;
wire n4107_1;
wire n4108;
wire n41080;
wire n41081;
wire n41082;
wire n41083;
wire n41084;
wire n41085;
wire n41087;
wire n41089;
wire n4109;
wire n41090;
wire n41091;
wire n41092;
wire n41093;
wire n41094;
wire n41095;
wire n41096;
wire n41097;
wire n41098;
wire n41099;
wire n4110;
wire n41100;
wire n41101;
wire n41102;
wire n41103;
wire n41105;
wire n41106;
wire n41107;
wire n41109;
wire n4111;
wire n41110;
wire n41111;
wire n41112;
wire n41113;
wire n41115;
wire n41116;
wire n41117;
wire n41118;
wire n4112;
wire n41120;
wire n41121;
wire n41122;
wire n41123;
wire n41124;
wire n41125;
wire n41126;
wire n41127;
wire n41128;
wire n41129;
wire n4112_1;
wire n4113;
wire n41130;
wire n41131;
wire n41132;
wire n41133;
wire n41135;
wire n41136;
wire n41137;
wire n41138;
wire n41139;
wire n4114;
wire n41140;
wire n41141;
wire n41142;
wire n41144;
wire n41145;
wire n41146;
wire n41147;
wire n41148;
wire n41149;
wire n4115;
wire n41150;
wire n41151;
wire n41152;
wire n41154;
wire n41155;
wire n41156;
wire n41157;
wire n41158;
wire n41159;
wire n4116;
wire n41160;
wire n41161;
wire n41162;
wire n41164;
wire n41165;
wire n41166;
wire n41167;
wire n41168;
wire n41169;
wire n4116_1;
wire n4117;
wire n41170;
wire n41171;
wire n41172;
wire n41173;
wire n41174;
wire n41175;
wire n41176;
wire n41177;
wire n41178;
wire n4118;
wire n41180;
wire n41181;
wire n41182;
wire n41183;
wire n41184;
wire n41185;
wire n41186;
wire n41187;
wire n41188;
wire n41189;
wire n4119;
wire n41190;
wire n41191;
wire n41192;
wire n41193;
wire n41194;
wire n41195;
wire n41196;
wire n41197;
wire n41198;
wire n41199;
wire n4120;
wire n41200;
wire n41201;
wire n41202;
wire n41203;
wire n41204;
wire n41205;
wire n41206;
wire n41207;
wire n41208;
wire n41209;
wire n4121;
wire n41210;
wire n41211;
wire n41212;
wire n41213;
wire n41214;
wire n41215;
wire n41217;
wire n41218;
wire n41219;
wire n4121_1;
wire n4122;
wire n41220;
wire n41221;
wire n41222;
wire n41223;
wire n41224;
wire n41225;
wire n41226;
wire n41227;
wire n41228;
wire n41229;
wire n4123;
wire n41230;
wire n41231;
wire n41232;
wire n41233;
wire n41234;
wire n41235;
wire n41236;
wire n41237;
wire n41238;
wire n41239;
wire n4124;
wire n41240;
wire n41241;
wire n41242;
wire n41243;
wire n41244;
wire n41245;
wire n41246;
wire n41247;
wire n41248;
wire n41249;
wire n4125;
wire n41250;
wire n41251;
wire n41252;
wire n41253;
wire n41254;
wire n41255;
wire n41257;
wire n41258;
wire n41259;
wire n4126;
wire n41260;
wire n41261;
wire n41262;
wire n41264;
wire n41266;
wire n41267;
wire n41268;
wire n41269;
wire n4126_1;
wire n4127;
wire n41270;
wire n41271;
wire n41272;
wire n41273;
wire n41274;
wire n41275;
wire n41276;
wire n41277;
wire n41278;
wire n41279;
wire n4128;
wire n41280;
wire n41281;
wire n41282;
wire n41283;
wire n41284;
wire n41285;
wire n41286;
wire n41287;
wire n41288;
wire n41289;
wire n4129;
wire n41290;
wire n41291;
wire n41292;
wire n41293;
wire n41294;
wire n41295;
wire n41296;
wire n41297;
wire n41298;
wire n41299;
wire n413;
wire n4130;
wire n41300;
wire n41301;
wire n41302;
wire n41303;
wire n41304;
wire n41305;
wire n41306;
wire n41307;
wire n41308;
wire n41309;
wire n4131;
wire n41310;
wire n41311;
wire n41312;
wire n41313;
wire n41314;
wire n41315;
wire n41316;
wire n41317;
wire n41318;
wire n41319;
wire n4131_1;
wire n4132;
wire n41320;
wire n41321;
wire n41322;
wire n41323;
wire n41324;
wire n41325;
wire n41326;
wire n41327;
wire n41328;
wire n41329;
wire n4133;
wire n41330;
wire n41331;
wire n41332;
wire n41333;
wire n41334;
wire n41335;
wire n41336;
wire n41337;
wire n41338;
wire n41339;
wire n4134;
wire n41340;
wire n41341;
wire n41342;
wire n41343;
wire n41344;
wire n41345;
wire n41346;
wire n41347;
wire n41348;
wire n41349;
wire n4135;
wire n41350;
wire n41351;
wire n41352;
wire n41353;
wire n41354;
wire n41355;
wire n41356;
wire n41357;
wire n41358;
wire n41359;
wire n4136;
wire n41360;
wire n41361;
wire n41362;
wire n41363;
wire n41364;
wire n41365;
wire n41366;
wire n41367;
wire n41368;
wire n41369;
wire n4136_1;
wire n4137;
wire n41370;
wire n41371;
wire n41372;
wire n41373;
wire n41374;
wire n41375;
wire n41376;
wire n41378;
wire n41379;
wire n4138;
wire n41380;
wire n41381;
wire n41382;
wire n41383;
wire n41384;
wire n41385;
wire n41386;
wire n41387;
wire n41388;
wire n41389;
wire n4139;
wire n41390;
wire n41391;
wire n41392;
wire n41393;
wire n41394;
wire n41395;
wire n41396;
wire n41397;
wire n41399;
wire n4140;
wire n41401;
wire n41402;
wire n41404;
wire n41405;
wire n41406;
wire n41407;
wire n41408;
wire n41409;
wire n4141;
wire n41410;
wire n41411;
wire n41412;
wire n41414;
wire n41415;
wire n41416;
wire n41418;
wire n41419;
wire n4141_1;
wire n4142;
wire n41420;
wire n41421;
wire n41422;
wire n41423;
wire n41424;
wire n41425;
wire n41427;
wire n41428;
wire n41429;
wire n4143;
wire n41430;
wire n41431;
wire n41432;
wire n41434;
wire n41435;
wire n41437;
wire n41439;
wire n4144;
wire n41440;
wire n41442;
wire n41443;
wire n41444;
wire n41445;
wire n41446;
wire n41447;
wire n41448;
wire n41449;
wire n4145;
wire n41450;
wire n41451;
wire n41452;
wire n41454;
wire n41455;
wire n41456;
wire n41457;
wire n41458;
wire n41459;
wire n4146;
wire n41460;
wire n41461;
wire n41463;
wire n41465;
wire n41466;
wire n41468;
wire n41469;
wire n4146_1;
wire n4147;
wire n41470;
wire n41471;
wire n41472;
wire n41473;
wire n41474;
wire n41475;
wire n41476;
wire n41477;
wire n41478;
wire n41479;
wire n4148;
wire n41480;
wire n41481;
wire n41482;
wire n41483;
wire n41484;
wire n41485;
wire n41486;
wire n41487;
wire n41488;
wire n41489;
wire n4149;
wire n41490;
wire n41491;
wire n41492;
wire n41493;
wire n41494;
wire n41495;
wire n41496;
wire n41497;
wire n41498;
wire n41499;
wire n4150;
wire n41500;
wire n41501;
wire n41503;
wire n41504;
wire n41506;
wire n41507;
wire n41508;
wire n41509;
wire n4151;
wire n41510;
wire n41511;
wire n41512;
wire n41513;
wire n41514;
wire n41515;
wire n41516;
wire n41517;
wire n41518;
wire n4151_1;
wire n4152;
wire n41520;
wire n41521;
wire n41522;
wire n41523;
wire n41524;
wire n41525;
wire n41527;
wire n41529;
wire n4153;
wire n41530;
wire n41531;
wire n41532;
wire n41533;
wire n41534;
wire n41535;
wire n41536;
wire n41537;
wire n41538;
wire n41539;
wire n4154;
wire n41540;
wire n41541;
wire n41542;
wire n41543;
wire n41544;
wire n41545;
wire n41546;
wire n41547;
wire n41548;
wire n41549;
wire n4155;
wire n41550;
wire n41551;
wire n41552;
wire n41553;
wire n41554;
wire n41555;
wire n41556;
wire n41557;
wire n41558;
wire n41559;
wire n4156;
wire n41560;
wire n41561;
wire n41562;
wire n41563;
wire n41564;
wire n41565;
wire n41566;
wire n41567;
wire n41568;
wire n41569;
wire n4156_1;
wire n4157;
wire n41570;
wire n41571;
wire n41572;
wire n41573;
wire n41574;
wire n41575;
wire n41576;
wire n41577;
wire n41578;
wire n41579;
wire n4158;
wire n41580;
wire n41581;
wire n41582;
wire n41583;
wire n41584;
wire n41585;
wire n41586;
wire n41587;
wire n41588;
wire n41589;
wire n4159;
wire n41590;
wire n41591;
wire n41592;
wire n41593;
wire n41594;
wire n41595;
wire n41596;
wire n41597;
wire n41598;
wire n41599;
wire n4160;
wire n41600;
wire n41601;
wire n41602;
wire n41603;
wire n41604;
wire n41605;
wire n41606;
wire n41607;
wire n41608;
wire n41609;
wire n4161;
wire n41610;
wire n41611;
wire n41612;
wire n41613;
wire n41614;
wire n41615;
wire n41616;
wire n41617;
wire n41618;
wire n41619;
wire n4161_1;
wire n4162;
wire n41620;
wire n41621;
wire n41622;
wire n41623;
wire n41624;
wire n41625;
wire n41626;
wire n41627;
wire n41628;
wire n41629;
wire n4163;
wire n41630;
wire n41631;
wire n41632;
wire n41633;
wire n41634;
wire n41635;
wire n41636;
wire n41637;
wire n41638;
wire n41639;
wire n4164;
wire n41640;
wire n41641;
wire n41642;
wire n41643;
wire n41644;
wire n41645;
wire n41646;
wire n41647;
wire n41649;
wire n4165;
wire n41650;
wire n41651;
wire n41652;
wire n41653;
wire n41654;
wire n41655;
wire n41656;
wire n41657;
wire n41658;
wire n41659;
wire n4166;
wire n41661;
wire n41662;
wire n41664;
wire n41665;
wire n41666;
wire n41667;
wire n41668;
wire n41669;
wire n4166_1;
wire n4167;
wire n41670;
wire n41671;
wire n41672;
wire n41674;
wire n41675;
wire n41676;
wire n41677;
wire n41678;
wire n41679;
wire n4168;
wire n41680;
wire n41681;
wire n41682;
wire n41683;
wire n41684;
wire n41685;
wire n41686;
wire n41687;
wire n41688;
wire n41689;
wire n4169;
wire n41690;
wire n41691;
wire n41692;
wire n41693;
wire n41694;
wire n41695;
wire n41696;
wire n41697;
wire n41698;
wire n41699;
wire n4170;
wire n41700;
wire n41701;
wire n41702;
wire n41703;
wire n41704;
wire n41705;
wire n41706;
wire n41707;
wire n41708;
wire n41709;
wire n4171;
wire n41710;
wire n41712;
wire n41713;
wire n41714;
wire n41715;
wire n41716;
wire n41718;
wire n41719;
wire n4171_1;
wire n4172;
wire n41720;
wire n41721;
wire n41722;
wire n41723;
wire n41724;
wire n41725;
wire n41726;
wire n41727;
wire n41728;
wire n41729;
wire n4173;
wire n41730;
wire n41731;
wire n41732;
wire n41733;
wire n41734;
wire n41735;
wire n41736;
wire n41737;
wire n41738;
wire n41739;
wire n4174;
wire n41740;
wire n41741;
wire n41742;
wire n41743;
wire n41744;
wire n41745;
wire n41746;
wire n41747;
wire n41749;
wire n4175;
wire n41750;
wire n41751;
wire n41752;
wire n41753;
wire n41755;
wire n41756;
wire n41757;
wire n41758;
wire n41759;
wire n4176;
wire n41761;
wire n41762;
wire n41763;
wire n41764;
wire n41765;
wire n41766;
wire n41767;
wire n41768;
wire n41769;
wire n4176_1;
wire n4177;
wire n41770;
wire n41771;
wire n41772;
wire n41773;
wire n41775;
wire n41776;
wire n41777;
wire n41778;
wire n41779;
wire n4178;
wire n41780;
wire n41781;
wire n41783;
wire n41785;
wire n41786;
wire n41787;
wire n41788;
wire n41789;
wire n4179;
wire n41790;
wire n41791;
wire n41792;
wire n41794;
wire n41795;
wire n41797;
wire n41798;
wire n41799;
wire n418;
wire n4180;
wire n41800;
wire n41801;
wire n41802;
wire n41803;
wire n41804;
wire n41805;
wire n41806;
wire n41807;
wire n41808;
wire n41809;
wire n4181;
wire n41810;
wire n41811;
wire n41812;
wire n41813;
wire n41814;
wire n41815;
wire n41817;
wire n41818;
wire n41819;
wire n4181_1;
wire n4182;
wire n41820;
wire n41822;
wire n41823;
wire n41824;
wire n41825;
wire n41826;
wire n41828;
wire n41829;
wire n4183;
wire n41830;
wire n41831;
wire n41832;
wire n41833;
wire n41834;
wire n41835;
wire n41836;
wire n41837;
wire n41838;
wire n41839;
wire n4184;
wire n41841;
wire n41843;
wire n41844;
wire n41845;
wire n41846;
wire n41847;
wire n41848;
wire n41849;
wire n4185;
wire n41850;
wire n41851;
wire n41852;
wire n41853;
wire n41854;
wire n41856;
wire n41857;
wire n41858;
wire n41859;
wire n4186;
wire n41860;
wire n41861;
wire n41862;
wire n41863;
wire n41865;
wire n41866;
wire n41867;
wire n41868;
wire n41869;
wire n4186_1;
wire n4187;
wire n41871;
wire n41872;
wire n41873;
wire n41874;
wire n41875;
wire n41876;
wire n41877;
wire n41878;
wire n41879;
wire n4188;
wire n41880;
wire n41881;
wire n41882;
wire n41884;
wire n41885;
wire n41886;
wire n41887;
wire n41888;
wire n41889;
wire n4189;
wire n41890;
wire n41891;
wire n41892;
wire n41893;
wire n41894;
wire n41895;
wire n41897;
wire n41898;
wire n41899;
wire n4190;
wire n41900;
wire n41901;
wire n41902;
wire n41903;
wire n41905;
wire n41906;
wire n41907;
wire n41908;
wire n41909;
wire n4191;
wire n41910;
wire n41911;
wire n41913;
wire n41915;
wire n41916;
wire n41917;
wire n41918;
wire n41919;
wire n4191_1;
wire n4192;
wire n41920;
wire n41921;
wire n41922;
wire n41923;
wire n41924;
wire n41925;
wire n41927;
wire n41928;
wire n41929;
wire n4193;
wire n41930;
wire n41932;
wire n41933;
wire n41934;
wire n41935;
wire n41936;
wire n41938;
wire n41939;
wire n4194;
wire n41940;
wire n41941;
wire n41942;
wire n41943;
wire n41944;
wire n41945;
wire n41946;
wire n41948;
wire n41949;
wire n4195;
wire n41950;
wire n41951;
wire n41952;
wire n41953;
wire n41954;
wire n41955;
wire n41956;
wire n41958;
wire n41959;
wire n4196;
wire n41960;
wire n41961;
wire n41962;
wire n41963;
wire n41964;
wire n41965;
wire n41966;
wire n41967;
wire n41969;
wire n4196_1;
wire n4197;
wire n41970;
wire n41971;
wire n41972;
wire n41973;
wire n41974;
wire n41975;
wire n41976;
wire n41977;
wire n41978;
wire n41979;
wire n4198;
wire n41980;
wire n41981;
wire n41982;
wire n41983;
wire n41984;
wire n41985;
wire n41987;
wire n41988;
wire n41989;
wire n4199;
wire n41990;
wire n41991;
wire n41992;
wire n41993;
wire n41994;
wire n41995;
wire n41996;
wire n41997;
wire n41998;
wire n41999;
wire n4200;
wire n42000;
wire n42001;
wire n42002;
wire n42003;
wire n42004;
wire n42005;
wire n42006;
wire n42007;
wire n42008;
wire n42009;
wire n4201;
wire n42010;
wire n42011;
wire n42012;
wire n42013;
wire n42014;
wire n42015;
wire n42016;
wire n42017;
wire n42018;
wire n42019;
wire n4201_1;
wire n4202;
wire n42020;
wire n42021;
wire n42022;
wire n42023;
wire n42024;
wire n42025;
wire n42026;
wire n42027;
wire n42028;
wire n42029;
wire n4203;
wire n42030;
wire n42032;
wire n42033;
wire n42034;
wire n42035;
wire n42036;
wire n42037;
wire n42038;
wire n4204;
wire n42040;
wire n42041;
wire n42043;
wire n42044;
wire n42045;
wire n42046;
wire n42047;
wire n42048;
wire n42049;
wire n4205;
wire n42050;
wire n42052;
wire n42053;
wire n42054;
wire n42055;
wire n42056;
wire n42058;
wire n42059;
wire n4206;
wire n42060;
wire n42061;
wire n42062;
wire n42063;
wire n42064;
wire n42065;
wire n42067;
wire n42068;
wire n4206_1;
wire n4207;
wire n42070;
wire n42071;
wire n42072;
wire n42073;
wire n42074;
wire n42075;
wire n42076;
wire n42077;
wire n42078;
wire n42079;
wire n4208;
wire n42080;
wire n42081;
wire n42084;
wire n42085;
wire n42087;
wire n42088;
wire n42089;
wire n4209;
wire n42090;
wire n42091;
wire n42092;
wire n42094;
wire n42095;
wire n42097;
wire n42098;
wire n42099;
wire n4210;
wire n42100;
wire n42101;
wire n42102;
wire n42103;
wire n42104;
wire n42106;
wire n42107;
wire n42109;
wire n4211;
wire n42110;
wire n42111;
wire n42112;
wire n42113;
wire n42114;
wire n42115;
wire n42116;
wire n42118;
wire n42119;
wire n4211_1;
wire n4212;
wire n42120;
wire n42121;
wire n42122;
wire n42123;
wire n42124;
wire n42125;
wire n42126;
wire n42128;
wire n42129;
wire n4213;
wire n42130;
wire n42131;
wire n42132;
wire n42134;
wire n42135;
wire n42136;
wire n42137;
wire n42138;
wire n42139;
wire n4214;
wire n42140;
wire n42141;
wire n42142;
wire n42144;
wire n42145;
wire n42146;
wire n42147;
wire n42148;
wire n42149;
wire n4215;
wire n42150;
wire n42151;
wire n42152;
wire n42153;
wire n42154;
wire n42156;
wire n42158;
wire n42159;
wire n4216;
wire n42160;
wire n42161;
wire n42162;
wire n42163;
wire n42165;
wire n42167;
wire n42168;
wire n42169;
wire n4216_1;
wire n4217;
wire n42170;
wire n42172;
wire n42173;
wire n42174;
wire n42175;
wire n42176;
wire n42177;
wire n42178;
wire n42179;
wire n4218;
wire n42181;
wire n42182;
wire n42183;
wire n42184;
wire n42185;
wire n42186;
wire n42187;
wire n42189;
wire n4219;
wire n42190;
wire n42191;
wire n42192;
wire n42193;
wire n42194;
wire n42195;
wire n42197;
wire n42198;
wire n42199;
wire n422;
wire n4220;
wire n42200;
wire n42201;
wire n42202;
wire n42204;
wire n42206;
wire n42207;
wire n42208;
wire n42209;
wire n4221;
wire n42210;
wire n42211;
wire n42212;
wire n42214;
wire n42215;
wire n42216;
wire n42217;
wire n42218;
wire n42219;
wire n4221_1;
wire n4222;
wire n42220;
wire n42221;
wire n42222;
wire n42224;
wire n42225;
wire n42226;
wire n42227;
wire n42228;
wire n42229;
wire n4223;
wire n42231;
wire n42233;
wire n42234;
wire n42235;
wire n42236;
wire n42237;
wire n42238;
wire n42239;
wire n4224;
wire n42240;
wire n42241;
wire n42242;
wire n42243;
wire n42244;
wire n42246;
wire n42247;
wire n42248;
wire n42249;
wire n4225;
wire n42250;
wire n42251;
wire n42253;
wire n42254;
wire n42255;
wire n42256;
wire n42257;
wire n42259;
wire n4226;
wire n42260;
wire n42261;
wire n42262;
wire n42263;
wire n42264;
wire n42266;
wire n42267;
wire n42268;
wire n42269;
wire n4226_1;
wire n4227;
wire n42270;
wire n42271;
wire n42272;
wire n42273;
wire n42275;
wire n42276;
wire n42277;
wire n42278;
wire n42279;
wire n4228;
wire n42280;
wire n42281;
wire n42283;
wire n42284;
wire n42285;
wire n42286;
wire n42287;
wire n42288;
wire n42289;
wire n4229;
wire n42290;
wire n42291;
wire n42292;
wire n42293;
wire n42294;
wire n42295;
wire n42296;
wire n42297;
wire n42298;
wire n42299;
wire n4230;
wire n42300;
wire n42301;
wire n42303;
wire n42304;
wire n42305;
wire n42306;
wire n42307;
wire n42308;
wire n42309;
wire n4231;
wire n42311;
wire n42312;
wire n42313;
wire n42314;
wire n42315;
wire n42316;
wire n42317;
wire n42318;
wire n42319;
wire n4231_1;
wire n4232;
wire n42320;
wire n42322;
wire n42323;
wire n42325;
wire n42326;
wire n42327;
wire n42328;
wire n42329;
wire n4233;
wire n42331;
wire n42332;
wire n42334;
wire n42335;
wire n42337;
wire n42338;
wire n42339;
wire n4234;
wire n42340;
wire n42341;
wire n42342;
wire n42343;
wire n42344;
wire n42345;
wire n42346;
wire n42347;
wire n42348;
wire n4235;
wire n42350;
wire n42351;
wire n42352;
wire n42353;
wire n42354;
wire n42355;
wire n42356;
wire n42357;
wire n42358;
wire n42359;
wire n4236;
wire n42360;
wire n42361;
wire n42362;
wire n42364;
wire n42365;
wire n42366;
wire n42367;
wire n42368;
wire n42369;
wire n4236_1;
wire n4237;
wire n42370;
wire n42371;
wire n42372;
wire n42373;
wire n42376;
wire n42377;
wire n42378;
wire n42379;
wire n4238;
wire n42380;
wire n42381;
wire n42382;
wire n42383;
wire n42384;
wire n42385;
wire n42386;
wire n42387;
wire n42388;
wire n42389;
wire n4239;
wire n42390;
wire n42391;
wire n42393;
wire n42394;
wire n42395;
wire n42396;
wire n42397;
wire n42398;
wire n42399;
wire n4240;
wire n42400;
wire n42401;
wire n42402;
wire n42403;
wire n42405;
wire n42406;
wire n42407;
wire n42408;
wire n42409;
wire n4241;
wire n42410;
wire n42411;
wire n42413;
wire n42414;
wire n42415;
wire n42416;
wire n42417;
wire n42419;
wire n4241_1;
wire n4242;
wire n42420;
wire n42421;
wire n42422;
wire n42423;
wire n42425;
wire n42426;
wire n42427;
wire n42428;
wire n42429;
wire n4243;
wire n42430;
wire n42431;
wire n42433;
wire n42434;
wire n42435;
wire n42436;
wire n42437;
wire n42438;
wire n42439;
wire n4244;
wire n42441;
wire n42442;
wire n42443;
wire n42444;
wire n42445;
wire n42446;
wire n42447;
wire n42448;
wire n42449;
wire n4245;
wire n42450;
wire n42451;
wire n42452;
wire n42453;
wire n42454;
wire n42455;
wire n42456;
wire n42457;
wire n42458;
wire n42459;
wire n4246;
wire n42461;
wire n42462;
wire n42463;
wire n42464;
wire n42465;
wire n42466;
wire n42467;
wire n42468;
wire n4246_1;
wire n4247;
wire n42470;
wire n42471;
wire n42472;
wire n42473;
wire n42474;
wire n42475;
wire n42476;
wire n42478;
wire n4248;
wire n42480;
wire n42481;
wire n42482;
wire n42483;
wire n42484;
wire n42485;
wire n42486;
wire n42487;
wire n42488;
wire n4249;
wire n42490;
wire n42492;
wire n42493;
wire n42494;
wire n42495;
wire n42496;
wire n42497;
wire n42498;
wire n42499;
wire n4250;
wire n42500;
wire n42501;
wire n42502;
wire n42504;
wire n42506;
wire n42507;
wire n42508;
wire n42509;
wire n4251;
wire n42510;
wire n42511;
wire n42512;
wire n42513;
wire n42514;
wire n42515;
wire n42517;
wire n42518;
wire n42519;
wire n4251_1;
wire n4252;
wire n42520;
wire n42521;
wire n42522;
wire n42523;
wire n42524;
wire n42525;
wire n42526;
wire n42527;
wire n42528;
wire n42529;
wire n4253;
wire n42530;
wire n42532;
wire n42533;
wire n42534;
wire n42535;
wire n42536;
wire n42538;
wire n42539;
wire n4254;
wire n42540;
wire n42541;
wire n42542;
wire n42543;
wire n42545;
wire n42546;
wire n42547;
wire n42548;
wire n42549;
wire n4255;
wire n42551;
wire n42552;
wire n42554;
wire n42555;
wire n42556;
wire n42557;
wire n42558;
wire n42559;
wire n4256;
wire n42560;
wire n42561;
wire n42562;
wire n42563;
wire n42564;
wire n42566;
wire n42567;
wire n42568;
wire n42569;
wire n4256_1;
wire n4257;
wire n42570;
wire n42571;
wire n42573;
wire n42574;
wire n42575;
wire n42576;
wire n42577;
wire n42579;
wire n4258;
wire n42580;
wire n42581;
wire n42582;
wire n42583;
wire n42584;
wire n42585;
wire n42586;
wire n42587;
wire n42588;
wire n42589;
wire n4259;
wire n42590;
wire n42591;
wire n42592;
wire n42594;
wire n42596;
wire n42597;
wire n42598;
wire n42599;
wire n4260;
wire n42600;
wire n42601;
wire n42603;
wire n42604;
wire n42605;
wire n42606;
wire n42607;
wire n42608;
wire n4261;
wire n42610;
wire n42611;
wire n42612;
wire n42613;
wire n42614;
wire n42615;
wire n42616;
wire n42618;
wire n42619;
wire n4261_1;
wire n4262;
wire n42620;
wire n42621;
wire n42622;
wire n42623;
wire n42625;
wire n42626;
wire n42627;
wire n42628;
wire n4263;
wire n42630;
wire n42631;
wire n42632;
wire n42633;
wire n42634;
wire n42635;
wire n42636;
wire n42637;
wire n42638;
wire n42639;
wire n4264;
wire n42640;
wire n42642;
wire n42643;
wire n42644;
wire n42645;
wire n42646;
wire n42647;
wire n42648;
wire n42649;
wire n4265;
wire n42650;
wire n42651;
wire n42652;
wire n42653;
wire n42655;
wire n42656;
wire n42657;
wire n42658;
wire n42659;
wire n4266;
wire n42660;
wire n42662;
wire n42663;
wire n42664;
wire n42665;
wire n42666;
wire n42667;
wire n42668;
wire n42669;
wire n4266_1;
wire n4267;
wire n42671;
wire n42672;
wire n42673;
wire n42674;
wire n42675;
wire n42676;
wire n42677;
wire n42678;
wire n4268;
wire n42680;
wire n42682;
wire n42683;
wire n42684;
wire n42685;
wire n42687;
wire n42688;
wire n42689;
wire n4269;
wire n42690;
wire n42691;
wire n42693;
wire n42694;
wire n42695;
wire n42696;
wire n42697;
wire n42698;
wire n42699;
wire n427;
wire n4270;
wire n42700;
wire n42701;
wire n42702;
wire n42703;
wire n42704;
wire n42705;
wire n42706;
wire n42707;
wire n42708;
wire n42709;
wire n4271;
wire n42711;
wire n42712;
wire n42713;
wire n42714;
wire n42716;
wire n42717;
wire n42718;
wire n42719;
wire n4271_1;
wire n4272;
wire n42720;
wire n42721;
wire n42722;
wire n42723;
wire n42724;
wire n42725;
wire n42726;
wire n42727;
wire n42728;
wire n42729;
wire n4273;
wire n42730;
wire n42732;
wire n42734;
wire n42735;
wire n42736;
wire n42737;
wire n42738;
wire n42739;
wire n4274;
wire n42740;
wire n42743;
wire n42744;
wire n42745;
wire n42746;
wire n42747;
wire n42748;
wire n42749;
wire n4275;
wire n42750;
wire n42751;
wire n42752;
wire n42753;
wire n42754;
wire n42755;
wire n42756;
wire n42758;
wire n42759;
wire n4275_1;
wire n4276;
wire n42760;
wire n42761;
wire n42762;
wire n42764;
wire n42765;
wire n42766;
wire n42767;
wire n42768;
wire n42769;
wire n4277;
wire n42771;
wire n42772;
wire n42773;
wire n42774;
wire n42775;
wire n42776;
wire n42777;
wire n42778;
wire n4278;
wire n42780;
wire n42781;
wire n42782;
wire n42783;
wire n42785;
wire n42787;
wire n42788;
wire n42789;
wire n4279;
wire n42790;
wire n42791;
wire n42792;
wire n42793;
wire n42795;
wire n42796;
wire n42797;
wire n42798;
wire n42799;
wire n4280;
wire n42800;
wire n42801;
wire n42803;
wire n42804;
wire n42805;
wire n42806;
wire n42807;
wire n42808;
wire n42809;
wire n4280_1;
wire n4281;
wire n42810;
wire n42811;
wire n42812;
wire n42814;
wire n42815;
wire n42816;
wire n42817;
wire n42818;
wire n42819;
wire n4282;
wire n42820;
wire n42821;
wire n42822;
wire n42823;
wire n42824;
wire n42825;
wire n42826;
wire n42827;
wire n42828;
wire n42829;
wire n4283;
wire n42830;
wire n42831;
wire n42832;
wire n42833;
wire n42834;
wire n42835;
wire n42836;
wire n42837;
wire n42838;
wire n42839;
wire n4284;
wire n42840;
wire n42841;
wire n42842;
wire n42843;
wire n42844;
wire n42845;
wire n42846;
wire n42847;
wire n42848;
wire n42849;
wire n4285;
wire n42850;
wire n42851;
wire n42852;
wire n42853;
wire n42854;
wire n42855;
wire n42856;
wire n42857;
wire n42858;
wire n42859;
wire n4285_1;
wire n4286;
wire n42860;
wire n42861;
wire n42862;
wire n42863;
wire n42864;
wire n42865;
wire n42866;
wire n42867;
wire n42868;
wire n42869;
wire n4287;
wire n42870;
wire n42871;
wire n42872;
wire n42873;
wire n42874;
wire n42875;
wire n42876;
wire n42877;
wire n42878;
wire n42879;
wire n4288;
wire n42880;
wire n42881;
wire n42882;
wire n42883;
wire n42884;
wire n42885;
wire n42886;
wire n42887;
wire n42888;
wire n42889;
wire n4289;
wire n42890;
wire n42891;
wire n42892;
wire n42893;
wire n42894;
wire n42896;
wire n42897;
wire n42898;
wire n42899;
wire n4290;
wire n42900;
wire n42901;
wire n42902;
wire n42904;
wire n42905;
wire n42906;
wire n42907;
wire n42908;
wire n42909;
wire n4290_1;
wire n4291;
wire n42910;
wire n42911;
wire n42912;
wire n42913;
wire n42914;
wire n42915;
wire n42916;
wire n42917;
wire n42918;
wire n42919;
wire n4292;
wire n42920;
wire n42921;
wire n42922;
wire n42923;
wire n42925;
wire n42926;
wire n42927;
wire n42928;
wire n42929;
wire n4293;
wire n42930;
wire n42931;
wire n42932;
wire n42933;
wire n42934;
wire n42936;
wire n42937;
wire n42938;
wire n42939;
wire n4294;
wire n42940;
wire n42941;
wire n42943;
wire n42945;
wire n42946;
wire n42947;
wire n42948;
wire n42949;
wire n4295;
wire n42950;
wire n42951;
wire n42952;
wire n42953;
wire n42954;
wire n42955;
wire n42957;
wire n42958;
wire n42959;
wire n4295_1;
wire n4296;
wire n42960;
wire n42961;
wire n42962;
wire n42963;
wire n42964;
wire n42966;
wire n42968;
wire n42969;
wire n4297;
wire n42970;
wire n42971;
wire n42972;
wire n42973;
wire n42974;
wire n42975;
wire n42976;
wire n42977;
wire n42978;
wire n42979;
wire n4298;
wire n42981;
wire n42982;
wire n42983;
wire n42984;
wire n42985;
wire n42986;
wire n42988;
wire n4299;
wire n42990;
wire n42991;
wire n42992;
wire n42993;
wire n42995;
wire n42996;
wire n42997;
wire n42998;
wire n42999;
wire n4300;
wire n43000;
wire n43001;
wire n43002;
wire n43003;
wire n43005;
wire n43006;
wire n43007;
wire n43008;
wire n43009;
wire n4300_1;
wire n4301;
wire n43010;
wire n43012;
wire n43013;
wire n43015;
wire n43016;
wire n43017;
wire n43018;
wire n43019;
wire n4302;
wire n43020;
wire n43021;
wire n43022;
wire n43023;
wire n43024;
wire n43025;
wire n43026;
wire n43028;
wire n43029;
wire n4303;
wire n43030;
wire n43031;
wire n43032;
wire n43034;
wire n43036;
wire n43037;
wire n43038;
wire n43039;
wire n4304;
wire n43040;
wire n43041;
wire n43042;
wire n43044;
wire n43045;
wire n43046;
wire n43047;
wire n43048;
wire n43049;
wire n4305;
wire n43050;
wire n43051;
wire n43052;
wire n43053;
wire n43055;
wire n43056;
wire n43057;
wire n43058;
wire n43059;
wire n4305_1;
wire n4306;
wire n43061;
wire n43062;
wire n43063;
wire n43064;
wire n43065;
wire n43067;
wire n43069;
wire n4307;
wire n43070;
wire n43071;
wire n43072;
wire n43073;
wire n43074;
wire n43075;
wire n43076;
wire n43077;
wire n43078;
wire n43079;
wire n4308;
wire n43081;
wire n43082;
wire n43083;
wire n43084;
wire n43085;
wire n43087;
wire n43088;
wire n43089;
wire n4309;
wire n43090;
wire n43092;
wire n43093;
wire n43094;
wire n43095;
wire n43096;
wire n43097;
wire n43098;
wire n43099;
wire n4310;
wire n43100;
wire n43101;
wire n43102;
wire n43103;
wire n43105;
wire n43106;
wire n43107;
wire n43108;
wire n43109;
wire n4310_1;
wire n4311;
wire n43110;
wire n43111;
wire n43112;
wire n43113;
wire n43114;
wire n43115;
wire n43116;
wire n43117;
wire n43118;
wire n43119;
wire n4312;
wire n43120;
wire n43121;
wire n43122;
wire n43123;
wire n43124;
wire n43125;
wire n43126;
wire n43127;
wire n43129;
wire n4313;
wire n43130;
wire n43131;
wire n43132;
wire n43133;
wire n43134;
wire n43135;
wire n43136;
wire n43137;
wire n43138;
wire n43139;
wire n4314;
wire n43140;
wire n43141;
wire n43142;
wire n43143;
wire n43145;
wire n43146;
wire n43148;
wire n43149;
wire n4315;
wire n43151;
wire n43152;
wire n43153;
wire n43154;
wire n43155;
wire n43156;
wire n43157;
wire n43158;
wire n43159;
wire n4315_1;
wire n4316;
wire n43160;
wire n43162;
wire n43163;
wire n43165;
wire n43166;
wire n43167;
wire n43168;
wire n43169;
wire n4317;
wire n43172;
wire n43173;
wire n43175;
wire n43176;
wire n43177;
wire n43178;
wire n4318;
wire n43180;
wire n43181;
wire n43182;
wire n43183;
wire n43184;
wire n43185;
wire n43186;
wire n43187;
wire n43188;
wire n43189;
wire n4319;
wire n43191;
wire n43192;
wire n43193;
wire n43194;
wire n43196;
wire n43197;
wire n43198;
wire n43199;
wire n432;
wire n4320;
wire n43200;
wire n43201;
wire n43203;
wire n43204;
wire n43205;
wire n43206;
wire n43207;
wire n43208;
wire n4320_1;
wire n4321;
wire n43210;
wire n43211;
wire n43212;
wire n43213;
wire n43214;
wire n43216;
wire n43217;
wire n43218;
wire n43219;
wire n4322;
wire n43220;
wire n43221;
wire n43222;
wire n43223;
wire n43225;
wire n43226;
wire n43228;
wire n43229;
wire n4323;
wire n43230;
wire n43231;
wire n43232;
wire n43233;
wire n43235;
wire n43236;
wire n43237;
wire n43238;
wire n43239;
wire n4324;
wire n43241;
wire n43242;
wire n43244;
wire n43245;
wire n43246;
wire n43248;
wire n43249;
wire n4325;
wire n43252;
wire n43253;
wire n43254;
wire n43255;
wire n43256;
wire n43257;
wire n43258;
wire n43259;
wire n4325_1;
wire n4326;
wire n43261;
wire n43262;
wire n43263;
wire n43264;
wire n43265;
wire n43266;
wire n43267;
wire n43268;
wire n43269;
wire n4327;
wire n43270;
wire n43272;
wire n43273;
wire n43275;
wire n43276;
wire n43277;
wire n43278;
wire n43279;
wire n4328;
wire n43280;
wire n43281;
wire n43282;
wire n43283;
wire n43284;
wire n43286;
wire n43287;
wire n43288;
wire n43289;
wire n4329;
wire n43291;
wire n43292;
wire n43294;
wire n43295;
wire n43296;
wire n43297;
wire n43298;
wire n43299;
wire n4330;
wire n43300;
wire n43301;
wire n43302;
wire n43304;
wire n43306;
wire n43307;
wire n43308;
wire n43309;
wire n4330_1;
wire n4331;
wire n43310;
wire n43311;
wire n43313;
wire n43314;
wire n43315;
wire n43316;
wire n43317;
wire n43318;
wire n4332;
wire n43320;
wire n43322;
wire n43323;
wire n43325;
wire n43326;
wire n43327;
wire n43328;
wire n43329;
wire n4333;
wire n43330;
wire n43332;
wire n43334;
wire n43335;
wire n43337;
wire n43338;
wire n43339;
wire n4334;
wire n43340;
wire n43342;
wire n43343;
wire n43344;
wire n43345;
wire n43347;
wire n43349;
wire n4334_1;
wire n4335;
wire n43350;
wire n43352;
wire n43353;
wire n43355;
wire n43356;
wire n43357;
wire n43358;
wire n43359;
wire n4336;
wire n43361;
wire n43362;
wire n43364;
wire n43365;
wire n43366;
wire n43367;
wire n43368;
wire n43369;
wire n4337;
wire n43370;
wire n43372;
wire n43373;
wire n43374;
wire n43375;
wire n43376;
wire n43377;
wire n43379;
wire n4338;
wire n43380;
wire n43381;
wire n43382;
wire n43383;
wire n43384;
wire n43385;
wire n43386;
wire n43387;
wire n43389;
wire n4339;
wire n43391;
wire n43393;
wire n43394;
wire n43395;
wire n43396;
wire n43397;
wire n43398;
wire n43399;
wire n4339_1;
wire n4340;
wire n43402;
wire n43403;
wire n43404;
wire n43405;
wire n43407;
wire n43408;
wire n43409;
wire n4341;
wire n43410;
wire n43411;
wire n43412;
wire n43413;
wire n43415;
wire n43416;
wire n43417;
wire n43418;
wire n43419;
wire n4342;
wire n43420;
wire n43421;
wire n43422;
wire n43423;
wire n43424;
wire n43425;
wire n43426;
wire n43427;
wire n43428;
wire n4343;
wire n43430;
wire n43431;
wire n43432;
wire n43433;
wire n43434;
wire n43435;
wire n43436;
wire n43437;
wire n43438;
wire n43439;
wire n4344;
wire n43441;
wire n43442;
wire n43443;
wire n43444;
wire n43445;
wire n43447;
wire n43448;
wire n43449;
wire n4344_1;
wire n4345;
wire n43450;
wire n43452;
wire n43453;
wire n43454;
wire n43456;
wire n43457;
wire n43458;
wire n43459;
wire n4346;
wire n43460;
wire n43462;
wire n43464;
wire n43465;
wire n43466;
wire n43467;
wire n43468;
wire n4347;
wire n43470;
wire n43472;
wire n43473;
wire n43474;
wire n43475;
wire n43476;
wire n43477;
wire n43478;
wire n43479;
wire n4348;
wire n43480;
wire n43481;
wire n43483;
wire n43484;
wire n43485;
wire n43486;
wire n43487;
wire n4349;
wire n43490;
wire n43491;
wire n43492;
wire n43493;
wire n43495;
wire n43497;
wire n43498;
wire n4349_1;
wire n4350;
wire n43500;
wire n43501;
wire n43502;
wire n43503;
wire n43505;
wire n43506;
wire n43507;
wire n43508;
wire n43509;
wire n4351;
wire n43510;
wire n43511;
wire n43513;
wire n43514;
wire n43515;
wire n43516;
wire n43518;
wire n43519;
wire n4352;
wire n43520;
wire n43521;
wire n43522;
wire n43523;
wire n43524;
wire n43525;
wire n43526;
wire n43527;
wire n43528;
wire n43529;
wire n4353;
wire n43530;
wire n43532;
wire n43533;
wire n43534;
wire n43535;
wire n43536;
wire n43538;
wire n43539;
wire n4354;
wire n43541;
wire n43542;
wire n43544;
wire n43545;
wire n43546;
wire n43547;
wire n43549;
wire n4354_1;
wire n4355;
wire n43550;
wire n43551;
wire n43552;
wire n43553;
wire n43554;
wire n43555;
wire n43557;
wire n43559;
wire n4356;
wire n43560;
wire n43561;
wire n43562;
wire n43563;
wire n43564;
wire n43565;
wire n43566;
wire n43567;
wire n4357;
wire n43570;
wire n43571;
wire n43572;
wire n43573;
wire n43574;
wire n43575;
wire n43576;
wire n43577;
wire n43579;
wire n4358;
wire n43580;
wire n43581;
wire n43582;
wire n43583;
wire n43585;
wire n43586;
wire n43587;
wire n43588;
wire n43589;
wire n4359;
wire n43590;
wire n43591;
wire n43592;
wire n43594;
wire n43595;
wire n43596;
wire n43597;
wire n43598;
wire n43599;
wire n4359_1;
wire n4360;
wire n43601;
wire n43602;
wire n43604;
wire n43606;
wire n43607;
wire n43608;
wire n43609;
wire n4361;
wire n43610;
wire n43611;
wire n43612;
wire n43613;
wire n43614;
wire n43616;
wire n43617;
wire n43618;
wire n43619;
wire n4362;
wire n43620;
wire n43621;
wire n43622;
wire n43623;
wire n43624;
wire n43625;
wire n43626;
wire n43627;
wire n43628;
wire n43629;
wire n4363;
wire n43631;
wire n43632;
wire n43633;
wire n43634;
wire n43635;
wire n43636;
wire n43637;
wire n43638;
wire n43639;
wire n4364;
wire n43640;
wire n43642;
wire n43644;
wire n43645;
wire n43647;
wire n43648;
wire n43649;
wire n4364_1;
wire n4365;
wire n43650;
wire n43651;
wire n43652;
wire n43653;
wire n43654;
wire n43655;
wire n43656;
wire n43657;
wire n43658;
wire n43659;
wire n4366;
wire n43660;
wire n43661;
wire n43662;
wire n43663;
wire n43665;
wire n43666;
wire n43667;
wire n43668;
wire n43669;
wire n4367;
wire n43670;
wire n43671;
wire n43672;
wire n43673;
wire n43675;
wire n43676;
wire n43677;
wire n43678;
wire n43679;
wire n4368;
wire n43681;
wire n43683;
wire n43684;
wire n43685;
wire n43686;
wire n43687;
wire n43688;
wire n43689;
wire n4369;
wire n43691;
wire n43692;
wire n43693;
wire n43694;
wire n43695;
wire n43696;
wire n43698;
wire n43699;
wire n4369_1;
wire n437;
wire n4370;
wire n43700;
wire n43701;
wire n43702;
wire n43703;
wire n43705;
wire n43706;
wire n43707;
wire n43708;
wire n43709;
wire n4371;
wire n43711;
wire n43712;
wire n43713;
wire n43715;
wire n43716;
wire n43717;
wire n43718;
wire n4372;
wire n43720;
wire n43722;
wire n43723;
wire n43724;
wire n43725;
wire n43726;
wire n43727;
wire n43729;
wire n4373;
wire n43730;
wire n43731;
wire n43732;
wire n43733;
wire n43734;
wire n43735;
wire n43736;
wire n43737;
wire n43738;
wire n4374;
wire n43740;
wire n43741;
wire n43742;
wire n43743;
wire n43744;
wire n43745;
wire n43747;
wire n43749;
wire n4374_1;
wire n4375;
wire n43750;
wire n43751;
wire n43752;
wire n43753;
wire n43754;
wire n43755;
wire n43756;
wire n43758;
wire n4376;
wire n43760;
wire n43761;
wire n43762;
wire n43763;
wire n43765;
wire n43766;
wire n43767;
wire n43768;
wire n43769;
wire n4377;
wire n43770;
wire n43771;
wire n43772;
wire n43773;
wire n43775;
wire n43777;
wire n43778;
wire n43779;
wire n4378;
wire n43780;
wire n43781;
wire n43782;
wire n43783;
wire n43784;
wire n43785;
wire n43786;
wire n43787;
wire n43788;
wire n43789;
wire n4379;
wire n43790;
wire n43791;
wire n43793;
wire n43794;
wire n43795;
wire n43796;
wire n43797;
wire n43799;
wire n4379_1;
wire n4380;
wire n43800;
wire n43801;
wire n43802;
wire n43803;
wire n43804;
wire n43806;
wire n43807;
wire n43808;
wire n43809;
wire n4381;
wire n43810;
wire n43811;
wire n43812;
wire n43813;
wire n43815;
wire n43816;
wire n43817;
wire n43818;
wire n43819;
wire n4382;
wire n43820;
wire n43821;
wire n43822;
wire n43823;
wire n43824;
wire n43826;
wire n43827;
wire n43829;
wire n4383;
wire n43830;
wire n43831;
wire n43832;
wire n43833;
wire n43834;
wire n43835;
wire n43836;
wire n43837;
wire n43838;
wire n4384;
wire n43840;
wire n43841;
wire n43842;
wire n43843;
wire n43844;
wire n43845;
wire n43846;
wire n43847;
wire n43848;
wire n43849;
wire n4384_1;
wire n4385;
wire n43850;
wire n43851;
wire n43852;
wire n43853;
wire n43854;
wire n43855;
wire n43857;
wire n43858;
wire n43859;
wire n4386;
wire n43860;
wire n43862;
wire n43863;
wire n43864;
wire n43865;
wire n43866;
wire n43867;
wire n43868;
wire n43869;
wire n4387;
wire n43870;
wire n43871;
wire n43872;
wire n43873;
wire n43874;
wire n43875;
wire n43876;
wire n43877;
wire n43878;
wire n43879;
wire n4388;
wire n43880;
wire n43881;
wire n43882;
wire n43883;
wire n43884;
wire n43885;
wire n43887;
wire n43888;
wire n4389;
wire n43890;
wire n43891;
wire n43892;
wire n43893;
wire n43895;
wire n43896;
wire n43897;
wire n43898;
wire n43899;
wire n4389_1;
wire n4390;
wire n43900;
wire n43901;
wire n43902;
wire n43903;
wire n43905;
wire n43906;
wire n43907;
wire n43908;
wire n43909;
wire n4391;
wire n43910;
wire n43911;
wire n43912;
wire n43913;
wire n43914;
wire n43916;
wire n43918;
wire n43919;
wire n4392;
wire n43920;
wire n43921;
wire n43922;
wire n43923;
wire n43924;
wire n43925;
wire n43927;
wire n43928;
wire n43929;
wire n4393;
wire n43930;
wire n43932;
wire n43933;
wire n43936;
wire n43937;
wire n43938;
wire n43939;
wire n4394;
wire n43940;
wire n43941;
wire n43942;
wire n43943;
wire n43944;
wire n43946;
wire n43947;
wire n43948;
wire n43949;
wire n4394_1;
wire n4395;
wire n43950;
wire n43951;
wire n43953;
wire n43954;
wire n43955;
wire n43956;
wire n43957;
wire n43959;
wire n4396;
wire n43960;
wire n43962;
wire n43963;
wire n43965;
wire n43966;
wire n43968;
wire n43969;
wire n4397;
wire n43970;
wire n43971;
wire n43972;
wire n43973;
wire n43974;
wire n43975;
wire n43976;
wire n43977;
wire n43979;
wire n4398;
wire n43980;
wire n43981;
wire n43982;
wire n43983;
wire n43985;
wire n43986;
wire n43987;
wire n43988;
wire n43989;
wire n4399;
wire n43990;
wire n43991;
wire n43992;
wire n43993;
wire n43994;
wire n43995;
wire n43996;
wire n43997;
wire n43999;
wire n4399_1;
wire n4400;
wire n44000;
wire n44001;
wire n44002;
wire n44003;
wire n44004;
wire n44005;
wire n44006;
wire n44007;
wire n44008;
wire n4401;
wire n44011;
wire n44012;
wire n44013;
wire n44014;
wire n44015;
wire n44016;
wire n44017;
wire n44018;
wire n44019;
wire n4402;
wire n44020;
wire n44021;
wire n44023;
wire n44024;
wire n44027;
wire n44028;
wire n44029;
wire n4403;
wire n44030;
wire n44031;
wire n44032;
wire n44033;
wire n44034;
wire n44036;
wire n44037;
wire n44038;
wire n44039;
wire n4404;
wire n44040;
wire n44041;
wire n44042;
wire n44043;
wire n44044;
wire n44045;
wire n44046;
wire n44047;
wire n44048;
wire n44049;
wire n4404_1;
wire n4405;
wire n44050;
wire n44052;
wire n44053;
wire n44055;
wire n44056;
wire n44058;
wire n44059;
wire n4406;
wire n44060;
wire n44061;
wire n44062;
wire n44063;
wire n44064;
wire n44065;
wire n44066;
wire n44068;
wire n44069;
wire n4407;
wire n44071;
wire n44073;
wire n44074;
wire n44076;
wire n44077;
wire n44078;
wire n44079;
wire n4408;
wire n44080;
wire n44081;
wire n44083;
wire n44084;
wire n44085;
wire n44086;
wire n44088;
wire n44089;
wire n4409;
wire n44090;
wire n44091;
wire n44093;
wire n44094;
wire n44096;
wire n44097;
wire n44098;
wire n44099;
wire n4409_1;
wire n4410;
wire n44100;
wire n44101;
wire n44102;
wire n44103;
wire n44104;
wire n44105;
wire n44106;
wire n44107;
wire n44108;
wire n44109;
wire n4411;
wire n44110;
wire n44111;
wire n44112;
wire n44114;
wire n44115;
wire n44116;
wire n44117;
wire n44118;
wire n44119;
wire n4412;
wire n44121;
wire n44122;
wire n44123;
wire n44124;
wire n44125;
wire n44126;
wire n44128;
wire n44129;
wire n4413;
wire n44130;
wire n44131;
wire n44132;
wire n44133;
wire n44134;
wire n44135;
wire n44136;
wire n44138;
wire n44139;
wire n4414;
wire n44140;
wire n44141;
wire n44142;
wire n44143;
wire n44144;
wire n44145;
wire n44146;
wire n44147;
wire n44148;
wire n44149;
wire n4414_1;
wire n4415;
wire n44150;
wire n44151;
wire n44153;
wire n44154;
wire n44155;
wire n44156;
wire n44157;
wire n44158;
wire n44159;
wire n4416;
wire n44160;
wire n44161;
wire n44162;
wire n44164;
wire n44165;
wire n44166;
wire n44167;
wire n44168;
wire n44169;
wire n4417;
wire n44170;
wire n44171;
wire n44172;
wire n44173;
wire n44174;
wire n44175;
wire n44176;
wire n44177;
wire n44178;
wire n44179;
wire n4418;
wire n44180;
wire n44181;
wire n44182;
wire n44183;
wire n44184;
wire n44185;
wire n44186;
wire n44187;
wire n44189;
wire n4419;
wire n44190;
wire n44191;
wire n44192;
wire n44193;
wire n44194;
wire n44195;
wire n44196;
wire n44198;
wire n44199;
wire n4419_1;
wire n442;
wire n4420;
wire n44200;
wire n44201;
wire n44202;
wire n44203;
wire n44204;
wire n44206;
wire n44208;
wire n44209;
wire n4421;
wire n44211;
wire n44212;
wire n44213;
wire n44214;
wire n44215;
wire n44216;
wire n44217;
wire n44219;
wire n4422;
wire n44220;
wire n44221;
wire n44222;
wire n44223;
wire n44224;
wire n44225;
wire n44227;
wire n4423;
wire n44230;
wire n44231;
wire n44232;
wire n44233;
wire n44234;
wire n44235;
wire n44237;
wire n44239;
wire n4424;
wire n44240;
wire n44241;
wire n44242;
wire n44243;
wire n44244;
wire n44245;
wire n44246;
wire n44248;
wire n44249;
wire n4424_1;
wire n4425;
wire n44250;
wire n44251;
wire n44252;
wire n44253;
wire n44254;
wire n44255;
wire n44256;
wire n44257;
wire n44258;
wire n44259;
wire n4426;
wire n44260;
wire n44261;
wire n44262;
wire n44264;
wire n44265;
wire n44267;
wire n44268;
wire n44269;
wire n4427;
wire n44270;
wire n44271;
wire n44273;
wire n44274;
wire n44276;
wire n44277;
wire n44279;
wire n4428;
wire n44280;
wire n44281;
wire n44282;
wire n44284;
wire n44285;
wire n44286;
wire n44287;
wire n44288;
wire n44289;
wire n4429;
wire n44291;
wire n44293;
wire n44294;
wire n44295;
wire n44296;
wire n44298;
wire n44299;
wire n4429_1;
wire n4430;
wire n44301;
wire n44302;
wire n44303;
wire n44304;
wire n44305;
wire n44306;
wire n44307;
wire n44309;
wire n4431;
wire n44310;
wire n44312;
wire n44313;
wire n44314;
wire n44315;
wire n44316;
wire n44317;
wire n44318;
wire n44319;
wire n4432;
wire n44320;
wire n44321;
wire n44322;
wire n44323;
wire n44325;
wire n44326;
wire n44327;
wire n44328;
wire n44329;
wire n4433;
wire n44330;
wire n44332;
wire n44333;
wire n44334;
wire n44336;
wire n44337;
wire n44338;
wire n44339;
wire n4434;
wire n44340;
wire n44341;
wire n44342;
wire n44343;
wire n44345;
wire n44347;
wire n44348;
wire n44349;
wire n4434_1;
wire n4435;
wire n44350;
wire n44351;
wire n44353;
wire n44354;
wire n44356;
wire n44357;
wire n44358;
wire n44359;
wire n4436;
wire n44361;
wire n44362;
wire n44363;
wire n44364;
wire n44365;
wire n44366;
wire n44367;
wire n44368;
wire n44369;
wire n4437;
wire n44370;
wire n44371;
wire n44373;
wire n44375;
wire n44376;
wire n44377;
wire n44378;
wire n44379;
wire n4438;
wire n44380;
wire n44382;
wire n44384;
wire n44385;
wire n44386;
wire n44387;
wire n44388;
wire n44389;
wire n4439;
wire n44390;
wire n44391;
wire n44392;
wire n44393;
wire n44394;
wire n44396;
wire n44397;
wire n44398;
wire n44399;
wire n4439_1;
wire n4440;
wire n44401;
wire n44403;
wire n44404;
wire n44406;
wire n44407;
wire n44408;
wire n44409;
wire n4441;
wire n44411;
wire n44412;
wire n44413;
wire n44414;
wire n44415;
wire n44417;
wire n44419;
wire n4442;
wire n44420;
wire n44421;
wire n44423;
wire n44424;
wire n44425;
wire n44426;
wire n44427;
wire n44428;
wire n44429;
wire n4443;
wire n44430;
wire n44432;
wire n44434;
wire n44435;
wire n44436;
wire n44437;
wire n44439;
wire n4443_1;
wire n4444;
wire n44440;
wire n44441;
wire n44442;
wire n44443;
wire n44445;
wire n44446;
wire n44447;
wire n44448;
wire n44449;
wire n4445;
wire n44450;
wire n44451;
wire n44452;
wire n44455;
wire n44457;
wire n44458;
wire n44459;
wire n4446;
wire n44460;
wire n44461;
wire n44463;
wire n44464;
wire n44465;
wire n44466;
wire n44468;
wire n44469;
wire n4447;
wire n44470;
wire n44471;
wire n44472;
wire n44473;
wire n44475;
wire n44476;
wire n44478;
wire n44479;
wire n4448;
wire n44480;
wire n44481;
wire n44484;
wire n44485;
wire n44486;
wire n44487;
wire n44488;
wire n44489;
wire n4448_1;
wire n4449;
wire n44490;
wire n44491;
wire n44492;
wire n44493;
wire n44494;
wire n44495;
wire n44496;
wire n44497;
wire n44498;
wire n44499;
wire n4450;
wire n44500;
wire n44501;
wire n44503;
wire n44504;
wire n44505;
wire n44506;
wire n44507;
wire n44508;
wire n44509;
wire n4451;
wire n44510;
wire n44511;
wire n44512;
wire n44513;
wire n44514;
wire n44516;
wire n44517;
wire n44518;
wire n44519;
wire n4452;
wire n44520;
wire n44521;
wire n44522;
wire n44523;
wire n44524;
wire n44525;
wire n44527;
wire n44528;
wire n44529;
wire n4453;
wire n44530;
wire n44531;
wire n44533;
wire n44536;
wire n44537;
wire n44538;
wire n44539;
wire n4453_1;
wire n4454;
wire n44540;
wire n44541;
wire n44542;
wire n44543;
wire n44544;
wire n44545;
wire n44546;
wire n44547;
wire n44548;
wire n44549;
wire n4455;
wire n44550;
wire n44551;
wire n44552;
wire n44553;
wire n44554;
wire n44555;
wire n44556;
wire n44557;
wire n44558;
wire n44559;
wire n4456;
wire n44560;
wire n44561;
wire n44562;
wire n44563;
wire n44564;
wire n44565;
wire n44566;
wire n44567;
wire n44568;
wire n44569;
wire n4457;
wire n44570;
wire n44572;
wire n44573;
wire n44574;
wire n44575;
wire n44577;
wire n44578;
wire n44579;
wire n4458;
wire n44580;
wire n44582;
wire n44583;
wire n44584;
wire n44585;
wire n44586;
wire n44587;
wire n44588;
wire n4458_1;
wire n4459;
wire n44590;
wire n44591;
wire n44592;
wire n44593;
wire n44594;
wire n44596;
wire n44597;
wire n44599;
wire n4460;
wire n44600;
wire n44601;
wire n44602;
wire n44603;
wire n44604;
wire n44605;
wire n44606;
wire n44607;
wire n44608;
wire n44609;
wire n4461;
wire n44610;
wire n44612;
wire n44613;
wire n44614;
wire n44615;
wire n44616;
wire n44617;
wire n44619;
wire n4462;
wire n44620;
wire n44621;
wire n44622;
wire n44623;
wire n44625;
wire n44626;
wire n44627;
wire n44628;
wire n44629;
wire n4463;
wire n44630;
wire n44631;
wire n44632;
wire n44633;
wire n44635;
wire n44636;
wire n44638;
wire n44639;
wire n4463_1;
wire n4464;
wire n44641;
wire n44642;
wire n44643;
wire n44644;
wire n44645;
wire n44646;
wire n44647;
wire n44648;
wire n44649;
wire n4465;
wire n44650;
wire n44652;
wire n44653;
wire n44654;
wire n44655;
wire n44656;
wire n44657;
wire n44658;
wire n44659;
wire n4466;
wire n44660;
wire n44662;
wire n44663;
wire n44664;
wire n44665;
wire n44666;
wire n44667;
wire n44668;
wire n44669;
wire n4467;
wire n44670;
wire n44671;
wire n44672;
wire n44673;
wire n44675;
wire n44676;
wire n44677;
wire n44678;
wire n44679;
wire n4468;
wire n44680;
wire n44681;
wire n44682;
wire n44683;
wire n44684;
wire n44685;
wire n44686;
wire n44687;
wire n44688;
wire n44689;
wire n4468_1;
wire n4469;
wire n44691;
wire n44692;
wire n44693;
wire n44694;
wire n44695;
wire n44696;
wire n44697;
wire n44698;
wire n447;
wire n4470;
wire n44700;
wire n44701;
wire n44702;
wire n44703;
wire n44704;
wire n44705;
wire n44706;
wire n44707;
wire n44708;
wire n44709;
wire n4471;
wire n44710;
wire n44711;
wire n44713;
wire n44714;
wire n44715;
wire n44716;
wire n44717;
wire n44718;
wire n44719;
wire n4472;
wire n44720;
wire n44722;
wire n44724;
wire n44725;
wire n44728;
wire n4473;
wire n44730;
wire n44731;
wire n44732;
wire n44733;
wire n44734;
wire n44735;
wire n44736;
wire n44737;
wire n44738;
wire n4473_1;
wire n4474;
wire n44740;
wire n44741;
wire n44743;
wire n44744;
wire n44745;
wire n44746;
wire n44747;
wire n44749;
wire n4475;
wire n44750;
wire n44751;
wire n44752;
wire n44754;
wire n44755;
wire n44756;
wire n44757;
wire n44758;
wire n44759;
wire n4476;
wire n44760;
wire n44761;
wire n44762;
wire n44763;
wire n44764;
wire n44765;
wire n44767;
wire n44768;
wire n44769;
wire n4477;
wire n44770;
wire n44771;
wire n44772;
wire n44774;
wire n44775;
wire n44777;
wire n44778;
wire n44779;
wire n4478;
wire n44780;
wire n44781;
wire n44782;
wire n44783;
wire n44785;
wire n44786;
wire n44787;
wire n44788;
wire n44789;
wire n4478_1;
wire n4479;
wire n44790;
wire n44791;
wire n44792;
wire n44793;
wire n44794;
wire n44795;
wire n44796;
wire n44797;
wire n44798;
wire n44799;
wire n4480;
wire n44800;
wire n44801;
wire n44802;
wire n44803;
wire n44804;
wire n44805;
wire n44806;
wire n44807;
wire n44808;
wire n44809;
wire n4481;
wire n44810;
wire n44811;
wire n44812;
wire n44813;
wire n44814;
wire n44815;
wire n44816;
wire n44817;
wire n44818;
wire n44819;
wire n4482;
wire n44820;
wire n44821;
wire n44822;
wire n44823;
wire n44824;
wire n44825;
wire n44827;
wire n44828;
wire n44829;
wire n4483;
wire n44830;
wire n44831;
wire n44833;
wire n44834;
wire n44836;
wire n44837;
wire n44838;
wire n44839;
wire n4483_1;
wire n4484;
wire n44840;
wire n44842;
wire n44844;
wire n44845;
wire n44847;
wire n44848;
wire n44849;
wire n4485;
wire n44850;
wire n44851;
wire n44852;
wire n44854;
wire n44855;
wire n44857;
wire n44858;
wire n44859;
wire n4486;
wire n44860;
wire n44861;
wire n44862;
wire n44863;
wire n44865;
wire n44866;
wire n44867;
wire n44868;
wire n4487;
wire n44870;
wire n44872;
wire n44873;
wire n44874;
wire n44875;
wire n44876;
wire n44877;
wire n44879;
wire n4488;
wire n44880;
wire n44882;
wire n44883;
wire n44884;
wire n44885;
wire n44886;
wire n44887;
wire n44888;
wire n4488_1;
wire n4489;
wire n44891;
wire n44892;
wire n44894;
wire n44895;
wire n44896;
wire n44897;
wire n44898;
wire n44899;
wire n4490;
wire n44901;
wire n44902;
wire n44903;
wire n44904;
wire n44905;
wire n44907;
wire n44908;
wire n4491;
wire n44910;
wire n44911;
wire n44912;
wire n44913;
wire n44914;
wire n44915;
wire n44916;
wire n44918;
wire n4492;
wire n44920;
wire n44921;
wire n44922;
wire n44923;
wire n44924;
wire n44925;
wire n44926;
wire n44928;
wire n44929;
wire n4493;
wire n44930;
wire n44931;
wire n44932;
wire n44933;
wire n44934;
wire n44936;
wire n44937;
wire n44939;
wire n4493_1;
wire n4494;
wire n44940;
wire n44941;
wire n44942;
wire n44943;
wire n44944;
wire n44946;
wire n44947;
wire n44948;
wire n44949;
wire n4495;
wire n44950;
wire n44951;
wire n44952;
wire n44953;
wire n44955;
wire n44956;
wire n44957;
wire n44958;
wire n44959;
wire n4496;
wire n44960;
wire n44961;
wire n44962;
wire n44963;
wire n44964;
wire n44966;
wire n44967;
wire n44968;
wire n4497;
wire n44970;
wire n44971;
wire n44972;
wire n44973;
wire n44974;
wire n44976;
wire n44977;
wire n44978;
wire n44979;
wire n4498;
wire n44980;
wire n44981;
wire n44982;
wire n44983;
wire n44985;
wire n44986;
wire n44987;
wire n44988;
wire n44989;
wire n4498_1;
wire n4499;
wire n44990;
wire n44992;
wire n44993;
wire n44995;
wire n44996;
wire n44997;
wire n44998;
wire n44999;
wire n4500;
wire n45000;
wire n45002;
wire n45003;
wire n45004;
wire n45005;
wire n45007;
wire n45008;
wire n45009;
wire n4501;
wire n45010;
wire n45012;
wire n45013;
wire n45015;
wire n45016;
wire n45017;
wire n45018;
wire n45019;
wire n4502;
wire n45020;
wire n45022;
wire n45023;
wire n45024;
wire n45025;
wire n45026;
wire n45027;
wire n45029;
wire n4503;
wire n45030;
wire n45032;
wire n45033;
wire n45035;
wire n45036;
wire n45037;
wire n45038;
wire n45039;
wire n4503_1;
wire n4504;
wire n45040;
wire n45041;
wire n45042;
wire n45043;
wire n45044;
wire n45045;
wire n45047;
wire n45048;
wire n45049;
wire n4505;
wire n45050;
wire n45051;
wire n45052;
wire n45053;
wire n45054;
wire n45056;
wire n45057;
wire n45058;
wire n45059;
wire n4506;
wire n45060;
wire n45061;
wire n45062;
wire n45064;
wire n45065;
wire n45067;
wire n45068;
wire n45069;
wire n4507;
wire n45070;
wire n45071;
wire n45072;
wire n45073;
wire n45074;
wire n45075;
wire n45076;
wire n45077;
wire n45078;
wire n45079;
wire n4508;
wire n45080;
wire n45082;
wire n45083;
wire n45084;
wire n45085;
wire n45086;
wire n45087;
wire n45088;
wire n45089;
wire n4508_1;
wire n4509;
wire n45090;
wire n45091;
wire n45092;
wire n45093;
wire n45094;
wire n45096;
wire n45097;
wire n45098;
wire n45099;
wire n4510;
wire n45100;
wire n45101;
wire n45102;
wire n45103;
wire n45104;
wire n45105;
wire n45106;
wire n45107;
wire n45108;
wire n45109;
wire n4511;
wire n45110;
wire n45112;
wire n45113;
wire n45114;
wire n45115;
wire n45116;
wire n45118;
wire n45119;
wire n4512;
wire n45120;
wire n45121;
wire n45122;
wire n45126;
wire n45127;
wire n45129;
wire n4513;
wire n45130;
wire n45131;
wire n45132;
wire n45133;
wire n45134;
wire n45136;
wire n45138;
wire n45139;
wire n4513_1;
wire n4514;
wire n45140;
wire n45141;
wire n45142;
wire n45143;
wire n45144;
wire n45146;
wire n45147;
wire n45149;
wire n4515;
wire n45150;
wire n45151;
wire n45152;
wire n45153;
wire n45154;
wire n45155;
wire n45156;
wire n45157;
wire n45159;
wire n4516;
wire n45160;
wire n45161;
wire n45162;
wire n45163;
wire n45164;
wire n45165;
wire n45166;
wire n45167;
wire n45169;
wire n4517;
wire n45170;
wire n45172;
wire n45173;
wire n45175;
wire n45176;
wire n45177;
wire n45178;
wire n45179;
wire n4518;
wire n45180;
wire n45181;
wire n45182;
wire n45183;
wire n45184;
wire n45185;
wire n45186;
wire n45187;
wire n45189;
wire n4518_1;
wire n4519;
wire n45190;
wire n45191;
wire n45192;
wire n45193;
wire n45194;
wire n45195;
wire n45196;
wire n45197;
wire n45198;
wire n45199;
wire n452;
wire n4520;
wire n45201;
wire n45202;
wire n45203;
wire n45204;
wire n45205;
wire n45206;
wire n45207;
wire n45209;
wire n4521;
wire n45210;
wire n45211;
wire n45212;
wire n45213;
wire n45214;
wire n45216;
wire n45217;
wire n45218;
wire n45219;
wire n4522;
wire n45220;
wire n45221;
wire n45222;
wire n45223;
wire n45224;
wire n45226;
wire n45227;
wire n45229;
wire n4523;
wire n45230;
wire n45231;
wire n45232;
wire n45233;
wire n45234;
wire n45235;
wire n45236;
wire n45237;
wire n45238;
wire n45239;
wire n4523_1;
wire n4524;
wire n45241;
wire n45243;
wire n45244;
wire n45245;
wire n45246;
wire n45247;
wire n45248;
wire n4525;
wire n45250;
wire n45251;
wire n45252;
wire n45253;
wire n45255;
wire n45256;
wire n45257;
wire n45258;
wire n45259;
wire n4526;
wire n45260;
wire n45261;
wire n45262;
wire n45263;
wire n45264;
wire n45265;
wire n45266;
wire n45267;
wire n45269;
wire n4527;
wire n45270;
wire n45271;
wire n45272;
wire n45274;
wire n45275;
wire n45276;
wire n45277;
wire n45278;
wire n4528;
wire n45280;
wire n45281;
wire n45282;
wire n45283;
wire n45285;
wire n45286;
wire n45287;
wire n45288;
wire n45289;
wire n4528_1;
wire n4529;
wire n45290;
wire n45292;
wire n45293;
wire n45294;
wire n45295;
wire n45296;
wire n45297;
wire n45298;
wire n45299;
wire n4530;
wire n45301;
wire n45302;
wire n45303;
wire n45304;
wire n45305;
wire n45306;
wire n45308;
wire n4531;
wire n45310;
wire n45311;
wire n45313;
wire n45315;
wire n45316;
wire n45317;
wire n45318;
wire n45319;
wire n4532;
wire n45320;
wire n45322;
wire n45324;
wire n45325;
wire n45326;
wire n45327;
wire n45328;
wire n45329;
wire n4533;
wire n45331;
wire n45332;
wire n45333;
wire n45334;
wire n45336;
wire n45337;
wire n45338;
wire n45339;
wire n4533_1;
wire n4534;
wire n45340;
wire n45341;
wire n45342;
wire n45343;
wire n45344;
wire n45346;
wire n45347;
wire n45348;
wire n45349;
wire n4535;
wire n45350;
wire n45351;
wire n45352;
wire n45353;
wire n45354;
wire n45356;
wire n45357;
wire n45358;
wire n4536;
wire n45360;
wire n45361;
wire n45362;
wire n45363;
wire n45365;
wire n45366;
wire n45367;
wire n45368;
wire n45369;
wire n4537;
wire n45370;
wire n45371;
wire n45372;
wire n45373;
wire n45375;
wire n45377;
wire n45378;
wire n45379;
wire n4538;
wire n45380;
wire n45382;
wire n45383;
wire n45384;
wire n45385;
wire n45386;
wire n45387;
wire n45388;
wire n45389;
wire n4538_1;
wire n4539;
wire n45390;
wire n45391;
wire n45392;
wire n45394;
wire n45395;
wire n45396;
wire n45397;
wire n45398;
wire n45399;
wire n4540;
wire n45401;
wire n45402;
wire n45403;
wire n45404;
wire n45405;
wire n45406;
wire n45408;
wire n45409;
wire n4541;
wire n45410;
wire n45411;
wire n45413;
wire n45414;
wire n45415;
wire n45416;
wire n45417;
wire n45418;
wire n45419;
wire n4542;
wire n45420;
wire n45421;
wire n45423;
wire n45424;
wire n45425;
wire n45426;
wire n45427;
wire n45428;
wire n45429;
wire n4543;
wire n45430;
wire n45431;
wire n45432;
wire n45433;
wire n45434;
wire n45435;
wire n45437;
wire n45438;
wire n45439;
wire n4543_1;
wire n4544;
wire n45440;
wire n45441;
wire n45442;
wire n45443;
wire n45444;
wire n45445;
wire n45446;
wire n45447;
wire n45448;
wire n45449;
wire n4545;
wire n45450;
wire n45452;
wire n45453;
wire n45454;
wire n45455;
wire n45456;
wire n45458;
wire n45459;
wire n4546;
wire n45460;
wire n45461;
wire n45462;
wire n45464;
wire n45466;
wire n45467;
wire n45468;
wire n45469;
wire n4547;
wire n45470;
wire n45472;
wire n45473;
wire n45475;
wire n45476;
wire n45478;
wire n45479;
wire n4548;
wire n45480;
wire n45481;
wire n45482;
wire n45484;
wire n45485;
wire n45487;
wire n45488;
wire n4548_1;
wire n4549;
wire n45490;
wire n45491;
wire n45493;
wire n45494;
wire n45495;
wire n45496;
wire n45497;
wire n45498;
wire n45499;
wire n4550;
wire n45500;
wire n45501;
wire n45502;
wire n45503;
wire n45505;
wire n45506;
wire n45507;
wire n45508;
wire n45509;
wire n4551;
wire n45510;
wire n45511;
wire n45512;
wire n45513;
wire n45515;
wire n45516;
wire n45517;
wire n45518;
wire n4552;
wire n45520;
wire n45521;
wire n45524;
wire n45525;
wire n45526;
wire n45527;
wire n45529;
wire n4553;
wire n45530;
wire n45532;
wire n45533;
wire n45534;
wire n45535;
wire n45537;
wire n45538;
wire n45539;
wire n4553_1;
wire n4554;
wire n45540;
wire n45542;
wire n45543;
wire n45544;
wire n45545;
wire n45546;
wire n45548;
wire n45549;
wire n4555;
wire n45550;
wire n45551;
wire n45553;
wire n45554;
wire n45555;
wire n45556;
wire n45557;
wire n45558;
wire n45559;
wire n4556;
wire n45560;
wire n45561;
wire n45562;
wire n45563;
wire n45564;
wire n45565;
wire n45567;
wire n45568;
wire n4557;
wire n45570;
wire n45571;
wire n45572;
wire n45573;
wire n45574;
wire n45575;
wire n45577;
wire n45578;
wire n45579;
wire n4558;
wire n45580;
wire n45581;
wire n45582;
wire n45584;
wire n45585;
wire n45586;
wire n45588;
wire n45589;
wire n4558_1;
wire n4559;
wire n45590;
wire n45591;
wire n45592;
wire n45595;
wire n45596;
wire n45597;
wire n45598;
wire n45599;
wire n4560;
wire n45600;
wire n45602;
wire n45603;
wire n45605;
wire n45606;
wire n45608;
wire n45609;
wire n4561;
wire n45610;
wire n45611;
wire n45612;
wire n45613;
wire n45614;
wire n45616;
wire n45617;
wire n45618;
wire n45619;
wire n4562;
wire n45620;
wire n45621;
wire n45622;
wire n45623;
wire n45624;
wire n45626;
wire n45627;
wire n45628;
wire n45629;
wire n4563;
wire n45630;
wire n45631;
wire n45632;
wire n45633;
wire n45635;
wire n45636;
wire n45638;
wire n45639;
wire n4563_1;
wire n4564;
wire n45640;
wire n45641;
wire n45642;
wire n45644;
wire n45645;
wire n45646;
wire n45647;
wire n45648;
wire n45649;
wire n4565;
wire n45650;
wire n45651;
wire n45653;
wire n45655;
wire n45656;
wire n45657;
wire n45658;
wire n45659;
wire n4566;
wire n45660;
wire n45661;
wire n45662;
wire n45663;
wire n45664;
wire n45666;
wire n45667;
wire n45668;
wire n45669;
wire n4567;
wire n45671;
wire n45672;
wire n45673;
wire n45674;
wire n45675;
wire n45676;
wire n45677;
wire n45678;
wire n45679;
wire n4568;
wire n45681;
wire n45682;
wire n45683;
wire n45684;
wire n45685;
wire n45686;
wire n45687;
wire n45688;
wire n4568_1;
wire n4569;
wire n45690;
wire n45691;
wire n45692;
wire n45693;
wire n45694;
wire n45695;
wire n45696;
wire n45697;
wire n45698;
wire n45699;
wire n457;
wire n4570;
wire n45701;
wire n45702;
wire n45704;
wire n45705;
wire n45707;
wire n45708;
wire n4571;
wire n45710;
wire n45711;
wire n45713;
wire n45714;
wire n45716;
wire n45717;
wire n45718;
wire n45719;
wire n4572;
wire n45720;
wire n45724;
wire n45725;
wire n45727;
wire n45728;
wire n4573;
wire n45730;
wire n45731;
wire n45733;
wire n45734;
wire n45736;
wire n45737;
wire n45738;
wire n45739;
wire n4573_1;
wire n4574;
wire n45740;
wire n45741;
wire n45742;
wire n45743;
wire n45744;
wire n45745;
wire n45747;
wire n45748;
wire n45749;
wire n4575;
wire n45750;
wire n45751;
wire n45752;
wire n45753;
wire n45754;
wire n45755;
wire n45756;
wire n45758;
wire n45759;
wire n4576;
wire n45761;
wire n45762;
wire n45763;
wire n45764;
wire n45765;
wire n45766;
wire n45767;
wire n4577;
wire n45771;
wire n45772;
wire n45773;
wire n45774;
wire n45775;
wire n45776;
wire n45777;
wire n45778;
wire n45779;
wire n4578;
wire n45780;
wire n45782;
wire n45783;
wire n45784;
wire n45785;
wire n45786;
wire n45787;
wire n45788;
wire n4578_1;
wire n4579;
wire n45790;
wire n45791;
wire n45793;
wire n45794;
wire n45795;
wire n45796;
wire n45797;
wire n45798;
wire n45799;
wire n4580;
wire n45800;
wire n45802;
wire n45803;
wire n45805;
wire n45806;
wire n45808;
wire n45809;
wire n4581;
wire n45810;
wire n45811;
wire n45812;
wire n45813;
wire n45814;
wire n45815;
wire n45816;
wire n45817;
wire n45818;
wire n45819;
wire n4582;
wire n45820;
wire n45823;
wire n45824;
wire n45827;
wire n45828;
wire n45829;
wire n4583;
wire n45830;
wire n45831;
wire n45832;
wire n45833;
wire n45834;
wire n45835;
wire n45838;
wire n45839;
wire n4583_1;
wire n4584;
wire n45840;
wire n45841;
wire n45842;
wire n45843;
wire n45844;
wire n45845;
wire n45846;
wire n45847;
wire n4585;
wire n45850;
wire n45851;
wire n45853;
wire n45854;
wire n45855;
wire n45856;
wire n45857;
wire n45858;
wire n45859;
wire n4586;
wire n45861;
wire n45862;
wire n45863;
wire n45864;
wire n45865;
wire n45866;
wire n45868;
wire n45869;
wire n4587;
wire n45870;
wire n45871;
wire n45872;
wire n45875;
wire n45876;
wire n4588;
wire n45880;
wire n45881;
wire n45882;
wire n45883;
wire n45884;
wire n45885;
wire n45887;
wire n45889;
wire n4588_1;
wire n4589;
wire n45890;
wire n45891;
wire n45892;
wire n45893;
wire n45894;
wire n45895;
wire n45896;
wire n45897;
wire n45899;
wire n4590;
wire n45900;
wire n45901;
wire n45902;
wire n45903;
wire n45905;
wire n45906;
wire n45907;
wire n45908;
wire n45909;
wire n4591;
wire n45910;
wire n45911;
wire n45912;
wire n45914;
wire n45915;
wire n45917;
wire n45918;
wire n4592;
wire n45920;
wire n45921;
wire n45922;
wire n45923;
wire n45924;
wire n45925;
wire n45926;
wire n45927;
wire n45928;
wire n45929;
wire n4593;
wire n45931;
wire n45932;
wire n45933;
wire n45934;
wire n45935;
wire n45936;
wire n45937;
wire n45938;
wire n45939;
wire n4593_1;
wire n4594;
wire n45941;
wire n45942;
wire n45944;
wire n45945;
wire n45946;
wire n45947;
wire n45948;
wire n45949;
wire n4595;
wire n45950;
wire n45951;
wire n45952;
wire n45953;
wire n45954;
wire n45955;
wire n45956;
wire n45958;
wire n45959;
wire n4596;
wire n45960;
wire n45961;
wire n45962;
wire n45963;
wire n45964;
wire n45965;
wire n45967;
wire n45968;
wire n45969;
wire n4597;
wire n45971;
wire n45972;
wire n45973;
wire n45974;
wire n45975;
wire n45976;
wire n45978;
wire n45979;
wire n4598;
wire n45980;
wire n45981;
wire n45983;
wire n45984;
wire n45985;
wire n45987;
wire n45988;
wire n45989;
wire n4598_1;
wire n4599;
wire n45990;
wire n45991;
wire n45992;
wire n45994;
wire n45995;
wire n45996;
wire n45997;
wire n45998;
wire n45999;
wire n4600;
wire n46000;
wire n46001;
wire n46003;
wire n46004;
wire n46005;
wire n46006;
wire n46008;
wire n46009;
wire n4601;
wire n46010;
wire n46011;
wire n46012;
wire n46013;
wire n46014;
wire n46015;
wire n46017;
wire n46018;
wire n46019;
wire n4602;
wire n46020;
wire n46021;
wire n46023;
wire n46024;
wire n46026;
wire n46027;
wire n46029;
wire n4603;
wire n46030;
wire n46031;
wire n46032;
wire n46033;
wire n46034;
wire n46035;
wire n46037;
wire n46038;
wire n46039;
wire n4603_1;
wire n4604;
wire n46040;
wire n46041;
wire n46042;
wire n46043;
wire n46045;
wire n46046;
wire n46048;
wire n46049;
wire n4605;
wire n46050;
wire n46051;
wire n46052;
wire n46053;
wire n46054;
wire n46055;
wire n46056;
wire n46058;
wire n46059;
wire n4606;
wire n46061;
wire n46062;
wire n46063;
wire n46064;
wire n46065;
wire n46068;
wire n46069;
wire n4607;
wire n46070;
wire n46071;
wire n46073;
wire n46074;
wire n46075;
wire n46076;
wire n46078;
wire n46079;
wire n4608;
wire n46080;
wire n46081;
wire n46082;
wire n46083;
wire n46084;
wire n46085;
wire n46086;
wire n46088;
wire n46089;
wire n4608_1;
wire n4609;
wire n46090;
wire n46091;
wire n46093;
wire n46095;
wire n46096;
wire n46097;
wire n46098;
wire n46099;
wire n4610;
wire n46102;
wire n46103;
wire n46104;
wire n46105;
wire n46106;
wire n46107;
wire n46109;
wire n4611;
wire n46110;
wire n46111;
wire n46112;
wire n46113;
wire n46114;
wire n46115;
wire n46117;
wire n46118;
wire n46119;
wire n4612;
wire n46120;
wire n46122;
wire n46123;
wire n46124;
wire n46125;
wire n46126;
wire n46127;
wire n46128;
wire n46129;
wire n4613;
wire n46130;
wire n46133;
wire n46134;
wire n46135;
wire n46136;
wire n46137;
wire n46138;
wire n46139;
wire n4613_1;
wire n4614;
wire n46140;
wire n46141;
wire n46143;
wire n46144;
wire n46145;
wire n46146;
wire n46147;
wire n46148;
wire n46149;
wire n4615;
wire n46151;
wire n46152;
wire n46153;
wire n46154;
wire n46156;
wire n46157;
wire n46158;
wire n46159;
wire n4616;
wire n46160;
wire n46161;
wire n46163;
wire n46164;
wire n46166;
wire n46167;
wire n46169;
wire n4617;
wire n46170;
wire n46171;
wire n46172;
wire n46173;
wire n46174;
wire n46175;
wire n46176;
wire n46177;
wire n46178;
wire n46179;
wire n4618;
wire n46181;
wire n46182;
wire n46184;
wire n46185;
wire n46186;
wire n46187;
wire n46189;
wire n4618_1;
wire n4619;
wire n46190;
wire n46192;
wire n46193;
wire n46195;
wire n46196;
wire n46197;
wire n46198;
wire n462;
wire n4620;
wire n46200;
wire n46201;
wire n46202;
wire n46203;
wire n46204;
wire n46205;
wire n46206;
wire n46208;
wire n46209;
wire n4621;
wire n46210;
wire n46211;
wire n46213;
wire n46214;
wire n46215;
wire n46216;
wire n46218;
wire n46219;
wire n4622;
wire n46220;
wire n46221;
wire n46223;
wire n46224;
wire n46225;
wire n46226;
wire n46227;
wire n46228;
wire n46229;
wire n4623;
wire n46230;
wire n46231;
wire n46232;
wire n46233;
wire n46235;
wire n46236;
wire n46237;
wire n46239;
wire n4623_1;
wire n4624;
wire n46240;
wire n46241;
wire n46242;
wire n46243;
wire n46244;
wire n46245;
wire n46246;
wire n46247;
wire n46249;
wire n4625;
wire n46250;
wire n46251;
wire n46252;
wire n46253;
wire n46254;
wire n46256;
wire n46258;
wire n46259;
wire n4626;
wire n46261;
wire n46262;
wire n46263;
wire n46264;
wire n46266;
wire n46267;
wire n46268;
wire n46269;
wire n4627;
wire n46270;
wire n46272;
wire n46273;
wire n46274;
wire n46275;
wire n46276;
wire n46278;
wire n46279;
wire n4628;
wire n46281;
wire n46284;
wire n46285;
wire n46286;
wire n46287;
wire n46288;
wire n46289;
wire n4628_1;
wire n4629;
wire n46290;
wire n46293;
wire n46294;
wire n46295;
wire n46296;
wire n46297;
wire n46298;
wire n4630;
wire n46300;
wire n46301;
wire n46302;
wire n46303;
wire n46304;
wire n46305;
wire n46306;
wire n46307;
wire n46308;
wire n46309;
wire n4631;
wire n46310;
wire n46311;
wire n46312;
wire n46313;
wire n46314;
wire n46315;
wire n46316;
wire n46317;
wire n46318;
wire n46319;
wire n4632;
wire n46320;
wire n46321;
wire n46322;
wire n46324;
wire n46325;
wire n46326;
wire n46327;
wire n46329;
wire n4633;
wire n46330;
wire n46332;
wire n46333;
wire n46335;
wire n46336;
wire n46337;
wire n46338;
wire n46339;
wire n4633_1;
wire n4634;
wire n46340;
wire n46341;
wire n46342;
wire n46344;
wire n46345;
wire n46347;
wire n46348;
wire n4635;
wire n46350;
wire n46351;
wire n46352;
wire n46353;
wire n46354;
wire n46355;
wire n46356;
wire n46357;
wire n46359;
wire n4636;
wire n46360;
wire n46361;
wire n46362;
wire n46364;
wire n46365;
wire n46366;
wire n46367;
wire n46369;
wire n4637;
wire n46371;
wire n46372;
wire n46374;
wire n46375;
wire n46377;
wire n46378;
wire n4638;
wire n46380;
wire n46381;
wire n46382;
wire n46383;
wire n46384;
wire n46385;
wire n46388;
wire n46389;
wire n4638_1;
wire n4639;
wire n46390;
wire n46391;
wire n46393;
wire n46394;
wire n46395;
wire n46396;
wire n46397;
wire n46398;
wire n46399;
wire n4640;
wire n46400;
wire n46401;
wire n46404;
wire n46405;
wire n46407;
wire n46408;
wire n46409;
wire n4641;
wire n46410;
wire n46411;
wire n46412;
wire n46413;
wire n46414;
wire n46415;
wire n46417;
wire n46418;
wire n46419;
wire n4642;
wire n46420;
wire n46421;
wire n46422;
wire n46424;
wire n46425;
wire n46426;
wire n46427;
wire n46428;
wire n46429;
wire n4643;
wire n46431;
wire n46432;
wire n46433;
wire n46434;
wire n46435;
wire n46437;
wire n46438;
wire n4643_1;
wire n4644;
wire n46440;
wire n46441;
wire n46443;
wire n46444;
wire n46445;
wire n46446;
wire n46449;
wire n4645;
wire n46450;
wire n46451;
wire n46452;
wire n46453;
wire n46454;
wire n46455;
wire n46456;
wire n46457;
wire n46459;
wire n4646;
wire n46460;
wire n46462;
wire n46463;
wire n46465;
wire n46466;
wire n46467;
wire n46468;
wire n46469;
wire n4647;
wire n46470;
wire n46471;
wire n46472;
wire n46474;
wire n46475;
wire n46476;
wire n46477;
wire n46478;
wire n46479;
wire n4648;
wire n46481;
wire n46482;
wire n46483;
wire n46484;
wire n46486;
wire n46487;
wire n46489;
wire n4648_1;
wire n4649;
wire n46490;
wire n46491;
wire n46493;
wire n46494;
wire n46495;
wire n46496;
wire n46497;
wire n46498;
wire n46499;
wire n4650;
wire n46500;
wire n46501;
wire n46502;
wire n46503;
wire n46504;
wire n46506;
wire n46507;
wire n46508;
wire n46509;
wire n4651;
wire n46510;
wire n46511;
wire n46513;
wire n46515;
wire n46516;
wire n46517;
wire n46518;
wire n4652;
wire n46520;
wire n46521;
wire n46522;
wire n46523;
wire n46524;
wire n46525;
wire n46526;
wire n46528;
wire n46529;
wire n4652_1;
wire n4653;
wire n46530;
wire n46531;
wire n46532;
wire n46534;
wire n46535;
wire n46536;
wire n46537;
wire n46538;
wire n46539;
wire n4654;
wire n46540;
wire n46541;
wire n46542;
wire n46544;
wire n46546;
wire n46547;
wire n46548;
wire n46549;
wire n4655;
wire n46551;
wire n46552;
wire n46554;
wire n46555;
wire n46557;
wire n46558;
wire n46559;
wire n4656;
wire n46560;
wire n46561;
wire n46563;
wire n46564;
wire n46565;
wire n46566;
wire n46567;
wire n46568;
wire n46569;
wire n4657;
wire n46570;
wire n46571;
wire n46573;
wire n46575;
wire n46576;
wire n46578;
wire n46579;
wire n4657_1;
wire n4658;
wire n46580;
wire n46581;
wire n46582;
wire n46584;
wire n46586;
wire n46587;
wire n46588;
wire n46589;
wire n4659;
wire n46591;
wire n46592;
wire n46594;
wire n46595;
wire n46596;
wire n46597;
wire n46598;
wire n46599;
wire n4660;
wire n46600;
wire n46601;
wire n46603;
wire n46604;
wire n46606;
wire n46607;
wire n46608;
wire n46609;
wire n4661;
wire n46610;
wire n46611;
wire n46612;
wire n46614;
wire n46615;
wire n46617;
wire n46618;
wire n46619;
wire n4662;
wire n46620;
wire n46621;
wire n46622;
wire n46623;
wire n46624;
wire n46625;
wire n46627;
wire n46628;
wire n46629;
wire n4662_1;
wire n4663;
wire n46630;
wire n46631;
wire n46632;
wire n46633;
wire n46634;
wire n46636;
wire n46637;
wire n46639;
wire n4664;
wire n46640;
wire n46642;
wire n46643;
wire n46644;
wire n46645;
wire n46646;
wire n46648;
wire n4665;
wire n46650;
wire n46651;
wire n46653;
wire n46654;
wire n46655;
wire n46656;
wire n46658;
wire n46659;
wire n4666;
wire n46660;
wire n46661;
wire n46663;
wire n46664;
wire n46665;
wire n46666;
wire n46668;
wire n46669;
wire n4667;
wire n46670;
wire n46671;
wire n46672;
wire n46673;
wire n46674;
wire n46675;
wire n46676;
wire n46677;
wire n46678;
wire n46679;
wire n4667_1;
wire n4668;
wire n46681;
wire n46682;
wire n46684;
wire n46685;
wire n46686;
wire n46687;
wire n46688;
wire n46689;
wire n4669;
wire n46690;
wire n46691;
wire n46692;
wire n46693;
wire n46694;
wire n46695;
wire n46696;
wire n46698;
wire n46699;
wire n467;
wire n4670;
wire n46700;
wire n46701;
wire n46702;
wire n46703;
wire n46704;
wire n46706;
wire n46707;
wire n46708;
wire n46709;
wire n4671;
wire n46710;
wire n46712;
wire n46713;
wire n46715;
wire n46716;
wire n46718;
wire n46719;
wire n4672;
wire n46720;
wire n46721;
wire n46722;
wire n46723;
wire n46724;
wire n46726;
wire n46727;
wire n46728;
wire n46729;
wire n4672_1;
wire n4673;
wire n46731;
wire n46732;
wire n46733;
wire n46734;
wire n46735;
wire n46736;
wire n46738;
wire n46739;
wire n4674;
wire n46741;
wire n46743;
wire n46744;
wire n46745;
wire n46746;
wire n46747;
wire n46748;
wire n4675;
wire n46750;
wire n46751;
wire n46753;
wire n46754;
wire n46755;
wire n46756;
wire n46757;
wire n46758;
wire n4676;
wire n46760;
wire n46761;
wire n46763;
wire n46764;
wire n46766;
wire n46767;
wire n46768;
wire n46769;
wire n4677;
wire n46770;
wire n46771;
wire n46772;
wire n46773;
wire n46775;
wire n46776;
wire n46778;
wire n46779;
wire n4677_1;
wire n4678;
wire n46780;
wire n46781;
wire n46783;
wire n46785;
wire n46786;
wire n46788;
wire n46789;
wire n4679;
wire n46791;
wire n46792;
wire n46793;
wire n46794;
wire n46795;
wire n46796;
wire n46797;
wire n46798;
wire n46799;
wire n4680;
wire n46802;
wire n46803;
wire n46805;
wire n46806;
wire n46807;
wire n46808;
wire n46809;
wire n4681;
wire n46810;
wire n46812;
wire n46813;
wire n46814;
wire n46815;
wire n46817;
wire n46818;
wire n46819;
wire n4682;
wire n46820;
wire n46821;
wire n46822;
wire n46824;
wire n46825;
wire n46826;
wire n46827;
wire n46828;
wire n46829;
wire n4682_1;
wire n4683;
wire n46830;
wire n46831;
wire n46832;
wire n46833;
wire n46834;
wire n46835;
wire n46836;
wire n46837;
wire n46839;
wire n4684;
wire n46840;
wire n46842;
wire n46843;
wire n46844;
wire n46845;
wire n46846;
wire n46849;
wire n4685;
wire n46850;
wire n46851;
wire n46852;
wire n46853;
wire n46854;
wire n46855;
wire n46856;
wire n46859;
wire n4686;
wire n46860;
wire n46861;
wire n46863;
wire n46864;
wire n46865;
wire n46866;
wire n46868;
wire n46869;
wire n4687;
wire n46871;
wire n46872;
wire n46874;
wire n46875;
wire n46876;
wire n46877;
wire n46879;
wire n4687_1;
wire n4688;
wire n46880;
wire n46881;
wire n46882;
wire n46883;
wire n46884;
wire n46885;
wire n46886;
wire n46887;
wire n46889;
wire n4689;
wire n46890;
wire n46891;
wire n46892;
wire n46893;
wire n46894;
wire n46895;
wire n46896;
wire n46897;
wire n46899;
wire n4690;
wire n46900;
wire n46901;
wire n46902;
wire n46903;
wire n46906;
wire n46907;
wire n46908;
wire n46909;
wire n4691;
wire n46910;
wire n46911;
wire n46912;
wire n46913;
wire n46914;
wire n46915;
wire n46916;
wire n46918;
wire n46919;
wire n4692;
wire n46920;
wire n46921;
wire n46922;
wire n46923;
wire n46924;
wire n46925;
wire n46926;
wire n46927;
wire n46929;
wire n4692_1;
wire n4693;
wire n46930;
wire n46931;
wire n46932;
wire n46933;
wire n46934;
wire n46935;
wire n46936;
wire n46938;
wire n46939;
wire n4694;
wire n46941;
wire n46942;
wire n46943;
wire n46944;
wire n46945;
wire n46946;
wire n46947;
wire n46949;
wire n4695;
wire n46950;
wire n46951;
wire n46952;
wire n46954;
wire n46955;
wire n46956;
wire n46957;
wire n46958;
wire n46959;
wire n4696;
wire n46961;
wire n46962;
wire n46963;
wire n46964;
wire n46966;
wire n46967;
wire n46969;
wire n4697;
wire n46970;
wire n46971;
wire n46972;
wire n46973;
wire n46974;
wire n46975;
wire n46976;
wire n46977;
wire n46978;
wire n46979;
wire n4697_1;
wire n4698;
wire n46980;
wire n46981;
wire n46982;
wire n46983;
wire n46984;
wire n46985;
wire n46986;
wire n46987;
wire n46988;
wire n46989;
wire n4699;
wire n46991;
wire n46992;
wire n46993;
wire n46994;
wire n46995;
wire n46996;
wire n46997;
wire n46998;
wire n46999;
wire n4700;
wire n47000;
wire n47001;
wire n47003;
wire n47004;
wire n47006;
wire n47007;
wire n47009;
wire n4701;
wire n47010;
wire n47011;
wire n47013;
wire n47014;
wire n47016;
wire n47017;
wire n47018;
wire n47019;
wire n4702;
wire n47021;
wire n47022;
wire n47023;
wire n47024;
wire n47026;
wire n47027;
wire n47028;
wire n4702_1;
wire n4703;
wire n47031;
wire n47032;
wire n47033;
wire n47034;
wire n47036;
wire n47037;
wire n47038;
wire n4704;
wire n47040;
wire n47041;
wire n47042;
wire n47043;
wire n47045;
wire n47046;
wire n47048;
wire n47049;
wire n4705;
wire n47051;
wire n47052;
wire n47053;
wire n47054;
wire n47055;
wire n47057;
wire n47058;
wire n47059;
wire n4706;
wire n47060;
wire n47062;
wire n47063;
wire n47065;
wire n47066;
wire n47067;
wire n47068;
wire n47069;
wire n4707;
wire n47071;
wire n47072;
wire n47073;
wire n47074;
wire n47075;
wire n47077;
wire n47078;
wire n47079;
wire n4707_1;
wire n4708;
wire n47080;
wire n47081;
wire n47082;
wire n47083;
wire n47085;
wire n47086;
wire n47088;
wire n47089;
wire n4709;
wire n47090;
wire n47091;
wire n47092;
wire n47093;
wire n47094;
wire n47096;
wire n47097;
wire n47098;
wire n47099;
wire n4710;
wire n47100;
wire n47101;
wire n47102;
wire n47103;
wire n47104;
wire n47106;
wire n47107;
wire n47108;
wire n47109;
wire n4711;
wire n47110;
wire n47111;
wire n47113;
wire n47114;
wire n47115;
wire n47116;
wire n47117;
wire n47118;
wire n47119;
wire n4712;
wire n47120;
wire n47122;
wire n47123;
wire n47125;
wire n47126;
wire n47128;
wire n47129;
wire n4712_1;
wire n4713;
wire n47131;
wire n47132;
wire n47133;
wire n47134;
wire n47135;
wire n47136;
wire n47138;
wire n47139;
wire n4714;
wire n47142;
wire n47143;
wire n47145;
wire n47146;
wire n47147;
wire n47148;
wire n47149;
wire n4715;
wire n47150;
wire n47151;
wire n47152;
wire n47154;
wire n47155;
wire n47156;
wire n47157;
wire n47158;
wire n47159;
wire n4716;
wire n47160;
wire n47162;
wire n47163;
wire n47165;
wire n47166;
wire n47168;
wire n47169;
wire n4717;
wire n47172;
wire n47173;
wire n47174;
wire n47175;
wire n47177;
wire n47178;
wire n47179;
wire n4717_1;
wire n4718;
wire n47180;
wire n47181;
wire n47182;
wire n47183;
wire n47184;
wire n47185;
wire n47186;
wire n47187;
wire n47189;
wire n4719;
wire n47191;
wire n47192;
wire n47193;
wire n47194;
wire n47196;
wire n47197;
wire n47198;
wire n47199;
wire n472;
wire n4720;
wire n47200;
wire n47201;
wire n47203;
wire n47204;
wire n47205;
wire n47206;
wire n47208;
wire n47209;
wire n4721;
wire n47210;
wire n47211;
wire n47213;
wire n47214;
wire n47215;
wire n47216;
wire n47218;
wire n47219;
wire n4722;
wire n47221;
wire n47222;
wire n47223;
wire n47224;
wire n47226;
wire n47227;
wire n47228;
wire n47229;
wire n4722_1;
wire n4723;
wire n47232;
wire n47233;
wire n47234;
wire n47235;
wire n47236;
wire n47238;
wire n47239;
wire n4724;
wire n47240;
wire n47241;
wire n47242;
wire n47243;
wire n47244;
wire n47246;
wire n47247;
wire n47248;
wire n47249;
wire n4725;
wire n47250;
wire n47251;
wire n47252;
wire n47256;
wire n47257;
wire n47259;
wire n4726;
wire n47260;
wire n47261;
wire n47262;
wire n47264;
wire n47265;
wire n47266;
wire n47267;
wire n47268;
wire n47269;
wire n4727;
wire n47270;
wire n47271;
wire n47272;
wire n47273;
wire n47274;
wire n47276;
wire n47277;
wire n47278;
wire n47279;
wire n4727_1;
wire n4728;
wire n47280;
wire n47281;
wire n47282;
wire n47283;
wire n47284;
wire n47286;
wire n47287;
wire n47288;
wire n47289;
wire n4729;
wire n47290;
wire n47291;
wire n47292;
wire n47293;
wire n47294;
wire n47295;
wire n47296;
wire n47298;
wire n4730;
wire n47300;
wire n47301;
wire n47303;
wire n47304;
wire n47305;
wire n47306;
wire n47308;
wire n47309;
wire n4731;
wire n47311;
wire n47312;
wire n47314;
wire n47315;
wire n47317;
wire n47318;
wire n4732;
wire n47320;
wire n47321;
wire n47323;
wire n47325;
wire n47326;
wire n47327;
wire n47328;
wire n4732_1;
wire n4733;
wire n47330;
wire n47331;
wire n47332;
wire n47333;
wire n47334;
wire n47335;
wire n47337;
wire n47338;
wire n4734;
wire n47340;
wire n47341;
wire n47342;
wire n47343;
wire n47345;
wire n47346;
wire n47347;
wire n47348;
wire n47349;
wire n4735;
wire n47351;
wire n47352;
wire n47354;
wire n47355;
wire n47357;
wire n47358;
wire n47359;
wire n4736;
wire n47360;
wire n47361;
wire n47363;
wire n47364;
wire n47365;
wire n47366;
wire n47367;
wire n47368;
wire n47369;
wire n4736_1;
wire n4737;
wire n47370;
wire n47372;
wire n47373;
wire n47374;
wire n47375;
wire n47376;
wire n47378;
wire n47379;
wire n4738;
wire n47380;
wire n47381;
wire n47382;
wire n47384;
wire n47386;
wire n47387;
wire n47388;
wire n47389;
wire n4739;
wire n47390;
wire n47391;
wire n47393;
wire n47394;
wire n47396;
wire n47397;
wire n47398;
wire n4740;
wire n47400;
wire n47401;
wire n47402;
wire n47403;
wire n47404;
wire n47405;
wire n47406;
wire n47407;
wire n47409;
wire n4741;
wire n47410;
wire n47411;
wire n47412;
wire n47413;
wire n47414;
wire n47415;
wire n47417;
wire n47418;
wire n4741_1;
wire n4742;
wire n47421;
wire n47422;
wire n47423;
wire n47424;
wire n47425;
wire n47426;
wire n47427;
wire n47428;
wire n4743;
wire n47430;
wire n47431;
wire n47432;
wire n47433;
wire n47434;
wire n47435;
wire n47437;
wire n47438;
wire n4744;
wire n47440;
wire n47441;
wire n47443;
wire n47444;
wire n47446;
wire n47447;
wire n47448;
wire n47449;
wire n4745;
wire n47450;
wire n47451;
wire n47453;
wire n47454;
wire n47455;
wire n47456;
wire n47457;
wire n47458;
wire n47459;
wire n4746;
wire n47460;
wire n47461;
wire n47462;
wire n47464;
wire n47465;
wire n47467;
wire n47468;
wire n47469;
wire n4746_1;
wire n4747;
wire n47470;
wire n47471;
wire n47472;
wire n47473;
wire n47474;
wire n47475;
wire n47476;
wire n47477;
wire n47478;
wire n47479;
wire n4748;
wire n47480;
wire n47481;
wire n47484;
wire n47485;
wire n47486;
wire n47487;
wire n47488;
wire n47489;
wire n4749;
wire n47491;
wire n47492;
wire n47493;
wire n47494;
wire n47495;
wire n47496;
wire n47497;
wire n47498;
wire n4750;
wire n47500;
wire n47501;
wire n47502;
wire n47503;
wire n47504;
wire n47506;
wire n47507;
wire n47509;
wire n4751;
wire n47510;
wire n47511;
wire n47512;
wire n47514;
wire n47515;
wire n47516;
wire n47517;
wire n47519;
wire n4751_1;
wire n4752;
wire n47520;
wire n47521;
wire n47522;
wire n47523;
wire n47524;
wire n47526;
wire n47527;
wire n47528;
wire n47529;
wire n4753;
wire n47530;
wire n47531;
wire n47532;
wire n47533;
wire n47534;
wire n47537;
wire n47538;
wire n47539;
wire n4754;
wire n47540;
wire n47542;
wire n47543;
wire n47545;
wire n47546;
wire n47548;
wire n47549;
wire n4755;
wire n47550;
wire n47551;
wire n47552;
wire n47553;
wire n47554;
wire n47555;
wire n47557;
wire n47558;
wire n4756;
wire n47560;
wire n47561;
wire n47562;
wire n47563;
wire n47564;
wire n47566;
wire n47567;
wire n4756_1;
wire n4757;
wire n4758;
wire n4759;
wire n476;
wire n4760;
wire n4761;
wire n4761_1;
wire n4762;
wire n4763;
wire n4764;
wire n4765;
wire n4766;
wire n4766_1;
wire n4767;
wire n4768;
wire n4769;
wire n4770;
wire n4771;
wire n4771_1;
wire n4772;
wire n4773;
wire n4774;
wire n4775;
wire n4776;
wire n4776_1;
wire n4777;
wire n4778;
wire n4779;
wire n4780;
wire n4781;
wire n4781_1;
wire n4782;
wire n4783;
wire n4784;
wire n4785;
wire n4786;
wire n4786_1;
wire n4787;
wire n4788;
wire n4789;
wire n4790;
wire n4791;
wire n4791_1;
wire n4792;
wire n4793;
wire n4794;
wire n4795;
wire n4796;
wire n4796_1;
wire n4797;
wire n4798;
wire n4799;
wire n4800;
wire n4801;
wire n4801_1;
wire n4802;
wire n4803;
wire n4804;
wire n4805;
wire n4806;
wire n4806_1;
wire n4807;
wire n4808;
wire n4809;
wire n481;
wire n4810;
wire n4810_1;
wire n4811;
wire n4812;
wire n4813;
wire n4814;
wire n4815;
wire n4815_1;
wire n4816;
wire n4817;
wire n4818;
wire n4819;
wire n4820;
wire n4820_1;
wire n4821;
wire n4822;
wire n4823;
wire n4824;
wire n4825;
wire n4825_1;
wire n4826;
wire n4827;
wire n4828;
wire n4829;
wire n4829_1;
wire n4830;
wire n4831;
wire n4832;
wire n4833;
wire n4834;
wire n4834_1;
wire n4835;
wire n4836;
wire n4837;
wire n4838;
wire n4839;
wire n4839_1;
wire n4840;
wire n4841;
wire n4842;
wire n4843;
wire n4843_1;
wire n4844;
wire n4845;
wire n4846;
wire n4847;
wire n4848;
wire n4848_1;
wire n4849;
wire n485;
wire n4850;
wire n4851;
wire n4852;
wire n4853;
wire n4853_1;
wire n4854;
wire n4855;
wire n4856;
wire n4857;
wire n4858;
wire n4858_1;
wire n4859;
wire n4860;
wire n4861;
wire n4862;
wire n4863;
wire n4863_1;
wire n4864;
wire n4865;
wire n4866;
wire n4867;
wire n4868;
wire n4868_1;
wire n4869;
wire n4870;
wire n4871;
wire n4872;
wire n4873;
wire n4873_1;
wire n4874;
wire n4875;
wire n4876;
wire n4877;
wire n4878;
wire n4878_1;
wire n4879;
wire n4880;
wire n4881;
wire n4882;
wire n4883;
wire n4883_1;
wire n4884;
wire n4885;
wire n4886;
wire n4887;
wire n4888;
wire n4888_1;
wire n4889;
wire n4890;
wire n4891;
wire n4892;
wire n4893;
wire n4893_1;
wire n4894;
wire n4895;
wire n4896;
wire n4897;
wire n4897_1;
wire n4898;
wire n4899;
wire n490;
wire n4900;
wire n4901;
wire n4902;
wire n4902_1;
wire n4903;
wire n4904;
wire n4905;
wire n4906;
wire n4907;
wire n4907_1;
wire n4908;
wire n4909;
wire n4910;
wire n4911;
wire n4912;
wire n4912_1;
wire n4913;
wire n4914;
wire n4915;
wire n4916;
wire n4917;
wire n4917_1;
wire n4918;
wire n4919;
wire n4920;
wire n4921;
wire n4922;
wire n4922_1;
wire n4923;
wire n4924;
wire n4925;
wire n4926;
wire n4927;
wire n4927_1;
wire n4928;
wire n4929;
wire n4930;
wire n4931;
wire n4932;
wire n4932_1;
wire n4933;
wire n4934;
wire n4935;
wire n4936;
wire n4937;
wire n4937_1;
wire n4938;
wire n4939;
wire n4940;
wire n4941;
wire n4942;
wire n4942_1;
wire n4943;
wire n4944;
wire n4945;
wire n4946;
wire n4947;
wire n4947_1;
wire n4948;
wire n4949;
wire n495;
wire n4950;
wire n4951;
wire n4952;
wire n4952_1;
wire n4953;
wire n4954;
wire n4955;
wire n4956;
wire n4957;
wire n4957_1;
wire n4958;
wire n4959;
wire n4960;
wire n4961;
wire n4962;
wire n4962_1;
wire n4963;
wire n4964;
wire n4965;
wire n4966;
wire n4967;
wire n4967_1;
wire n4968;
wire n4969;
wire n4970;
wire n4971;
wire n4972;
wire n4972_1;
wire n4973;
wire n4974;
wire n4975;
wire n4976;
wire n4977;
wire n4977_1;
wire n4978;
wire n4979;
wire n4980;
wire n4981;
wire n4982;
wire n4982_1;
wire n4983;
wire n4984;
wire n4985;
wire n4986;
wire n4987;
wire n4987_1;
wire n4988;
wire n4989;
wire n4990;
wire n4991;
wire n4992;
wire n4992_1;
wire n4993;
wire n4994;
wire n4995;
wire n4997;
wire n4997_1;
wire n4998;
wire n4999;
wire n500;
wire n5000;
wire n5001;
wire n5001_1;
wire n5002;
wire n5003;
wire n5004;
wire n5005;
wire n5006;
wire n5006_1;
wire n5007;
wire n5008;
wire n5009;
wire n5010;
wire n5011;
wire n5011_1;
wire n5012;
wire n5013;
wire n5014;
wire n5015;
wire n5016;
wire n5016_1;
wire n5017;
wire n5018;
wire n5019;
wire n5020;
wire n5021;
wire n5021_1;
wire n5022;
wire n5023;
wire n5024;
wire n5025;
wire n5026;
wire n5026_1;
wire n5027;
wire n5028;
wire n5029;
wire n5030;
wire n5031;
wire n5031_1;
wire n5032;
wire n5033;
wire n5034;
wire n5035;
wire n5036;
wire n5036_1;
wire n5037;
wire n5038;
wire n5039;
wire n5040;
wire n5041;
wire n5041_1;
wire n5042;
wire n5043;
wire n5044;
wire n5045;
wire n5046;
wire n5046_1;
wire n5047;
wire n5048;
wire n5049;
wire n505;
wire n5050;
wire n5051;
wire n5051_1;
wire n5052;
wire n5053;
wire n5054;
wire n5055;
wire n5056;
wire n5056_1;
wire n5057;
wire n5058;
wire n5059;
wire n5060;
wire n5061;
wire n5061_1;
wire n5062;
wire n5063;
wire n5064;
wire n5065;
wire n5066;
wire n5066_1;
wire n5067;
wire n5068;
wire n5069;
wire n5070;
wire n5070_1;
wire n5071;
wire n5072;
wire n5073;
wire n5074;
wire n5075;
wire n5075_1;
wire n5076;
wire n5077;
wire n5078;
wire n5079;
wire n5080;
wire n5080_1;
wire n5081;
wire n5082;
wire n5083;
wire n5084;
wire n5085;
wire n5085_1;
wire n5086;
wire n5087;
wire n5088;
wire n5089;
wire n509;
wire n5090;
wire n5090_1;
wire n5091;
wire n5092;
wire n5093;
wire n5094;
wire n5095;
wire n5095_1;
wire n5096;
wire n5097;
wire n5098;
wire n5099;
wire n5100;
wire n5100_1;
wire n5101;
wire n5102;
wire n5103;
wire n5104;
wire n5105;
wire n5105_1;
wire n5106;
wire n5107;
wire n5108;
wire n5109;
wire n5110;
wire n5110_1;
wire n5111;
wire n5112;
wire n5113;
wire n5114;
wire n5115;
wire n5115_1;
wire n5116;
wire n5117;
wire n5118;
wire n5119;
wire n5120;
wire n5120_1;
wire n5121;
wire n5122;
wire n5123;
wire n5124;
wire n5125;
wire n5125_1;
wire n5126;
wire n5127;
wire n5128;
wire n5129;
wire n5130;
wire n5130_1;
wire n5131;
wire n5132;
wire n5133;
wire n5134;
wire n5135;
wire n5135_1;
wire n5136;
wire n5137;
wire n5138;
wire n5139;
wire n514;
wire n5140;
wire n5140_1;
wire n5141;
wire n5142;
wire n5143;
wire n5144;
wire n5145;
wire n5145_1;
wire n5146;
wire n5147;
wire n5148;
wire n5149;
wire n5150;
wire n5150_1;
wire n5151;
wire n5152;
wire n5153;
wire n5154;
wire n5155;
wire n5155_1;
wire n5156;
wire n5157;
wire n5158;
wire n5159;
wire n5160;
wire n5160_1;
wire n5161;
wire n5162;
wire n5163;
wire n5164;
wire n5165;
wire n5165_1;
wire n5166;
wire n5167;
wire n5168;
wire n5169;
wire n5170;
wire n5170_1;
wire n5171;
wire n5172;
wire n5173;
wire n5174;
wire n5175;
wire n5175_1;
wire n5176;
wire n5177;
wire n5178;
wire n5179;
wire n5180;
wire n5180_1;
wire n5181;
wire n5182;
wire n5183;
wire n5184;
wire n5185;
wire n5185_1;
wire n5186;
wire n5187;
wire n5188;
wire n5189;
wire n519;
wire n5190;
wire n5190_1;
wire n5191;
wire n5192;
wire n5193;
wire n5194;
wire n5195;
wire n5195_1;
wire n5196;
wire n5197;
wire n5198;
wire n5199;
wire n5200;
wire n5200_1;
wire n5201;
wire n5202;
wire n5203;
wire n5204;
wire n5205;
wire n5205_1;
wire n5206;
wire n5207;
wire n5208;
wire n5209;
wire n5210;
wire n5210_1;
wire n5211;
wire n5212;
wire n5213;
wire n5214;
wire n5215;
wire n5215_1;
wire n5216;
wire n5217;
wire n5218;
wire n5219;
wire n5220;
wire n5220_1;
wire n5221;
wire n5222;
wire n5223;
wire n5224;
wire n5225;
wire n5225_1;
wire n5226;
wire n5227;
wire n5228;
wire n5229;
wire n5230;
wire n5230_1;
wire n5231;
wire n5232;
wire n5233;
wire n5234;
wire n5235;
wire n5235_1;
wire n5236;
wire n5237;
wire n5238;
wire n5239;
wire n524;
wire n5240;
wire n5240_1;
wire n5241;
wire n5242;
wire n5243;
wire n5244;
wire n5245;
wire n5245_1;
wire n5246;
wire n5247;
wire n5248;
wire n5249;
wire n5250;
wire n5250_1;
wire n5251;
wire n5252;
wire n5253;
wire n5254;
wire n5255;
wire n5255_1;
wire n5256;
wire n5257;
wire n5258;
wire n5259;
wire n5260;
wire n5260_1;
wire n5261;
wire n5262;
wire n5263;
wire n5264;
wire n5265;
wire n5265_1;
wire n5266;
wire n5267;
wire n5268;
wire n5269;
wire n5270;
wire n5270_1;
wire n5271;
wire n5272;
wire n5273;
wire n5274;
wire n5275;
wire n5275_1;
wire n5276;
wire n5277;
wire n5278;
wire n5279;
wire n5280;
wire n5280_1;
wire n5281;
wire n5282;
wire n5283;
wire n5284;
wire n5285;
wire n5285_1;
wire n5286;
wire n5287;
wire n5288;
wire n5289;
wire n529;
wire n5290;
wire n5290_1;
wire n5291;
wire n5292;
wire n5293;
wire n5294;
wire n5295;
wire n5295_1;
wire n5296;
wire n5297;
wire n5298;
wire n5299;
wire n5300;
wire n5300_1;
wire n5301;
wire n5302;
wire n5303;
wire n5304;
wire n5305;
wire n5305_1;
wire n5306;
wire n5307;
wire n5308;
wire n5309;
wire n5310;
wire n5310_1;
wire n5311;
wire n5312;
wire n5313;
wire n5314;
wire n5315;
wire n5315_1;
wire n5316;
wire n5317;
wire n5318;
wire n5319;
wire n5320;
wire n5320_1;
wire n5321;
wire n5322;
wire n5323;
wire n5324;
wire n5325;
wire n5325_1;
wire n5326;
wire n5327;
wire n5328;
wire n5329;
wire n5330;
wire n5330_1;
wire n5331;
wire n5332;
wire n5333;
wire n5334;
wire n5335;
wire n5335_1;
wire n5336;
wire n5337;
wire n5338;
wire n5339;
wire n534;
wire n5340;
wire n5340_1;
wire n5341;
wire n5342;
wire n5343;
wire n5344;
wire n5345;
wire n5345_1;
wire n5346;
wire n5347;
wire n5348;
wire n5349;
wire n5350;
wire n5350_1;
wire n5351;
wire n5352;
wire n5353;
wire n5354;
wire n5355;
wire n5355_1;
wire n5356;
wire n5357;
wire n5358;
wire n5359;
wire n5360;
wire n5360_1;
wire n5361;
wire n5362;
wire n5363;
wire n5364;
wire n5365;
wire n5365_1;
wire n5366;
wire n5367;
wire n5368;
wire n5369;
wire n5370;
wire n5370_1;
wire n5371;
wire n5372;
wire n5373;
wire n5374;
wire n5375;
wire n5375_1;
wire n5376;
wire n5377;
wire n5378;
wire n5379;
wire n5380;
wire n5380_1;
wire n5381;
wire n5382;
wire n5383;
wire n5384;
wire n5385;
wire n5385_1;
wire n5386;
wire n5387;
wire n5388;
wire n5389;
wire n539;
wire n5390;
wire n5390_1;
wire n5391;
wire n5392;
wire n5393;
wire n5394;
wire n5395;
wire n5395_1;
wire n5396;
wire n5397;
wire n5398;
wire n5399;
wire n5400;
wire n5400_1;
wire n5401;
wire n5402;
wire n5403;
wire n5404;
wire n5405;
wire n5405_1;
wire n5406;
wire n5407;
wire n5408;
wire n5409;
wire n5410;
wire n5410_1;
wire n5411;
wire n5412;
wire n5413;
wire n5414;
wire n5415;
wire n5415_1;
wire n5416;
wire n5417;
wire n5418;
wire n5419;
wire n5420;
wire n5420_1;
wire n5421;
wire n5422;
wire n5423;
wire n5424;
wire n5425;
wire n5425_1;
wire n5426;
wire n5427;
wire n5428;
wire n5429;
wire n5430;
wire n5430_1;
wire n5431;
wire n5432;
wire n5433;
wire n5434;
wire n5435;
wire n5435_1;
wire n5436;
wire n5437;
wire n5438;
wire n5439;
wire n544;
wire n5440;
wire n5440_1;
wire n5441;
wire n5442;
wire n5443;
wire n5444;
wire n5445;
wire n5445_1;
wire n5446;
wire n5447;
wire n5448;
wire n5449;
wire n5450;
wire n5450_1;
wire n5451;
wire n5452;
wire n5453;
wire n5454;
wire n5455;
wire n5455_1;
wire n5456;
wire n5457;
wire n5458;
wire n5459;
wire n5459_1;
wire n5460;
wire n5461;
wire n5462;
wire n5463;
wire n5464;
wire n5464_1;
wire n5465;
wire n5466;
wire n5467;
wire n5468;
wire n5469;
wire n5469_1;
wire n5470;
wire n5471;
wire n5472;
wire n5473;
wire n5474;
wire n5474_1;
wire n5475;
wire n5476;
wire n5477;
wire n5478;
wire n5479;
wire n5479_1;
wire n5480;
wire n5481;
wire n5482;
wire n5483;
wire n5483_1;
wire n5484;
wire n5485;
wire n5486;
wire n5487;
wire n5488;
wire n5488_1;
wire n5489;
wire n549;
wire n5490;
wire n5491;
wire n5492;
wire n5493;
wire n5493_1;
wire n5494;
wire n5495;
wire n5496;
wire n5497;
wire n5498;
wire n5498_1;
wire n5499;
wire n5500;
wire n5501;
wire n5502;
wire n5503;
wire n5503_1;
wire n5504;
wire n5505;
wire n5506;
wire n5507;
wire n5508;
wire n5508_1;
wire n5509;
wire n5510;
wire n5511;
wire n5512;
wire n5513;
wire n5513_1;
wire n5514;
wire n5515;
wire n5516;
wire n5517;
wire n5518;
wire n5518_1;
wire n5519;
wire n5520;
wire n5521;
wire n5522;
wire n5523;
wire n5523_1;
wire n5524;
wire n5525;
wire n5526;
wire n5527;
wire n5528;
wire n5528_1;
wire n5529;
wire n5530;
wire n5531;
wire n5532;
wire n5533;
wire n5533_1;
wire n5534;
wire n5535;
wire n5536;
wire n5537;
wire n5538;
wire n5538_1;
wire n5539;
wire n554;
wire n5540;
wire n5541;
wire n5542;
wire n5543;
wire n5543_1;
wire n5544;
wire n5545;
wire n5546;
wire n5547;
wire n5548;
wire n5548_1;
wire n5549;
wire n5550;
wire n5551;
wire n5552;
wire n5553;
wire n5553_1;
wire n5554;
wire n5555;
wire n5556;
wire n5557;
wire n5558;
wire n5558_1;
wire n5559;
wire n5560;
wire n5561;
wire n5562;
wire n5563;
wire n5563_1;
wire n5564;
wire n5565;
wire n5566;
wire n5567;
wire n5568;
wire n5568_1;
wire n5569;
wire n5570;
wire n5571;
wire n5572;
wire n5573;
wire n5573_1;
wire n5574;
wire n5575;
wire n5576;
wire n5577;
wire n5578;
wire n5578_1;
wire n5579;
wire n5580;
wire n5581;
wire n5582;
wire n5583;
wire n5583_1;
wire n5584;
wire n5585;
wire n5586;
wire n5587;
wire n5588;
wire n5588_1;
wire n5589;
wire n559;
wire n5590;
wire n5591;
wire n5592;
wire n5593;
wire n5593_1;
wire n5594;
wire n5595;
wire n5596;
wire n5597;
wire n5598;
wire n5598_1;
wire n5599;
wire n5600;
wire n5601;
wire n5602;
wire n5603;
wire n5603_1;
wire n5604;
wire n5605;
wire n5606;
wire n5607;
wire n5608;
wire n5608_1;
wire n5609;
wire n5610;
wire n5611;
wire n5612;
wire n5613;
wire n5613_1;
wire n5614;
wire n5615;
wire n5616;
wire n5617;
wire n5618;
wire n5618_1;
wire n5619;
wire n5620;
wire n5621;
wire n5622;
wire n5623;
wire n5623_1;
wire n5624;
wire n5625;
wire n5626;
wire n5627;
wire n5628;
wire n5628_1;
wire n5629;
wire n5630;
wire n5631;
wire n5632;
wire n5633;
wire n5633_1;
wire n5634;
wire n5635;
wire n5636;
wire n5637;
wire n5638;
wire n5638_1;
wire n5639;
wire n564;
wire n5640;
wire n5641;
wire n5642;
wire n5643;
wire n5643_1;
wire n5644;
wire n5645;
wire n5646;
wire n5647;
wire n5648;
wire n5648_1;
wire n5649;
wire n5650;
wire n5651;
wire n5652;
wire n5653;
wire n5653_1;
wire n5654;
wire n5655;
wire n5656;
wire n5657;
wire n5657_1;
wire n5658;
wire n5659;
wire n5660;
wire n5661;
wire n5662;
wire n5662_1;
wire n5663;
wire n5664;
wire n5665;
wire n5666;
wire n5667;
wire n5667_1;
wire n5668;
wire n5669;
wire n5670;
wire n5671;
wire n5672;
wire n5672_1;
wire n5673;
wire n5674;
wire n5675;
wire n5676;
wire n5677;
wire n5677_1;
wire n5678;
wire n5679;
wire n5680;
wire n5681;
wire n5682;
wire n5682_1;
wire n5683;
wire n5684;
wire n5685;
wire n5686;
wire n5687;
wire n5687_1;
wire n5688;
wire n5689;
wire n569;
wire n5690;
wire n5691;
wire n5692;
wire n5692_1;
wire n5693;
wire n5694;
wire n5695;
wire n5696;
wire n5697;
wire n5697_1;
wire n5698;
wire n5699;
wire n5700;
wire n5701;
wire n5701_1;
wire n5702;
wire n5703;
wire n5704;
wire n5705;
wire n5706;
wire n5706_1;
wire n5707;
wire n5708;
wire n5709;
wire n5710;
wire n5711;
wire n5711_1;
wire n5712;
wire n5713;
wire n5714;
wire n5715;
wire n5716;
wire n5716_1;
wire n5717;
wire n5718;
wire n5719;
wire n5720;
wire n5721;
wire n5721_1;
wire n5722;
wire n5723;
wire n5724;
wire n5725;
wire n5726;
wire n5726_1;
wire n5727;
wire n5728;
wire n5729;
wire n5730;
wire n5730_1;
wire n5731;
wire n5732;
wire n5733;
wire n5734;
wire n5735;
wire n5735_1;
wire n5736;
wire n5737;
wire n5738;
wire n5739;
wire n574;
wire n5740;
wire n5740_1;
wire n5741;
wire n5742;
wire n5743;
wire n5744;
wire n5745;
wire n5745_1;
wire n5746;
wire n5747;
wire n5748;
wire n5749;
wire n5750;
wire n5750_1;
wire n5751;
wire n5752;
wire n5753;
wire n5754;
wire n5755;
wire n5755_1;
wire n5756;
wire n5757;
wire n5758;
wire n5759;
wire n5760;
wire n5760_1;
wire n5761;
wire n5762;
wire n5763;
wire n5764;
wire n5765;
wire n5765_1;
wire n5766;
wire n5767;
wire n5768;
wire n5769;
wire n5769_1;
wire n5770;
wire n5771;
wire n5772;
wire n5773;
wire n5774;
wire n5774_1;
wire n5775;
wire n5776;
wire n5777;
wire n5778;
wire n5779;
wire n5779_1;
wire n5780;
wire n5781;
wire n5782;
wire n5783;
wire n5784;
wire n5784_1;
wire n5785;
wire n5786;
wire n5787;
wire n5788;
wire n5789;
wire n5789_1;
wire n579;
wire n5790;
wire n5791;
wire n5792;
wire n5793;
wire n5794;
wire n5794_1;
wire n5795;
wire n5796;
wire n5797;
wire n5798;
wire n5799;
wire n5799_1;
wire n5800;
wire n5801;
wire n5802;
wire n5803;
wire n5804;
wire n5804_1;
wire n5805;
wire n5806;
wire n5807;
wire n5808;
wire n5809;
wire n5809_1;
wire n5810;
wire n5811;
wire n5812;
wire n5813;
wire n5814;
wire n5814_1;
wire n5815;
wire n5816;
wire n5817;
wire n5818;
wire n5819;
wire n5819_1;
wire n5820;
wire n5821;
wire n5822;
wire n5823;
wire n5824;
wire n5824_1;
wire n5825;
wire n5826;
wire n5827;
wire n5828;
wire n5829;
wire n5829_1;
wire n5830;
wire n5831;
wire n5832;
wire n5833;
wire n5834;
wire n5834_1;
wire n5835;
wire n5836;
wire n5837;
wire n5838;
wire n5839;
wire n5839_1;
wire n584;
wire n5840;
wire n5841;
wire n5842;
wire n5843;
wire n5844;
wire n5844_1;
wire n5845;
wire n5846;
wire n5847;
wire n5848;
wire n5849;
wire n5849_1;
wire n5850;
wire n5851;
wire n5852;
wire n5853;
wire n5854;
wire n5854_1;
wire n5855;
wire n5856;
wire n5857;
wire n5858;
wire n5859;
wire n5859_1;
wire n5860;
wire n5861;
wire n5862;
wire n5863;
wire n5864;
wire n5864_1;
wire n5865;
wire n5866;
wire n5867;
wire n5868;
wire n5869;
wire n5869_1;
wire n5870;
wire n5871;
wire n5872;
wire n5873;
wire n5874;
wire n5875;
wire n5876;
wire n5877;
wire n5878;
wire n5878_1;
wire n5879;
wire n5880;
wire n5881;
wire n5882;
wire n5883;
wire n5883_1;
wire n5884;
wire n5885;
wire n5886;
wire n5887;
wire n5888;
wire n5888_1;
wire n5889;
wire n589;
wire n5890;
wire n5891;
wire n5892;
wire n5893;
wire n5893_1;
wire n5894;
wire n5895;
wire n5896;
wire n5897;
wire n5898;
wire n5898_1;
wire n5899;
wire n5900;
wire n5901;
wire n5902;
wire n5903;
wire n5903_1;
wire n5904;
wire n5905;
wire n5906;
wire n5907;
wire n5908;
wire n5908_1;
wire n5909;
wire n5910;
wire n5911;
wire n5912;
wire n5913;
wire n5913_1;
wire n5914;
wire n5915;
wire n5916;
wire n5917;
wire n5918;
wire n5918_1;
wire n5919;
wire n5920;
wire n5921;
wire n5922;
wire n5923;
wire n5923_1;
wire n5924;
wire n5925;
wire n5926;
wire n5927;
wire n5928;
wire n5928_1;
wire n5929;
wire n5930;
wire n5931;
wire n5932;
wire n5933;
wire n5933_1;
wire n5934;
wire n5935;
wire n5936;
wire n5937;
wire n5938;
wire n5938_1;
wire n5939;
wire n594;
wire n5940;
wire n5941;
wire n5942;
wire n5943;
wire n5943_1;
wire n5944;
wire n5945;
wire n5946;
wire n5947;
wire n5948;
wire n5948_1;
wire n5949;
wire n5950;
wire n5951;
wire n5952;
wire n5953;
wire n5953_1;
wire n5954;
wire n5955;
wire n5956;
wire n5957;
wire n5958;
wire n5958_1;
wire n5959;
wire n5960;
wire n5961;
wire n5962;
wire n5963;
wire n5963_1;
wire n5964;
wire n5965;
wire n5966;
wire n5967;
wire n5968;
wire n5968_1;
wire n5969;
wire n5970;
wire n5971;
wire n5972;
wire n5973;
wire n5973_1;
wire n5974;
wire n5975;
wire n5976;
wire n5977;
wire n5978;
wire n5978_1;
wire n5979;
wire n5980;
wire n5981;
wire n5982;
wire n5983;
wire n5983_1;
wire n5984;
wire n5985;
wire n5986;
wire n5987;
wire n5988;
wire n5988_1;
wire n5989;
wire n599;
wire n5990;
wire n5991;
wire n5992;
wire n5993;
wire n5993_1;
wire n5994;
wire n5995;
wire n5996;
wire n5997;
wire n5998;
wire n5998_1;
wire n5999;
wire n6000;
wire n6001;
wire n6002;
wire n6003;
wire n6003_1;
wire n6004;
wire n6005;
wire n6006;
wire n6007;
wire n6007_1;
wire n6008;
wire n6009;
wire n6010;
wire n6011;
wire n6012;
wire n6012_1;
wire n6013;
wire n6014;
wire n6015;
wire n6016;
wire n6017;
wire n6017_1;
wire n6018;
wire n6019;
wire n6020;
wire n6021;
wire n6022;
wire n6022_1;
wire n6023;
wire n6024;
wire n6025;
wire n6026;
wire n6027;
wire n6027_1;
wire n6028;
wire n6029;
wire n6030;
wire n6031;
wire n6032;
wire n6032_1;
wire n6033;
wire n6034;
wire n6035;
wire n6036;
wire n6037;
wire n6037_1;
wire n6038;
wire n6039;
wire n604;
wire n6040;
wire n6041;
wire n6042;
wire n6042_1;
wire n6043;
wire n6044;
wire n6045;
wire n6046;
wire n6047;
wire n6047_1;
wire n6048;
wire n6049;
wire n6050;
wire n6051;
wire n6051_1;
wire n6052;
wire n6053;
wire n6054;
wire n6055;
wire n6056;
wire n6056_1;
wire n6057;
wire n6058;
wire n6059;
wire n6060;
wire n6061;
wire n6061_1;
wire n6062;
wire n6063;
wire n6064;
wire n6065;
wire n6066;
wire n6066_1;
wire n6067;
wire n6068;
wire n6069;
wire n6070;
wire n6071;
wire n6071_1;
wire n6072;
wire n6073;
wire n6075;
wire n6076;
wire n6076_1;
wire n6077;
wire n6078;
wire n6079;
wire n6080;
wire n6081;
wire n6081_1;
wire n6082;
wire n6083;
wire n6084;
wire n6085;
wire n6086;
wire n6086_1;
wire n6087;
wire n6088;
wire n6089;
wire n609;
wire n6090;
wire n6091;
wire n6091_1;
wire n6092;
wire n6093;
wire n6094;
wire n6095;
wire n6096;
wire n6096_1;
wire n6097;
wire n6098;
wire n6099;
wire n6100;
wire n6101;
wire n6101_1;
wire n6102;
wire n6103;
wire n6104;
wire n6105;
wire n6106;
wire n6106_1;
wire n6107;
wire n6108;
wire n6109;
wire n6110;
wire n6111;
wire n6111_1;
wire n6112;
wire n6113;
wire n6114;
wire n6115;
wire n6116;
wire n6116_1;
wire n6117;
wire n6118;
wire n6119;
wire n6120;
wire n6121;
wire n6121_1;
wire n6122;
wire n6123;
wire n6124;
wire n6125;
wire n6125_1;
wire n6126;
wire n6127;
wire n6128;
wire n6129;
wire n6130;
wire n6130_1;
wire n6131;
wire n6132;
wire n6133;
wire n6134;
wire n6135;
wire n6135_1;
wire n6136;
wire n6137;
wire n6138;
wire n6139;
wire n614;
wire n6140;
wire n6140_1;
wire n6141;
wire n6142;
wire n6143;
wire n6144;
wire n6145;
wire n6145_1;
wire n6146;
wire n6147;
wire n6148;
wire n6149;
wire n6149_1;
wire n6150;
wire n6151;
wire n6152;
wire n6153;
wire n6154;
wire n6154_1;
wire n6155;
wire n6156;
wire n6157;
wire n6158;
wire n6159;
wire n6159_1;
wire n6160;
wire n6161;
wire n6162;
wire n6163;
wire n6163_1;
wire n6164;
wire n6165;
wire n6166;
wire n6167;
wire n6168;
wire n6168_1;
wire n6169;
wire n6170;
wire n6171;
wire n6172;
wire n6172_1;
wire n6173;
wire n6174;
wire n6175;
wire n6176;
wire n6177;
wire n6177_1;
wire n6178;
wire n6179;
wire n6180;
wire n6181;
wire n6182;
wire n6182_1;
wire n6183;
wire n6184;
wire n6185;
wire n6186;
wire n6187;
wire n6187_1;
wire n6188;
wire n6189;
wire n619;
wire n6190;
wire n6191;
wire n6192;
wire n6192_1;
wire n6193;
wire n6194;
wire n6195;
wire n6196;
wire n6197;
wire n6197_1;
wire n6198;
wire n6199;
wire n6200;
wire n6201;
wire n6202;
wire n6202_1;
wire n6203;
wire n6205;
wire n6206;
wire n6207;
wire n6207_1;
wire n6208;
wire n6209;
wire n6210;
wire n6211;
wire n6212;
wire n6212_1;
wire n6213;
wire n6214;
wire n6215;
wire n6216;
wire n6217;
wire n6217_1;
wire n6218;
wire n6219;
wire n6220;
wire n6221;
wire n6222;
wire n6222_1;
wire n6223;
wire n6224;
wire n6225;
wire n6226;
wire n6227;
wire n6227_1;
wire n6228;
wire n6229;
wire n6230;
wire n6231;
wire n6231_1;
wire n6232;
wire n6233;
wire n6234;
wire n6235;
wire n6236;
wire n6236_1;
wire n6237;
wire n6238;
wire n6239;
wire n624;
wire n6240;
wire n6241;
wire n6241_1;
wire n6242;
wire n6243;
wire n6244;
wire n6245;
wire n6246;
wire n6246_1;
wire n6247;
wire n6248;
wire n6249;
wire n6250;
wire n6251;
wire n6251_1;
wire n6252;
wire n6253;
wire n6254;
wire n6255;
wire n6256;
wire n6256_1;
wire n6257;
wire n6258;
wire n6259;
wire n6260;
wire n6260_1;
wire n6261;
wire n6262;
wire n6263;
wire n6264;
wire n6265;
wire n6265_1;
wire n6266;
wire n6267;
wire n6268;
wire n6269;
wire n6270;
wire n6271;
wire n6272;
wire n6273;
wire n6274;
wire n6275;
wire n6276;
wire n6277;
wire n6278;
wire n6279;
wire n6280;
wire n6281;
wire n6282;
wire n6283;
wire n6284;
wire n6285;
wire n6286;
wire n6287;
wire n6288;
wire n6289;
wire n629;
wire n6290;
wire n6291;
wire n6292;
wire n6293;
wire n6294;
wire n6295;
wire n6296;
wire n6297;
wire n6298;
wire n6299;
wire n6300;
wire n6301;
wire n6302;
wire n6303;
wire n6304;
wire n6305;
wire n6306;
wire n6307;
wire n6308;
wire n6309;
wire n6310;
wire n6311;
wire n6312;
wire n6313;
wire n6314;
wire n6315;
wire n6316;
wire n6317;
wire n6318;
wire n6319;
wire n6320;
wire n6321;
wire n6322;
wire n6323;
wire n6324;
wire n6325;
wire n6326;
wire n6327;
wire n6328;
wire n6329;
wire n6330;
wire n6331;
wire n6332;
wire n6333;
wire n6334;
wire n6335;
wire n6336;
wire n6337;
wire n6338;
wire n6339;
wire n634;
wire n6340;
wire n6341;
wire n6342;
wire n6343;
wire n6344;
wire n6345;
wire n6346;
wire n6347;
wire n6348;
wire n6349;
wire n6350;
wire n6351;
wire n6352;
wire n6353;
wire n6354;
wire n6355;
wire n6356;
wire n6357;
wire n6358;
wire n6359;
wire n6360;
wire n6361;
wire n6362;
wire n6363;
wire n6364;
wire n6365;
wire n6366;
wire n6367;
wire n6368;
wire n6369;
wire n6370;
wire n6371;
wire n6372;
wire n6373;
wire n6374;
wire n6375;
wire n6376;
wire n6377;
wire n6378;
wire n6379;
wire n6380;
wire n6381;
wire n6382;
wire n6383;
wire n6384;
wire n6385;
wire n6386;
wire n6387;
wire n6388;
wire n6389;
wire n639;
wire n6390;
wire n6391;
wire n6392;
wire n6393;
wire n6394;
wire n6395;
wire n6396;
wire n6397;
wire n6398;
wire n6399;
wire n6400;
wire n6401;
wire n6402;
wire n6403;
wire n6404;
wire n6405;
wire n6406;
wire n6407;
wire n6408;
wire n6409;
wire n6410;
wire n6411;
wire n6412;
wire n6413;
wire n6414;
wire n6415;
wire n6416;
wire n6417;
wire n6418;
wire n6419;
wire n6420;
wire n6421;
wire n6422;
wire n6423;
wire n6424;
wire n6425;
wire n6426;
wire n6427;
wire n6428;
wire n6429;
wire n6430;
wire n6431;
wire n6432;
wire n6433;
wire n6434;
wire n6435;
wire n6436;
wire n6437;
wire n6438;
wire n6439;
wire n644;
wire n6440;
wire n6441;
wire n6442;
wire n6443;
wire n6444;
wire n6445;
wire n6446;
wire n6447;
wire n6448;
wire n6449;
wire n6450;
wire n6451;
wire n6452;
wire n6453;
wire n6454;
wire n6455;
wire n6456;
wire n6457;
wire n6458;
wire n6459;
wire n6460;
wire n6461;
wire n6462;
wire n6463;
wire n6464;
wire n6465;
wire n6466;
wire n6467;
wire n6468;
wire n6469;
wire n6470;
wire n6471;
wire n6472;
wire n6473;
wire n6474;
wire n6475;
wire n6476;
wire n6477;
wire n6478;
wire n6479;
wire n6480;
wire n6481;
wire n6482;
wire n6483;
wire n6484;
wire n6485;
wire n6486;
wire n6487;
wire n6488;
wire n6489;
wire n649;
wire n6490;
wire n6491;
wire n6492;
wire n6493;
wire n6494;
wire n6495;
wire n6496;
wire n6497;
wire n6498;
wire n6499;
wire n6500;
wire n6501;
wire n6502;
wire n6503;
wire n6504;
wire n6505;
wire n6506;
wire n6507;
wire n6508;
wire n6509;
wire n6510;
wire n6511;
wire n6512;
wire n6513;
wire n6514;
wire n6515;
wire n6516;
wire n6517;
wire n6518;
wire n6519;
wire n6520;
wire n6521;
wire n6522;
wire n6523;
wire n6524;
wire n6525;
wire n6526;
wire n6527;
wire n6528;
wire n6529;
wire n653;
wire n6530;
wire n6531;
wire n6532;
wire n6533;
wire n6534;
wire n6535;
wire n6536;
wire n6537;
wire n6538;
wire n6539;
wire n6540;
wire n6541;
wire n6542;
wire n6543;
wire n6544;
wire n6545;
wire n6546;
wire n6547;
wire n6548;
wire n6549;
wire n6550;
wire n6551;
wire n6552;
wire n6553;
wire n6554;
wire n6555;
wire n6556;
wire n6557;
wire n6558;
wire n6559;
wire n6560;
wire n6561;
wire n6562;
wire n6563;
wire n6564;
wire n6565;
wire n6567;
wire n6568;
wire n6569;
wire n6570;
wire n6571;
wire n6572;
wire n6573;
wire n6574;
wire n6575;
wire n6576;
wire n6577;
wire n6578;
wire n6579;
wire n658;
wire n6580;
wire n6581;
wire n6582;
wire n6583;
wire n6584;
wire n6585;
wire n6586;
wire n6587;
wire n6588;
wire n6589;
wire n6590;
wire n6591;
wire n6592;
wire n6593;
wire n6594;
wire n6595;
wire n6596;
wire n6597;
wire n6598;
wire n6599;
wire n6600;
wire n6601;
wire n6602;
wire n6603;
wire n6604;
wire n6605;
wire n6606;
wire n6607;
wire n6608;
wire n6609;
wire n6610;
wire n6611;
wire n6612;
wire n6613;
wire n6614;
wire n6615;
wire n6616;
wire n6617;
wire n6618;
wire n6619;
wire n6620;
wire n6621;
wire n6622;
wire n6623;
wire n6624;
wire n6625;
wire n6626;
wire n6627;
wire n6628;
wire n6629;
wire n663;
wire n6630;
wire n6631;
wire n6632;
wire n6633;
wire n6634;
wire n6635;
wire n6636;
wire n6637;
wire n6638;
wire n6639;
wire n6640;
wire n6641;
wire n6642;
wire n6643;
wire n6644;
wire n6645;
wire n6646;
wire n6647;
wire n6648;
wire n6649;
wire n6650;
wire n6651;
wire n6652;
wire n6653;
wire n6654;
wire n6655;
wire n6656;
wire n6657;
wire n6658;
wire n6659;
wire n6660;
wire n6661;
wire n6662;
wire n6663;
wire n6664;
wire n6665;
wire n6666;
wire n6667;
wire n6668;
wire n6669;
wire n6670;
wire n6671;
wire n6672;
wire n6673;
wire n6674;
wire n6675;
wire n6676;
wire n6677;
wire n6678;
wire n6679;
wire n668;
wire n6680;
wire n6681;
wire n6682;
wire n6683;
wire n6684;
wire n6685;
wire n6686;
wire n6687;
wire n6688;
wire n6689;
wire n6690;
wire n6691;
wire n6692;
wire n6693;
wire n6694;
wire n6695;
wire n6696;
wire n6697;
wire n6698;
wire n6699;
wire n6700;
wire n6701;
wire n6702;
wire n6703;
wire n6704;
wire n6705;
wire n6706;
wire n6707;
wire n6708;
wire n6709;
wire n6710;
wire n6711;
wire n6712;
wire n6713;
wire n6714;
wire n6715;
wire n6716;
wire n6717;
wire n6718;
wire n6719;
wire n6720;
wire n6721;
wire n6722;
wire n6723;
wire n6724;
wire n6725;
wire n6726;
wire n6727;
wire n6728;
wire n6729;
wire n673;
wire n6730;
wire n6731;
wire n6732;
wire n6733;
wire n6734;
wire n6735;
wire n6736;
wire n6737;
wire n6738;
wire n6739;
wire n6740;
wire n6741;
wire n6742;
wire n6743;
wire n6744;
wire n6745;
wire n6746;
wire n6747;
wire n6748;
wire n6749;
wire n6750;
wire n6751;
wire n6752;
wire n6753;
wire n6754;
wire n6755;
wire n6756;
wire n6757;
wire n6758;
wire n6759;
wire n6760;
wire n6761;
wire n6762;
wire n6763;
wire n6764;
wire n6765;
wire n6766;
wire n6767;
wire n6768;
wire n6769;
wire n6770;
wire n6771;
wire n6772;
wire n6773;
wire n6774;
wire n6775;
wire n6776;
wire n6777;
wire n6778;
wire n6779;
wire n678;
wire n6780;
wire n6781;
wire n6782;
wire n6783;
wire n6784;
wire n6785;
wire n6786;
wire n6787;
wire n6788;
wire n6789;
wire n6790;
wire n6791;
wire n6792;
wire n6793;
wire n6794;
wire n6795;
wire n6796;
wire n6797;
wire n6798;
wire n6799;
wire n6800;
wire n6801;
wire n6802;
wire n6803;
wire n6804;
wire n6805;
wire n6806;
wire n6807;
wire n6808;
wire n6809;
wire n6810;
wire n6811;
wire n6812;
wire n6813;
wire n6814;
wire n6815;
wire n6816;
wire n6817;
wire n6818;
wire n6819;
wire n6820;
wire n6821;
wire n6822;
wire n6823;
wire n6824;
wire n6825;
wire n6826;
wire n6827;
wire n6828;
wire n6829;
wire n683;
wire n6830;
wire n6831;
wire n6832;
wire n6833;
wire n6834;
wire n6835;
wire n6836;
wire n6837;
wire n6838;
wire n6839;
wire n6840;
wire n6841;
wire n6842;
wire n6843;
wire n6844;
wire n6845;
wire n6846;
wire n6847;
wire n6848;
wire n6849;
wire n6850;
wire n6851;
wire n6852;
wire n6853;
wire n6854;
wire n6855;
wire n6856;
wire n6857;
wire n6858;
wire n6859;
wire n6860;
wire n6861;
wire n6862;
wire n6863;
wire n6864;
wire n6865;
wire n6866;
wire n6867;
wire n6868;
wire n6869;
wire n6870;
wire n6871;
wire n6872;
wire n6873;
wire n6874;
wire n6875;
wire n6876;
wire n6877;
wire n6878;
wire n6879;
wire n688;
wire n6880;
wire n6881;
wire n6882;
wire n6883;
wire n6884;
wire n6885;
wire n6886;
wire n6887;
wire n6888;
wire n6889;
wire n6890;
wire n6891;
wire n6892;
wire n6893;
wire n6894;
wire n6895;
wire n6896;
wire n6897;
wire n6898;
wire n6899;
wire n6900;
wire n6901;
wire n6902;
wire n6903;
wire n6905;
wire n6906;
wire n6907;
wire n6908;
wire n6909;
wire n6910;
wire n6911;
wire n6912;
wire n6913;
wire n6914;
wire n6915;
wire n6916;
wire n6917;
wire n6918;
wire n6919;
wire n6920;
wire n6921;
wire n6922;
wire n6923;
wire n6924;
wire n6925;
wire n6926;
wire n6927;
wire n6928;
wire n6929;
wire n693;
wire n6930;
wire n6931;
wire n6932;
wire n6933;
wire n6934;
wire n6935;
wire n6936;
wire n6937;
wire n6938;
wire n6939;
wire n6940;
wire n6941;
wire n6942;
wire n6943;
wire n6944;
wire n6945;
wire n6946;
wire n6947;
wire n6948;
wire n6949;
wire n6950;
wire n6951;
wire n6952;
wire n6953;
wire n6954;
wire n6955;
wire n6956;
wire n6957;
wire n6958;
wire n6959;
wire n6960;
wire n6961;
wire n6962;
wire n6963;
wire n6964;
wire n6965;
wire n6966;
wire n6967;
wire n6968;
wire n6969;
wire n6970;
wire n6971;
wire n6972;
wire n6973;
wire n6974;
wire n6975;
wire n6976;
wire n6977;
wire n6978;
wire n6979;
wire n698;
wire n6980;
wire n6981;
wire n6982;
wire n6983;
wire n6984;
wire n6985;
wire n6986;
wire n6987;
wire n6988;
wire n6989;
wire n6990;
wire n6991;
wire n6992;
wire n6993;
wire n6994;
wire n6995;
wire n6996;
wire n6997;
wire n6998;
wire n6999;
wire n7000;
wire n7001;
wire n7002;
wire n7003;
wire n7004;
wire n7005;
wire n7006;
wire n7007;
wire n7008;
wire n7009;
wire n7010;
wire n7011;
wire n7012;
wire n7013;
wire n7014;
wire n7015;
wire n7016;
wire n7017;
wire n7018;
wire n7019;
wire n7020;
wire n7021;
wire n7022;
wire n7023;
wire n7024;
wire n7025;
wire n7026;
wire n7027;
wire n7028;
wire n7029;
wire n703;
wire n7030;
wire n7031;
wire n7033;
wire n7034;
wire n7035;
wire n7036;
wire n7037;
wire n7038;
wire n7039;
wire n7040;
wire n7041;
wire n7042;
wire n7043;
wire n7044;
wire n7045;
wire n7046;
wire n7047;
wire n7048;
wire n7049;
wire n7050;
wire n7051;
wire n7052;
wire n7053;
wire n7054;
wire n7055;
wire n7056;
wire n7057;
wire n7058;
wire n7059;
wire n7060;
wire n7061;
wire n7062;
wire n7063;
wire n7064;
wire n7065;
wire n7066;
wire n7067;
wire n7068;
wire n7069;
wire n7070;
wire n7071;
wire n7072;
wire n7073;
wire n7074;
wire n7075;
wire n7076;
wire n7077;
wire n7078;
wire n7079;
wire n708;
wire n7080;
wire n7081;
wire n7082;
wire n7083;
wire n7084;
wire n7085;
wire n7086;
wire n7087;
wire n7088;
wire n7089;
wire n7090;
wire n7091;
wire n7092;
wire n7093;
wire n7094;
wire n7095;
wire n7096;
wire n7097;
wire n7098;
wire n7099;
wire n7100;
wire n7101;
wire n7102;
wire n7103;
wire n7104;
wire n7105;
wire n7106;
wire n7107;
wire n7108;
wire n7109;
wire n7110;
wire n7111;
wire n7112;
wire n7113;
wire n7114;
wire n7115;
wire n7116;
wire n7117;
wire n7118;
wire n7119;
wire n7120;
wire n7121;
wire n7122;
wire n7123;
wire n7124;
wire n7125;
wire n7126;
wire n7127;
wire n7128;
wire n7129;
wire n713;
wire n7130;
wire n7131;
wire n7132;
wire n7133;
wire n7134;
wire n7135;
wire n7136;
wire n7137;
wire n7138;
wire n7139;
wire n7140;
wire n7141;
wire n7142;
wire n7143;
wire n7144;
wire n7145;
wire n7146;
wire n7147;
wire n7148;
wire n7149;
wire n7150;
wire n7151;
wire n7152;
wire n7153;
wire n7154;
wire n7155;
wire n7156;
wire n7157;
wire n7158;
wire n7159;
wire n7160;
wire n7161;
wire n7162;
wire n7163;
wire n7164;
wire n7165;
wire n7166;
wire n7167;
wire n7168;
wire n7169;
wire n7170;
wire n7171;
wire n7172;
wire n7173;
wire n7174;
wire n7175;
wire n7176;
wire n7177;
wire n7178;
wire n7179;
wire n718;
wire n7180;
wire n7181;
wire n7182;
wire n7183;
wire n7184;
wire n7185;
wire n7186;
wire n7187;
wire n7188;
wire n7189;
wire n7190;
wire n7191;
wire n7192;
wire n7193;
wire n7194;
wire n7195;
wire n7196;
wire n7197;
wire n7198;
wire n7199;
wire n7200;
wire n7201;
wire n7202;
wire n7203;
wire n7204;
wire n7205;
wire n7206;
wire n7207;
wire n7208;
wire n7209;
wire n7210;
wire n7211;
wire n7212;
wire n7213;
wire n7214;
wire n7215;
wire n7216;
wire n7217;
wire n7218;
wire n7219;
wire n7220;
wire n7221;
wire n7222;
wire n7223;
wire n7224;
wire n7225;
wire n7226;
wire n7227;
wire n7228;
wire n7229;
wire n723;
wire n7230;
wire n7231;
wire n7232;
wire n7233;
wire n7234;
wire n7235;
wire n7236;
wire n7237;
wire n7238;
wire n7239;
wire n7240;
wire n7241;
wire n7242;
wire n7243;
wire n7244;
wire n7245;
wire n7246;
wire n7247;
wire n7248;
wire n7249;
wire n7250;
wire n7251;
wire n7252;
wire n7253;
wire n7254;
wire n7255;
wire n7256;
wire n7257;
wire n7258;
wire n7259;
wire n7260;
wire n7261;
wire n7262;
wire n7263;
wire n7264;
wire n7265;
wire n7266;
wire n7267;
wire n7268;
wire n7269;
wire n727;
wire n7270;
wire n7271;
wire n7272;
wire n7273;
wire n7274;
wire n7275;
wire n7276;
wire n7277;
wire n7278;
wire n7279;
wire n7280;
wire n7281;
wire n7282;
wire n7283;
wire n7284;
wire n7285;
wire n7286;
wire n7287;
wire n7288;
wire n7289;
wire n7290;
wire n7291;
wire n7292;
wire n7293;
wire n7294;
wire n7295;
wire n7296;
wire n7297;
wire n7298;
wire n7299;
wire n7300;
wire n7301;
wire n7302;
wire n7303;
wire n7304;
wire n7305;
wire n7306;
wire n7307;
wire n7308;
wire n7309;
wire n7310;
wire n7311;
wire n7312;
wire n7313;
wire n7314;
wire n7315;
wire n7316;
wire n7317;
wire n7318;
wire n7319;
wire n732;
wire n7320;
wire n7321;
wire n7322;
wire n7323;
wire n7324;
wire n7325;
wire n7326;
wire n7327;
wire n7328;
wire n7329;
wire n7330;
wire n7331;
wire n7332;
wire n7333;
wire n7334;
wire n7335;
wire n7336;
wire n7337;
wire n7338;
wire n7339;
wire n7340;
wire n7341;
wire n7342;
wire n7343;
wire n7344;
wire n7345;
wire n7346;
wire n7347;
wire n7348;
wire n7349;
wire n7350;
wire n7351;
wire n7352;
wire n7353;
wire n7354;
wire n7355;
wire n7356;
wire n7357;
wire n7358;
wire n7359;
wire n7360;
wire n7361;
wire n7362;
wire n7363;
wire n7364;
wire n7365;
wire n7366;
wire n7367;
wire n7368;
wire n7369;
wire n737;
wire n7370;
wire n7371;
wire n7372;
wire n7373;
wire n7374;
wire n7375;
wire n7376;
wire n7377;
wire n7378;
wire n7379;
wire n7380;
wire n7381;
wire n7382;
wire n7383;
wire n7384;
wire n7385;
wire n7386;
wire n7387;
wire n7388;
wire n7389;
wire n7390;
wire n7391;
wire n7392;
wire n7393;
wire n7394;
wire n7395;
wire n7396;
wire n7397;
wire n7398;
wire n7399;
wire n7400;
wire n7401;
wire n7402;
wire n7403;
wire n7404;
wire n7405;
wire n7406;
wire n7407;
wire n7408;
wire n7409;
wire n7410;
wire n7411;
wire n7412;
wire n7413;
wire n7414;
wire n7415;
wire n7416;
wire n7417;
wire n7418;
wire n7419;
wire n742;
wire n7420;
wire n7421;
wire n7422;
wire n7423;
wire n7424;
wire n7425;
wire n7426;
wire n7427;
wire n7428;
wire n7429;
wire n7430;
wire n7431;
wire n7432;
wire n7433;
wire n7434;
wire n7435;
wire n7436;
wire n7437;
wire n7438;
wire n7439;
wire n7440;
wire n7441;
wire n7442;
wire n7443;
wire n7444;
wire n7445;
wire n7446;
wire n7447;
wire n7448;
wire n7449;
wire n7450;
wire n7451;
wire n7452;
wire n7453;
wire n7454;
wire n7455;
wire n7456;
wire n7457;
wire n7458;
wire n7459;
wire n7460;
wire n7461;
wire n7462;
wire n7463;
wire n7464;
wire n7465;
wire n7466;
wire n7467;
wire n7468;
wire n7469;
wire n747;
wire n7470;
wire n7471;
wire n7472;
wire n7473;
wire n7474;
wire n7475;
wire n7476;
wire n7477;
wire n7478;
wire n7479;
wire n7480;
wire n7481;
wire n7482;
wire n7483;
wire n7484;
wire n7485;
wire n7486;
wire n7487;
wire n7488;
wire n7489;
wire n7490;
wire n7491;
wire n7492;
wire n7493;
wire n7494;
wire n7495;
wire n7496;
wire n7497;
wire n7498;
wire n7499;
wire n7500;
wire n7501;
wire n7502;
wire n7503;
wire n7504;
wire n7505;
wire n7506;
wire n7507;
wire n7508;
wire n7509;
wire n7510;
wire n7511;
wire n7512;
wire n7513;
wire n7514;
wire n7515;
wire n7516;
wire n7517;
wire n7518;
wire n7519;
wire n752;
wire n7520;
wire n7521;
wire n7522;
wire n7523;
wire n7524;
wire n7525;
wire n7526;
wire n7527;
wire n7528;
wire n7529;
wire n7530;
wire n7531;
wire n7532;
wire n7533;
wire n7534;
wire n7535;
wire n7536;
wire n7537;
wire n7538;
wire n7539;
wire n7540;
wire n7541;
wire n7542;
wire n7543;
wire n7544;
wire n7545;
wire n7546;
wire n7547;
wire n7548;
wire n7550;
wire n7551;
wire n7552;
wire n7553;
wire n7554;
wire n7555;
wire n7556;
wire n7557;
wire n7558;
wire n7559;
wire n756;
wire n7560;
wire n7561;
wire n7562;
wire n7563;
wire n7564;
wire n7565;
wire n7566;
wire n7567;
wire n7568;
wire n7569;
wire n7570;
wire n7571;
wire n7572;
wire n7573;
wire n7574;
wire n7575;
wire n7576;
wire n7577;
wire n7578;
wire n7579;
wire n7580;
wire n7581;
wire n7582;
wire n7583;
wire n7584;
wire n7585;
wire n7586;
wire n7587;
wire n7588;
wire n7589;
wire n7590;
wire n7591;
wire n7592;
wire n7593;
wire n7594;
wire n7595;
wire n7596;
wire n7597;
wire n7598;
wire n7599;
wire n7600;
wire n7601;
wire n7602;
wire n7603;
wire n7604;
wire n7605;
wire n7606;
wire n7607;
wire n7608;
wire n7609;
wire n761;
wire n7610;
wire n7611;
wire n7612;
wire n7613;
wire n7614;
wire n7615;
wire n7616;
wire n7617;
wire n7618;
wire n7619;
wire n7620;
wire n7621;
wire n7622;
wire n7623;
wire n7624;
wire n7625;
wire n7626;
wire n7627;
wire n7628;
wire n7629;
wire n7630;
wire n7631;
wire n7632;
wire n7633;
wire n7634;
wire n7635;
wire n7636;
wire n7637;
wire n7638;
wire n7639;
wire n7640;
wire n7641;
wire n7642;
wire n7643;
wire n7644;
wire n7645;
wire n7646;
wire n7647;
wire n7648;
wire n7649;
wire n765;
wire n7650;
wire n7651;
wire n7652;
wire n7653;
wire n7654;
wire n7655;
wire n7656;
wire n7657;
wire n7658;
wire n7659;
wire n7660;
wire n7661;
wire n7662;
wire n7663;
wire n7664;
wire n7665;
wire n7666;
wire n7667;
wire n7668;
wire n7669;
wire n7670;
wire n7671;
wire n7672;
wire n7673;
wire n7674;
wire n7675;
wire n7676;
wire n7677;
wire n7678;
wire n7679;
wire n7680;
wire n7681;
wire n7682;
wire n7683;
wire n7684;
wire n7685;
wire n7686;
wire n7687;
wire n7688;
wire n7689;
wire n7690;
wire n7691;
wire n7692;
wire n7693;
wire n7694;
wire n7695;
wire n7696;
wire n7697;
wire n7698;
wire n7699;
wire n770;
wire n7700;
wire n7701;
wire n7702;
wire n7703;
wire n7704;
wire n7705;
wire n7706;
wire n7707;
wire n7708;
wire n7709;
wire n7710;
wire n7711;
wire n7712;
wire n7713;
wire n7714;
wire n7715;
wire n7716;
wire n7717;
wire n7718;
wire n7719;
wire n7720;
wire n7721;
wire n7722;
wire n7723;
wire n7724;
wire n7725;
wire n7726;
wire n7727;
wire n7728;
wire n7729;
wire n7730;
wire n7731;
wire n7732;
wire n7733;
wire n7734;
wire n7735;
wire n7736;
wire n7737;
wire n7738;
wire n7739;
wire n7740;
wire n7741;
wire n7742;
wire n7743;
wire n7744;
wire n7745;
wire n7746;
wire n7747;
wire n7748;
wire n7749;
wire n775;
wire n7750;
wire n7751;
wire n7752;
wire n7753;
wire n7754;
wire n7755;
wire n7756;
wire n7757;
wire n7758;
wire n7759;
wire n7760;
wire n7761;
wire n7762;
wire n7763;
wire n7764;
wire n7765;
wire n7766;
wire n7767;
wire n7768;
wire n7769;
wire n7770;
wire n7771;
wire n7772;
wire n7773;
wire n7774;
wire n7775;
wire n7776;
wire n7777;
wire n7778;
wire n7779;
wire n7780;
wire n7781;
wire n7782;
wire n7783;
wire n7784;
wire n7785;
wire n7786;
wire n7787;
wire n7788;
wire n7789;
wire n7790;
wire n7791;
wire n7792;
wire n7793;
wire n7794;
wire n7795;
wire n7796;
wire n7797;
wire n7798;
wire n7799;
wire n780;
wire n7800;
wire n7801;
wire n7802;
wire n7803;
wire n7804;
wire n7805;
wire n7806;
wire n7807;
wire n7808;
wire n7809;
wire n7810;
wire n7811;
wire n7812;
wire n7813;
wire n7814;
wire n7815;
wire n7816;
wire n7817;
wire n7818;
wire n7819;
wire n7820;
wire n7821;
wire n7822;
wire n7823;
wire n7824;
wire n7825;
wire n7826;
wire n7827;
wire n7828;
wire n7829;
wire n7830;
wire n7831;
wire n7832;
wire n7833;
wire n7834;
wire n7835;
wire n7836;
wire n7837;
wire n7838;
wire n7839;
wire n7840;
wire n7841;
wire n7842;
wire n7843;
wire n7844;
wire n7845;
wire n7846;
wire n7847;
wire n7848;
wire n7849;
wire n785;
wire n7850;
wire n7851;
wire n7852;
wire n7853;
wire n7854;
wire n7855;
wire n7856;
wire n7857;
wire n7858;
wire n7859;
wire n7860;
wire n7861;
wire n7862;
wire n7863;
wire n7864;
wire n7865;
wire n7866;
wire n7867;
wire n7868;
wire n7869;
wire n7870;
wire n7871;
wire n7872;
wire n7873;
wire n7874;
wire n7875;
wire n7876;
wire n7877;
wire n7878;
wire n7879;
wire n7880;
wire n7881;
wire n7882;
wire n7883;
wire n7884;
wire n7885;
wire n7886;
wire n7887;
wire n7888;
wire n7889;
wire n7890;
wire n7891;
wire n7892;
wire n7893;
wire n7894;
wire n7895;
wire n7896;
wire n7897;
wire n7898;
wire n7899;
wire n790;
wire n7900;
wire n7901;
wire n7902;
wire n7903;
wire n7904;
wire n7905;
wire n7906;
wire n7907;
wire n7908;
wire n7909;
wire n7910;
wire n7911;
wire n7912;
wire n7913;
wire n7914;
wire n7915;
wire n7916;
wire n7917;
wire n7918;
wire n7919;
wire n7920;
wire n7921;
wire n7922;
wire n7923;
wire n7924;
wire n7925;
wire n7926;
wire n7927;
wire n7928;
wire n7929;
wire n7930;
wire n7931;
wire n7932;
wire n7933;
wire n7934;
wire n7935;
wire n7936;
wire n7937;
wire n7938;
wire n7939;
wire n794;
wire n7940;
wire n7941;
wire n7942;
wire n7943;
wire n7944;
wire n7945;
wire n7946;
wire n7947;
wire n7948;
wire n7949;
wire n7950;
wire n7951;
wire n7952;
wire n7953;
wire n7954;
wire n7955;
wire n7956;
wire n7957;
wire n7958;
wire n7959;
wire n7960;
wire n7961;
wire n7962;
wire n7963;
wire n7964;
wire n7965;
wire n7966;
wire n7967;
wire n7968;
wire n7969;
wire n7970;
wire n7971;
wire n7972;
wire n7973;
wire n7974;
wire n7975;
wire n7976;
wire n7977;
wire n7978;
wire n7979;
wire n7980;
wire n7981;
wire n7982;
wire n7983;
wire n7984;
wire n7985;
wire n7986;
wire n7987;
wire n7988;
wire n7989;
wire n799;
wire n7990;
wire n7991;
wire n7992;
wire n7993;
wire n7994;
wire n7995;
wire n7996;
wire n7997;
wire n7998;
wire n7999;
wire n8000;
wire n8001;
wire n8002;
wire n8003;
wire n8004;
wire n8005;
wire n8006;
wire n8007;
wire n8008;
wire n8009;
wire n8010;
wire n8011;
wire n8012;
wire n8013;
wire n8014;
wire n8015;
wire n8016;
wire n8017;
wire n8018;
wire n8019;
wire n8020;
wire n8021;
wire n8022;
wire n8023;
wire n8024;
wire n8025;
wire n8026;
wire n8027;
wire n8028;
wire n8029;
wire n8030;
wire n8031;
wire n8032;
wire n8033;
wire n8034;
wire n8035;
wire n8036;
wire n8037;
wire n8038;
wire n8039;
wire n804;
wire n8040;
wire n8041;
wire n8042;
wire n8043;
wire n8044;
wire n8045;
wire n8046;
wire n8047;
wire n8048;
wire n8049;
wire n8050;
wire n8051;
wire n8052;
wire n8053;
wire n8054;
wire n8055;
wire n8056;
wire n8057;
wire n8058;
wire n8059;
wire n8060;
wire n8061;
wire n8062;
wire n8063;
wire n8064;
wire n8065;
wire n8066;
wire n8068;
wire n8069;
wire n8070;
wire n8071;
wire n8072;
wire n8073;
wire n8074;
wire n8075;
wire n8076;
wire n8077;
wire n8078;
wire n8079;
wire n8080;
wire n8081;
wire n8082;
wire n8083;
wire n8084;
wire n8085;
wire n8086;
wire n8087;
wire n8088;
wire n8089;
wire n809;
wire n8090;
wire n8091;
wire n8092;
wire n8093;
wire n8094;
wire n8095;
wire n8096;
wire n8097;
wire n8098;
wire n8099;
wire n8100;
wire n8101;
wire n8102;
wire n8103;
wire n8104;
wire n8105;
wire n8106;
wire n8107;
wire n8108;
wire n8109;
wire n8110;
wire n8111;
wire n8112;
wire n8113;
wire n8114;
wire n8115;
wire n8116;
wire n8117;
wire n8118;
wire n8119;
wire n8120;
wire n8121;
wire n8122;
wire n8123;
wire n8124;
wire n8125;
wire n8126;
wire n8127;
wire n8128;
wire n8129;
wire n8130;
wire n8131;
wire n8132;
wire n8133;
wire n8134;
wire n8135;
wire n8136;
wire n8137;
wire n8138;
wire n8139;
wire n814;
wire n8140;
wire n8141;
wire n8142;
wire n8143;
wire n8144;
wire n8145;
wire n8146;
wire n8147;
wire n8148;
wire n8149;
wire n8150;
wire n8151;
wire n8152;
wire n8153;
wire n8154;
wire n8155;
wire n8156;
wire n8157;
wire n8158;
wire n8159;
wire n8160;
wire n8161;
wire n8162;
wire n8163;
wire n8164;
wire n8165;
wire n8166;
wire n8167;
wire n8168;
wire n8169;
wire n8170;
wire n8171;
wire n8172;
wire n8173;
wire n8174;
wire n8175;
wire n8176;
wire n8177;
wire n8178;
wire n8179;
wire n818;
wire n8180;
wire n8181;
wire n8182;
wire n8183;
wire n8184;
wire n8185;
wire n8186;
wire n8187;
wire n8188;
wire n8189;
wire n8190;
wire n8191;
wire n8192;
wire n8193;
wire n8194;
wire n8195;
wire n8196;
wire n8197;
wire n8198;
wire n8199;
wire n8200;
wire n8201;
wire n8202;
wire n8203;
wire n8204;
wire n8205;
wire n8206;
wire n8207;
wire n8208;
wire n8209;
wire n8210;
wire n8211;
wire n8212;
wire n8213;
wire n8214;
wire n8215;
wire n8216;
wire n8217;
wire n8218;
wire n8219;
wire n8220;
wire n8221;
wire n8222;
wire n8223;
wire n8224;
wire n8225;
wire n8226;
wire n8227;
wire n8228;
wire n8229;
wire n823;
wire n8230;
wire n8231;
wire n8232;
wire n8233;
wire n8234;
wire n8235;
wire n8236;
wire n8237;
wire n8238;
wire n8239;
wire n8240;
wire n8241;
wire n8242;
wire n8243;
wire n8244;
wire n8245;
wire n8246;
wire n8247;
wire n8248;
wire n8249;
wire n8250;
wire n8251;
wire n8252;
wire n8253;
wire n8254;
wire n8255;
wire n8256;
wire n8257;
wire n8258;
wire n8259;
wire n8260;
wire n8261;
wire n8262;
wire n8263;
wire n8264;
wire n8265;
wire n8266;
wire n8267;
wire n8268;
wire n8269;
wire n8270;
wire n8271;
wire n8272;
wire n8273;
wire n8274;
wire n8275;
wire n8276;
wire n8277;
wire n8278;
wire n8279;
wire n828;
wire n8280;
wire n8281;
wire n8282;
wire n8283;
wire n8284;
wire n8285;
wire n8286;
wire n8287;
wire n8288;
wire n8289;
wire n8290;
wire n8291;
wire n8292;
wire n8293;
wire n8294;
wire n8295;
wire n8296;
wire n8297;
wire n8298;
wire n8299;
wire n8300;
wire n8301;
wire n8302;
wire n8303;
wire n8304;
wire n8305;
wire n8306;
wire n8307;
wire n8308;
wire n8309;
wire n8310;
wire n8311;
wire n8312;
wire n8313;
wire n8314;
wire n8315;
wire n8316;
wire n8317;
wire n8318;
wire n8319;
wire n8320;
wire n8321;
wire n8322;
wire n8323;
wire n8324;
wire n8325;
wire n8326;
wire n8327;
wire n8328;
wire n8329;
wire n833;
wire n8330;
wire n8331;
wire n8332;
wire n8333;
wire n8334;
wire n8335;
wire n8336;
wire n8337;
wire n8338;
wire n8339;
wire n8340;
wire n8341;
wire n8342;
wire n8343;
wire n8344;
wire n8345;
wire n8346;
wire n8347;
wire n8348;
wire n8349;
wire n8350;
wire n8351;
wire n8352;
wire n8353;
wire n8354;
wire n8355;
wire n8356;
wire n8357;
wire n8358;
wire n8359;
wire n8360;
wire n8361;
wire n8362;
wire n8363;
wire n8364;
wire n8365;
wire n8366;
wire n8367;
wire n8368;
wire n8369;
wire n8370;
wire n8371;
wire n8372;
wire n8373;
wire n8374;
wire n8375;
wire n8376;
wire n8377;
wire n8378;
wire n8379;
wire n838;
wire n8380;
wire n8381;
wire n8382;
wire n8383;
wire n8384;
wire n8385;
wire n8386;
wire n8387;
wire n8388;
wire n8389;
wire n8390;
wire n8391;
wire n8392;
wire n8393;
wire n8394;
wire n8395;
wire n8396;
wire n8397;
wire n8398;
wire n8399;
wire n8400;
wire n8401;
wire n8402;
wire n8403;
wire n8404;
wire n8405;
wire n8406;
wire n8407;
wire n8408;
wire n8409;
wire n8410;
wire n8411;
wire n8412;
wire n8414;
wire n8415;
wire n8416;
wire n8417;
wire n8418;
wire n8419;
wire n8420;
wire n8421;
wire n8422;
wire n8423;
wire n8424;
wire n8425;
wire n8426;
wire n8427;
wire n8428;
wire n8429;
wire n843;
wire n8430;
wire n8431;
wire n8432;
wire n8433;
wire n8434;
wire n8435;
wire n8436;
wire n8437;
wire n8438;
wire n8439;
wire n8440;
wire n8441;
wire n8442;
wire n8443;
wire n8444;
wire n8445;
wire n8446;
wire n8447;
wire n8448;
wire n8449;
wire n8450;
wire n8451;
wire n8452;
wire n8453;
wire n8454;
wire n8455;
wire n8456;
wire n8457;
wire n8458;
wire n8459;
wire n8460;
wire n8461;
wire n8462;
wire n8463;
wire n8464;
wire n8465;
wire n8466;
wire n8467;
wire n8468;
wire n8469;
wire n847;
wire n8470;
wire n8471;
wire n8472;
wire n8473;
wire n8474;
wire n8475;
wire n8476;
wire n8477;
wire n8478;
wire n8479;
wire n8480;
wire n8481;
wire n8482;
wire n8483;
wire n8484;
wire n8485;
wire n8486;
wire n8487;
wire n8488;
wire n8489;
wire n8490;
wire n8491;
wire n8492;
wire n8493;
wire n8494;
wire n8495;
wire n8496;
wire n8497;
wire n8498;
wire n8499;
wire n8500;
wire n8501;
wire n8502;
wire n8503;
wire n8504;
wire n8505;
wire n8506;
wire n8507;
wire n8508;
wire n8509;
wire n8510;
wire n8511;
wire n8512;
wire n8513;
wire n8514;
wire n8515;
wire n8516;
wire n8517;
wire n8518;
wire n8519;
wire n852;
wire n8520;
wire n8521;
wire n8522;
wire n8523;
wire n8524;
wire n8525;
wire n8526;
wire n8527;
wire n8528;
wire n8529;
wire n8530;
wire n8531;
wire n8532;
wire n8533;
wire n8534;
wire n8535;
wire n8536;
wire n8537;
wire n8538;
wire n8539;
wire n8540;
wire n8541;
wire n8542;
wire n8543;
wire n8544;
wire n8545;
wire n8546;
wire n8547;
wire n8548;
wire n8549;
wire n8550;
wire n8551;
wire n8552;
wire n8553;
wire n8554;
wire n8555;
wire n8556;
wire n8557;
wire n8558;
wire n8559;
wire n8560;
wire n8561;
wire n8562;
wire n8563;
wire n8564;
wire n8565;
wire n8566;
wire n8567;
wire n8568;
wire n8569;
wire n857;
wire n8570;
wire n8571;
wire n8572;
wire n8573;
wire n8574;
wire n8575;
wire n8576;
wire n8577;
wire n8578;
wire n8579;
wire n8580;
wire n8581;
wire n8582;
wire n8583;
wire n8584;
wire n8585;
wire n8586;
wire n8587;
wire n8588;
wire n8589;
wire n8590;
wire n8591;
wire n8592;
wire n8593;
wire n8594;
wire n8595;
wire n8596;
wire n8597;
wire n8598;
wire n8599;
wire n8600;
wire n8601;
wire n8602;
wire n8603;
wire n8604;
wire n8605;
wire n8606;
wire n8607;
wire n8608;
wire n8609;
wire n8610;
wire n8611;
wire n8612;
wire n8613;
wire n8614;
wire n8615;
wire n8616;
wire n8617;
wire n8618;
wire n8619;
wire n862;
wire n8620;
wire n8621;
wire n8622;
wire n8623;
wire n8624;
wire n8625;
wire n8626;
wire n8627;
wire n8628;
wire n8629;
wire n8630;
wire n8631;
wire n8632;
wire n8633;
wire n8634;
wire n8635;
wire n8636;
wire n8637;
wire n8638;
wire n8639;
wire n8640;
wire n8641;
wire n8642;
wire n8643;
wire n8644;
wire n8645;
wire n8646;
wire n8647;
wire n8648;
wire n8649;
wire n8650;
wire n8651;
wire n8652;
wire n8653;
wire n8654;
wire n8655;
wire n8656;
wire n8657;
wire n8658;
wire n8659;
wire n8660;
wire n8661;
wire n8662;
wire n8663;
wire n8664;
wire n8665;
wire n8666;
wire n8667;
wire n8668;
wire n8669;
wire n867;
wire n8670;
wire n8671;
wire n8672;
wire n8673;
wire n8674;
wire n8675;
wire n8676;
wire n8677;
wire n8678;
wire n8679;
wire n8680;
wire n8681;
wire n8682;
wire n8683;
wire n8684;
wire n8685;
wire n8686;
wire n8687;
wire n8688;
wire n8689;
wire n8690;
wire n8691;
wire n8692;
wire n8693;
wire n8694;
wire n8695;
wire n8696;
wire n8697;
wire n8698;
wire n8699;
wire n8700;
wire n8701;
wire n8702;
wire n8703;
wire n8704;
wire n8705;
wire n8706;
wire n8707;
wire n8708;
wire n8709;
wire n8710;
wire n8711;
wire n8712;
wire n8713;
wire n8714;
wire n8715;
wire n8716;
wire n8717;
wire n8718;
wire n8719;
wire n872;
wire n8720;
wire n8721;
wire n8722;
wire n8723;
wire n8724;
wire n8725;
wire n8726;
wire n8727;
wire n8728;
wire n8729;
wire n8730;
wire n8731;
wire n8732;
wire n8733;
wire n8734;
wire n8735;
wire n8736;
wire n8737;
wire n8738;
wire n8739;
wire n8740;
wire n8741;
wire n8742;
wire n8743;
wire n8744;
wire n8745;
wire n8746;
wire n8747;
wire n8748;
wire n8749;
wire n8750;
wire n8751;
wire n8752;
wire n8753;
wire n8754;
wire n8755;
wire n8756;
wire n8757;
wire n8758;
wire n8759;
wire n876;
wire n8760;
wire n8761;
wire n8764;
wire n8765;
wire n8766;
wire n8767;
wire n8768;
wire n8769;
wire n8770;
wire n8771;
wire n8772;
wire n8773;
wire n8774;
wire n8775;
wire n8776;
wire n8777;
wire n8778;
wire n8779;
wire n8780;
wire n8781;
wire n8782;
wire n8783;
wire n8784;
wire n8785;
wire n8786;
wire n8787;
wire n8788;
wire n8789;
wire n8790;
wire n8791;
wire n8792;
wire n8793;
wire n8794;
wire n8795;
wire n8796;
wire n8797;
wire n8798;
wire n8799;
wire n8800;
wire n8801;
wire n8802;
wire n8803;
wire n8804;
wire n8805;
wire n8806;
wire n8807;
wire n8808;
wire n8809;
wire n881;
wire n8810;
wire n8811;
wire n8812;
wire n8813;
wire n8814;
wire n8815;
wire n8816;
wire n8817;
wire n8818;
wire n8819;
wire n8820;
wire n8821;
wire n8822;
wire n8823;
wire n8824;
wire n8825;
wire n8826;
wire n8827;
wire n8828;
wire n8829;
wire n8830;
wire n8831;
wire n8832;
wire n8833;
wire n8834;
wire n8835;
wire n8836;
wire n8837;
wire n8838;
wire n8839;
wire n8840;
wire n8841;
wire n8842;
wire n8843;
wire n8844;
wire n8845;
wire n8846;
wire n8847;
wire n8848;
wire n8849;
wire n8850;
wire n8851;
wire n8852;
wire n8853;
wire n8854;
wire n8855;
wire n8856;
wire n8857;
wire n8858;
wire n8859;
wire n886;
wire n8860;
wire n8861;
wire n8862;
wire n8863;
wire n8864;
wire n8865;
wire n8866;
wire n8867;
wire n8868;
wire n8869;
wire n8870;
wire n8871;
wire n8872;
wire n8873;
wire n8874;
wire n8875;
wire n8876;
wire n8877;
wire n8878;
wire n8879;
wire n8880;
wire n8881;
wire n8882;
wire n8883;
wire n8884;
wire n8885;
wire n8886;
wire n8887;
wire n8888;
wire n8889;
wire n8890;
wire n8891;
wire n8892;
wire n8893;
wire n8894;
wire n8895;
wire n8896;
wire n8897;
wire n8898;
wire n8899;
wire n8900;
wire n8901;
wire n8902;
wire n8903;
wire n8904;
wire n8905;
wire n8906;
wire n8907;
wire n8908;
wire n8909;
wire n891;
wire n8910;
wire n8911;
wire n8912;
wire n8913;
wire n8914;
wire n8915;
wire n8916;
wire n8917;
wire n8918;
wire n8919;
wire n8920;
wire n8921;
wire n8922;
wire n8923;
wire n8924;
wire n8925;
wire n8926;
wire n8927;
wire n8928;
wire n8929;
wire n8930;
wire n8931;
wire n8932;
wire n8933;
wire n8934;
wire n8935;
wire n8936;
wire n8937;
wire n8938;
wire n8939;
wire n8940;
wire n8941;
wire n8942;
wire n8943;
wire n8944;
wire n8945;
wire n8946;
wire n8947;
wire n8948;
wire n8949;
wire n8950;
wire n8951;
wire n8952;
wire n8953;
wire n8954;
wire n8955;
wire n8956;
wire n8957;
wire n8958;
wire n8959;
wire n896;
wire n8960;
wire n8961;
wire n8962;
wire n8963;
wire n8964;
wire n8965;
wire n8966;
wire n8967;
wire n8968;
wire n8969;
wire n8970;
wire n8971;
wire n8972;
wire n8974;
wire n8975;
wire n8976;
wire n8977;
wire n8978;
wire n8979;
wire n8980;
wire n8981;
wire n8982;
wire n8983;
wire n8984;
wire n8985;
wire n8986;
wire n8987;
wire n8988;
wire n8989;
wire n8990;
wire n8991;
wire n8992;
wire n8993;
wire n8994;
wire n8995;
wire n8996;
wire n8997;
wire n8998;
wire n8999;
wire n9000;
wire n9001;
wire n9002;
wire n9003;
wire n9004;
wire n9005;
wire n9006;
wire n9007;
wire n9008;
wire n9009;
wire n901;
wire n9010;
wire n9011;
wire n9012;
wire n9013;
wire n9014;
wire n9015;
wire n9016;
wire n9017;
wire n9018;
wire n9019;
wire n9020;
wire n9021;
wire n9022;
wire n9023;
wire n9024;
wire n9025;
wire n9026;
wire n9027;
wire n9028;
wire n9029;
wire n9030;
wire n9031;
wire n9032;
wire n9033;
wire n9034;
wire n9035;
wire n9036;
wire n9037;
wire n9038;
wire n9039;
wire n9040;
wire n9041;
wire n9042;
wire n9043;
wire n9044;
wire n9045;
wire n9046;
wire n9047;
wire n9048;
wire n9049;
wire n9050;
wire n9051;
wire n9052;
wire n9053;
wire n9054;
wire n9055;
wire n9056;
wire n9057;
wire n9058;
wire n9059;
wire n906;
wire n9060;
wire n9061;
wire n9062;
wire n9063;
wire n9064;
wire n9065;
wire n9066;
wire n9067;
wire n9068;
wire n9069;
wire n9070;
wire n9071;
wire n9072;
wire n9073;
wire n9074;
wire n9075;
wire n9076;
wire n9077;
wire n9078;
wire n9079;
wire n9080;
wire n9081;
wire n9082;
wire n9083;
wire n9084;
wire n9085;
wire n9086;
wire n9087;
wire n9088;
wire n9089;
wire n9090;
wire n9091;
wire n9092;
wire n9093;
wire n9094;
wire n9095;
wire n9096;
wire n9097;
wire n9098;
wire n9099;
wire n9100;
wire n9101;
wire n9102;
wire n9103;
wire n9104;
wire n9105;
wire n9106;
wire n9107;
wire n9108;
wire n9109;
wire n911;
wire n9110;
wire n9111;
wire n9112;
wire n9113;
wire n9114;
wire n9115;
wire n9116;
wire n9117;
wire n9118;
wire n9119;
wire n9120;
wire n9121;
wire n9122;
wire n9123;
wire n9124;
wire n9125;
wire n9126;
wire n9127;
wire n9128;
wire n9129;
wire n9130;
wire n9131;
wire n9132;
wire n9133;
wire n9134;
wire n9135;
wire n9136;
wire n9137;
wire n9138;
wire n9139;
wire n9140;
wire n9141;
wire n9142;
wire n9143;
wire n9144;
wire n9145;
wire n9146;
wire n9147;
wire n9148;
wire n9149;
wire n9150;
wire n9151;
wire n9152;
wire n9153;
wire n9154;
wire n9155;
wire n9156;
wire n9157;
wire n9158;
wire n9159;
wire n916;
wire n9160;
wire n9161;
wire n9162;
wire n9163;
wire n9164;
wire n9165;
wire n9166;
wire n9167;
wire n9168;
wire n9169;
wire n9170;
wire n9171;
wire n9172;
wire n9173;
wire n9174;
wire n9175;
wire n9176;
wire n9177;
wire n9178;
wire n9179;
wire n9180;
wire n9181;
wire n9182;
wire n9183;
wire n9184;
wire n9185;
wire n9186;
wire n9187;
wire n9188;
wire n9189;
wire n9190;
wire n9191;
wire n9192;
wire n9193;
wire n9194;
wire n9195;
wire n9196;
wire n9197;
wire n9198;
wire n9199;
wire n9200;
wire n9201;
wire n9202;
wire n9203;
wire n9204;
wire n9205;
wire n9206;
wire n9207;
wire n9208;
wire n9209;
wire n921;
wire n9210;
wire n9211;
wire n9212;
wire n9213;
wire n9214;
wire n9215;
wire n9216;
wire n9217;
wire n9218;
wire n9219;
wire n9220;
wire n9221;
wire n9222;
wire n9223;
wire n9224;
wire n9225;
wire n9226;
wire n9227;
wire n9228;
wire n9229;
wire n9230;
wire n9231;
wire n9232;
wire n9233;
wire n9234;
wire n9236;
wire n9238;
wire n9239;
wire n9240;
wire n9241;
wire n9242;
wire n9243;
wire n9245;
wire n9246;
wire n9247;
wire n9248;
wire n9249;
wire n9250;
wire n9251;
wire n9252;
wire n9253;
wire n9254;
wire n9255;
wire n9256;
wire n9257;
wire n9258;
wire n9259;
wire n926;
wire n9260;
wire n9261;
wire n9262;
wire n9263;
wire n9264;
wire n9265;
wire n9266;
wire n9267;
wire n9268;
wire n9269;
wire n9270;
wire n9271;
wire n9272;
wire n9273;
wire n9274;
wire n9275;
wire n9276;
wire n9277;
wire n9278;
wire n9279;
wire n9280;
wire n9281;
wire n9282;
wire n9283;
wire n9284;
wire n9285;
wire n9286;
wire n9287;
wire n9288;
wire n9289;
wire n9290;
wire n9291;
wire n9292;
wire n9293;
wire n9294;
wire n9295;
wire n9296;
wire n9297;
wire n9298;
wire n9299;
wire n9300;
wire n9301;
wire n9302;
wire n9303;
wire n9304;
wire n9305;
wire n9306;
wire n9307;
wire n9308;
wire n9309;
wire n931;
wire n9310;
wire n9311;
wire n9312;
wire n9313;
wire n9314;
wire n9315;
wire n9316;
wire n9317;
wire n9318;
wire n9319;
wire n9320;
wire n9321;
wire n9322;
wire n9323;
wire n9324;
wire n9325;
wire n9326;
wire n9327;
wire n9328;
wire n9329;
wire n9330;
wire n9331;
wire n9332;
wire n9333;
wire n9334;
wire n9335;
wire n9336;
wire n9337;
wire n9338;
wire n9339;
wire n9340;
wire n9341;
wire n9342;
wire n9343;
wire n9344;
wire n9345;
wire n9346;
wire n9347;
wire n9348;
wire n9350;
wire n9351;
wire n9352;
wire n9353;
wire n9354;
wire n9355;
wire n9356;
wire n9357;
wire n9358;
wire n9359;
wire n936;
wire n9360;
wire n9361;
wire n9362;
wire n9363;
wire n9364;
wire n9365;
wire n9366;
wire n9367;
wire n9368;
wire n9369;
wire n9370;
wire n9371;
wire n9372;
wire n9373;
wire n9374;
wire n9375;
wire n9376;
wire n9377;
wire n9378;
wire n9379;
wire n9380;
wire n9381;
wire n9382;
wire n9383;
wire n9384;
wire n9385;
wire n9386;
wire n9387;
wire n9388;
wire n9389;
wire n9390;
wire n9391;
wire n9392;
wire n9393;
wire n9394;
wire n9395;
wire n9396;
wire n9397;
wire n9398;
wire n9399;
wire n9400;
wire n9401;
wire n9402;
wire n9403;
wire n9404;
wire n9405;
wire n9406;
wire n9407;
wire n9408;
wire n9409;
wire n941;
wire n9410;
wire n9411;
wire n9412;
wire n9413;
wire n9414;
wire n9415;
wire n9416;
wire n9417;
wire n9418;
wire n9419;
wire n9420;
wire n9421;
wire n9422;
wire n9423;
wire n9424;
wire n9425;
wire n9426;
wire n9427;
wire n9428;
wire n9429;
wire n9430;
wire n9431;
wire n9432;
wire n9433;
wire n9434;
wire n9435;
wire n9436;
wire n9437;
wire n9438;
wire n9439;
wire n9440;
wire n9441;
wire n9442;
wire n9443;
wire n9444;
wire n9445;
wire n9446;
wire n9447;
wire n9448;
wire n9449;
wire n9450;
wire n9451;
wire n9452;
wire n9453;
wire n9454;
wire n9455;
wire n9456;
wire n9457;
wire n9458;
wire n9459;
wire n946;
wire n9460;
wire n9461;
wire n9462;
wire n9463;
wire n9464;
wire n9465;
wire n9466;
wire n9467;
wire n9468;
wire n9469;
wire n9470;
wire n9471;
wire n9472;
wire n9473;
wire n9474;
wire n9475;
wire n9476;
wire n9477;
wire n9478;
wire n9479;
wire n9480;
wire n9481;
wire n9482;
wire n9483;
wire n9484;
wire n9485;
wire n9486;
wire n9487;
wire n9488;
wire n9489;
wire n9490;
wire n9491;
wire n9492;
wire n9493;
wire n9494;
wire n9495;
wire n9496;
wire n9497;
wire n9498;
wire n9499;
wire n9500;
wire n9501;
wire n9502;
wire n9503;
wire n9504;
wire n9505;
wire n9506;
wire n9507;
wire n9508;
wire n9509;
wire n951;
wire n9510;
wire n9511;
wire n9512;
wire n9513;
wire n9514;
wire n9515;
wire n9516;
wire n9517;
wire n9518;
wire n9519;
wire n9520;
wire n9521;
wire n9522;
wire n9523;
wire n9524;
wire n9525;
wire n9526;
wire n9527;
wire n9528;
wire n9529;
wire n9530;
wire n9531;
wire n9532;
wire n9533;
wire n9534;
wire n9535;
wire n9536;
wire n9537;
wire n9538;
wire n9539;
wire n9540;
wire n9541;
wire n9542;
wire n9543;
wire n9544;
wire n9545;
wire n9546;
wire n9547;
wire n9548;
wire n9549;
wire n9550;
wire n9551;
wire n9552;
wire n9553;
wire n9554;
wire n9555;
wire n9556;
wire n9557;
wire n9558;
wire n9559;
wire n956;
wire n9560;
wire n9561;
wire n9562;
wire n9563;
wire n9564;
wire n9565;
wire n9566;
wire n9567;
wire n9568;
wire n9569;
wire n9570;
wire n9571;
wire n9572;
wire n9573;
wire n9574;
wire n9575;
wire n9576;
wire n9577;
wire n9578;
wire n9579;
wire n9580;
wire n9581;
wire n9582;
wire n9583;
wire n9584;
wire n9585;
wire n9586;
wire n9587;
wire n9588;
wire n9589;
wire n9590;
wire n9591;
wire n9592;
wire n9593;
wire n9594;
wire n9595;
wire n9596;
wire n9597;
wire n9598;
wire n9599;
wire n9600;
wire n9601;
wire n9602;
wire n9603;
wire n9604;
wire n9605;
wire n9606;
wire n9607;
wire n9608;
wire n9609;
wire n961;
wire n9610;
wire n9611;
wire n9612;
wire n9613;
wire n9614;
wire n9615;
wire n9616;
wire n9617;
wire n9618;
wire n9619;
wire n9620;
wire n9621;
wire n9622;
wire n9623;
wire n9624;
wire n9625;
wire n9626;
wire n9627;
wire n9628;
wire n9629;
wire n9630;
wire n9631;
wire n9632;
wire n9633;
wire n9634;
wire n9635;
wire n9636;
wire n9637;
wire n9638;
wire n9639;
wire n9640;
wire n9641;
wire n9642;
wire n9643;
wire n9644;
wire n9645;
wire n9646;
wire n9648;
wire n9650;
wire n9651;
wire n9652;
wire n9653;
wire n9654;
wire n9655;
wire n9656;
wire n9657;
wire n9658;
wire n9659;
wire n966;
wire n9660;
wire n9661;
wire n9662;
wire n9663;
wire n9664;
wire n9665;
wire n9666;
wire n9667;
wire n9668;
wire n9669;
wire n9670;
wire n9671;
wire n9672;
wire n9673;
wire n9674;
wire n9675;
wire n9676;
wire n9677;
wire n9678;
wire n9679;
wire n9680;
wire n9681;
wire n9682;
wire n9683;
wire n9684;
wire n9685;
wire n9686;
wire n9687;
wire n9688;
wire n9689;
wire n9690;
wire n9691;
wire n9692;
wire n9693;
wire n9694;
wire n9695;
wire n9696;
wire n9697;
wire n9698;
wire n9699;
wire n9700;
wire n9701;
wire n9702;
wire n9703;
wire n9704;
wire n9705;
wire n9706;
wire n9707;
wire n9708;
wire n9709;
wire n971;
wire n9710;
wire n9711;
wire n9712;
wire n9713;
wire n9714;
wire n9715;
wire n9716;
wire n9717;
wire n9718;
wire n9719;
wire n9720;
wire n9721;
wire n9722;
wire n9723;
wire n9724;
wire n9725;
wire n9726;
wire n9727;
wire n9728;
wire n9729;
wire n9730;
wire n9731;
wire n9732;
wire n9733;
wire n9734;
wire n9735;
wire n9736;
wire n9737;
wire n9738;
wire n9739;
wire n9740;
wire n9741;
wire n9742;
wire n9743;
wire n9744;
wire n9745;
wire n9746;
wire n9747;
wire n9748;
wire n9749;
wire n9750;
wire n9751;
wire n9752;
wire n9753;
wire n9754;
wire n9755;
wire n9756;
wire n9757;
wire n9758;
wire n9759;
wire n976;
wire n9760;
wire n9761;
wire n9762;
wire n9763;
wire n9764;
wire n9765;
wire n9766;
wire n9767;
wire n9768;
wire n9769;
wire n9770;
wire n9771;
wire n9772;
wire n9773;
wire n9774;
wire n9775;
wire n9776;
wire n9777;
wire n9778;
wire n9779;
wire n9780;
wire n9781;
wire n9782;
wire n9783;
wire n9784;
wire n9785;
wire n9786;
wire n9787;
wire n9788;
wire n9789;
wire n9790;
wire n9791;
wire n9792;
wire n9793;
wire n9794;
wire n9795;
wire n9796;
wire n9797;
wire n9798;
wire n9799;
wire n9800;
wire n9801;
wire n9802;
wire n9803;
wire n9804;
wire n9805;
wire n9806;
wire n9807;
wire n9808;
wire n9809;
wire n981;
wire n9810;
wire n9811;
wire n9812;
wire n9813;
wire n9814;
wire n9815;
wire n9816;
wire n9817;
wire n9818;
wire n9819;
wire n9820;
wire n9821;
wire n9822;
wire n9823;
wire n9824;
wire n9825;
wire n9826;
wire n9827;
wire n9828;
wire n9829;
wire n9830;
wire n9831;
wire n9832;
wire n9833;
wire n9834;
wire n9835;
wire n9836;
wire n9837;
wire n9838;
wire n9839;
wire n9840;
wire n9841;
wire n9842;
wire n9843;
wire n9844;
wire n9845;
wire n9846;
wire n9847;
wire n9848;
wire n9849;
wire n9850;
wire n9851;
wire n9852;
wire n9853;
wire n9854;
wire n9855;
wire n9856;
wire n9857;
wire n9858;
wire n9859;
wire n986;
wire n9860;
wire n9861;
wire n9862;
wire n9863;
wire n9864;
wire n9865;
wire n9866;
wire n9867;
wire n9868;
wire n9869;
wire n9870;
wire n9871;
wire n9872;
wire n9873;
wire n9874;
wire n9875;
wire n9876;
wire n9877;
wire n9878;
wire n9879;
wire n9880;
wire n9881;
wire n9882;
wire n9883;
wire n9884;
wire n9885;
wire n9886;
wire n9887;
wire n9888;
wire n9889;
wire n9890;
wire n9891;
wire n9892;
wire n9893;
wire n9894;
wire n9895;
wire n9896;
wire n9897;
wire n9898;
wire n9899;
wire n9900;
wire n9901;
wire n9903;
wire n9904;
wire n9905;
wire n9906;
wire n9907;
wire n9908;
wire n9909;
wire n991;
wire n9910;
wire n9911;
wire n9912;
wire n9913;
wire n9914;
wire n9915;
wire n9916;
wire n9917;
wire n9918;
wire n9919;
wire n9920;
wire n9921;
wire n9922;
wire n9923;
wire n9924;
wire n9925;
wire n9926;
wire n9927;
wire n9928;
wire n9929;
wire n9930;
wire n9931;
wire n9932;
wire n9933;
wire n9934;
wire n9935;
wire n9936;
wire n9937;
wire n9938;
wire n9939;
wire n9940;
wire n9941;
wire n9942;
wire n9943;
wire n9944;
wire n9945;
wire n9946;
wire n9947;
wire n9948;
wire n9949;
wire n9950;
wire n9951;
wire n9952;
wire n9953;
wire n9954;
wire n9955;
wire n9956;
wire n9957;
wire n9958;
wire n9959;
wire n996;
wire n9960;
wire n9961;
wire n9962;
wire n9963;
wire n9964;
wire n9965;
wire n9966;
wire n9967;
wire n9968;
wire n9969;
wire n9970;
wire n9971;
wire n9972;
wire n9973;
wire n9974;
wire n9975;
wire n9976;
wire n9977;
wire n9978;
wire n9979;
wire n9980;
wire n9981;
wire n9982;
wire n9983;
wire n9984;
wire n9985;
wire n9986;
wire n9987;
wire n9988;
wire n9989;
wire n9990;
wire n9991;
wire n9992;
wire n9993;
wire n9994;
wire n9995;
wire n9996;
wire n9997;
wire n9998;
wire n9999;
wire n_17093;
wire n_186;
wire n_22641;
wire n_25834;
wire n_27014;
wire n_27923;
wire n_44061;
wire n_44365;
wire n_44422;
wire n_44610;
wire n_44695;
wire n_44721;
wire n_44722;
wire n_44847;
wire n_44962;
wire n_45202;
wire n_45204;
wire n_45209;
wire n_45224;
wire n_45622;
wire n_46254;
wire state_cordic_1_;

// Start cells
in01f01 g00000 ( .a(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n3789) );
in01f01 g00001 ( .a(n_44962), .o(n3790) );
no02f01 g00002 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_6_), .b(n3790), .o(n3791) );
no02f01 g00003 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_5_), .b(n3790), .o(n3792_1) );
no02f01 g00004 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_2_), .b(n3790), .o(n3793) );
in01f01 g00005 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_1_), .o(n3794) );
na02f01 g00006 ( .a(n3794), .b(n_44962), .o(n3795) );
in01f01 g00007 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_0_), .o(n3796) );
na02f01 g00008 ( .a(n3796), .b(n_44962), .o(n3797_1) );
na02f01 g00009 ( .a(n3797_1), .b(n3795), .o(n3798) );
no02f01 g00010 ( .a(n3798), .b(n3793), .o(n3799) );
no02f01 g00011 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_3_), .b(n3790), .o(n3800) );
no02f01 g00012 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_4_), .b(n3790), .o(n3801) );
no02f01 g00013 ( .a(n3801), .b(n3800), .o(n3802_1) );
na02f01 g00014 ( .a(n3802_1), .b(n3799), .o(n3803) );
no02f01 g00015 ( .a(n3803), .b(n3792_1), .o(n3804) );
in01f01 g00016 ( .a(n3804), .o(n3805) );
no02f01 g00017 ( .a(n3805), .b(n3791), .o(n3806_1) );
no02f01 g00018 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_9_), .b(n3790), .o(n3807) );
no02f01 g00019 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_8_), .b(n3790), .o(n3808) );
no02f01 g00020 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_7_), .b(n3790), .o(n3809) );
no03f01 g00021 ( .a(n3809), .b(n3808), .c(n3807), .o(n3810) );
na02f01 g00022 ( .a(n3810), .b(n3806_1), .o(n3811_1) );
in01f01 g00023 ( .a(n3811_1), .o(n3812) );
in01f01 g00024 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_10_), .o(n3813) );
no02f01 g00025 ( .a(n3813), .b(n_44962), .o(n3814) );
in01f01 g00026 ( .a(n3814), .o(n3815) );
no03f01 g00027 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_8_), .b(delay_xor_ln22_unr21_stage8_stallmux_q_9_), .c(n_44962), .o(n3816_1) );
no02f01 g00028 ( .a(n3816_1), .b(delay_xor_ln22_unr21_stage8_stallmux_q_10_), .o(n3817) );
ao12f01 g00029 ( .a(n3817), .b(n3815), .c(n3812), .o(n3818) );
no02f01 g00030 ( .a(n3818), .b(delay_add_ln22_unr20_stage8_stallmux_q_23_), .o(n3819) );
in01f01 g00031 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_23_), .o(n3820) );
in01f01 g00032 ( .a(n3818), .o(n3821_1) );
no02f01 g00033 ( .a(n3821_1), .b(n3820), .o(n3822) );
no02f01 g00034 ( .a(n3822), .b(n3819), .o(n3823) );
in01f01 g00035 ( .a(n3823), .o(n3824) );
ao12f01 g00036 ( .a(n3818), .b(delay_add_ln22_unr20_stage8_stallmux_q_16_), .c(delay_add_ln22_unr20_stage8_stallmux_q_17_), .o(n3825) );
in01f01 g00037 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_14_), .o(n3826_1) );
in01f01 g00038 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_15_), .o(n3827) );
ao12f01 g00039 ( .a(n3821_1), .b(n3827), .c(n3826_1), .o(n3828) );
no03f01 g00040 ( .a(n3809), .b(n3792_1), .c(n3791), .o(n3829) );
na03f01 g00041 ( .a(n3829), .b(n3802_1), .c(n3799), .o(n3830) );
no02f01 g00042 ( .a(n3830), .b(n3808), .o(n3831_1) );
in01f01 g00043 ( .a(n3831_1), .o(n3832) );
na02f01 g00044 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_9_), .b(n3790), .o(n3833) );
in01f01 g00045 ( .a(n3833), .o(n3834) );
no02f01 g00046 ( .a(n3834), .b(n3807), .o(n3835) );
no02f01 g00047 ( .a(n3835), .b(n3832), .o(n3836_1) );
na02f01 g00048 ( .a(n3835), .b(n3832), .o(n3837) );
in01f01 g00049 ( .a(n3837), .o(n3838) );
no02f01 g00050 ( .a(n3838), .b(n3836_1), .o(n3839) );
in01f01 g00051 ( .a(n3839), .o(n3840) );
no02f01 g00052 ( .a(n3840), .b(delay_add_ln22_unr20_stage8_stallmux_q_9_), .o(n3841_1) );
in01f01 g00053 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_8_), .o(n3842) );
in01f01 g00054 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_8_), .o(n3843) );
no02f01 g00055 ( .a(n3843), .b(n_44962), .o(n3844) );
no02f01 g00056 ( .a(n3844), .b(n3808), .o(n3845) );
no02f01 g00057 ( .a(n3845), .b(n3830), .o(n3846_1) );
na02f01 g00058 ( .a(n3845), .b(n3830), .o(n3847) );
in01f01 g00059 ( .a(n3847), .o(n3848) );
no02f01 g00060 ( .a(n3848), .b(n3846_1), .o(n3849) );
no02f01 g00061 ( .a(n3849), .b(n3842), .o(n3850_1) );
in01f01 g00062 ( .a(n3806_1), .o(n3851) );
na02f01 g00063 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_7_), .b(n3790), .o(n3852) );
in01f01 g00064 ( .a(n3852), .o(n3853) );
no02f01 g00065 ( .a(n3853), .b(n3809), .o(n3854) );
no02f01 g00066 ( .a(n3854), .b(n3851), .o(n3855_1) );
na02f01 g00067 ( .a(n3854), .b(n3851), .o(n3856) );
in01f01 g00068 ( .a(n3856), .o(n3857) );
no02f01 g00069 ( .a(n3857), .b(n3855_1), .o(n3858) );
in01f01 g00070 ( .a(n3858), .o(n3859) );
no02f01 g00071 ( .a(n3859), .b(delay_add_ln22_unr20_stage8_stallmux_q_7_), .o(n3860_1) );
in01f01 g00072 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_6_), .o(n3861) );
na02f01 g00073 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_6_), .b(n3790), .o(n3862) );
in01f01 g00074 ( .a(n3862), .o(n3863) );
no02f01 g00075 ( .a(n3863), .b(n3791), .o(n3864) );
in01f01 g00076 ( .a(n3864), .o(n3865_1) );
no02f01 g00077 ( .a(n3865_1), .b(n3804), .o(n3866) );
no02f01 g00078 ( .a(n3864), .b(n3805), .o(n3867) );
no02f01 g00079 ( .a(n3867), .b(n3866), .o(n3868) );
no02f01 g00080 ( .a(n3868), .b(n3861), .o(n3869) );
in01f01 g00081 ( .a(n3869), .o(n3870_1) );
na02f01 g00082 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_5_), .b(n3790), .o(n3871) );
in01f01 g00083 ( .a(n3871), .o(n3872) );
no02f01 g00084 ( .a(n3872), .b(n3792_1), .o(n3873) );
no02f01 g00085 ( .a(n3873), .b(n3803), .o(n3874) );
na02f01 g00086 ( .a(n3873), .b(n3803), .o(n3875_1) );
in01f01 g00087 ( .a(n3875_1), .o(n3876) );
no02f01 g00088 ( .a(n3876), .b(n3874), .o(n3877) );
in01f01 g00089 ( .a(n3877), .o(n3878) );
no02f01 g00090 ( .a(n3878), .b(delay_add_ln22_unr20_stage8_stallmux_q_5_), .o(n3879) );
in01f01 g00091 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_4_), .o(n3880_1) );
na02f01 g00092 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_4_), .b(n3790), .o(n3881) );
in01f01 g00093 ( .a(n3881), .o(n3882) );
no02f01 g00094 ( .a(n3882), .b(n3801), .o(n3883) );
in01f01 g00095 ( .a(n3883), .o(n3884) );
in01f01 g00096 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_2_), .o(n3885_1) );
na02f01 g00097 ( .a(n3885_1), .b(n_44962), .o(n3886) );
no02f01 g00098 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_1_), .b(n3790), .o(n3887) );
no02f01 g00099 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_0_), .b(n3790), .o(n3888) );
no02f01 g00100 ( .a(n3888), .b(n3887), .o(n3889) );
na02f01 g00101 ( .a(n3889), .b(n3886), .o(n3890_1) );
no02f01 g00102 ( .a(n3800), .b(n3890_1), .o(n3891) );
no02f01 g00103 ( .a(n3891), .b(n3884), .o(n3892) );
na02f01 g00104 ( .a(n3891), .b(n3884), .o(n3893) );
in01f01 g00105 ( .a(n3893), .o(n3894) );
no02f01 g00106 ( .a(n3894), .b(n3892), .o(n3895_1) );
no02f01 g00107 ( .a(n3895_1), .b(n3880_1), .o(n3896) );
in01f01 g00108 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_3_), .o(n3897) );
na02f01 g00109 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_3_), .b(n3790), .o(n3898) );
in01f01 g00110 ( .a(n3898), .o(n3899) );
no02f01 g00111 ( .a(n3899), .b(n3800), .o(n3900_1) );
no02f01 g00112 ( .a(n3900_1), .b(n3890_1), .o(n3901) );
no03f01 g00113 ( .a(n3899), .b(n3800), .c(n3799), .o(n3902) );
no02f01 g00114 ( .a(n3902), .b(n3901), .o(n3903) );
no02f01 g00115 ( .a(n3903), .b(n3897), .o(n3904) );
in01f01 g00116 ( .a(n3904), .o(n3905_1) );
in01f01 g00117 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_2_), .o(n3906) );
na02f01 g00118 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_2_), .b(n3790), .o(n3907) );
na02f01 g00119 ( .a(n3907), .b(n3886), .o(n3908) );
no02f01 g00120 ( .a(n3908), .b(n3889), .o(n3909) );
ao12f01 g00121 ( .a(n3798), .b(n3907), .c(n3886), .o(n3910_1) );
no02f01 g00122 ( .a(n3910_1), .b(n3909), .o(n3911) );
no02f01 g00123 ( .a(n3911), .b(n3906), .o(n3912) );
na02f01 g00124 ( .a(n3911), .b(n3906), .o(n3913) );
in01f01 g00125 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_0_), .o(n3914) );
na02f01 g00126 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_0_), .b(n_44962), .o(n3915_1) );
no02f01 g00127 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_0_), .b(n_44962), .o(n3916) );
in01f01 g00128 ( .a(n3916), .o(n3917) );
na02f01 g00129 ( .a(n3917), .b(n3915_1), .o(n3918) );
no02f01 g00130 ( .a(n3918), .b(n3914), .o(n3919) );
na02f01 g00131 ( .a(n3919), .b(delay_add_ln22_unr20_stage8_stallmux_q_1_), .o(n3920_1) );
na02f01 g00132 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_1_), .b(n3790), .o(n3921) );
na02f01 g00133 ( .a(n3921), .b(n3795), .o(n3922) );
no02f01 g00134 ( .a(n3922), .b(n3797_1), .o(n3923) );
ao12f01 g00135 ( .a(n3888), .b(n3921), .c(n3795), .o(n3924) );
no02f01 g00136 ( .a(n3924), .b(n3923), .o(n3925_1) );
no02f01 g00137 ( .a(n3919), .b(delay_add_ln22_unr20_stage8_stallmux_q_1_), .o(n3926) );
oa12f01 g00138 ( .a(n3920_1), .b(n3926), .c(n3925_1), .o(n3927) );
ao12f01 g00139 ( .a(n3912), .b(n3927), .c(n3913), .o(n3928) );
no03f01 g00140 ( .a(n3902), .b(n3901), .c(delay_add_ln22_unr20_stage8_stallmux_q_3_), .o(n3929) );
oa12f01 g00141 ( .a(n3905_1), .b(n3929), .c(n3928), .o(n3930_1) );
no03f01 g00142 ( .a(n3894), .b(n3892), .c(delay_add_ln22_unr20_stage8_stallmux_q_4_), .o(n3931) );
in01f01 g00143 ( .a(n3931), .o(n3932) );
ao12f01 g00144 ( .a(n3896), .b(n3932), .c(n3930_1), .o(n3933) );
na02f01 g00145 ( .a(n3878), .b(delay_add_ln22_unr20_stage8_stallmux_q_5_), .o(n3934) );
ao12f01 g00146 ( .a(n3879), .b(n3934), .c(n3933), .o(n3935_1) );
na02f01 g00147 ( .a(n3868), .b(n3861), .o(n3936) );
na02f01 g00148 ( .a(n3936), .b(n3935_1), .o(n3937) );
na02f01 g00149 ( .a(n3937), .b(n3870_1), .o(n3938) );
na02f01 g00150 ( .a(n3859), .b(delay_add_ln22_unr20_stage8_stallmux_q_7_), .o(n3939) );
in01f01 g00151 ( .a(n3939), .o(n3940_1) );
no02f01 g00152 ( .a(n3940_1), .b(n3938), .o(n3941) );
no02f01 g00153 ( .a(n3941), .b(n3860_1), .o(n3942) );
in01f01 g00154 ( .a(n3942), .o(n3943) );
na02f01 g00155 ( .a(n3849), .b(n3842), .o(n3944) );
in01f01 g00156 ( .a(n3944), .o(n3945_1) );
no02f01 g00157 ( .a(n3945_1), .b(n3943), .o(n3946) );
no02f01 g00158 ( .a(n3946), .b(n3850_1), .o(n3947) );
na02f01 g00159 ( .a(n3840), .b(delay_add_ln22_unr20_stage8_stallmux_q_9_), .o(n3948) );
ao12f01 g00160 ( .a(n3841_1), .b(n3948), .c(n3947), .o(n3949) );
in01f01 g00161 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_10_), .o(n3950_1) );
no02f01 g00162 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_10_), .b(n3790), .o(n3951) );
no02f01 g00163 ( .a(n3951), .b(n3814), .o(n3952) );
no02f01 g00164 ( .a(n3952), .b(n3811_1), .o(n3953) );
na02f01 g00165 ( .a(n3952), .b(n3811_1), .o(n3954) );
in01f01 g00166 ( .a(n3954), .o(n3955_1) );
no02f01 g00167 ( .a(n3955_1), .b(n3953), .o(n3956) );
no02f01 g00168 ( .a(n3956), .b(n3950_1), .o(n3957) );
in01f01 g00169 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_11_), .o(n3958) );
no02f01 g00170 ( .a(n3821_1), .b(n3958), .o(n3959) );
no02f01 g00171 ( .a(n3959), .b(n3957), .o(n3960_1) );
in01f01 g00172 ( .a(n3960_1), .o(n3961) );
na02f01 g00173 ( .a(n3956), .b(n3950_1), .o(n3962) );
in01f01 g00174 ( .a(n3962), .o(n3963) );
no02f01 g00175 ( .a(n3818), .b(delay_add_ln22_unr20_stage8_stallmux_q_11_), .o(n3964) );
no02f01 g00176 ( .a(n3964), .b(n3963), .o(n3965_1) );
oa12f01 g00177 ( .a(n3965_1), .b(n3961), .c(n3949), .o(n3966) );
in01f01 g00178 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_13_), .o(n3967) );
in01f01 g00179 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_12_), .o(n3968) );
ao12f01 g00180 ( .a(n3821_1), .b(n3968), .c(n3967), .o(n3969) );
in01f01 g00181 ( .a(n3969), .o(n3970_1) );
na02f01 g00182 ( .a(n3970_1), .b(n3966), .o(n3971) );
no02f01 g00183 ( .a(n3818), .b(delay_add_ln22_unr20_stage8_stallmux_q_14_), .o(n3972) );
no02f01 g00184 ( .a(n3818), .b(delay_add_ln22_unr20_stage8_stallmux_q_15_), .o(n3973) );
ao12f01 g00185 ( .a(n3818), .b(delay_add_ln22_unr20_stage8_stallmux_q_12_), .c(delay_add_ln22_unr20_stage8_stallmux_q_13_), .o(n3974) );
no03f01 g00186 ( .a(n3974), .b(n3973), .c(n3972), .o(n3975_1) );
oa12f01 g00187 ( .a(n3975_1), .b(n3971), .c(n3828), .o(n3976) );
no02f01 g00188 ( .a(n3976), .b(n3825), .o(n3977) );
no02f01 g00189 ( .a(n3818), .b(delay_add_ln22_unr20_stage8_stallmux_q_18_), .o(n3978) );
no02f01 g00190 ( .a(n3818), .b(delay_add_ln22_unr20_stage8_stallmux_q_19_), .o(n3979) );
no02f01 g00191 ( .a(n3979), .b(n3978), .o(n3980_1) );
no02f01 g00192 ( .a(n3818), .b(delay_add_ln22_unr20_stage8_stallmux_q_20_), .o(n3981) );
no02f01 g00193 ( .a(n3818), .b(delay_add_ln22_unr20_stage8_stallmux_q_21_), .o(n3982) );
no02f01 g00194 ( .a(n3982), .b(n3981), .o(n3983) );
na03f01 g00195 ( .a(n3983), .b(n3980_1), .c(n3977), .o(n3984) );
no02f01 g00196 ( .a(n3818), .b(delay_add_ln22_unr20_stage8_stallmux_q_22_), .o(n3985_1) );
no02f01 g00197 ( .a(n3985_1), .b(n3984), .o(n3986) );
in01f01 g00198 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_17_), .o(n3987) );
in01f01 g00199 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_16_), .o(n3988) );
ao12f01 g00200 ( .a(n3821_1), .b(n3988), .c(n3987), .o(n3989) );
in01f01 g00201 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_18_), .o(n3990_1) );
in01f01 g00202 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_19_), .o(n3991) );
ao12f01 g00203 ( .a(n3821_1), .b(n3991), .c(n3990_1), .o(n3992) );
no02f01 g00204 ( .a(n3992), .b(n3989), .o(n3993) );
in01f01 g00205 ( .a(n3993), .o(n3994_1) );
in01f01 g00206 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_21_), .o(n3995) );
in01f01 g00207 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_20_), .o(n3996) );
ao12f01 g00208 ( .a(n3821_1), .b(n3996), .c(n3995), .o(n3997) );
no02f01 g00209 ( .a(n3997), .b(n3994_1), .o(n3998) );
in01f01 g00210 ( .a(n3998), .o(n3999_1) );
in01f01 g00211 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_22_), .o(n4000) );
no02f01 g00212 ( .a(n3821_1), .b(n4000), .o(n4001) );
no02f01 g00213 ( .a(n4001), .b(n3999_1), .o(n4002) );
in01f01 g00214 ( .a(n4002), .o(n4003) );
no03f01 g00215 ( .a(n4003), .b(n3986), .c(n3824), .o(n4004_1) );
in01f01 g00216 ( .a(n4004_1), .o(n4005) );
oa12f01 g00217 ( .a(n3824), .b(n4003), .c(n3986), .o(n4006) );
na02f01 g00218 ( .a(n4006), .b(n4005), .o(n4007) );
in01f01 g00219 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_10_), .o(n4008) );
in01f01 g00220 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_9_), .o(n4009_1) );
in01f01 g00221 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_8_), .o(n4010) );
in01f01 g00222 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_1_), .o(n4011) );
na02f01 g00223 ( .a(n4011), .b(n_44962), .o(n4012) );
in01f01 g00224 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_0_), .o(n4013) );
na02f01 g00225 ( .a(n4013), .b(n_44962), .o(n4014_1) );
na02f01 g00226 ( .a(n4014_1), .b(n4012), .o(n4015) );
no02f01 g00227 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_4_), .b(n3790), .o(n4016) );
no02f01 g00228 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_3_), .b(n3790), .o(n4017) );
no02f01 g00229 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_2_), .b(n3790), .o(n4018) );
no02f01 g00230 ( .a(n4018), .b(n4017), .o(n4019_1) );
in01f01 g00231 ( .a(n4019_1), .o(n4020) );
no03f01 g00232 ( .a(n4020), .b(n4016), .c(n4015), .o(n4021) );
no02f01 g00233 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_5_), .b(n3790), .o(n4022) );
no02f01 g00234 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_7_), .b(n3790), .o(n4023) );
no02f01 g00235 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_6_), .b(n3790), .o(n4024_1) );
no02f01 g00236 ( .a(n4024_1), .b(n4023), .o(n4025) );
in01f01 g00237 ( .a(n4025), .o(n4026) );
no02f01 g00238 ( .a(n4026), .b(n4022), .o(n4027) );
na02f01 g00239 ( .a(n4027), .b(n4021), .o(n4028_1) );
no04f01 g00240 ( .a(n4028_1), .b(n4010), .c(n4009_1), .d(n3790), .o(n4029) );
no02f01 g00241 ( .a(n4029), .b(n4008), .o(n4030) );
in01f01 g00242 ( .a(n4030), .o(n4031) );
no02f01 g00243 ( .a(n4031), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_11_), .o(n4032) );
in01f01 g00244 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_9_), .o(n4033_1) );
in01f01 g00245 ( .a(n4021), .o(n4034) );
no02f01 g00246 ( .a(n4022), .b(n4034), .o(n4035) );
in01f01 g00247 ( .a(n4035), .o(n4036) );
no02f01 g00248 ( .a(n4036), .b(n4024_1), .o(n4037) );
no02f01 g00249 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_9_), .b(n3790), .o(n4038_1) );
no02f01 g00250 ( .a(n4009_1), .b(n_44962), .o(n4039) );
no02f01 g00251 ( .a(n4039), .b(n4038_1), .o(n4040) );
no02f01 g00252 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_8_), .b(n3790), .o(n4041) );
no03f01 g00253 ( .a(n4040), .b(n4041), .c(n4023), .o(n4042) );
in01f01 g00254 ( .a(n4028_1), .o(n4043_1) );
in01f01 g00255 ( .a(n4041), .o(n4044) );
na02f01 g00256 ( .a(n4044), .b(n4043_1), .o(n4045) );
ao22f01 g00257 ( .a(n4045), .b(n4040), .c(n4042), .d(n4037), .o(n4046) );
in01f01 g00258 ( .a(n4046), .o(n4047) );
no02f01 g00259 ( .a(n4047), .b(n4033_1), .o(n4048_1) );
in01f01 g00260 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_8_), .o(n4049) );
no02f01 g00261 ( .a(n4010), .b(n_44962), .o(n4050) );
no02f01 g00262 ( .a(n4050), .b(n4041), .o(n4051) );
no03f01 g00263 ( .a(n4051), .b(n4036), .c(n4026), .o(n4052) );
ao12f01 g00264 ( .a(n4052), .b(n4051), .c(n4028_1), .o(n4053_1) );
in01f01 g00265 ( .a(n4053_1), .o(n4054) );
no02f01 g00266 ( .a(n4054), .b(n4049), .o(n4055) );
in01f01 g00267 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_7_), .o(n4056) );
in01f01 g00268 ( .a(n4023), .o(n4057) );
na02f01 g00269 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_7_), .b(n3790), .o(n4058_1) );
na02f01 g00270 ( .a(n4058_1), .b(n4057), .o(n4059) );
no02f01 g00271 ( .a(n4059), .b(n4037), .o(n4060) );
in01f01 g00272 ( .a(n4022), .o(n4061) );
in01f01 g00273 ( .a(n4024_1), .o(n4062) );
na04f01 g00274 ( .a(n4059), .b(n4062), .c(n4061), .d(n4021), .o(n4063_1) );
in01f01 g00275 ( .a(n4063_1), .o(n4064) );
no03f01 g00276 ( .a(n4064), .b(n4060), .c(n4056), .o(n4065) );
na02f01 g00277 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_6_), .b(n3790), .o(n4066) );
na02f01 g00278 ( .a(n4066), .b(n4062), .o(n4067) );
no02f01 g00279 ( .a(n4067), .b(n4035), .o(n4068_1) );
in01f01 g00280 ( .a(n4068_1), .o(n4069) );
in01f01 g00281 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_6_), .o(n4070) );
no02f01 g00282 ( .a(n4020), .b(n4015), .o(n4071) );
in01f01 g00283 ( .a(n4071), .o(n4072) );
in01f01 g00284 ( .a(n4016), .o(n4073_1) );
na03f01 g00285 ( .a(n4067), .b(n4061), .c(n4073_1), .o(n4074) );
no02f01 g00286 ( .a(n4074), .b(n4072), .o(n4075) );
no02f01 g00287 ( .a(n4075), .b(n4070), .o(n4076) );
na02f01 g00288 ( .a(n4076), .b(n4069), .o(n4077) );
in01f01 g00289 ( .a(n4077), .o(n4078_1) );
na02f01 g00290 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_5_), .b(n3790), .o(n4079) );
na02f01 g00291 ( .a(n4079), .b(n4061), .o(n4080) );
in01f01 g00292 ( .a(n4080), .o(n4081) );
no02f01 g00293 ( .a(n4018), .b(n4015), .o(n4082) );
no03f01 g00294 ( .a(n4081), .b(n4017), .c(n4016), .o(n4083_1) );
ao22f01 g00295 ( .a(n4083_1), .b(n4082), .c(n4081), .d(n4034), .o(n4084) );
no02f01 g00296 ( .a(n4084), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_5_), .o(n4085) );
na02f01 g00297 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_4_), .b(n3790), .o(n4086) );
na02f01 g00298 ( .a(n4086), .b(n4073_1), .o(n4087) );
in01f01 g00299 ( .a(n4087), .o(n4088_1) );
no02f01 g00300 ( .a(n4088_1), .b(n4072), .o(n4089) );
no02f01 g00301 ( .a(n4087), .b(n4071), .o(n4090) );
no02f01 g00302 ( .a(n4090), .b(n4089), .o(n4091) );
no02f01 g00303 ( .a(n4091), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_4_), .o(n4092) );
in01f01 g00304 ( .a(n4092), .o(n4093_1) );
in01f01 g00305 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_3_), .o(n4094) );
na02f01 g00306 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_3_), .b(n3790), .o(n4095) );
in01f01 g00307 ( .a(n4095), .o(n4096) );
no02f01 g00308 ( .a(n4096), .b(n4017), .o(n4097) );
oa12f01 g00309 ( .a(n4097), .b(n4018), .c(n4015), .o(n4098_1) );
oa12f01 g00310 ( .a(n4082), .b(n4096), .c(n4017), .o(n4099) );
na02f01 g00311 ( .a(n4099), .b(n4098_1), .o(n4100) );
no02f01 g00312 ( .a(n4100), .b(n4094), .o(n4101) );
in01f01 g00313 ( .a(n4101), .o(n4102) );
in01f01 g00314 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_2_), .o(n4103_1) );
in01f01 g00315 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_2_), .o(n4104) );
no02f01 g00316 ( .a(n4104), .b(n_44962), .o(n4105) );
no02f01 g00317 ( .a(n4105), .b(n4018), .o(n4106) );
na02f01 g00318 ( .a(n4106), .b(n4015), .o(n4107_1) );
no02f01 g00319 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_1_), .b(n3790), .o(n4108) );
no02f01 g00320 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_0_), .b(n3790), .o(n4109) );
no02f01 g00321 ( .a(n4109), .b(n4108), .o(n4110) );
oa12f01 g00322 ( .a(n4110), .b(n4105), .c(n4018), .o(n4111) );
na02f01 g00323 ( .a(n4111), .b(n4107_1), .o(n4112_1) );
no02f01 g00324 ( .a(n4112_1), .b(n4103_1), .o(n4113) );
na02f01 g00325 ( .a(n4112_1), .b(n4103_1), .o(n4114) );
in01f01 g00326 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_1_), .o(n4115) );
no02f01 g00327 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_0_), .b(n_44962), .o(n4116_1) );
no02f01 g00328 ( .a(n4013), .b(n3790), .o(n4117) );
no02f01 g00329 ( .a(n4117), .b(n4116_1), .o(n4118) );
in01f01 g00330 ( .a(n4118), .o(n4119) );
no02f01 g00331 ( .a(n4119), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_0_), .o(n4120) );
no03f01 g00332 ( .a(n4119), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_1_), .c(delay_sub_ln21_0_unr20_stage8_stallmux_q_0_), .o(n4121_1) );
na03f01 g00333 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_1_), .b(n4013), .c(n_44962), .o(n4122) );
no02f01 g00334 ( .a(n4011), .b(n_44962), .o(n4123) );
oa12f01 g00335 ( .a(n4014_1), .b(n4123), .c(n4108), .o(n4124) );
na02f01 g00336 ( .a(n4124), .b(n4122), .o(n4125) );
oa22f01 g00337 ( .a(n4125), .b(n4121_1), .c(n4120), .d(n4115), .o(n4126_1) );
ao12f01 g00338 ( .a(n4113), .b(n4126_1), .c(n4114), .o(n4127) );
ao12f01 g00339 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_3_), .b(n4099), .c(n4098_1), .o(n4128) );
oa12f01 g00340 ( .a(n4102), .b(n4128), .c(n4127), .o(n4129) );
na02f01 g00341 ( .a(n4129), .b(n4093_1), .o(n4130) );
na02f01 g00342 ( .a(n4084), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_5_), .o(n4131_1) );
na02f01 g00343 ( .a(n4091), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_4_), .o(n4132) );
na02f01 g00344 ( .a(n4132), .b(n4131_1), .o(n4133) );
in01f01 g00345 ( .a(n4133), .o(n4134) );
ao12f01 g00346 ( .a(n4085), .b(n4134), .c(n4130), .o(n4135) );
oa12f01 g00347 ( .a(n4070), .b(n4075), .c(n4068_1), .o(n4136_1) );
ao12f01 g00348 ( .a(n4078_1), .b(n4136_1), .c(n4135), .o(n4137) );
in01f01 g00349 ( .a(n4137), .o(n4138) );
oa12f01 g00350 ( .a(n4056), .b(n4064), .c(n4060), .o(n4139) );
ao12f01 g00351 ( .a(n4065), .b(n4139), .c(n4138), .o(n4140) );
no02f01 g00352 ( .a(n4053_1), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_8_), .o(n4141_1) );
no02f01 g00353 ( .a(n4141_1), .b(n4140), .o(n4142) );
no02f01 g00354 ( .a(n4142), .b(n4055), .o(n4143) );
in01f01 g00355 ( .a(n4143), .o(n4144) );
no02f01 g00356 ( .a(n4144), .b(n4048_1), .o(n4145) );
no02f01 g00357 ( .a(n4046), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_9_), .o(n4146_1) );
no02f01 g00358 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_10_), .b(n3790), .o(n4147) );
no02f01 g00359 ( .a(n4008), .b(n_44962), .o(n4148) );
no02f01 g00360 ( .a(n4148), .b(n4147), .o(n4149) );
no03f01 g00361 ( .a(n4038_1), .b(n4041), .c(n4023), .o(n4150) );
na02f01 g00362 ( .a(n4150), .b(n4037), .o(n4151_1) );
no03f01 g00363 ( .a(n4149), .b(n4038_1), .c(n4041), .o(n4152) );
ao22f01 g00364 ( .a(n4152), .b(n4043_1), .c(n4151_1), .d(n4149), .o(n4153) );
no02f01 g00365 ( .a(n4153), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_10_), .o(n4154) );
no02f01 g00366 ( .a(n4154), .b(n4146_1), .o(n4155) );
in01f01 g00367 ( .a(n4155), .o(n4156_1) );
no02f01 g00368 ( .a(n4156_1), .b(n4145), .o(n4157) );
in01f01 g00369 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_11_), .o(n4158) );
na02f01 g00370 ( .a(n4153), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_10_), .o(n4159) );
ao12f01 g00371 ( .a(n4030), .b(n4159), .c(n4158), .o(n4160) );
no02f01 g00372 ( .a(n4160), .b(n4157), .o(n4161_1) );
in01f01 g00373 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_14_), .o(n4162) );
in01f01 g00374 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_15_), .o(n4163) );
ao12f01 g00375 ( .a(n4030), .b(n4163), .c(n4162), .o(n4164) );
in01f01 g00376 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_13_), .o(n4165) );
in01f01 g00377 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_12_), .o(n4166_1) );
ao12f01 g00378 ( .a(n4030), .b(n4166_1), .c(n4165), .o(n4167) );
no02f01 g00379 ( .a(n4167), .b(n4164), .o(n4168) );
oa12f01 g00380 ( .a(n4168), .b(n4161_1), .c(n4032), .o(n4169) );
no02f01 g00381 ( .a(n4031), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_13_), .o(n4170) );
no02f01 g00382 ( .a(n4031), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_12_), .o(n4171_1) );
no02f01 g00383 ( .a(n4171_1), .b(n4170), .o(n4172) );
in01f01 g00384 ( .a(n4172), .o(n4173) );
no02f01 g00385 ( .a(n4031), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_15_), .o(n4174) );
no02f01 g00386 ( .a(n4031), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_14_), .o(n4175) );
no03f01 g00387 ( .a(n4175), .b(n4174), .c(n4173), .o(n4176_1) );
no02f01 g00388 ( .a(n4031), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_20_), .o(n4177) );
no02f01 g00389 ( .a(n4031), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_21_), .o(n4178) );
no02f01 g00390 ( .a(n4178), .b(n4177), .o(n4179) );
in01f01 g00391 ( .a(n4179), .o(n4180) );
ao12f01 g00392 ( .a(n4031), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_16_), .c(delay_sub_ln21_0_unr20_stage8_stallmux_q_17_), .o(n4181_1) );
no02f01 g00393 ( .a(n4031), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_19_), .o(n4182) );
no02f01 g00394 ( .a(n4182), .b(n4181_1), .o(n4183) );
in01f01 g00395 ( .a(n4183), .o(n4184) );
no02f01 g00396 ( .a(n4031), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_18_), .o(n4185) );
no02f01 g00397 ( .a(n4031), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_22_), .o(n4186_1) );
no04f01 g00398 ( .a(n4186_1), .b(n4185), .c(n4184), .d(n4180), .o(n4187) );
na03f01 g00399 ( .a(n4187), .b(n4176_1), .c(n4169), .o(n4188) );
no02f01 g00400 ( .a(n4031), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_23_), .o(n4189) );
no02f01 g00401 ( .a(n4189), .b(n4188), .o(n4190) );
no02f01 g00402 ( .a(n4031), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_24_), .o(n4191_1) );
in01f01 g00403 ( .a(n4191_1), .o(n4192) );
na02f01 g00404 ( .a(n4192), .b(n4190), .o(n4193) );
no02f01 g00405 ( .a(n4031), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_25_), .o(n4194) );
no02f01 g00406 ( .a(n4194), .b(n4193), .o(n4195) );
no02f01 g00407 ( .a(n4031), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_26_), .o(n4196_1) );
no02f01 g00408 ( .a(n4031), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_27_), .o(n4197) );
no02f01 g00409 ( .a(n4197), .b(n4196_1), .o(n4198) );
in01f01 g00410 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_19_), .o(n4199) );
in01f01 g00411 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_18_), .o(n4200) );
ao12f01 g00412 ( .a(n4030), .b(n4200), .c(n4199), .o(n4201_1) );
in01f01 g00413 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_17_), .o(n4202) );
in01f01 g00414 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_16_), .o(n4203) );
ao12f01 g00415 ( .a(n4030), .b(n4203), .c(n4202), .o(n4204) );
no02f01 g00416 ( .a(n4204), .b(n4201_1), .o(n4205) );
in01f01 g00417 ( .a(n4205), .o(n4206_1) );
in01f01 g00418 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_21_), .o(n4207) );
in01f01 g00419 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_20_), .o(n4208) );
ao12f01 g00420 ( .a(n4030), .b(n4208), .c(n4207), .o(n4209) );
no02f01 g00421 ( .a(n4209), .b(n4206_1), .o(n4210) );
in01f01 g00422 ( .a(n4210), .o(n4211_1) );
in01f01 g00423 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_22_), .o(n4212) );
in01f01 g00424 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_23_), .o(n4213) );
ao12f01 g00425 ( .a(n4030), .b(n4213), .c(n4212), .o(n4214) );
no02f01 g00426 ( .a(n4214), .b(n4211_1), .o(n4215) );
in01f01 g00427 ( .a(n4215), .o(n4216_1) );
in01f01 g00428 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_24_), .o(n4217) );
in01f01 g00429 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_25_), .o(n4218) );
ao12f01 g00430 ( .a(n4030), .b(n4218), .c(n4217), .o(n4219) );
no02f01 g00431 ( .a(n4219), .b(n4216_1), .o(n4220) );
in01f01 g00432 ( .a(n4220), .o(n4221_1) );
in01f01 g00433 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_27_), .o(n4222) );
in01f01 g00434 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_26_), .o(n4223) );
ao12f01 g00435 ( .a(n4030), .b(n4223), .c(n4222), .o(n4224) );
no02f01 g00436 ( .a(n4224), .b(n4221_1), .o(n4225) );
in01f01 g00437 ( .a(n4225), .o(n4226_1) );
ao12f01 g00438 ( .a(n4226_1), .b(n4198), .c(n4195), .o(n4227) );
in01f01 g00439 ( .a(n4227), .o(n4228) );
in01f01 g00440 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_28_), .o(n4229) );
no02f01 g00441 ( .a(n4030), .b(n4229), .o(n4230) );
no02f01 g00442 ( .a(n4031), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_28_), .o(n4231_1) );
no02f01 g00443 ( .a(n4031), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_29_), .o(n4232) );
no02f01 g00444 ( .a(n4232), .b(n4231_1), .o(n4233) );
oa12f01 g00445 ( .a(n4233), .b(n4230), .c(n4228), .o(n4234) );
na02f01 g00446 ( .a(n4031), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_29_), .o(n4235) );
na02f01 g00447 ( .a(n4235), .b(n4234), .o(n4236_1) );
no02f01 g00448 ( .a(n4236_1), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_30_), .o(n4237) );
na02f01 g00449 ( .a(n4233), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_30_), .o(n4238) );
oa22f01 g00450 ( .a(n4238), .b(n4227), .c(n4237), .d(n4030), .o(n4239) );
no02f01 g00451 ( .a(n4031), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_31_), .o(n4240) );
na02f01 g00452 ( .a(n4031), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_31_), .o(n4241_1) );
in01f01 g00453 ( .a(n4241_1), .o(n4242) );
no02f01 g00454 ( .a(n4242), .b(n4240), .o(n4243) );
in01f01 g00455 ( .a(n4243), .o(n4244) );
no02f01 g00456 ( .a(n4244), .b(n4239), .o(n4245) );
na02f01 g00457 ( .a(n4244), .b(n4239), .o(n4246_1) );
in01f01 g00458 ( .a(n4246_1), .o(n4247) );
no02f01 g00459 ( .a(n4247), .b(n4245), .o(n4248) );
in01f01 g00460 ( .a(delay_sub_ln23_0_unr21_stage8_stallmux_q), .o(n4249) );
no02f01 g00461 ( .a(n4248), .b(n4249), .o(n4250) );
in01f01 g00462 ( .a(n4231_1), .o(n4251_1) );
oa12f01 g00463 ( .a(n4251_1), .b(n4230), .c(n4228), .o(n4252) );
in01f01 g00464 ( .a(n4235), .o(n4253) );
no02f01 g00465 ( .a(n4253), .b(n4232), .o(n4254) );
na02f01 g00466 ( .a(n4254), .b(n4252), .o(n4255) );
in01f01 g00467 ( .a(n4255), .o(n4256_1) );
no02f01 g00468 ( .a(n4254), .b(n4252), .o(n4257) );
no02f01 g00469 ( .a(n4257), .b(n4256_1), .o(n4258) );
no02f01 g00470 ( .a(n4231_1), .b(n4230), .o(n4259) );
in01f01 g00471 ( .a(n4259), .o(n4260) );
no02f01 g00472 ( .a(n4260), .b(n4228), .o(n4261_1) );
no02f01 g00473 ( .a(n4259), .b(n4227), .o(n4262) );
no02f01 g00474 ( .a(n4262), .b(n4261_1), .o(n4263) );
no02f01 g00475 ( .a(n4263), .b(n4249), .o(n4264) );
no02f01 g00476 ( .a(n4030), .b(n4223), .o(n4265) );
no02f01 g00477 ( .a(n4221_1), .b(n4195), .o(n4266_1) );
in01f01 g00478 ( .a(n4266_1), .o(n4267) );
no02f01 g00479 ( .a(n4267), .b(n4265), .o(n4268) );
no02f01 g00480 ( .a(n4030), .b(n4222), .o(n4269) );
no02f01 g00481 ( .a(n4269), .b(n4197), .o(n4270) );
oa12f01 g00482 ( .a(n4270), .b(n4268), .c(n4196_1), .o(n4271_1) );
in01f01 g00483 ( .a(n4271_1), .o(n4272) );
no03f01 g00484 ( .a(n4270), .b(n4268), .c(n4196_1), .o(n4273) );
no02f01 g00485 ( .a(n4273), .b(n4272), .o(n4274) );
no02f01 g00486 ( .a(n4265), .b(n4196_1), .o(n4275_1) );
na02f01 g00487 ( .a(n4275_1), .b(n4266_1), .o(n4276) );
in01f01 g00488 ( .a(n4276), .o(n4277) );
no02f01 g00489 ( .a(n4275_1), .b(n4266_1), .o(n4278) );
no02f01 g00490 ( .a(n4278), .b(n4277), .o(n4279) );
no02f01 g00491 ( .a(n4030), .b(n4212), .o(n4280_1) );
no02f01 g00492 ( .a(n4280_1), .b(n4186_1), .o(n4281) );
in01f01 g00493 ( .a(n4281), .o(n4282) );
no02f01 g00494 ( .a(n4161_1), .b(n4032), .o(n4283) );
in01f01 g00495 ( .a(n4168), .o(n4284) );
no02f01 g00496 ( .a(n4284), .b(n4283), .o(n4285_1) );
in01f01 g00497 ( .a(n4176_1), .o(n4286) );
no02f01 g00498 ( .a(n4185), .b(n4184), .o(n4287) );
in01f01 g00499 ( .a(n4287), .o(n4288) );
no04f01 g00500 ( .a(n4288), .b(n4180), .c(n4286), .d(n4285_1), .o(n4289) );
no03f01 g00501 ( .a(n4289), .b(n4282), .c(n4211_1), .o(n4290_1) );
na04f01 g00502 ( .a(n4287), .b(n4179), .c(n4176_1), .d(n4169), .o(n4291) );
ao12f01 g00503 ( .a(n4281), .b(n4291), .c(n4210), .o(n4292) );
oa12f01 g00504 ( .a(delay_sub_ln23_0_unr21_stage8_stallmux_q), .b(n4292), .c(n4290_1), .o(n4293) );
no02f01 g00505 ( .a(n4030), .b(n4213), .o(n4294) );
no02f01 g00506 ( .a(n4294), .b(n4189), .o(n4295_1) );
no02f01 g00507 ( .a(n4280_1), .b(n4211_1), .o(n4296) );
na03f01 g00508 ( .a(n4296), .b(n4295_1), .c(n4188), .o(n4297) );
in01f01 g00509 ( .a(n4295_1), .o(n4298) );
na02f01 g00510 ( .a(n4296), .b(n4188), .o(n4299) );
na02f01 g00511 ( .a(n4299), .b(n4298), .o(n4300_1) );
na02f01 g00512 ( .a(n4300_1), .b(n4297), .o(n4301) );
na02f01 g00513 ( .a(n4301), .b(delay_sub_ln23_0_unr21_stage8_stallmux_q), .o(n4302) );
na02f01 g00514 ( .a(n4302), .b(n4293), .o(n4303) );
in01f01 g00515 ( .a(n4187), .o(n4304) );
no03f01 g00516 ( .a(n4304), .b(n4286), .c(n4285_1), .o(n4305_1) );
in01f01 g00517 ( .a(n4189), .o(n4306) );
na02f01 g00518 ( .a(n4306), .b(n4305_1), .o(n4307) );
no02f01 g00519 ( .a(n4030), .b(n4217), .o(n4308) );
no02f01 g00520 ( .a(n4308), .b(n4191_1), .o(n4309) );
ao12f01 g00521 ( .a(n4309), .b(n4215), .c(n4307), .o(n4310_1) );
in01f01 g00522 ( .a(n4309), .o(n4311) );
no03f01 g00523 ( .a(n4311), .b(n4216_1), .c(n4190), .o(n4312) );
no02f01 g00524 ( .a(n4312), .b(n4310_1), .o(n4313) );
no02f01 g00525 ( .a(n4313), .b(n4249), .o(n4314) );
no02f01 g00526 ( .a(n4308), .b(n4216_1), .o(n4315_1) );
no02f01 g00527 ( .a(n4030), .b(n4218), .o(n4316) );
no02f01 g00528 ( .a(n4316), .b(n4194), .o(n4317) );
na03f01 g00529 ( .a(n4317), .b(n4315_1), .c(n4193), .o(n4318) );
na02f01 g00530 ( .a(n4315_1), .b(n4193), .o(n4319) );
in01f01 g00531 ( .a(n4317), .o(n4320_1) );
na02f01 g00532 ( .a(n4320_1), .b(n4319), .o(n4321) );
na02f01 g00533 ( .a(n4321), .b(n4318), .o(n4322) );
no03f01 g00534 ( .a(n4322), .b(n4314), .c(n4303), .o(n4323) );
ao12f01 g00535 ( .a(n4249), .b(n4323), .c(n4279), .o(n4324) );
in01f01 g00536 ( .a(n4324), .o(n4325_1) );
oa12f01 g00537 ( .a(n4325_1), .b(n4274), .c(n4249), .o(n4326) );
no02f01 g00538 ( .a(n4326), .b(n4264), .o(n4327) );
oa12f01 g00539 ( .a(n4327), .b(n4258), .c(n4249), .o(n4328) );
no02f01 g00540 ( .a(n4031), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_30_), .o(n4329) );
in01f01 g00541 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_30_), .o(n4330_1) );
no02f01 g00542 ( .a(n4030), .b(n4330_1), .o(n4331) );
no02f01 g00543 ( .a(n4331), .b(n4329), .o(n4332) );
in01f01 g00544 ( .a(n4332), .o(n4333) );
na02f01 g00545 ( .a(n4333), .b(n4236_1), .o(n4334_1) );
in01f01 g00546 ( .a(n4334_1), .o(n4335) );
no02f01 g00547 ( .a(n4333), .b(n4236_1), .o(n4336) );
no02f01 g00548 ( .a(n4336), .b(n4335), .o(n4337) );
in01f01 g00549 ( .a(n4337), .o(n4338) );
ao12f01 g00550 ( .a(n4328), .b(n4338), .c(delay_sub_ln23_0_unr21_stage8_stallmux_q), .o(n4339_1) );
ao12f01 g00551 ( .a(n4250), .b(n4339_1), .c(n4248), .o(n4340) );
no02f01 g00552 ( .a(n4340), .b(n4007), .o(n4341) );
in01f01 g00553 ( .a(n4006), .o(n4342) );
no02f01 g00554 ( .a(n4342), .b(n4004_1), .o(n4343) );
in01f01 g00555 ( .a(n4340), .o(n4344_1) );
no02f01 g00556 ( .a(n4344_1), .b(n4343), .o(n4345) );
no02f01 g00557 ( .a(n4345), .b(n4341), .o(n4346) );
in01f01 g00558 ( .a(n4346), .o(n4347) );
ao12f01 g00559 ( .a(n3994_1), .b(n3980_1), .c(n3977), .o(n4348) );
no02f01 g00560 ( .a(n3821_1), .b(n3996), .o(n4349_1) );
no02f01 g00561 ( .a(n4349_1), .b(n3981), .o(n4350) );
no02f01 g00562 ( .a(n4350), .b(n4348), .o(n4351) );
na02f01 g00563 ( .a(n4350), .b(n4348), .o(n4352) );
in01f01 g00564 ( .a(n4352), .o(n4353) );
no02f01 g00565 ( .a(n4353), .b(n4351), .o(n4354_1) );
in01f01 g00566 ( .a(n4354_1), .o(n4355) );
in01f01 g00567 ( .a(n3977), .o(n4356) );
in01f01 g00568 ( .a(n3980_1), .o(n4357) );
no03f01 g00569 ( .a(n3981), .b(n4357), .c(n4356), .o(n4358) );
no03f01 g00570 ( .a(n4358), .b(n4349_1), .c(n3994_1), .o(n4359_1) );
in01f01 g00571 ( .a(n4359_1), .o(n4360) );
no02f01 g00572 ( .a(n3821_1), .b(n3995), .o(n4361) );
no02f01 g00573 ( .a(n4361), .b(n3982), .o(n4362) );
in01f01 g00574 ( .a(n4362), .o(n4363) );
no02f01 g00575 ( .a(n4363), .b(n4360), .o(n4364_1) );
no02f01 g00576 ( .a(n4362), .b(n4359_1), .o(n4365) );
no02f01 g00577 ( .a(n4365), .b(n4364_1), .o(n4366) );
in01f01 g00578 ( .a(n4366), .o(n4367) );
ao12f01 g00579 ( .a(n4340), .b(n4367), .c(n4355), .o(n4368) );
in01f01 g00580 ( .a(n4368), .o(n4369_1) );
in01f01 g00581 ( .a(n4258), .o(n4370) );
in01f01 g00582 ( .a(n4264), .o(n4371) );
in01f01 g00583 ( .a(n4273), .o(n4372) );
na02f01 g00584 ( .a(n4372), .b(n4271_1), .o(n4373) );
ao12f01 g00585 ( .a(n4324), .b(n4373), .c(delay_sub_ln23_0_unr21_stage8_stallmux_q), .o(n4374_1) );
na02f01 g00586 ( .a(n4374_1), .b(n4371), .o(n4375) );
ao12f01 g00587 ( .a(n4375), .b(n4370), .c(delay_sub_ln23_0_unr21_stage8_stallmux_q), .o(n4376) );
oa12f01 g00588 ( .a(n4376), .b(n4337), .c(n4249), .o(n4377) );
na02f01 g00589 ( .a(n4377), .b(n4248), .o(n4378) );
in01f01 g00590 ( .a(n4248), .o(n4379_1) );
na02f01 g00591 ( .a(n4339_1), .b(n4379_1), .o(n4380) );
na02f01 g00592 ( .a(n4380), .b(n4378), .o(n4381) );
in01f01 g00593 ( .a(n3948), .o(n4382) );
no02f01 g00594 ( .a(n4382), .b(n3841_1), .o(n4383) );
in01f01 g00595 ( .a(n4383), .o(n4384_1) );
no03f01 g00596 ( .a(n4384_1), .b(n3946), .c(n3850_1), .o(n4385) );
no02f01 g00597 ( .a(n4383), .b(n3947), .o(n4386) );
no02f01 g00598 ( .a(n4386), .b(n4385), .o(n4387) );
in01f01 g00599 ( .a(n4387), .o(n4388) );
no02f01 g00600 ( .a(n4388), .b(n4381), .o(n4389_1) );
no02f01 g00601 ( .a(n4338), .b(n4376), .o(n4390) );
no02f01 g00602 ( .a(n4337), .b(n4328), .o(n4391) );
no02f01 g00603 ( .a(n4391), .b(n4390), .o(n4392) );
no02f01 g00604 ( .a(n3945_1), .b(n3850_1), .o(n4393) );
no02f01 g00605 ( .a(n4393), .b(n3943), .o(n4394_1) );
na02f01 g00606 ( .a(n4393), .b(n3943), .o(n4395) );
in01f01 g00607 ( .a(n4395), .o(n4396) );
no02f01 g00608 ( .a(n4396), .b(n4394_1), .o(n4397) );
no02f01 g00609 ( .a(n4397), .b(n4392), .o(n4398) );
no02f01 g00610 ( .a(n4264), .b(n4258), .o(n4399_1) );
ao22f01 g00611 ( .a(n4399_1), .b(n4374_1), .c(n4375), .d(n4258), .o(n4400) );
no02f01 g00612 ( .a(n3940_1), .b(n3860_1), .o(n4401) );
in01f01 g00613 ( .a(n4401), .o(n4402) );
no02f01 g00614 ( .a(n4402), .b(n3938), .o(n4403) );
na02f01 g00615 ( .a(n4402), .b(n3938), .o(n4404_1) );
in01f01 g00616 ( .a(n4404_1), .o(n4405) );
no02f01 g00617 ( .a(n4405), .b(n4403), .o(n4406) );
no02f01 g00618 ( .a(n4406), .b(n4400), .o(n4407) );
in01f01 g00619 ( .a(n4407), .o(n4408) );
na02f01 g00620 ( .a(n4399_1), .b(n4374_1), .o(n4409_1) );
oa12f01 g00621 ( .a(n4409_1), .b(n4327), .c(n4370), .o(n4410) );
in01f01 g00622 ( .a(n4406), .o(n4411) );
in01f01 g00623 ( .a(n4263), .o(n4412) );
na02f01 g00624 ( .a(n4374_1), .b(n4412), .o(n4413) );
na02f01 g00625 ( .a(n4326), .b(n4263), .o(n4414_1) );
na02f01 g00626 ( .a(n3936), .b(n3870_1), .o(n4415) );
no02f01 g00627 ( .a(n4415), .b(n3935_1), .o(n4416) );
na02f01 g00628 ( .a(n4415), .b(n3935_1), .o(n4417) );
in01f01 g00629 ( .a(n4417), .o(n4418) );
no02f01 g00630 ( .a(n4418), .b(n4416), .o(n4419_1) );
ao12f01 g00631 ( .a(n4419_1), .b(n4414_1), .c(n4413), .o(n4420) );
na02f01 g00632 ( .a(n4324), .b(n4274), .o(n4421) );
na02f01 g00633 ( .a(n4325_1), .b(n4373), .o(n4422) );
in01f01 g00634 ( .a(n3933), .o(n4423) );
in01f01 g00635 ( .a(n3934), .o(n4424_1) );
no03f01 g00636 ( .a(n4424_1), .b(n4423), .c(n3879), .o(n4425) );
in01f01 g00637 ( .a(n3879), .o(n4426) );
ao12f01 g00638 ( .a(n3933), .b(n3934), .c(n4426), .o(n4427) );
no02f01 g00639 ( .a(n4427), .b(n4425), .o(n4428) );
ao12f01 g00640 ( .a(n4428), .b(n4422), .c(n4421), .o(n4429_1) );
in01f01 g00641 ( .a(n4429_1), .o(n4430) );
no02f01 g00642 ( .a(n4323), .b(n4249), .o(n4431) );
na02f01 g00643 ( .a(n4431), .b(n4279), .o(n4432) );
in01f01 g00644 ( .a(n4278), .o(n4433) );
na02f01 g00645 ( .a(n4433), .b(n4276), .o(n4434_1) );
oa12f01 g00646 ( .a(n4434_1), .b(n4323), .c(n4249), .o(n4435) );
no03f01 g00647 ( .a(n3931), .b(n3930_1), .c(n3896), .o(n4436) );
in01f01 g00648 ( .a(n3930_1), .o(n4437) );
no02f01 g00649 ( .a(n3931), .b(n3896), .o(n4438) );
no02f01 g00650 ( .a(n4438), .b(n4437), .o(n4439_1) );
no02f01 g00651 ( .a(n4439_1), .b(n4436), .o(n4440) );
ao12f01 g00652 ( .a(n4440), .b(n4435), .c(n4432), .o(n4441) );
no03f01 g00653 ( .a(n4323), .b(n4434_1), .c(n4249), .o(n4442) );
no02f01 g00654 ( .a(n4431), .b(n4279), .o(n4443_1) );
in01f01 g00655 ( .a(n4440), .o(n4444) );
no03f01 g00656 ( .a(n4444), .b(n4443_1), .c(n4442), .o(n4445) );
in01f01 g00657 ( .a(n4318), .o(n4446) );
ao12f01 g00658 ( .a(n4317), .b(n4315_1), .c(n4193), .o(n4447) );
no02f01 g00659 ( .a(n4447), .b(n4446), .o(n4448_1) );
oa12f01 g00660 ( .a(n4448_1), .b(n4314), .c(n4303), .o(n4449) );
no02f01 g00661 ( .a(n4292), .b(n4290_1), .o(n4450) );
no02f01 g00662 ( .a(n4450), .b(n4249), .o(n4451) );
in01f01 g00663 ( .a(n4297), .o(n4452) );
ao12f01 g00664 ( .a(n4295_1), .b(n4296), .c(n4188), .o(n4453_1) );
no02f01 g00665 ( .a(n4453_1), .b(n4452), .o(n4454) );
no02f01 g00666 ( .a(n4454), .b(n4249), .o(n4455) );
no02f01 g00667 ( .a(n4455), .b(n4451), .o(n4456) );
oa12f01 g00668 ( .a(n4311), .b(n4216_1), .c(n4190), .o(n4457) );
in01f01 g00669 ( .a(n4312), .o(n4458_1) );
na02f01 g00670 ( .a(n4458_1), .b(n4457), .o(n4459) );
na02f01 g00671 ( .a(n4459), .b(delay_sub_ln23_0_unr21_stage8_stallmux_q), .o(n4460) );
na03f01 g00672 ( .a(n4322), .b(n4460), .c(n4456), .o(n4461) );
no02f01 g00673 ( .a(n3929), .b(n3904), .o(n4462) );
no02f01 g00674 ( .a(n4462), .b(n3928), .o(n4463_1) );
na02f01 g00675 ( .a(n4462), .b(n3928), .o(n4464) );
in01f01 g00676 ( .a(n4464), .o(n4465) );
no02f01 g00677 ( .a(n4465), .b(n4463_1), .o(n4466) );
ao12f01 g00678 ( .a(n4466), .b(n4461), .c(n4449), .o(n4467) );
in01f01 g00679 ( .a(n4467), .o(n4468_1) );
ao12f01 g00680 ( .a(n4459), .b(n4302), .c(n4293), .o(n4469) );
no03f01 g00681 ( .a(n4313), .b(n4455), .c(n4451), .o(n4470) );
no02f01 g00682 ( .a(n4470), .b(n4469), .o(n4471) );
in01f01 g00683 ( .a(n3927), .o(n4472) );
in01f01 g00684 ( .a(n3913), .o(n4473_1) );
no02f01 g00685 ( .a(n4473_1), .b(n3912), .o(n4474) );
no02f01 g00686 ( .a(n4474), .b(n4472), .o(n4475) );
na02f01 g00687 ( .a(n4474), .b(n4472), .o(n4476) );
in01f01 g00688 ( .a(n4476), .o(n4477) );
no02f01 g00689 ( .a(n4477), .b(n4475), .o(n4478_1) );
no02f01 g00690 ( .a(n4478_1), .b(n4471), .o(n4479) );
no02f01 g00691 ( .a(n3918), .b(delay_add_ln22_unr20_stage8_stallmux_q_0_), .o(n4480) );
ao12f01 g00692 ( .a(n3914), .b(n3917), .c(n3915_1), .o(n4481) );
no02f01 g00693 ( .a(n4481), .b(n4480), .o(n4482) );
no02f01 g00694 ( .a(n4482), .b(n4450), .o(n4483_1) );
in01f01 g00695 ( .a(n4483_1), .o(n4484) );
no03f01 g00696 ( .a(n3924), .b(n3923), .c(delay_add_ln22_unr20_stage8_stallmux_q_1_), .o(n4485) );
in01f01 g00697 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_1_), .o(n4486) );
no02f01 g00698 ( .a(n3925_1), .b(n4486), .o(n4487) );
no03f01 g00699 ( .a(n4487), .b(n4485), .c(n3919), .o(n4488_1) );
in01f01 g00700 ( .a(n3919), .o(n4489) );
no02f01 g00701 ( .a(n4487), .b(n4485), .o(n4490) );
no02f01 g00702 ( .a(n4490), .b(n4489), .o(n4491) );
no02f01 g00703 ( .a(n4491), .b(n4488_1), .o(n4492) );
no02f01 g00704 ( .a(n4492), .b(n4484), .o(n4493_1) );
in01f01 g00705 ( .a(n4493_1), .o(n4494) );
in01f01 g00706 ( .a(n4492), .o(n4495) );
na03f01 g00707 ( .a(n4291), .b(n4281), .c(n4210), .o(n4496) );
in01f01 g00708 ( .a(n4292), .o(n4497) );
na02f01 g00709 ( .a(n4497), .b(n4496), .o(n4498_1) );
ao12f01 g00710 ( .a(n4454), .b(n4498_1), .c(delay_sub_ln23_0_unr21_stage8_stallmux_q), .o(n4499) );
no02f01 g00711 ( .a(n4301), .b(n4293), .o(n4500) );
oa22f01 g00712 ( .a(n4500), .b(n4499), .c(n4495), .d(n4483_1), .o(n4501) );
ao22f01 g00713 ( .a(n4501), .b(n4494), .c(n4478_1), .d(n4471), .o(n4502) );
na03f01 g00714 ( .a(n4466), .b(n4461), .c(n4449), .o(n4503_1) );
oa12f01 g00715 ( .a(n4503_1), .b(n4502), .c(n4479), .o(n4504) );
ao12f01 g00716 ( .a(n4445), .b(n4504), .c(n4468_1), .o(n4505) );
na03f01 g00717 ( .a(n4428), .b(n4422), .c(n4421), .o(n4506) );
oa12f01 g00718 ( .a(n4506), .b(n4505), .c(n4441), .o(n4507) );
no02f01 g00719 ( .a(n4326), .b(n4263), .o(n4508_1) );
no02f01 g00720 ( .a(n4374_1), .b(n4412), .o(n4509) );
in01f01 g00721 ( .a(n4419_1), .o(n4510) );
no03f01 g00722 ( .a(n4510), .b(n4509), .c(n4508_1), .o(n4511) );
ao12f01 g00723 ( .a(n4511), .b(n4507), .c(n4430), .o(n4512) );
oa22f01 g00724 ( .a(n4512), .b(n4420), .c(n4411), .d(n4410), .o(n4513_1) );
in01f01 g00725 ( .a(n4397), .o(n4514) );
no03f01 g00726 ( .a(n4514), .b(n4391), .c(n4390), .o(n4515) );
ao12f01 g00727 ( .a(n4515), .b(n4513_1), .c(n4408), .o(n4516) );
ao12f01 g00728 ( .a(n4387), .b(n4380), .c(n4378), .o(n4517) );
no03f01 g00729 ( .a(n4517), .b(n4516), .c(n4398), .o(n4518_1) );
ao12f01 g00730 ( .a(n3957), .b(n3962), .c(n3949), .o(n4519) );
in01f01 g00731 ( .a(n4519), .o(n4520) );
no02f01 g00732 ( .a(n3964), .b(n3959), .o(n4521) );
in01f01 g00733 ( .a(n4521), .o(n4522) );
no02f01 g00734 ( .a(n4522), .b(n4520), .o(n4523_1) );
no02f01 g00735 ( .a(n4521), .b(n4519), .o(n4524) );
no02f01 g00736 ( .a(n4524), .b(n4523_1), .o(n4525) );
in01f01 g00737 ( .a(n4525), .o(n4526) );
in01f01 g00738 ( .a(n3949), .o(n4527) );
no02f01 g00739 ( .a(n3963), .b(n3957), .o(n4528_1) );
no02f01 g00740 ( .a(n4528_1), .b(n4527), .o(n4529) );
na02f01 g00741 ( .a(n4528_1), .b(n4527), .o(n4530) );
in01f01 g00742 ( .a(n4530), .o(n4531) );
no02f01 g00743 ( .a(n4531), .b(n4529), .o(n4532) );
in01f01 g00744 ( .a(n4532), .o(n4533_1) );
oa12f01 g00745 ( .a(n4340), .b(n4533_1), .c(n4526), .o(n4534) );
oa12f01 g00746 ( .a(n4534), .b(n4518_1), .c(n4389_1), .o(n4535) );
no02f01 g00747 ( .a(n4533_1), .b(n4340), .o(n4536) );
no02f01 g00748 ( .a(n4526), .b(n4340), .o(n4537) );
no02f01 g00749 ( .a(n4537), .b(n4536), .o(n4538_1) );
no02f01 g00750 ( .a(n3821_1), .b(n3968), .o(n4539) );
no02f01 g00751 ( .a(n3818), .b(delay_add_ln22_unr20_stage8_stallmux_q_12_), .o(n4540) );
no02f01 g00752 ( .a(n4540), .b(n4539), .o(n4541) );
no02f01 g00753 ( .a(n4541), .b(n3966), .o(n4542) );
na02f01 g00754 ( .a(n4541), .b(n3966), .o(n4543_1) );
in01f01 g00755 ( .a(n4543_1), .o(n4544) );
no02f01 g00756 ( .a(n4544), .b(n4542), .o(n4545) );
in01f01 g00757 ( .a(n4545), .o(n4546) );
no02f01 g00758 ( .a(n4546), .b(n4340), .o(n4547) );
in01f01 g00759 ( .a(n4547), .o(n4548_1) );
in01f01 g00760 ( .a(n3974), .o(n4549) );
no02f01 g00761 ( .a(n3821_1), .b(n3826_1), .o(n4550) );
no02f01 g00762 ( .a(n3972), .b(n4550), .o(n4551) );
in01f01 g00763 ( .a(n4551), .o(n4552) );
ao12f01 g00764 ( .a(n4552), .b(n4549), .c(n3971), .o(n4553_1) );
na02f01 g00765 ( .a(n4549), .b(n3971), .o(n4554) );
no02f01 g00766 ( .a(n4551), .b(n4554), .o(n4555) );
no02f01 g00767 ( .a(n4555), .b(n4553_1), .o(n4556) );
in01f01 g00768 ( .a(n4556), .o(n4557) );
no02f01 g00769 ( .a(n4557), .b(n4340), .o(n4558_1) );
in01f01 g00770 ( .a(n4539), .o(n4559) );
ao12f01 g00771 ( .a(n4540), .b(n4559), .c(n3966), .o(n4560) );
no02f01 g00772 ( .a(n3818), .b(delay_add_ln22_unr20_stage8_stallmux_q_13_), .o(n4561) );
no02f01 g00773 ( .a(n3821_1), .b(n3967), .o(n4562) );
no02f01 g00774 ( .a(n4562), .b(n4561), .o(n4563_1) );
in01f01 g00775 ( .a(n4563_1), .o(n4564) );
no02f01 g00776 ( .a(n4564), .b(n4560), .o(n4565) );
na02f01 g00777 ( .a(n4564), .b(n4560), .o(n4566) );
in01f01 g00778 ( .a(n4566), .o(n4567) );
no02f01 g00779 ( .a(n4567), .b(n4565), .o(n4568_1) );
in01f01 g00780 ( .a(n4568_1), .o(n4569) );
no02f01 g00781 ( .a(n4569), .b(n4340), .o(n4570) );
no03f01 g00782 ( .a(n3974), .b(n3972), .c(n3966), .o(n4571) );
no03f01 g00783 ( .a(n4571), .b(n3969), .c(n4550), .o(n4572) );
in01f01 g00784 ( .a(n4572), .o(n4573_1) );
no02f01 g00785 ( .a(n3821_1), .b(n3827), .o(n4574) );
no02f01 g00786 ( .a(n4574), .b(n3973), .o(n4575) );
in01f01 g00787 ( .a(n4575), .o(n4576) );
no02f01 g00788 ( .a(n4576), .b(n4573_1), .o(n4577) );
no02f01 g00789 ( .a(n4575), .b(n4572), .o(n4578_1) );
no02f01 g00790 ( .a(n4578_1), .b(n4577), .o(n4579) );
in01f01 g00791 ( .a(n4579), .o(n4580) );
no02f01 g00792 ( .a(n4580), .b(n4340), .o(n4581) );
no03f01 g00793 ( .a(n4581), .b(n4570), .c(n4558_1), .o(n4582) );
na04f01 g00794 ( .a(n4582), .b(n4548_1), .c(n4538_1), .d(n4535), .o(n4583_1) );
ao12f01 g00795 ( .a(n4344_1), .b(n4579), .c(n4556), .o(n4584) );
ao12f01 g00796 ( .a(n4344_1), .b(n4568_1), .c(n4545), .o(n4585) );
no02f01 g00797 ( .a(n4585), .b(n4584), .o(n4586) );
na02f01 g00798 ( .a(n4586), .b(n4583_1), .o(n4587) );
in01f01 g00799 ( .a(n3976), .o(n4588_1) );
no02f01 g00800 ( .a(n3821_1), .b(n3988), .o(n4589) );
no02f01 g00801 ( .a(n3818), .b(delay_add_ln22_unr20_stage8_stallmux_q_16_), .o(n4590) );
in01f01 g00802 ( .a(n4590), .o(n4591) );
ao12f01 g00803 ( .a(n4589), .b(n4591), .c(n4588_1), .o(n4592) );
in01f01 g00804 ( .a(n4592), .o(n4593_1) );
no02f01 g00805 ( .a(n3818), .b(delay_add_ln22_unr20_stage8_stallmux_q_17_), .o(n4594) );
no02f01 g00806 ( .a(n3821_1), .b(n3987), .o(n4595) );
no02f01 g00807 ( .a(n4595), .b(n4594), .o(n4596) );
in01f01 g00808 ( .a(n4596), .o(n4597) );
no02f01 g00809 ( .a(n4597), .b(n4593_1), .o(n4598_1) );
no02f01 g00810 ( .a(n4596), .b(n4592), .o(n4599) );
no02f01 g00811 ( .a(n4599), .b(n4598_1), .o(n4600) );
in01f01 g00812 ( .a(n4600), .o(n4601) );
no02f01 g00813 ( .a(n4601), .b(n4340), .o(n4602) );
no02f01 g00814 ( .a(n4590), .b(n4589), .o(n4603_1) );
no02f01 g00815 ( .a(n4603_1), .b(n3976), .o(n4604) );
na02f01 g00816 ( .a(n4603_1), .b(n3976), .o(n4605) );
in01f01 g00817 ( .a(n4605), .o(n4606) );
no02f01 g00818 ( .a(n4606), .b(n4604), .o(n4607) );
in01f01 g00819 ( .a(n4607), .o(n4608_1) );
no02f01 g00820 ( .a(n4608_1), .b(n4340), .o(n4609) );
no02f01 g00821 ( .a(n4609), .b(n4602), .o(n4610) );
no02f01 g00822 ( .a(n3821_1), .b(n3990_1), .o(n4611) );
no02f01 g00823 ( .a(n3978), .b(n4356), .o(n4612) );
no03f01 g00824 ( .a(n4612), .b(n4611), .c(n3989), .o(n4613_1) );
no02f01 g00825 ( .a(n3821_1), .b(n3991), .o(n4614) );
no02f01 g00826 ( .a(n4614), .b(n3979), .o(n4615) );
no02f01 g00827 ( .a(n4615), .b(n4613_1), .o(n4616) );
na02f01 g00828 ( .a(n4615), .b(n4613_1), .o(n4617) );
in01f01 g00829 ( .a(n4617), .o(n4618_1) );
no02f01 g00830 ( .a(n4618_1), .b(n4616), .o(n4619) );
in01f01 g00831 ( .a(n4619), .o(n4620) );
no02f01 g00832 ( .a(n4620), .b(n4340), .o(n4621) );
no02f01 g00833 ( .a(n4611), .b(n3978), .o(n4622) );
in01f01 g00834 ( .a(n4622), .o(n4623_1) );
no03f01 g00835 ( .a(n4623_1), .b(n3989), .c(n3977), .o(n4624) );
no02f01 g00836 ( .a(n3989), .b(n3977), .o(n4625) );
no02f01 g00837 ( .a(n4622), .b(n4625), .o(n4626) );
no02f01 g00838 ( .a(n4626), .b(n4624), .o(n4627) );
in01f01 g00839 ( .a(n4627), .o(n4628_1) );
no02f01 g00840 ( .a(n4628_1), .b(n4340), .o(n4629) );
no02f01 g00841 ( .a(n4629), .b(n4621), .o(n4630) );
na04f01 g00842 ( .a(n4630), .b(n4610), .c(n4587), .d(n4369_1), .o(n4631) );
ao12f01 g00843 ( .a(n4344_1), .b(n4627), .c(n4619), .o(n4632) );
ao12f01 g00844 ( .a(n4344_1), .b(n4607), .c(n4600), .o(n4633_1) );
no02f01 g00845 ( .a(n4633_1), .b(n4632), .o(n4634) );
in01f01 g00846 ( .a(n4634), .o(n4635) );
ao12f01 g00847 ( .a(n4344_1), .b(n4366), .c(n4354_1), .o(n4636) );
no02f01 g00848 ( .a(n4636), .b(n4635), .o(n4637) );
no02f01 g00849 ( .a(n4001), .b(n3985_1), .o(n4638_1) );
ao12f01 g00850 ( .a(n4638_1), .b(n3998), .c(n3984), .o(n4639) );
na03f01 g00851 ( .a(n4638_1), .b(n3998), .c(n3984), .o(n4640) );
in01f01 g00852 ( .a(n4640), .o(n4641) );
no02f01 g00853 ( .a(n4641), .b(n4639), .o(n4642) );
no02f01 g00854 ( .a(n4642), .b(n4344_1), .o(n4643_1) );
in01f01 g00855 ( .a(n4643_1), .o(n4644) );
na03f01 g00856 ( .a(n4644), .b(n4637), .c(n4631), .o(n4645) );
in01f01 g00857 ( .a(n4642), .o(n4646) );
no02f01 g00858 ( .a(n4646), .b(n4340), .o(n4647) );
in01f01 g00859 ( .a(n4647), .o(n4648_1) );
ao12f01 g00860 ( .a(n4347), .b(n4648_1), .c(n4645), .o(n4649) );
in01f01 g00861 ( .a(n4389_1), .o(n4650) );
in01f01 g00862 ( .a(n4398), .o(n4651) );
in01f01 g00863 ( .a(n4420), .o(n4652_1) );
in01f01 g00864 ( .a(n4441), .o(n4653) );
na03f01 g00865 ( .a(n4440), .b(n4435), .c(n4432), .o(n4654) );
oa12f01 g00866 ( .a(n4313), .b(n4455), .c(n4451), .o(n4655) );
na03f01 g00867 ( .a(n4459), .b(n4302), .c(n4293), .o(n4656) );
na02f01 g00868 ( .a(n4656), .b(n4655), .o(n4657_1) );
in01f01 g00869 ( .a(n4478_1), .o(n4658) );
na02f01 g00870 ( .a(n4658), .b(n4657_1), .o(n4659) );
na02f01 g00871 ( .a(n4301), .b(n4293), .o(n4660) );
na02f01 g00872 ( .a(n4454), .b(n4451), .o(n4661) );
ao22f01 g00873 ( .a(n4661), .b(n4660), .c(n4492), .d(n4484), .o(n4662_1) );
oa22f01 g00874 ( .a(n4662_1), .b(n4493_1), .c(n4658), .d(n4657_1), .o(n4663) );
ao12f01 g00875 ( .a(n4322), .b(n4460), .c(n4456), .o(n4664) );
no03f01 g00876 ( .a(n4448_1), .b(n4314), .c(n4303), .o(n4665) );
in01f01 g00877 ( .a(n4466), .o(n4666) );
no03f01 g00878 ( .a(n4666), .b(n4665), .c(n4664), .o(n4667_1) );
ao12f01 g00879 ( .a(n4667_1), .b(n4663), .c(n4659), .o(n4668) );
oa12f01 g00880 ( .a(n4654), .b(n4668), .c(n4467), .o(n4669) );
no02f01 g00881 ( .a(n4325_1), .b(n4373), .o(n4670) );
no02f01 g00882 ( .a(n4324), .b(n4274), .o(n4671) );
in01f01 g00883 ( .a(n4428), .o(n4672_1) );
no03f01 g00884 ( .a(n4672_1), .b(n4671), .c(n4670), .o(n4673) );
ao12f01 g00885 ( .a(n4673), .b(n4669), .c(n4653), .o(n4674) );
na03f01 g00886 ( .a(n4419_1), .b(n4414_1), .c(n4413), .o(n4675) );
oa12f01 g00887 ( .a(n4675), .b(n4674), .c(n4429_1), .o(n4676) );
no02f01 g00888 ( .a(n4411), .b(n4410), .o(n4677_1) );
ao12f01 g00889 ( .a(n4677_1), .b(n4676), .c(n4652_1), .o(n4678) );
in01f01 g00890 ( .a(n4515), .o(n4679) );
oa12f01 g00891 ( .a(n4679), .b(n4678), .c(n4407), .o(n4680) );
in01f01 g00892 ( .a(n4517), .o(n4681) );
na03f01 g00893 ( .a(n4681), .b(n4680), .c(n4651), .o(n4682_1) );
in01f01 g00894 ( .a(n4534), .o(n4683) );
ao12f01 g00895 ( .a(n4683), .b(n4682_1), .c(n4650), .o(n4684) );
in01f01 g00896 ( .a(n4538_1), .o(n4685) );
in01f01 g00897 ( .a(n4582), .o(n4686) );
no04f01 g00898 ( .a(n4686), .b(n4547), .c(n4685), .d(n4684), .o(n4687_1) );
in01f01 g00899 ( .a(n4586), .o(n4688) );
no02f01 g00900 ( .a(n4688), .b(n4687_1), .o(n4689) );
in01f01 g00901 ( .a(n4610), .o(n4690) );
in01f01 g00902 ( .a(n4630), .o(n4691) );
no04f01 g00903 ( .a(n4691), .b(n4690), .c(n4689), .d(n4368), .o(n4692_1) );
in01f01 g00904 ( .a(n4637), .o(n4693) );
no03f01 g00905 ( .a(n4643_1), .b(n4693), .c(n4692_1), .o(n4694) );
no03f01 g00906 ( .a(n4647), .b(n4694), .c(n4346), .o(n4695) );
no02f01 g00907 ( .a(n4695), .b(n4649), .o(n4696) );
ao12f01 g00908 ( .a(n4690), .b(n4586), .c(n4583_1), .o(n4697_1) );
no02f01 g00909 ( .a(n4647), .b(n4341), .o(n4698) );
na04f01 g00910 ( .a(n4698), .b(n4630), .c(n4697_1), .d(n4369_1), .o(n4699) );
ao12f01 g00911 ( .a(n4344_1), .b(n4642), .c(n4343), .o(n4700) );
no02f01 g00912 ( .a(n4700), .b(n4693), .o(n4701) );
na02f01 g00913 ( .a(n4701), .b(n4699), .o(n4702_1) );
in01f01 g00914 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_24_), .o(n4703) );
no02f01 g00915 ( .a(n3821_1), .b(n4703), .o(n4704) );
no02f01 g00916 ( .a(n3818), .b(delay_add_ln22_unr20_stage8_stallmux_q_24_), .o(n4705) );
no02f01 g00917 ( .a(n4705), .b(n4704), .o(n4706) );
no03f01 g00918 ( .a(n3985_1), .b(n3984), .c(n3819), .o(n4707_1) );
ao12f01 g00919 ( .a(n3821_1), .b(n4000), .c(n3820), .o(n4708) );
no02f01 g00920 ( .a(n4708), .b(n3999_1), .o(n4709) );
in01f01 g00921 ( .a(n4709), .o(n4710) );
no02f01 g00922 ( .a(n4710), .b(n4707_1), .o(n4711) );
na02f01 g00923 ( .a(n4711), .b(n4706), .o(n4712_1) );
no02f01 g00924 ( .a(n4711), .b(n4706), .o(n4713) );
in01f01 g00925 ( .a(n4713), .o(n4714) );
na02f01 g00926 ( .a(n4714), .b(n4712_1), .o(n4715) );
no02f01 g00927 ( .a(n4715), .b(n4340), .o(n4716) );
in01f01 g00928 ( .a(n4712_1), .o(n4717_1) );
no02f01 g00929 ( .a(n4713), .b(n4717_1), .o(n4718) );
no02f01 g00930 ( .a(n4718), .b(n4344_1), .o(n4719) );
no02f01 g00931 ( .a(n4719), .b(n4716), .o(n4720) );
in01f01 g00932 ( .a(n4720), .o(n4721) );
no02f01 g00933 ( .a(n4721), .b(n4702_1), .o(n4722_1) );
oa12f01 g00934 ( .a(n4610), .b(n4688), .c(n4687_1), .o(n4723) );
in01f01 g00935 ( .a(n4698), .o(n4724) );
no04f01 g00936 ( .a(n4724), .b(n4691), .c(n4723), .d(n4368), .o(n4725) );
in01f01 g00937 ( .a(n4701), .o(n4726) );
no02f01 g00938 ( .a(n4726), .b(n4725), .o(n4727_1) );
no02f01 g00939 ( .a(n4720), .b(n4727_1), .o(n4728) );
no02f01 g00940 ( .a(n4728), .b(n4722_1), .o(n4729) );
ao12f01 g00941 ( .a(n3789), .b(n4729), .c(n4696), .o(n4730) );
no02f01 g00942 ( .a(n3818), .b(delay_add_ln22_unr20_stage8_stallmux_q_25_), .o(n4731) );
in01f01 g00943 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_25_), .o(n4732_1) );
no02f01 g00944 ( .a(n3821_1), .b(n4732_1), .o(n4733) );
no02f01 g00945 ( .a(n4733), .b(n4731), .o(n4734) );
in01f01 g00946 ( .a(n4734), .o(n4735) );
in01f01 g00947 ( .a(n4705), .o(n4736_1) );
na02f01 g00948 ( .a(n4707_1), .b(n4736_1), .o(n4737) );
no02f01 g00949 ( .a(n4710), .b(n4704), .o(n4738) );
na02f01 g00950 ( .a(n4738), .b(n4737), .o(n4739) );
no02f01 g00951 ( .a(n4739), .b(n4735), .o(n4740) );
in01f01 g00952 ( .a(n4740), .o(n4741_1) );
na02f01 g00953 ( .a(n4739), .b(n4735), .o(n4742) );
na02f01 g00954 ( .a(n4742), .b(n4741_1), .o(n4743) );
no02f01 g00955 ( .a(n4743), .b(n4340), .o(n4744) );
in01f01 g00956 ( .a(n4742), .o(n4745) );
no02f01 g00957 ( .a(n4745), .b(n4740), .o(n4746_1) );
no02f01 g00958 ( .a(n4746_1), .b(n4344_1), .o(n4747) );
no02f01 g00959 ( .a(n4747), .b(n4744), .o(n4748) );
in01f01 g00960 ( .a(n4748), .o(n4749) );
ao12f01 g00961 ( .a(n4716), .b(n4701), .c(n4699), .o(n4750) );
no03f01 g00962 ( .a(n4750), .b(n4749), .c(n4719), .o(n4751_1) );
in01f01 g00963 ( .a(n4751_1), .o(n4752) );
oa12f01 g00964 ( .a(n4749), .b(n4750), .c(n4719), .o(n4753) );
ao12f01 g00965 ( .a(n3789), .b(n4753), .c(n4752), .o(n4754) );
no02f01 g00966 ( .a(n4754), .b(n4730), .o(n4755) );
ao12f01 g00967 ( .a(n4340), .b(n4743), .c(n4715), .o(n4756_1) );
ao12f01 g00968 ( .a(n4344_1), .b(n4746_1), .c(n4718), .o(n4757) );
no02f01 g00969 ( .a(n4757), .b(n4726), .o(n4758) );
oa12f01 g00970 ( .a(n4758), .b(n4756_1), .c(n4699), .o(n4759) );
in01f01 g00971 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_26_), .o(n4760) );
no02f01 g00972 ( .a(n3821_1), .b(n4760), .o(n4761_1) );
no02f01 g00973 ( .a(n3818), .b(delay_add_ln22_unr20_stage8_stallmux_q_26_), .o(n4762) );
no02f01 g00974 ( .a(n4762), .b(n4761_1), .o(n4763) );
in01f01 g00975 ( .a(n4763), .o(n4764) );
no02f01 g00976 ( .a(n4737), .b(n4731), .o(n4765) );
ao12f01 g00977 ( .a(n3821_1), .b(n4732_1), .c(n4703), .o(n4766_1) );
no02f01 g00978 ( .a(n4766_1), .b(n4710), .o(n4767) );
in01f01 g00979 ( .a(n4767), .o(n4768) );
no02f01 g00980 ( .a(n4768), .b(n4765), .o(n4769) );
in01f01 g00981 ( .a(n4769), .o(n4770) );
no02f01 g00982 ( .a(n4770), .b(n4764), .o(n4771_1) );
no02f01 g00983 ( .a(n4769), .b(n4763), .o(n4772) );
no02f01 g00984 ( .a(n4772), .b(n4771_1), .o(n4773) );
in01f01 g00985 ( .a(n4773), .o(n4774) );
no02f01 g00986 ( .a(n4774), .b(n4340), .o(n4775) );
no02f01 g00987 ( .a(n4773), .b(n4344_1), .o(n4776_1) );
no02f01 g00988 ( .a(n4776_1), .b(n4775), .o(n4777) );
in01f01 g00989 ( .a(n4777), .o(n4778) );
na02f01 g00990 ( .a(n4778), .b(n4759), .o(n4779) );
no02f01 g00991 ( .a(n4778), .b(n4759), .o(n4780) );
in01f01 g00992 ( .a(n4780), .o(n4781_1) );
na02f01 g00993 ( .a(n4781_1), .b(n4779), .o(n4782) );
na02f01 g00994 ( .a(n4782), .b(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n4783) );
in01f01 g00995 ( .a(n4779), .o(n4784) );
no02f01 g00996 ( .a(n4780), .b(n4784), .o(n4785) );
no02f01 g00997 ( .a(n4785), .b(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n4786_1) );
ao12f01 g00998 ( .a(n4786_1), .b(n4783), .c(n4755), .o(n4787) );
in01f01 g00999 ( .a(n4761_1), .o(n4788) );
na02f01 g01000 ( .a(n4769), .b(n4788), .o(n4789) );
in01f01 g01001 ( .a(n4762), .o(n4790) );
na02f01 g01002 ( .a(n4789), .b(n4790), .o(n4791_1) );
no02f01 g01003 ( .a(n3818), .b(delay_add_ln22_unr20_stage8_stallmux_q_27_), .o(n4792) );
in01f01 g01004 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_27_), .o(n4793) );
no02f01 g01005 ( .a(n3821_1), .b(n4793), .o(n4794) );
no02f01 g01006 ( .a(n4794), .b(n4792), .o(n4795) );
no02f01 g01007 ( .a(n4795), .b(n4762), .o(n4796_1) );
ao22f01 g01008 ( .a(n4796_1), .b(n4789), .c(n4795), .d(n4791_1), .o(n4797) );
in01f01 g01009 ( .a(n4797), .o(n4798) );
no02f01 g01010 ( .a(n4798), .b(n4340), .o(n4799) );
no02f01 g01011 ( .a(n4797), .b(n4344_1), .o(n4800) );
no02f01 g01012 ( .a(n4800), .b(n4799), .o(n4801_1) );
in01f01 g01013 ( .a(n4775), .o(n4802) );
oa12f01 g01014 ( .a(n4802), .b(n4776_1), .c(n4759), .o(n4803) );
no02f01 g01015 ( .a(n4803), .b(n4801_1), .o(n4804) );
na02f01 g01016 ( .a(n4803), .b(n4801_1), .o(n4805) );
in01f01 g01017 ( .a(n4805), .o(n4806_1) );
no02f01 g01018 ( .a(n4806_1), .b(n4804), .o(n4807) );
no02f01 g01019 ( .a(n4807), .b(n3789), .o(n4808) );
no02f01 g01020 ( .a(n4807), .b(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n4809) );
no02f01 g01021 ( .a(n4809), .b(n4808), .o(n4810_1) );
no02f01 g01022 ( .a(n4810_1), .b(n4787), .o(n4811) );
in01f01 g01023 ( .a(n4787), .o(n4812) );
in01f01 g01024 ( .a(n4804), .o(n4813) );
na02f01 g01025 ( .a(n4805), .b(n4813), .o(n4814) );
na02f01 g01026 ( .a(n4814), .b(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n4815_1) );
na02f01 g01027 ( .a(n4814), .b(n3789), .o(n4816) );
na02f01 g01028 ( .a(n4816), .b(n4815_1), .o(n4817) );
no02f01 g01029 ( .a(n4817), .b(n4812), .o(n4818) );
in01f01 g01030 ( .a(n4639), .o(n4819) );
ao12f01 g01031 ( .a(n4249), .b(n4640), .c(n4819), .o(n4820_1) );
no03f01 g01032 ( .a(n4820_1), .b(n4342), .c(n4004_1), .o(n4821) );
no02f01 g01033 ( .a(n4821), .b(n4249), .o(n4822) );
no02f01 g01034 ( .a(n4718), .b(n4249), .o(n4823) );
no02f01 g01035 ( .a(n4823), .b(n4822), .o(n4824) );
oa12f01 g01036 ( .a(n4824), .b(n4746_1), .c(n4249), .o(n4825_1) );
na02f01 g01037 ( .a(n4825_1), .b(n4773), .o(n4826) );
oa12f01 g01038 ( .a(delay_sub_ln23_0_unr21_stage8_stallmux_q), .b(n4641), .c(n4639), .o(n4827) );
na03f01 g01039 ( .a(n4827), .b(n4006), .c(n4005), .o(n4828) );
na02f01 g01040 ( .a(n4828), .b(delay_sub_ln23_0_unr21_stage8_stallmux_q), .o(n4829_1) );
na02f01 g01041 ( .a(n4715), .b(delay_sub_ln23_0_unr21_stage8_stallmux_q), .o(n4830) );
na02f01 g01042 ( .a(n4830), .b(n4829_1), .o(n4831) );
ao12f01 g01043 ( .a(n4831), .b(n4743), .c(delay_sub_ln23_0_unr21_stage8_stallmux_q), .o(n4832) );
na02f01 g01044 ( .a(n4832), .b(n4774), .o(n4833) );
in01f01 g01045 ( .a(n4132), .o(n4834_1) );
no03f01 g01046 ( .a(n4834_1), .b(n4129), .c(n4092), .o(n4835) );
in01f01 g01047 ( .a(n4129), .o(n4836) );
ao12f01 g01048 ( .a(n4836), .b(n4132), .c(n4093_1), .o(n4837) );
no02f01 g01049 ( .a(n4837), .b(n4835), .o(n4838) );
in01f01 g01050 ( .a(n4838), .o(n4839_1) );
ao12f01 g01051 ( .a(n4839_1), .b(n4833), .c(n4826), .o(n4840) );
no02f01 g01052 ( .a(n4832), .b(n4774), .o(n4841) );
no02f01 g01053 ( .a(n4825_1), .b(n4773), .o(n4842) );
no03f01 g01054 ( .a(n4838), .b(n4842), .c(n4841), .o(n4843_1) );
no02f01 g01055 ( .a(n4843_1), .b(n4840), .o(n4844) );
ao12f01 g01056 ( .a(n4743), .b(n4830), .c(n4829_1), .o(n4845) );
no03f01 g01057 ( .a(n4823), .b(n4822), .c(n4746_1), .o(n4846) );
in01f01 g01058 ( .a(n4127), .o(n4847) );
no03f01 g01059 ( .a(n4128), .b(n4847), .c(n4101), .o(n4848_1) );
no02f01 g01060 ( .a(n4128), .b(n4101), .o(n4849) );
no02f01 g01061 ( .a(n4849), .b(n4127), .o(n4850) );
no02f01 g01062 ( .a(n4850), .b(n4848_1), .o(n4851) );
no03f01 g01063 ( .a(n4851), .b(n4846), .c(n4845), .o(n4852) );
oa12f01 g01064 ( .a(n4715), .b(n4821), .c(n4249), .o(n4853_1) );
na03f01 g01065 ( .a(n4828), .b(n4718), .c(delay_sub_ln23_0_unr21_stage8_stallmux_q), .o(n4854) );
in01f01 g01066 ( .a(n4126_1), .o(n4855) );
in01f01 g01067 ( .a(n4114), .o(n4856) );
no02f01 g01068 ( .a(n4856), .b(n4113), .o(n4857) );
no02f01 g01069 ( .a(n4857), .b(n4855), .o(n4858_1) );
na02f01 g01070 ( .a(n4857), .b(n4855), .o(n4859) );
in01f01 g01071 ( .a(n4859), .o(n4860) );
no02f01 g01072 ( .a(n4860), .b(n4858_1), .o(n4861) );
in01f01 g01073 ( .a(n4861), .o(n4862) );
na03f01 g01074 ( .a(n4862), .b(n4854), .c(n4853_1), .o(n4863_1) );
ao12f01 g01075 ( .a(n4862), .b(n4854), .c(n4853_1), .o(n4864) );
in01f01 g01076 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_0_), .o(n4865) );
no02f01 g01077 ( .a(n4119), .b(n4865), .o(n4866) );
no02f01 g01078 ( .a(n4118), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_0_), .o(n4867) );
no02f01 g01079 ( .a(n4867), .b(n4866), .o(n4868_1) );
no02f01 g01080 ( .a(n4868_1), .b(n4642), .o(n4869) );
in01f01 g01081 ( .a(n4120), .o(n4870) );
no02f01 g01082 ( .a(n4125), .b(n4115), .o(n4871) );
na02f01 g01083 ( .a(n4125), .b(n4115), .o(n4872) );
in01f01 g01084 ( .a(n4872), .o(n4873_1) );
no03f01 g01085 ( .a(n4873_1), .b(n4871), .c(n4870), .o(n4874) );
in01f01 g01086 ( .a(n4871), .o(n4875) );
ao12f01 g01087 ( .a(n4120), .b(n4872), .c(n4875), .o(n4876) );
no02f01 g01088 ( .a(n4876), .b(n4874), .o(n4877) );
no02f01 g01089 ( .a(n4877), .b(n4869), .o(n4878_1) );
no02f01 g01090 ( .a(n4827), .b(n4007), .o(n4879) );
no02f01 g01091 ( .a(n4820_1), .b(n4343), .o(n4880) );
no02f01 g01092 ( .a(n4880), .b(n4879), .o(n4881) );
na02f01 g01093 ( .a(n4877), .b(n4869), .o(n4882) );
ao12f01 g01094 ( .a(n4878_1), .b(n4882), .c(n4881), .o(n4883_1) );
oa12f01 g01095 ( .a(n4863_1), .b(n4883_1), .c(n4864), .o(n4884) );
oa12f01 g01096 ( .a(n4851), .b(n4846), .c(n4845), .o(n4885) );
ao12f01 g01097 ( .a(n4852), .b(n4885), .c(n4884), .o(n4886) );
no02f01 g01098 ( .a(n4886), .b(n4844), .o(n4887) );
na02f01 g01099 ( .a(n4886), .b(n4844), .o(n4888_1) );
in01f01 g01100 ( .a(n4888_1), .o(n4889) );
no02f01 g01101 ( .a(n4889), .b(n4887), .o(n4890) );
no03f01 g01102 ( .a(n4890), .b(n4818), .c(n4811), .o(n4891) );
na02f01 g01103 ( .a(n4817), .b(n4812), .o(n4892) );
na02f01 g01104 ( .a(n4810_1), .b(n4787), .o(n4893_1) );
in01f01 g01105 ( .a(n4890), .o(n4894) );
ao12f01 g01106 ( .a(n4894), .b(n4893_1), .c(n4892), .o(n4895) );
na02f01 g01107 ( .a(n4782), .b(n3789), .o(n4896) );
na02f01 g01108 ( .a(n4896), .b(n4783), .o(n4897_1) );
na02f01 g01109 ( .a(n4897_1), .b(n4755), .o(n4898) );
in01f01 g01110 ( .a(n4755), .o(n4899) );
no02f01 g01111 ( .a(n4785), .b(n3789), .o(n4900) );
no02f01 g01112 ( .a(n4786_1), .b(n4900), .o(n4901) );
na02f01 g01113 ( .a(n4901), .b(n4899), .o(n4902_1) );
ao12f01 g01114 ( .a(n4718), .b(n4828), .c(delay_sub_ln23_0_unr21_stage8_stallmux_q), .o(n4903) );
no03f01 g01115 ( .a(n4821), .b(n4715), .c(n4249), .o(n4904) );
no03f01 g01116 ( .a(n4861), .b(n4904), .c(n4903), .o(n4905) );
oa12f01 g01117 ( .a(n4861), .b(n4904), .c(n4903), .o(n4906) );
in01f01 g01118 ( .a(n4878_1), .o(n4907_1) );
na02f01 g01119 ( .a(n4820_1), .b(n4343), .o(n4908) );
na02f01 g01120 ( .a(n4827), .b(n4007), .o(n4909) );
na02f01 g01121 ( .a(n4909), .b(n4908), .o(n4910) );
in01f01 g01122 ( .a(n4882), .o(n4911) );
oa12f01 g01123 ( .a(n4907_1), .b(n4911), .c(n4910), .o(n4912_1) );
ao12f01 g01124 ( .a(n4905), .b(n4912_1), .c(n4906), .o(n4913) );
oa12f01 g01125 ( .a(n4746_1), .b(n4823), .c(n4822), .o(n4914) );
na03f01 g01126 ( .a(n4830), .b(n4829_1), .c(n4743), .o(n4915) );
in01f01 g01127 ( .a(n4851), .o(n4916) );
ao12f01 g01128 ( .a(n4916), .b(n4915), .c(n4914), .o(n4917_1) );
no02f01 g01129 ( .a(n4917_1), .b(n4852), .o(n4918) );
no02f01 g01130 ( .a(n4918), .b(n4913), .o(n4919) );
na02f01 g01131 ( .a(n4918), .b(n4913), .o(n4920) );
in01f01 g01132 ( .a(n4920), .o(n4921) );
no02f01 g01133 ( .a(n4921), .b(n4919), .o(n4922_1) );
in01f01 g01134 ( .a(n4922_1), .o(n4923) );
na03f01 g01135 ( .a(n4923), .b(n4902_1), .c(n4898), .o(n4924) );
oa12f01 g01136 ( .a(n4346), .b(n4647), .c(n4694), .o(n4925) );
na03f01 g01137 ( .a(n4648_1), .b(n4645), .c(n4347), .o(n4926) );
na02f01 g01138 ( .a(n4926), .b(n4925), .o(n4927_1) );
na02f01 g01139 ( .a(n4720), .b(n4727_1), .o(n4928) );
na02f01 g01140 ( .a(n4721), .b(n4702_1), .o(n4929) );
na02f01 g01141 ( .a(n4929), .b(n4928), .o(n4930) );
oa12f01 g01142 ( .a(delay_sub_ln23_0_unr22_stage8_stallmux_q), .b(n4930), .c(n4927_1), .o(n4931) );
ao12f01 g01143 ( .a(delay_sub_ln23_0_unr22_stage8_stallmux_q), .b(n4753), .c(n4752), .o(n4932_1) );
no03f01 g01144 ( .a(n4932_1), .b(n4754), .c(n4931), .o(n4933) );
in01f01 g01145 ( .a(n4719), .o(n4934) );
in01f01 g01146 ( .a(n4716), .o(n4935) );
oa12f01 g01147 ( .a(n4935), .b(n4726), .c(n4725), .o(n4936) );
ao12f01 g01148 ( .a(n4748), .b(n4936), .c(n4934), .o(n4937_1) );
oa12f01 g01149 ( .a(delay_sub_ln23_0_unr22_stage8_stallmux_q), .b(n4937_1), .c(n4751_1), .o(n4938) );
oa12f01 g01150 ( .a(n3789), .b(n4937_1), .c(n4751_1), .o(n4939) );
ao12f01 g01151 ( .a(n4730), .b(n4939), .c(n4938), .o(n4940) );
no02f01 g01152 ( .a(n4864), .b(n4905), .o(n4941) );
no02f01 g01153 ( .a(n4941), .b(n4883_1), .o(n4942_1) );
na02f01 g01154 ( .a(n4941), .b(n4883_1), .o(n4943) );
in01f01 g01155 ( .a(n4943), .o(n4944) );
no02f01 g01156 ( .a(n4944), .b(n4942_1), .o(n4945) );
no03f01 g01157 ( .a(n4945), .b(n4940), .c(n4933), .o(n4946) );
oa12f01 g01158 ( .a(n4945), .b(n4940), .c(n4933), .o(n4947_1) );
na03f01 g01159 ( .a(n4729), .b(n4927_1), .c(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n4948) );
oa12f01 g01160 ( .a(n4930), .b(n4696), .c(n3789), .o(n4949) );
in01f01 g01161 ( .a(n4877), .o(n4950) );
no02f01 g01162 ( .a(n4881), .b(n4950), .o(n4951) );
no02f01 g01163 ( .a(n4910), .b(n4877), .o(n4952_1) );
no02f01 g01164 ( .a(n4952_1), .b(n4951), .o(n4953) );
no02f01 g01165 ( .a(n4953), .b(n4869), .o(n4954) );
na02f01 g01166 ( .a(n4953), .b(n4869), .o(n4955) );
in01f01 g01167 ( .a(n4955), .o(n4956) );
no02f01 g01168 ( .a(n4956), .b(n4954), .o(n4957_1) );
in01f01 g01169 ( .a(n4957_1), .o(n4958) );
ao12f01 g01170 ( .a(n4958), .b(n4949), .c(n4948), .o(n4959) );
no02f01 g01171 ( .a(n4927_1), .b(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n4960) );
no02f01 g01172 ( .a(n4927_1), .b(n3789), .o(n4961) );
in01f01 g01173 ( .a(n4868_1), .o(n4962_1) );
no02f01 g01174 ( .a(n4962_1), .b(n4642), .o(n4963) );
no02f01 g01175 ( .a(n4868_1), .b(n4646), .o(n4964) );
no02f01 g01176 ( .a(n4964), .b(n4963), .o(n4965) );
no03f01 g01177 ( .a(n4965), .b(n4961), .c(n4960), .o(n4966) );
na03f01 g01178 ( .a(n4958), .b(n4949), .c(n4948), .o(n4967_1) );
oa12f01 g01179 ( .a(n4967_1), .b(n4966), .c(n4959), .o(n4968) );
ao12f01 g01180 ( .a(n4946), .b(n4968), .c(n4947_1), .o(n4969) );
ao12f01 g01181 ( .a(n4923), .b(n4902_1), .c(n4898), .o(n4970) );
oa12f01 g01182 ( .a(n4924), .b(n4970), .c(n4969), .o(n4971) );
oa12f01 g01183 ( .a(n4971), .b(n4895), .c(n4891), .o(n4972_1) );
na03f01 g01184 ( .a(n4894), .b(n4893_1), .c(n4892), .o(n4973) );
oa12f01 g01185 ( .a(n4890), .b(n4818), .c(n4811), .o(n4974) );
no02f01 g01186 ( .a(n4901), .b(n4899), .o(n4975) );
no02f01 g01187 ( .a(n4897_1), .b(n4755), .o(n4976) );
no03f01 g01188 ( .a(n4922_1), .b(n4976), .c(n4975), .o(n4977_1) );
na03f01 g01189 ( .a(n4939), .b(n4938), .c(n4730), .o(n4978) );
oa12f01 g01190 ( .a(n4931), .b(n4932_1), .c(n4754), .o(n4979) );
in01f01 g01191 ( .a(n4945), .o(n4980) );
na03f01 g01192 ( .a(n4980), .b(n4979), .c(n4978), .o(n4981) );
ao12f01 g01193 ( .a(n4980), .b(n4979), .c(n4978), .o(n4982_1) );
no03f01 g01194 ( .a(n4930), .b(n4696), .c(n3789), .o(n4983) );
ao12f01 g01195 ( .a(n4729), .b(n4927_1), .c(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n4984) );
oa12f01 g01196 ( .a(n4957_1), .b(n4984), .c(n4983), .o(n4985) );
na02f01 g01197 ( .a(n4696), .b(n3789), .o(n4986) );
na02f01 g01198 ( .a(n4696), .b(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n4987_1) );
in01f01 g01199 ( .a(n4965), .o(n4988) );
na03f01 g01200 ( .a(n4988), .b(n4987_1), .c(n4986), .o(n4989) );
no03f01 g01201 ( .a(n4957_1), .b(n4984), .c(n4983), .o(n4990) );
ao12f01 g01202 ( .a(n4990), .b(n4989), .c(n4985), .o(n4991) );
oa12f01 g01203 ( .a(n4981), .b(n4991), .c(n4982_1), .o(n4992_1) );
oa12f01 g01204 ( .a(n4922_1), .b(n4976), .c(n4975), .o(n4993) );
ao12f01 g01205 ( .a(n4977_1), .b(n4993), .c(n4992_1), .o(n4994) );
na03f01 g01206 ( .a(n4994), .b(n4974), .c(n4973), .o(n4995) );
na02f01 g01207 ( .a(n4995), .b(n4972_1), .o(n198) );
in01f01 g01208 ( .a(n_45224), .o(n4997_1) );
no02f01 g01209 ( .a(n4997_1), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_22_), .o(n4998) );
no02f01 g01210 ( .a(n4997_1), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_21_), .o(n4999) );
no02f01 g01211 ( .a(n4999), .b(n4998), .o(n5000) );
in01f01 g01212 ( .a(n5000), .o(n5001_1) );
in01f01 g01213 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_21_), .o(n5002) );
in01f01 g01214 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_22_), .o(n5003) );
ao12f01 g01215 ( .a(n_45224), .b(n5003), .c(n5002), .o(n5004) );
no02f01 g01216 ( .a(n4997_1), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_20_), .o(n5005) );
na02f01 g01217 ( .a(n4997_1), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_20_), .o(n5006_1) );
in01f01 g01218 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_19_), .o(n5007) );
no02f01 g01219 ( .a(n5007), .b(delay_sub_ln23_unr9_stage4_stallmux_q_3_), .o(n5008) );
in01f01 g01220 ( .a(n5008), .o(n5009) );
ao12f01 g01221 ( .a(n5005), .b(n5009), .c(n5006_1), .o(n5010) );
oa12f01 g01222 ( .a(n5000), .b(n5010), .c(n5004), .o(n5011_1) );
in01f01 g01223 ( .a(delay_sub_ln23_unr9_stage4_stallmux_q_3_), .o(n5012) );
ao12f01 g01224 ( .a(n5012), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_15_), .c(delay_sub_ln23_0_unr8_stage4_stallmux_q_16_), .o(n5013) );
in01f01 g01225 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_14_), .o(n5014) );
in01f01 g01226 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_0_), .o(n5015) );
na02f01 g01227 ( .a(n_45224), .b(n5015), .o(n5016_1) );
no02f01 g01228 ( .a(n_45224), .b(n5015), .o(n5017) );
ao12f01 g01229 ( .a(n5017), .b(n5016_1), .c(cordic_combinational_sub_ln23_0_unr12_z_0_), .o(n5018) );
no02f01 g01230 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_2_), .b(n5012), .o(n5019) );
no02f01 g01231 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_1_), .b(n5012), .o(n5020) );
no03f01 g01232 ( .a(n5020), .b(n5019), .c(n5018), .o(n5021_1) );
in01f01 g01233 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_2_), .o(n5022) );
no02f01 g01234 ( .a(n5022), .b(delay_sub_ln23_unr9_stage4_stallmux_q_3_), .o(n5023) );
in01f01 g01235 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_1_), .o(n5024) );
no02f01 g01236 ( .a(n5024), .b(delay_sub_ln23_unr9_stage4_stallmux_q_3_), .o(n5025) );
no03f01 g01237 ( .a(n5025), .b(n5023), .c(n5021_1), .o(n5026_1) );
ao12f01 g01238 ( .a(n5012), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_3_), .c(delay_sub_ln23_0_unr8_stage4_stallmux_q_4_), .o(n5027) );
no02f01 g01239 ( .a(n5027), .b(n5026_1), .o(n5028) );
no02f01 g01240 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_5_), .b(n5012), .o(n5029) );
no02f01 g01241 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_6_), .b(n5012), .o(n5030) );
no02f01 g01242 ( .a(n5030), .b(n5029), .o(n5031_1) );
in01f01 g01243 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_4_), .o(n5032) );
in01f01 g01244 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_3_), .o(n5033) );
ao12f01 g01245 ( .a(delay_sub_ln23_unr9_stage4_stallmux_q_3_), .b(n5033), .c(n5032), .o(n5034) );
na02f01 g01246 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_5_), .b(n5012), .o(n5035) );
in01f01 g01247 ( .a(n5035), .o(n5036_1) );
na02f01 g01248 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_6_), .b(n5012), .o(n5037) );
in01f01 g01249 ( .a(n5037), .o(n5038) );
no03f01 g01250 ( .a(n5038), .b(n5036_1), .c(n5034), .o(n5039) );
in01f01 g01251 ( .a(n5039), .o(n5040) );
ao12f01 g01252 ( .a(n5040), .b(n5031_1), .c(n5028), .o(n5041_1) );
in01f01 g01253 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_7_), .o(n5042) );
na02f01 g01254 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_8_), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_9_), .o(n5043) );
oa12f01 g01255 ( .a(delay_sub_ln23_unr9_stage4_stallmux_q_3_), .b(n5043), .c(n5042), .o(n5044) );
no02f01 g01256 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_10_), .b(n5012), .o(n5045) );
in01f01 g01257 ( .a(n5045), .o(n5046_1) );
na02f01 g01258 ( .a(n5046_1), .b(n5044), .o(n5047) );
no02f01 g01259 ( .a(n5047), .b(n5041_1), .o(n5048) );
no02f01 g01260 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_11_), .b(n5012), .o(n5049) );
no02f01 g01261 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_12_), .b(n5012), .o(n5050) );
no02f01 g01262 ( .a(n5050), .b(n5049), .o(n5051_1) );
in01f01 g01263 ( .a(n5051_1), .o(n5052) );
no02f01 g01264 ( .a(n5012), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_13_), .o(n5053) );
no02f01 g01265 ( .a(n5053), .b(n5052), .o(n5054) );
na02f01 g01266 ( .a(n5054), .b(n5048), .o(n5055) );
na02f01 g01267 ( .a(n5012), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_13_), .o(n5056_1) );
na03f01 g01268 ( .a(n5056_1), .b(n5055), .c(n5014), .o(n5057) );
in01f01 g01269 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_8_), .o(n5058) );
ao12f01 g01270 ( .a(delay_sub_ln23_unr9_stage4_stallmux_q_3_), .b(n5042), .c(n5058), .o(n5059) );
in01f01 g01271 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_9_), .o(n5060) );
no02f01 g01272 ( .a(n5060), .b(delay_sub_ln23_unr9_stage4_stallmux_q_3_), .o(n5061_1) );
no02f01 g01273 ( .a(n5061_1), .b(n5059), .o(n5062) );
in01f01 g01274 ( .a(n5062), .o(n5063) );
na02f01 g01275 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_10_), .b(n5012), .o(n5064) );
in01f01 g01276 ( .a(n5064), .o(n5065) );
no02f01 g01277 ( .a(n5065), .b(n5063), .o(n5066_1) );
in01f01 g01278 ( .a(n5066_1), .o(n5067) );
in01f01 g01279 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_12_), .o(n5068) );
in01f01 g01280 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_11_), .o(n5069) );
ao12f01 g01281 ( .a(delay_sub_ln23_unr9_stage4_stallmux_q_3_), .b(n5069), .c(n5068), .o(n5070_1) );
no02f01 g01282 ( .a(n5070_1), .b(n5067), .o(n5071) );
oa12f01 g01283 ( .a(n5071), .b(n5055), .c(n5014), .o(n5072) );
ao12f01 g01284 ( .a(n5072), .b(n5057), .c(n5012), .o(n5073) );
no02f01 g01285 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_18_), .b(n5012), .o(n5074) );
no02f01 g01286 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_17_), .b(n5012), .o(n5075_1) );
no02f01 g01287 ( .a(n5075_1), .b(n5074), .o(n5076) );
in01f01 g01288 ( .a(n5076), .o(n5077) );
no03f01 g01289 ( .a(n5077), .b(n5073), .c(n5013), .o(n5078) );
in01f01 g01290 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_16_), .o(n5079) );
in01f01 g01291 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_15_), .o(n5080_1) );
ao12f01 g01292 ( .a(delay_sub_ln23_unr9_stage4_stallmux_q_3_), .b(n5080_1), .c(n5079), .o(n5081) );
in01f01 g01293 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_18_), .o(n5082) );
in01f01 g01294 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_17_), .o(n5083) );
ao12f01 g01295 ( .a(delay_sub_ln23_unr9_stage4_stallmux_q_3_), .b(n5083), .c(n5082), .o(n5084) );
no02f01 g01296 ( .a(n5084), .b(n5081), .o(n5085_1) );
in01f01 g01297 ( .a(n5085_1), .o(n5086) );
no02f01 g01298 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_19_), .b(n5012), .o(n5087) );
no02f01 g01299 ( .a(n5087), .b(n5005), .o(n5088) );
oa12f01 g01300 ( .a(n5088), .b(n5086), .c(n5078), .o(n5089) );
oa12f01 g01301 ( .a(n5011_1), .b(n5089), .c(n5001_1), .o(n5090_1) );
in01f01 g01302 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_27_), .o(n5091) );
in01f01 g01303 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_28_), .o(n5092) );
ao12f01 g01304 ( .a(n_45224), .b(n5092), .c(n5091), .o(n5093) );
no02f01 g01305 ( .a(n5093), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_29_), .o(n5094) );
no02f01 g01306 ( .a(n5094), .b(n_45224), .o(n5095_1) );
in01f01 g01307 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_23_), .o(n5096) );
in01f01 g01308 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_24_), .o(n5097) );
ao12f01 g01309 ( .a(n_45224), .b(n5097), .c(n5096), .o(n5098) );
in01f01 g01310 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_26_), .o(n5099) );
in01f01 g01311 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_25_), .o(n5100_1) );
ao12f01 g01312 ( .a(n_45224), .b(n5100_1), .c(n5099), .o(n5101) );
no02f01 g01313 ( .a(n5101), .b(n5098), .o(n5102) );
in01f01 g01314 ( .a(n5102), .o(n5103) );
no02f01 g01315 ( .a(n5103), .b(n5095_1), .o(n5104) );
in01f01 g01316 ( .a(n5104), .o(n5105_1) );
no02f01 g01317 ( .a(n4997_1), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_23_), .o(n5106) );
no02f01 g01318 ( .a(n4997_1), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_24_), .o(n5107) );
no02f01 g01319 ( .a(n5107), .b(n5106), .o(n5108) );
no02f01 g01320 ( .a(n4997_1), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_26_), .o(n5109) );
no02f01 g01321 ( .a(n4997_1), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_25_), .o(n5110_1) );
no02f01 g01322 ( .a(n5110_1), .b(n5109), .o(n5111) );
na02f01 g01323 ( .a(n5111), .b(n5108), .o(n5112) );
no02f01 g01324 ( .a(n4997_1), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_29_), .o(n5113) );
no02f01 g01325 ( .a(n4997_1), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_27_), .o(n5114) );
no02f01 g01326 ( .a(n4997_1), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_28_), .o(n5115_1) );
no02f01 g01327 ( .a(n5115_1), .b(n5114), .o(n5116) );
in01f01 g01328 ( .a(n5116), .o(n5117) );
no03f01 g01329 ( .a(n5117), .b(n5113), .c(n5112), .o(n5118) );
oa12f01 g01330 ( .a(n5118), .b(n5105_1), .c(n5090_1), .o(n5119) );
no03f01 g01331 ( .a(n5029), .b(n5027), .c(n5026_1), .o(n5120_1) );
no03f01 g01332 ( .a(n5120_1), .b(n5036_1), .c(n5034), .o(n5121) );
in01f01 g01333 ( .a(n5121), .o(n5122) );
no02f01 g01334 ( .a(n5038), .b(n5030), .o(n5123) );
in01f01 g01335 ( .a(n5123), .o(n5124) );
no02f01 g01336 ( .a(n5124), .b(n5122), .o(n5125_1) );
no02f01 g01337 ( .a(n5123), .b(n5121), .o(n5126) );
no02f01 g01338 ( .a(n5126), .b(n5125_1), .o(n5127) );
in01f01 g01339 ( .a(n5127), .o(n5128) );
no02f01 g01340 ( .a(n5128), .b(n5119), .o(n5129) );
in01f01 g01341 ( .a(n5129), .o(n5130_1) );
in01f01 g01342 ( .a(n5018), .o(n5131) );
in01f01 g01343 ( .a(n5020), .o(n5132) );
ao12f01 g01344 ( .a(n5025), .b(n5132), .c(n5131), .o(n5133) );
in01f01 g01345 ( .a(n5133), .o(n5134) );
no02f01 g01346 ( .a(n5023), .b(n5019), .o(n5135_1) );
in01f01 g01347 ( .a(n5135_1), .o(n5136) );
no02f01 g01348 ( .a(n5136), .b(n5134), .o(n5137) );
no02f01 g01349 ( .a(n5135_1), .b(n5133), .o(n5138) );
no02f01 g01350 ( .a(n5138), .b(n5137), .o(n5139) );
in01f01 g01351 ( .a(n5139), .o(n5140_1) );
no02f01 g01352 ( .a(n5140_1), .b(n5119), .o(n5141) );
in01f01 g01353 ( .a(n5119), .o(n5142) );
no02f01 g01354 ( .a(n5025), .b(n5020), .o(n5143) );
in01f01 g01355 ( .a(n5143), .o(n5144) );
no02f01 g01356 ( .a(n5144), .b(n5131), .o(n5145_1) );
no02f01 g01357 ( .a(n5143), .b(n5018), .o(n5146) );
no02f01 g01358 ( .a(n5146), .b(n5145_1), .o(n5147) );
na02f01 g01359 ( .a(n5147), .b(n5142), .o(n5148) );
in01f01 g01360 ( .a(n5016_1), .o(n5149) );
no03f01 g01361 ( .a(n5017), .b(n5149), .c(cordic_combinational_sub_ln23_0_unr12_z_0_), .o(n5150_1) );
in01f01 g01362 ( .a(cordic_combinational_sub_ln23_0_unr12_z_0_), .o(n5151) );
in01f01 g01363 ( .a(n5017), .o(n5152) );
ao12f01 g01364 ( .a(n5151), .b(n5152), .c(n5016_1), .o(n5153) );
no02f01 g01365 ( .a(n5153), .b(n5150_1), .o(n5154) );
in01f01 g01366 ( .a(n5154), .o(n5155_1) );
na02f01 g01367 ( .a(n5155_1), .b(n5119), .o(n5156) );
no02f01 g01368 ( .a(n5155_1), .b(n5119), .o(n5157) );
oa12f01 g01369 ( .a(n5156), .b(n5157), .c(cordic_combinational_sub_ln23_0_unr12_z_0_), .o(n5158) );
na02f01 g01370 ( .a(n5158), .b(n5148), .o(n5159) );
no02f01 g01371 ( .a(n5139), .b(n5142), .o(n5160_1) );
no02f01 g01372 ( .a(n5147), .b(n5142), .o(n5161) );
no02f01 g01373 ( .a(n5161), .b(n5160_1), .o(n5162) );
oa12f01 g01374 ( .a(n5162), .b(n5159), .c(n5141), .o(n5163) );
in01f01 g01375 ( .a(n5026_1), .o(n5164) );
no02f01 g01376 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_3_), .b(n5012), .o(n5165_1) );
no02f01 g01377 ( .a(n5033), .b(delay_sub_ln23_unr9_stage4_stallmux_q_3_), .o(n5166) );
no02f01 g01378 ( .a(n5166), .b(n5165_1), .o(n5167) );
in01f01 g01379 ( .a(n5167), .o(n5168) );
no02f01 g01380 ( .a(n5168), .b(n5164), .o(n5169) );
no02f01 g01381 ( .a(n5167), .b(n5026_1), .o(n5170_1) );
no02f01 g01382 ( .a(n5170_1), .b(n5169), .o(n5171) );
in01f01 g01383 ( .a(n5171), .o(n5172) );
no02f01 g01384 ( .a(n5172), .b(n5119), .o(n5173) );
in01f01 g01385 ( .a(n5173), .o(n5174) );
na02f01 g01386 ( .a(n5174), .b(n5163), .o(n5175_1) );
no02f01 g01387 ( .a(n5034), .b(n5028), .o(n5176) );
no02f01 g01388 ( .a(n5036_1), .b(n5029), .o(n5177) );
no02f01 g01389 ( .a(n5177), .b(n5176), .o(n5178) );
na02f01 g01390 ( .a(n5177), .b(n5176), .o(n5179) );
in01f01 g01391 ( .a(n5179), .o(n5180_1) );
no02f01 g01392 ( .a(n5180_1), .b(n5178), .o(n5181) );
in01f01 g01393 ( .a(n5181), .o(n5182) );
no02f01 g01394 ( .a(n5182), .b(n5119), .o(n5183) );
in01f01 g01395 ( .a(n5165_1), .o(n5184) );
ao12f01 g01396 ( .a(n5166), .b(n5184), .c(n5164), .o(n5185_1) );
in01f01 g01397 ( .a(n5185_1), .o(n5186) );
no02f01 g01398 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_4_), .b(n5012), .o(n5187) );
no02f01 g01399 ( .a(n5032), .b(delay_sub_ln23_unr9_stage4_stallmux_q_3_), .o(n5188) );
no02f01 g01400 ( .a(n5188), .b(n5187), .o(n5189) );
in01f01 g01401 ( .a(n5189), .o(n5190_1) );
no02f01 g01402 ( .a(n5190_1), .b(n5186), .o(n5191) );
no02f01 g01403 ( .a(n5189), .b(n5185_1), .o(n5192) );
no02f01 g01404 ( .a(n5192), .b(n5191), .o(n5193) );
in01f01 g01405 ( .a(n5193), .o(n5194) );
no02f01 g01406 ( .a(n5194), .b(n5119), .o(n5195_1) );
no02f01 g01407 ( .a(n5195_1), .b(n5183), .o(n5196) );
in01f01 g01408 ( .a(n5196), .o(n5197) );
no02f01 g01409 ( .a(n5197), .b(n5175_1), .o(n5198) );
no02f01 g01410 ( .a(n5193), .b(n5142), .o(n5199) );
no02f01 g01411 ( .a(n5171), .b(n5142), .o(n5200_1) );
no02f01 g01412 ( .a(n5200_1), .b(n5199), .o(n5201) );
in01f01 g01413 ( .a(n5201), .o(n5202) );
no02f01 g01414 ( .a(n5127), .b(n5142), .o(n5203) );
no02f01 g01415 ( .a(n5181), .b(n5142), .o(n5204) );
no03f01 g01416 ( .a(n5204), .b(n5203), .c(n5202), .o(n5205_1) );
in01f01 g01417 ( .a(n5205_1), .o(n5206) );
ao12f01 g01418 ( .a(n5206), .b(n5198), .c(n5130_1), .o(n5207) );
no02f01 g01419 ( .a(n5042), .b(delay_sub_ln23_unr9_stage4_stallmux_q_3_), .o(n5208) );
no02f01 g01420 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_7_), .b(n5012), .o(n5209) );
no02f01 g01421 ( .a(n5209), .b(n5041_1), .o(n5210_1) );
no02f01 g01422 ( .a(n5210_1), .b(n5208), .o(n5211) );
no02f01 g01423 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_8_), .b(n5012), .o(n5212) );
no02f01 g01424 ( .a(n5058), .b(delay_sub_ln23_unr9_stage4_stallmux_q_3_), .o(n5213) );
no02f01 g01425 ( .a(n5213), .b(n5212), .o(n5214) );
no02f01 g01426 ( .a(n5214), .b(n5211), .o(n5215_1) );
na02f01 g01427 ( .a(n5214), .b(n5211), .o(n5216) );
in01f01 g01428 ( .a(n5216), .o(n5217) );
no02f01 g01429 ( .a(n5217), .b(n5215_1), .o(n5218) );
in01f01 g01430 ( .a(n5218), .o(n5219) );
no02f01 g01431 ( .a(n5219), .b(n5119), .o(n5220_1) );
in01f01 g01432 ( .a(n5041_1), .o(n5221) );
no02f01 g01433 ( .a(n5208), .b(n5209), .o(n5222) );
in01f01 g01434 ( .a(n5222), .o(n5223) );
no02f01 g01435 ( .a(n5223), .b(n5221), .o(n5224) );
no02f01 g01436 ( .a(n5222), .b(n5041_1), .o(n5225_1) );
no02f01 g01437 ( .a(n5225_1), .b(n5224), .o(n5226) );
in01f01 g01438 ( .a(n5226), .o(n5227) );
no02f01 g01439 ( .a(n5227), .b(n5119), .o(n5228) );
no02f01 g01440 ( .a(n5228), .b(n5220_1), .o(n5229) );
in01f01 g01441 ( .a(n5229), .o(n5230_1) );
no02f01 g01442 ( .a(n5230_1), .b(n5207), .o(n5231) );
oa12f01 g01443 ( .a(delay_sub_ln23_unr9_stage4_stallmux_q_3_), .b(n5042), .c(n5058), .o(n5232) );
na02f01 g01444 ( .a(n5232), .b(n5221), .o(n5233) );
in01f01 g01445 ( .a(n5233), .o(n5234) );
no02f01 g01446 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_9_), .b(n5012), .o(n5235_1) );
no02f01 g01447 ( .a(n5235_1), .b(n5061_1), .o(n5236) );
in01f01 g01448 ( .a(n5236), .o(n5237) );
no03f01 g01449 ( .a(n5237), .b(n5234), .c(n5059), .o(n5238) );
in01f01 g01450 ( .a(n5059), .o(n5239) );
ao12f01 g01451 ( .a(n5236), .b(n5233), .c(n5239), .o(n5240_1) );
no02f01 g01452 ( .a(n5240_1), .b(n5238), .o(n5241) );
in01f01 g01453 ( .a(n5241), .o(n5242) );
no02f01 g01454 ( .a(n5242), .b(n5119), .o(n5243) );
ao12f01 g01455 ( .a(n5063), .b(n5044), .c(n5221), .o(n5244) );
no02f01 g01456 ( .a(n5065), .b(n5045), .o(n5245_1) );
no02f01 g01457 ( .a(n5245_1), .b(n5244), .o(n5246) );
na02f01 g01458 ( .a(n5245_1), .b(n5244), .o(n5247) );
in01f01 g01459 ( .a(n5247), .o(n5248) );
no02f01 g01460 ( .a(n5248), .b(n5246), .o(n5249) );
in01f01 g01461 ( .a(n5249), .o(n5250_1) );
no02f01 g01462 ( .a(n5250_1), .b(n5119), .o(n5251) );
no02f01 g01463 ( .a(n5251), .b(n5243), .o(n5252) );
na02f01 g01464 ( .a(n5252), .b(n5231), .o(n5253) );
no02f01 g01465 ( .a(n5069), .b(delay_sub_ln23_unr9_stage4_stallmux_q_3_), .o(n5254) );
no02f01 g01466 ( .a(n5254), .b(n5049), .o(n5255_1) );
in01f01 g01467 ( .a(n5255_1), .o(n5256) );
no03f01 g01468 ( .a(n5256), .b(n5067), .c(n5048), .o(n5257) );
in01f01 g01469 ( .a(n5048), .o(n5258) );
ao12f01 g01470 ( .a(n5255_1), .b(n5066_1), .c(n5258), .o(n5259) );
no02f01 g01471 ( .a(n5259), .b(n5257), .o(n5260_1) );
in01f01 g01472 ( .a(n5260_1), .o(n5261) );
no02f01 g01473 ( .a(n5261), .b(n5119), .o(n5262) );
no02f01 g01474 ( .a(n5049), .b(n5258), .o(n5263) );
no03f01 g01475 ( .a(n5263), .b(n5254), .c(n5067), .o(n5264) );
no02f01 g01476 ( .a(n5068), .b(delay_sub_ln23_unr9_stage4_stallmux_q_3_), .o(n5265_1) );
no02f01 g01477 ( .a(n5265_1), .b(n5050), .o(n5266) );
no02f01 g01478 ( .a(n5266), .b(n5264), .o(n5267) );
na02f01 g01479 ( .a(n5266), .b(n5264), .o(n5268) );
in01f01 g01480 ( .a(n5268), .o(n5269) );
no02f01 g01481 ( .a(n5269), .b(n5267), .o(n5270_1) );
in01f01 g01482 ( .a(n5270_1), .o(n5271) );
no02f01 g01483 ( .a(n5271), .b(n5119), .o(n5272) );
no02f01 g01484 ( .a(n5272), .b(n5262), .o(n5273) );
in01f01 g01485 ( .a(n5273), .o(n5274) );
no02f01 g01486 ( .a(n5274), .b(n5253), .o(n5275_1) );
na03f01 g01487 ( .a(n5071), .b(n5056_1), .c(n5055), .o(n5276) );
in01f01 g01488 ( .a(n5276), .o(n5277) );
no02f01 g01489 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_14_), .b(n5012), .o(n5278) );
no02f01 g01490 ( .a(n5014), .b(delay_sub_ln23_unr9_stage4_stallmux_q_3_), .o(n5279) );
no02f01 g01491 ( .a(n5279), .b(n5278), .o(n5280_1) );
no02f01 g01492 ( .a(n5280_1), .b(n5277), .o(n5281) );
na02f01 g01493 ( .a(n5280_1), .b(n5277), .o(n5282) );
in01f01 g01494 ( .a(n5282), .o(n5283) );
no02f01 g01495 ( .a(n5283), .b(n5281), .o(n5284) );
in01f01 g01496 ( .a(n5284), .o(n5285_1) );
no02f01 g01497 ( .a(n5285_1), .b(n5119), .o(n5286) );
in01f01 g01498 ( .a(n5071), .o(n5287) );
ao12f01 g01499 ( .a(n5287), .b(n5051_1), .c(n5048), .o(n5288) );
in01f01 g01500 ( .a(n5056_1), .o(n5289) );
no02f01 g01501 ( .a(n5289), .b(n5053), .o(n5290_1) );
no02f01 g01502 ( .a(n5290_1), .b(n5288), .o(n5291) );
na02f01 g01503 ( .a(n5290_1), .b(n5288), .o(n5292) );
in01f01 g01504 ( .a(n5292), .o(n5293) );
no02f01 g01505 ( .a(n5293), .b(n5291), .o(n5294) );
in01f01 g01506 ( .a(n5294), .o(n5295_1) );
no02f01 g01507 ( .a(n5295_1), .b(n5119), .o(n5296) );
no02f01 g01508 ( .a(n5296), .b(n5286), .o(n5297) );
na02f01 g01509 ( .a(n5297), .b(n5275_1), .o(n5298) );
no02f01 g01510 ( .a(n5218), .b(n5142), .o(n5299) );
no02f01 g01511 ( .a(n5226), .b(n5142), .o(n5300_1) );
no02f01 g01512 ( .a(n5300_1), .b(n5299), .o(n5301) );
no02f01 g01513 ( .a(n5241), .b(n5142), .o(n5302) );
no02f01 g01514 ( .a(n5249), .b(n5142), .o(n5303) );
no02f01 g01515 ( .a(n5303), .b(n5302), .o(n5304) );
no02f01 g01516 ( .a(n5260_1), .b(n5142), .o(n5305_1) );
no02f01 g01517 ( .a(n5270_1), .b(n5142), .o(n5306) );
no02f01 g01518 ( .a(n5306), .b(n5305_1), .o(n5307) );
na03f01 g01519 ( .a(n5307), .b(n5304), .c(n5301), .o(n5308) );
no02f01 g01520 ( .a(n5294), .b(n5142), .o(n5309) );
no02f01 g01521 ( .a(n5284), .b(n5142), .o(n5310_1) );
no03f01 g01522 ( .a(n5310_1), .b(n5309), .c(n5308), .o(n5311) );
na02f01 g01523 ( .a(n5311), .b(n5298), .o(n5312) );
in01f01 g01524 ( .a(n5073), .o(n5313) );
no02f01 g01525 ( .a(n5080_1), .b(delay_sub_ln23_unr9_stage4_stallmux_q_3_), .o(n5314) );
no02f01 g01526 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_15_), .b(n5012), .o(n5315_1) );
in01f01 g01527 ( .a(n5315_1), .o(n5316) );
ao12f01 g01528 ( .a(n5314), .b(n5316), .c(n5313), .o(n5317) );
in01f01 g01529 ( .a(n5317), .o(n5318) );
no02f01 g01530 ( .a(n5012), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_16_), .o(n5319) );
no02f01 g01531 ( .a(delay_sub_ln23_unr9_stage4_stallmux_q_3_), .b(n5079), .o(n5320_1) );
no02f01 g01532 ( .a(n5320_1), .b(n5319), .o(n5321) );
in01f01 g01533 ( .a(n5321), .o(n5322) );
no02f01 g01534 ( .a(n5322), .b(n5318), .o(n5323) );
no02f01 g01535 ( .a(n5321), .b(n5317), .o(n5324) );
no02f01 g01536 ( .a(n5324), .b(n5323), .o(n5325_1) );
in01f01 g01537 ( .a(n5325_1), .o(n5326) );
no02f01 g01538 ( .a(n5326), .b(n5119), .o(n5327) );
no02f01 g01539 ( .a(n5315_1), .b(n5314), .o(n5328) );
in01f01 g01540 ( .a(n5328), .o(n5329) );
no02f01 g01541 ( .a(n5329), .b(n5313), .o(n5330_1) );
no02f01 g01542 ( .a(n5328), .b(n5073), .o(n5331) );
no02f01 g01543 ( .a(n5331), .b(n5330_1), .o(n5332) );
in01f01 g01544 ( .a(n5332), .o(n5333) );
no02f01 g01545 ( .a(n5333), .b(n5119), .o(n5334) );
no02f01 g01546 ( .a(n5334), .b(n5327), .o(n5335_1) );
in01f01 g01547 ( .a(n5335_1), .o(n5336) );
no02f01 g01548 ( .a(n5083), .b(delay_sub_ln23_unr9_stage4_stallmux_q_3_), .o(n5337) );
no03f01 g01549 ( .a(n5075_1), .b(n5073), .c(n5013), .o(n5338) );
no03f01 g01550 ( .a(n5338), .b(n5337), .c(n5081), .o(n5339) );
no02f01 g01551 ( .a(n5082), .b(delay_sub_ln23_unr9_stage4_stallmux_q_3_), .o(n5340_1) );
no02f01 g01552 ( .a(n5340_1), .b(n5074), .o(n5341) );
no02f01 g01553 ( .a(n5341), .b(n5339), .o(n5342) );
na02f01 g01554 ( .a(n5341), .b(n5339), .o(n5343) );
in01f01 g01555 ( .a(n5343), .o(n5344) );
no03f01 g01556 ( .a(n5344), .b(n5342), .c(n5119), .o(n5345_1) );
no02f01 g01557 ( .a(n5073), .b(n5013), .o(n5346) );
no02f01 g01558 ( .a(n5337), .b(n5075_1), .o(n5347) );
in01f01 g01559 ( .a(n5347), .o(n5348) );
no03f01 g01560 ( .a(n5348), .b(n5081), .c(n5346), .o(n5349) );
no02f01 g01561 ( .a(n5081), .b(n5346), .o(n5350_1) );
no02f01 g01562 ( .a(n5347), .b(n5350_1), .o(n5351) );
no02f01 g01563 ( .a(n5351), .b(n5349), .o(n5352) );
in01f01 g01564 ( .a(n5352), .o(n5353) );
no02f01 g01565 ( .a(n5353), .b(n5119), .o(n5354) );
no03f01 g01566 ( .a(n5354), .b(n5345_1), .c(n5336), .o(n5355_1) );
na02f01 g01567 ( .a(n5355_1), .b(n5312), .o(n5356) );
in01f01 g01568 ( .a(n5356), .o(n5357) );
in01f01 g01569 ( .a(n5087), .o(n5358) );
na02f01 g01570 ( .a(n5358), .b(n5078), .o(n5359) );
na03f01 g01571 ( .a(n5359), .b(n5085_1), .c(n5009), .o(n5360_1) );
in01f01 g01572 ( .a(n5006_1), .o(n5361) );
no02f01 g01573 ( .a(n5361), .b(n5005), .o(n5362) );
in01f01 g01574 ( .a(n5362), .o(n5363) );
no02f01 g01575 ( .a(n5363), .b(n5360_1), .o(n5364) );
na02f01 g01576 ( .a(n5363), .b(n5360_1), .o(n5365_1) );
in01f01 g01577 ( .a(n5365_1), .o(n5366) );
no03f01 g01578 ( .a(n5366), .b(n5364), .c(n5142), .o(n5367) );
no02f01 g01579 ( .a(n5086), .b(n5078), .o(n5368) );
no02f01 g01580 ( .a(n5087), .b(n5008), .o(n5369) );
no02f01 g01581 ( .a(n5369), .b(n5368), .o(n5370_1) );
na02f01 g01582 ( .a(n5369), .b(n5368), .o(n5371) );
in01f01 g01583 ( .a(n5371), .o(n5372) );
no02f01 g01584 ( .a(n5372), .b(n5370_1), .o(n5373) );
in01f01 g01585 ( .a(n5373), .o(n5374) );
no02f01 g01586 ( .a(n5374), .b(n5142), .o(n5375_1) );
no02f01 g01587 ( .a(n5375_1), .b(n5367), .o(n5376) );
in01f01 g01588 ( .a(n5376), .o(n5377) );
in01f01 g01589 ( .a(n5089), .o(n5378) );
no02f01 g01590 ( .a(n5378), .b(n5010), .o(n5379) );
no02f01 g01591 ( .a(n_45224), .b(n5002), .o(n5380_1) );
no02f01 g01592 ( .a(n5380_1), .b(n4999), .o(n5381) );
no02f01 g01593 ( .a(n5381), .b(n5379), .o(n5382) );
na02f01 g01594 ( .a(n5381), .b(n5379), .o(n5383) );
in01f01 g01595 ( .a(n5383), .o(n5384) );
no02f01 g01596 ( .a(n5384), .b(n5382), .o(n5385_1) );
in01f01 g01597 ( .a(n5385_1), .o(n5386) );
no02f01 g01598 ( .a(n5386), .b(n5142), .o(n5387) );
in01f01 g01599 ( .a(n5380_1), .o(n5388) );
ao12f01 g01600 ( .a(n4999), .b(n5379), .c(n5388), .o(n5389) );
no02f01 g01601 ( .a(n_45224), .b(n5003), .o(n5390_1) );
no02f01 g01602 ( .a(n5390_1), .b(n4998), .o(n5391) );
in01f01 g01603 ( .a(n5391), .o(n5392) );
no02f01 g01604 ( .a(n5392), .b(n5389), .o(n5393) );
na02f01 g01605 ( .a(n5392), .b(n5389), .o(n5394) );
in01f01 g01606 ( .a(n5394), .o(n5395_1) );
no03f01 g01607 ( .a(n5395_1), .b(n5393), .c(n5142), .o(n5396) );
no02f01 g01608 ( .a(n5396), .b(n5387), .o(n5397) );
in01f01 g01609 ( .a(n5397), .o(n5398) );
no02f01 g01610 ( .a(n5398), .b(n5377), .o(n5399) );
no02f01 g01611 ( .a(n5332), .b(n5142), .o(n5400_1) );
in01f01 g01612 ( .a(n5400_1), .o(n5401) );
no02f01 g01613 ( .a(n5352), .b(n5142), .o(n5402) );
no02f01 g01614 ( .a(n5325_1), .b(n5142), .o(n5403) );
no02f01 g01615 ( .a(n5403), .b(n5402), .o(n5404) );
na02f01 g01616 ( .a(n5404), .b(n5401), .o(n5405_1) );
no02f01 g01617 ( .a(n5344), .b(n5342), .o(n5406) );
no02f01 g01618 ( .a(n5406), .b(n5142), .o(n5407) );
no02f01 g01619 ( .a(n5407), .b(n5405_1), .o(n5408) );
no02f01 g01620 ( .a(n5408), .b(n5377), .o(n5409) );
na02f01 g01621 ( .a(n5409), .b(n5397), .o(n5410_1) );
no02f01 g01622 ( .a(n5373), .b(n5119), .o(n5411) );
in01f01 g01623 ( .a(n5411), .o(n5412) );
in01f01 g01624 ( .a(n5364), .o(n5413) );
ao12f01 g01625 ( .a(n5119), .b(n5365_1), .c(n5413), .o(n5414) );
no02f01 g01626 ( .a(n5385_1), .b(n5119), .o(n5415_1) );
no02f01 g01627 ( .a(n5415_1), .b(n5414), .o(n5416) );
na02f01 g01628 ( .a(n5416), .b(n5412), .o(n5417) );
in01f01 g01629 ( .a(n5393), .o(n5418) );
ao12f01 g01630 ( .a(n5119), .b(n5394), .c(n5418), .o(n5419) );
no02f01 g01631 ( .a(n5419), .b(n5417), .o(n5420_1) );
na02f01 g01632 ( .a(n5420_1), .b(n5410_1), .o(n5421) );
ao12f01 g01633 ( .a(n5421), .b(n5399), .c(n5357), .o(n5422) );
in01f01 g01634 ( .a(n5422), .o(n5423) );
no02f01 g01635 ( .a(n_45224), .b(n5096), .o(n5424) );
in01f01 g01636 ( .a(n5106), .o(n5425_1) );
ao12f01 g01637 ( .a(n5424), .b(n5425_1), .c(n5090_1), .o(n5426) );
in01f01 g01638 ( .a(n5426), .o(n5427) );
no02f01 g01639 ( .a(n_45224), .b(n5097), .o(n5428) );
no02f01 g01640 ( .a(n5428), .b(n5107), .o(n5429) );
in01f01 g01641 ( .a(n5429), .o(n5430_1) );
no02f01 g01642 ( .a(n5430_1), .b(n5427), .o(n5431) );
no02f01 g01643 ( .a(n5429), .b(n5426), .o(n5432) );
no02f01 g01644 ( .a(n5432), .b(n5431), .o(n5433) );
no02f01 g01645 ( .a(n5433), .b(n5119), .o(n5434) );
ao12f01 g01646 ( .a(n5098), .b(n5108), .c(n5090_1), .o(n5435_1) );
no02f01 g01647 ( .a(n_45224), .b(n5100_1), .o(n5436) );
no02f01 g01648 ( .a(n5110_1), .b(n5436), .o(n5437) );
no02f01 g01649 ( .a(n5437), .b(n5435_1), .o(n5438) );
na02f01 g01650 ( .a(n5437), .b(n5435_1), .o(n5439) );
in01f01 g01651 ( .a(n5439), .o(n5440_1) );
no02f01 g01652 ( .a(n5440_1), .b(n5438), .o(n5441) );
no02f01 g01653 ( .a(n5441), .b(n5119), .o(n5442) );
in01f01 g01654 ( .a(n5090_1), .o(n5443) );
no02f01 g01655 ( .a(n5106), .b(n5424), .o(n5444) );
no02f01 g01656 ( .a(n5444), .b(n5443), .o(n5445_1) );
na02f01 g01657 ( .a(n5444), .b(n5443), .o(n5446) );
in01f01 g01658 ( .a(n5446), .o(n5447) );
no02f01 g01659 ( .a(n5447), .b(n5445_1), .o(n5448) );
no02f01 g01660 ( .a(n5448), .b(n5119), .o(n5449) );
no03f01 g01661 ( .a(n5449), .b(n5442), .c(n5434), .o(n5450_1) );
in01f01 g01662 ( .a(n5108), .o(n5451) );
no03f01 g01663 ( .a(n5110_1), .b(n5451), .c(n5443), .o(n5452) );
no03f01 g01664 ( .a(n5452), .b(n5436), .c(n5098), .o(n5453) );
no02f01 g01665 ( .a(n_45224), .b(n5099), .o(n5454) );
no02f01 g01666 ( .a(n5454), .b(n5109), .o(n5455_1) );
no02f01 g01667 ( .a(n5455_1), .b(n5453), .o(n5456) );
na02f01 g01668 ( .a(n5455_1), .b(n5453), .o(n5457) );
in01f01 g01669 ( .a(n5457), .o(n5458) );
no02f01 g01670 ( .a(n5458), .b(n5456), .o(n5459_1) );
no02f01 g01671 ( .a(n5459_1), .b(n5119), .o(n5460) );
no02f01 g01672 ( .a(n5112), .b(n5443), .o(n5461) );
no02f01 g01673 ( .a(n5461), .b(n5103), .o(n5462) );
no02f01 g01674 ( .a(n_45224), .b(n5091), .o(n5463) );
no02f01 g01675 ( .a(n5114), .b(n5463), .o(n5464_1) );
no02f01 g01676 ( .a(n5464_1), .b(n5462), .o(n5465) );
na02f01 g01677 ( .a(n5464_1), .b(n5462), .o(n5466) );
in01f01 g01678 ( .a(n5466), .o(n5467) );
no02f01 g01679 ( .a(n5467), .b(n5465), .o(n5468) );
no02f01 g01680 ( .a(n5468), .b(n5119), .o(n5469_1) );
no02f01 g01681 ( .a(n5469_1), .b(n5460), .o(n5470) );
na02f01 g01682 ( .a(n5470), .b(n5450_1), .o(n5471) );
no02f01 g01683 ( .a(n5471), .b(n5423), .o(n5472) );
in01f01 g01684 ( .a(n5472), .o(n5473) );
in01f01 g01685 ( .a(n5461), .o(n5474_1) );
no02f01 g01686 ( .a(n5474_1), .b(n5114), .o(n5475) );
no03f01 g01687 ( .a(n5475), .b(n5103), .c(n5463), .o(n5476) );
no02f01 g01688 ( .a(n_45224), .b(n5092), .o(n5477) );
no02f01 g01689 ( .a(n5477), .b(n5115_1), .o(n5478) );
no02f01 g01690 ( .a(n5478), .b(n5476), .o(n5479_1) );
na02f01 g01691 ( .a(n5478), .b(n5476), .o(n5480) );
in01f01 g01692 ( .a(n5480), .o(n5481) );
no02f01 g01693 ( .a(n5481), .b(n5479_1), .o(n5482) );
no02f01 g01694 ( .a(n5482), .b(n5119), .o(n5483_1) );
na02f01 g01695 ( .a(n5433), .b(n5119), .o(n5484) );
in01f01 g01696 ( .a(n5484), .o(n5485) );
na02f01 g01697 ( .a(n5448), .b(n5119), .o(n5486) );
in01f01 g01698 ( .a(n5486), .o(n5487) );
no02f01 g01699 ( .a(n5487), .b(n5485), .o(n5488_1) );
in01f01 g01700 ( .a(n5488_1), .o(n5489) );
na02f01 g01701 ( .a(n5441), .b(n5119), .o(n5490) );
in01f01 g01702 ( .a(n5490), .o(n5491) );
no02f01 g01703 ( .a(n5491), .b(n5489), .o(n5492) );
in01f01 g01704 ( .a(n5492), .o(n5493_1) );
na02f01 g01705 ( .a(n5459_1), .b(n5119), .o(n5494) );
in01f01 g01706 ( .a(n5494), .o(n5495) );
no02f01 g01707 ( .a(n5495), .b(n5493_1), .o(n5496) );
in01f01 g01708 ( .a(n5496), .o(n5497) );
na02f01 g01709 ( .a(n5482), .b(n5119), .o(n5498_1) );
in01f01 g01710 ( .a(n5498_1), .o(n5499) );
na02f01 g01711 ( .a(n5468), .b(n5119), .o(n5500) );
in01f01 g01712 ( .a(n5500), .o(n5501) );
no02f01 g01713 ( .a(n5501), .b(n5499), .o(n5502) );
in01f01 g01714 ( .a(n5502), .o(n5503_1) );
no02f01 g01715 ( .a(n5503_1), .b(n5497), .o(n5504) );
oa12f01 g01716 ( .a(n5504), .b(n5483_1), .c(n5473), .o(n5505) );
in01f01 g01717 ( .a(n5505), .o(n5506) );
no02f01 g01718 ( .a(n5474_1), .b(n5117), .o(n5507) );
no03f01 g01719 ( .a(n5507), .b(n5103), .c(n5093), .o(n5508_1) );
in01f01 g01720 ( .a(n5508_1), .o(n5509) );
in01f01 g01721 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_29_), .o(n5510) );
no02f01 g01722 ( .a(n_45224), .b(n5510), .o(n5511) );
no02f01 g01723 ( .a(n5511), .b(n5113), .o(n5512) );
in01f01 g01724 ( .a(n5512), .o(n5513_1) );
no02f01 g01725 ( .a(n5513_1), .b(n5509), .o(n5514) );
no02f01 g01726 ( .a(n5512), .b(n5508_1), .o(n5515) );
no02f01 g01727 ( .a(n5515), .b(n5514), .o(n5516) );
no02f01 g01728 ( .a(n5516), .b(n5119), .o(n5517) );
na02f01 g01729 ( .a(n5516), .b(n5119), .o(n5518_1) );
in01f01 g01730 ( .a(n5518_1), .o(n5519) );
no02f01 g01731 ( .a(n5519), .b(n5517), .o(n5520) );
in01f01 g01732 ( .a(n5520), .o(n5521) );
no02f01 g01733 ( .a(n5521), .b(n5506), .o(n5522) );
no02f01 g01734 ( .a(n5520), .b(n5505), .o(n5523_1) );
no03f01 g01735 ( .a(n5519), .b(n5503_1), .c(n5497), .o(n5524) );
in01f01 g01736 ( .a(n5524), .o(n5525) );
no03f01 g01737 ( .a(n5517), .b(n5483_1), .c(n5471), .o(n5526) );
oa12f01 g01738 ( .a(n5526), .b(n5525), .c(n5422), .o(n5527) );
no03f01 g01739 ( .a(n5527), .b(n5523_1), .c(n5522), .o(n5528_1) );
in01f01 g01740 ( .a(n5527), .o(n5529) );
ao12f01 g01741 ( .a(n5449), .b(n5486), .c(n5423), .o(n5530) );
in01f01 g01742 ( .a(n5530), .o(n5531) );
no02f01 g01743 ( .a(n5485), .b(n5434), .o(n5532) );
in01f01 g01744 ( .a(n5532), .o(n5533_1) );
no02f01 g01745 ( .a(n5533_1), .b(n5531), .o(n5534) );
no02f01 g01746 ( .a(n5532), .b(n5530), .o(n5535) );
no02f01 g01747 ( .a(n5535), .b(n5534), .o(n5536) );
no02f01 g01748 ( .a(n5536), .b(n5529), .o(n5537) );
no02f01 g01749 ( .a(n5487), .b(n5449), .o(n5538_1) );
in01f01 g01750 ( .a(n5538_1), .o(n5539) );
no02f01 g01751 ( .a(n5539), .b(n5423), .o(n5540) );
no02f01 g01752 ( .a(n5538_1), .b(n5422), .o(n5541) );
no02f01 g01753 ( .a(n5541), .b(n5540), .o(n5542) );
no02f01 g01754 ( .a(n5542), .b(n5529), .o(n5543_1) );
no02f01 g01755 ( .a(n5543_1), .b(n5537), .o(n5544) );
in01f01 g01756 ( .a(n5544), .o(n5545) );
no02f01 g01757 ( .a(n5449), .b(n5434), .o(n5546) );
oa12f01 g01758 ( .a(n5546), .b(n5489), .c(n5422), .o(n5547) );
in01f01 g01759 ( .a(n5547), .o(n5548_1) );
no02f01 g01760 ( .a(n5491), .b(n5442), .o(n5549) );
no02f01 g01761 ( .a(n5549), .b(n5548_1), .o(n5550) );
na02f01 g01762 ( .a(n5549), .b(n5548_1), .o(n5551) );
in01f01 g01763 ( .a(n5551), .o(n5552) );
no02f01 g01764 ( .a(n5552), .b(n5550), .o(n5553_1) );
no02f01 g01765 ( .a(n5553_1), .b(n5529), .o(n5554) );
ao12f01 g01766 ( .a(n5493_1), .b(n5450_1), .c(n5422), .o(n5555) );
no02f01 g01767 ( .a(n5495), .b(n5460), .o(n5556) );
in01f01 g01768 ( .a(n5556), .o(n5557) );
no02f01 g01769 ( .a(n5557), .b(n5555), .o(n5558_1) );
na02f01 g01770 ( .a(n5557), .b(n5555), .o(n5559) );
in01f01 g01771 ( .a(n5559), .o(n5560) );
no02f01 g01772 ( .a(n5560), .b(n5558_1), .o(n5561) );
no02f01 g01773 ( .a(n5561), .b(n5529), .o(n5562) );
no03f01 g01774 ( .a(n5562), .b(n5554), .c(n5545), .o(n5563_1) );
na03f01 g01775 ( .a(n5500), .b(n5496), .c(n5473), .o(n5564) );
no02f01 g01776 ( .a(n5499), .b(n5483_1), .o(n5565) );
no02f01 g01777 ( .a(n5565), .b(n5564), .o(n5566) );
na02f01 g01778 ( .a(n5565), .b(n5564), .o(n5567) );
in01f01 g01779 ( .a(n5567), .o(n5568_1) );
no03f01 g01780 ( .a(n5568_1), .b(n5566), .c(n5527), .o(n5569) );
in01f01 g01781 ( .a(n5450_1), .o(n5570) );
no02f01 g01782 ( .a(n5460), .b(n5570), .o(n5571) );
oa12f01 g01783 ( .a(n5571), .b(n5497), .c(n5422), .o(n5572) );
in01f01 g01784 ( .a(n5572), .o(n5573_1) );
no02f01 g01785 ( .a(n5501), .b(n5469_1), .o(n5574) );
no02f01 g01786 ( .a(n5574), .b(n5573_1), .o(n5575) );
na02f01 g01787 ( .a(n5574), .b(n5573_1), .o(n5576) );
in01f01 g01788 ( .a(n5576), .o(n5577) );
no03f01 g01789 ( .a(n5577), .b(n5575), .c(n5527), .o(n5578_1) );
no02f01 g01790 ( .a(n5578_1), .b(n5569), .o(n5579) );
in01f01 g01791 ( .a(n5579), .o(n5580) );
no02f01 g01792 ( .a(n5580), .b(n5563_1), .o(n5581) );
in01f01 g01793 ( .a(n5566), .o(n5582) );
ao12f01 g01794 ( .a(n5529), .b(n5567), .c(n5582), .o(n5583_1) );
no02f01 g01795 ( .a(n5577), .b(n5575), .o(n5584) );
no02f01 g01796 ( .a(n5584), .b(n5529), .o(n5585) );
no02f01 g01797 ( .a(n5585), .b(n5583_1), .o(n5586) );
in01f01 g01798 ( .a(n5586), .o(n5587) );
no02f01 g01799 ( .a(n5523_1), .b(n5522), .o(n5588_1) );
no02f01 g01800 ( .a(n5529), .b(n5588_1), .o(n5589) );
no03f01 g01801 ( .a(n5589), .b(n5587), .c(n5581), .o(n5590) );
no02f01 g01802 ( .a(n5590), .b(n5528_1), .o(n5591) );
in01f01 g01803 ( .a(n5591), .o(n5592) );
no03f01 g01804 ( .a(n5204), .b(n5202), .c(n5198), .o(n5593_1) );
no02f01 g01805 ( .a(n5203), .b(n5129), .o(n5594) );
no02f01 g01806 ( .a(n5594), .b(n5593_1), .o(n5595) );
na02f01 g01807 ( .a(n5594), .b(n5593_1), .o(n5596) );
in01f01 g01808 ( .a(n5596), .o(n5597) );
no02f01 g01809 ( .a(n5597), .b(n5595), .o(n5598_1) );
in01f01 g01810 ( .a(n5598_1), .o(n5599) );
no02f01 g01811 ( .a(n5599), .b(n5529), .o(n5600) );
in01f01 g01812 ( .a(n5159), .o(n5601) );
no02f01 g01813 ( .a(n5160_1), .b(n5141), .o(n5602) );
in01f01 g01814 ( .a(n5602), .o(n5603_1) );
no03f01 g01815 ( .a(n5603_1), .b(n5161), .c(n5601), .o(n5604) );
in01f01 g01816 ( .a(n5161), .o(n5605) );
ao12f01 g01817 ( .a(n5602), .b(n5605), .c(n5159), .o(n5606) );
no02f01 g01818 ( .a(n5606), .b(n5604), .o(n5607) );
in01f01 g01819 ( .a(n5607), .o(n5608_1) );
no02f01 g01820 ( .a(n5608_1), .b(n5529), .o(n5609) );
in01f01 g01821 ( .a(n5158), .o(n5610) );
in01f01 g01822 ( .a(n5148), .o(n5611) );
no02f01 g01823 ( .a(n5161), .b(n5611), .o(n5612) );
no02f01 g01824 ( .a(n5612), .b(n5610), .o(n5613_1) );
na02f01 g01825 ( .a(n5612), .b(n5610), .o(n5614) );
in01f01 g01826 ( .a(n5614), .o(n5615) );
no02f01 g01827 ( .a(n5615), .b(n5613_1), .o(n5616) );
in01f01 g01828 ( .a(n5616), .o(n5617) );
no02f01 g01829 ( .a(n5617), .b(n5529), .o(n5618_1) );
in01f01 g01830 ( .a(n5618_1), .o(n5619) );
in01f01 g01831 ( .a(n5156), .o(n5620) );
no03f01 g01832 ( .a(n5157), .b(n5620), .c(n5151), .o(n5621) );
in01f01 g01833 ( .a(n5157), .o(n5622) );
ao12f01 g01834 ( .a(cordic_combinational_sub_ln23_0_unr12_z_0_), .b(n5622), .c(n5156), .o(n5623_1) );
no02f01 g01835 ( .a(n5623_1), .b(n5621), .o(n5624) );
no02f01 g01836 ( .a(n5624), .b(n5527), .o(n5625) );
in01f01 g01837 ( .a(n5625), .o(n5626) );
na02f01 g01838 ( .a(n5624), .b(n5527), .o(n5627) );
na02f01 g01839 ( .a(n5627), .b(cordic_combinational_sub_ln23_0_unr12_z_0_), .o(n5628_1) );
na02f01 g01840 ( .a(n5628_1), .b(n5626), .o(n5629) );
na02f01 g01841 ( .a(n5629), .b(n5619), .o(n5630) );
no02f01 g01842 ( .a(n5616), .b(n5527), .o(n5631) );
no02f01 g01843 ( .a(n5607), .b(n5527), .o(n5632) );
no02f01 g01844 ( .a(n5632), .b(n5631), .o(n5633_1) );
oa12f01 g01845 ( .a(n5633_1), .b(n5630), .c(n5609), .o(n5634) );
in01f01 g01846 ( .a(n5634), .o(n5635) );
no02f01 g01847 ( .a(n5200_1), .b(n5173), .o(n5636) );
in01f01 g01848 ( .a(n5636), .o(n5637) );
no02f01 g01849 ( .a(n5637), .b(n5163), .o(n5638_1) );
in01f01 g01850 ( .a(n5163), .o(n5639) );
no02f01 g01851 ( .a(n5636), .b(n5639), .o(n5640) );
no02f01 g01852 ( .a(n5640), .b(n5638_1), .o(n5641) );
in01f01 g01853 ( .a(n5641), .o(n5642) );
no02f01 g01854 ( .a(n5642), .b(n5529), .o(n5643_1) );
no02f01 g01855 ( .a(n5643_1), .b(n5635), .o(n5644) );
in01f01 g01856 ( .a(n5175_1), .o(n5645) );
in01f01 g01857 ( .a(n5195_1), .o(n5646) );
ao12f01 g01858 ( .a(n5202), .b(n5646), .c(n5645), .o(n5647) );
in01f01 g01859 ( .a(n5647), .o(n5648_1) );
no02f01 g01860 ( .a(n5204), .b(n5183), .o(n5649) );
in01f01 g01861 ( .a(n5649), .o(n5650) );
no02f01 g01862 ( .a(n5650), .b(n5648_1), .o(n5651) );
no02f01 g01863 ( .a(n5649), .b(n5647), .o(n5652) );
no02f01 g01864 ( .a(n5652), .b(n5651), .o(n5653_1) );
in01f01 g01865 ( .a(n5653_1), .o(n5654) );
no02f01 g01866 ( .a(n5654), .b(n5529), .o(n5655) );
no02f01 g01867 ( .a(n5199), .b(n5195_1), .o(n5656) );
in01f01 g01868 ( .a(n5656), .o(n5657_1) );
no03f01 g01869 ( .a(n5657_1), .b(n5200_1), .c(n5645), .o(n5658) );
in01f01 g01870 ( .a(n5200_1), .o(n5659) );
ao12f01 g01871 ( .a(n5656), .b(n5659), .c(n5175_1), .o(n5660) );
no02f01 g01872 ( .a(n5660), .b(n5658), .o(n5661) );
in01f01 g01873 ( .a(n5661), .o(n5662_1) );
no02f01 g01874 ( .a(n5662_1), .b(n5529), .o(n5663) );
no02f01 g01875 ( .a(n5663), .b(n5655), .o(n5664) );
na02f01 g01876 ( .a(n5664), .b(n5644), .o(n5665) );
no02f01 g01877 ( .a(n5661), .b(n5527), .o(n5666) );
no02f01 g01878 ( .a(n5641), .b(n5527), .o(n5667_1) );
no02f01 g01879 ( .a(n5667_1), .b(n5666), .o(n5668) );
in01f01 g01880 ( .a(n5668), .o(n5669) );
no02f01 g01881 ( .a(n5598_1), .b(n5527), .o(n5670) );
no02f01 g01882 ( .a(n5653_1), .b(n5527), .o(n5671) );
no03f01 g01883 ( .a(n5671), .b(n5670), .c(n5669), .o(n5672_1) );
oa12f01 g01884 ( .a(n5672_1), .b(n5665), .c(n5600), .o(n5673) );
no02f01 g01885 ( .a(n5300_1), .b(n5228), .o(n5674) );
no02f01 g01886 ( .a(n5674), .b(n5207), .o(n5675) );
na02f01 g01887 ( .a(n5674), .b(n5207), .o(n5676) );
in01f01 g01888 ( .a(n5676), .o(n5677_1) );
no02f01 g01889 ( .a(n5677_1), .b(n5675), .o(n5678) );
in01f01 g01890 ( .a(n5678), .o(n5679) );
no02f01 g01891 ( .a(n5679), .b(n5529), .o(n5680) );
no02f01 g01892 ( .a(n5228), .b(n5207), .o(n5681) );
no02f01 g01893 ( .a(n5681), .b(n5300_1), .o(n5682_1) );
no02f01 g01894 ( .a(n5299), .b(n5220_1), .o(n5683) );
no02f01 g01895 ( .a(n5683), .b(n5682_1), .o(n5684) );
na02f01 g01896 ( .a(n5683), .b(n5682_1), .o(n5685) );
in01f01 g01897 ( .a(n5685), .o(n5686) );
no02f01 g01898 ( .a(n5686), .b(n5684), .o(n5687_1) );
in01f01 g01899 ( .a(n5687_1), .o(n5688) );
no02f01 g01900 ( .a(n5688), .b(n5529), .o(n5689) );
no02f01 g01901 ( .a(n5689), .b(n5680), .o(n5690) );
na02f01 g01902 ( .a(n5690), .b(n5673), .o(n5691) );
in01f01 g01903 ( .a(n5231), .o(n5692_1) );
in01f01 g01904 ( .a(n5301), .o(n5693) );
no02f01 g01905 ( .a(n5302), .b(n5693), .o(n5694) );
oa12f01 g01906 ( .a(n5694), .b(n5243), .c(n5692_1), .o(n5695) );
in01f01 g01907 ( .a(n5695), .o(n5696) );
no02f01 g01908 ( .a(n5303), .b(n5251), .o(n5697_1) );
no02f01 g01909 ( .a(n5697_1), .b(n5696), .o(n5698) );
na02f01 g01910 ( .a(n5697_1), .b(n5696), .o(n5699) );
in01f01 g01911 ( .a(n5699), .o(n5700) );
no02f01 g01912 ( .a(n5700), .b(n5698), .o(n5701_1) );
in01f01 g01913 ( .a(n5701_1), .o(n5702) );
no02f01 g01914 ( .a(n5702), .b(n5529), .o(n5703) );
no02f01 g01915 ( .a(n5693), .b(n5231), .o(n5704) );
no02f01 g01916 ( .a(n5302), .b(n5243), .o(n5705) );
no02f01 g01917 ( .a(n5705), .b(n5704), .o(n5706_1) );
na02f01 g01918 ( .a(n5705), .b(n5704), .o(n5707) );
in01f01 g01919 ( .a(n5707), .o(n5708) );
no02f01 g01920 ( .a(n5708), .b(n5706_1), .o(n5709) );
in01f01 g01921 ( .a(n5709), .o(n5710) );
no02f01 g01922 ( .a(n5710), .b(n5529), .o(n5711_1) );
no02f01 g01923 ( .a(n5711_1), .b(n5703), .o(n5712) );
in01f01 g01924 ( .a(n5712), .o(n5713) );
no02f01 g01925 ( .a(n5678), .b(n5527), .o(n5714) );
no02f01 g01926 ( .a(n5687_1), .b(n5527), .o(n5715) );
no02f01 g01927 ( .a(n5715), .b(n5714), .o(n5716_1) );
in01f01 g01928 ( .a(n5716_1), .o(n5717) );
no02f01 g01929 ( .a(n5709), .b(n5527), .o(n5718) );
no02f01 g01930 ( .a(n5701_1), .b(n5527), .o(n5719) );
no03f01 g01931 ( .a(n5719), .b(n5718), .c(n5717), .o(n5720) );
oa12f01 g01932 ( .a(n5720), .b(n5713), .c(n5691), .o(n5721_1) );
in01f01 g01933 ( .a(n5721_1), .o(n5722) );
in01f01 g01934 ( .a(n5253), .o(n5723) );
na02f01 g01935 ( .a(n5304), .b(n5301), .o(n5724) );
no02f01 g01936 ( .a(n5305_1), .b(n5262), .o(n5725) );
in01f01 g01937 ( .a(n5725), .o(n5726_1) );
no03f01 g01938 ( .a(n5726_1), .b(n5724), .c(n5723), .o(n5727) );
in01f01 g01939 ( .a(n5724), .o(n5728) );
ao12f01 g01940 ( .a(n5725), .b(n5728), .c(n5253), .o(n5729) );
no02f01 g01941 ( .a(n5729), .b(n5727), .o(n5730_1) );
in01f01 g01942 ( .a(n5730_1), .o(n5731) );
no02f01 g01943 ( .a(n5731), .b(n5529), .o(n5732) );
no02f01 g01944 ( .a(n5305_1), .b(n5724), .o(n5733) );
oa12f01 g01945 ( .a(n5733), .b(n5262), .c(n5253), .o(n5734) );
in01f01 g01946 ( .a(n5734), .o(n5735_1) );
no02f01 g01947 ( .a(n5306), .b(n5272), .o(n5736) );
no02f01 g01948 ( .a(n5736), .b(n5735_1), .o(n5737) );
na02f01 g01949 ( .a(n5736), .b(n5735_1), .o(n5738) );
in01f01 g01950 ( .a(n5738), .o(n5739) );
no02f01 g01951 ( .a(n5739), .b(n5737), .o(n5740_1) );
in01f01 g01952 ( .a(n5740_1), .o(n5741) );
no02f01 g01953 ( .a(n5741), .b(n5529), .o(n5742) );
no03f01 g01954 ( .a(n5742), .b(n5732), .c(n5722), .o(n5743) );
no02f01 g01955 ( .a(n5309), .b(n5296), .o(n5744) );
in01f01 g01956 ( .a(n5744), .o(n5745_1) );
no03f01 g01957 ( .a(n5745_1), .b(n5308), .c(n5275_1), .o(n5746) );
no02f01 g01958 ( .a(n5308), .b(n5275_1), .o(n5747) );
no02f01 g01959 ( .a(n5744), .b(n5747), .o(n5748) );
no02f01 g01960 ( .a(n5748), .b(n5746), .o(n5749) );
in01f01 g01961 ( .a(n5749), .o(n5750_1) );
no02f01 g01962 ( .a(n5750_1), .b(n5529), .o(n5751) );
in01f01 g01963 ( .a(n5751), .o(n5752) );
na02f01 g01964 ( .a(n5752), .b(n5743), .o(n5753) );
no02f01 g01965 ( .a(n5740_1), .b(n5527), .o(n5754) );
no02f01 g01966 ( .a(n5730_1), .b(n5527), .o(n5755_1) );
no02f01 g01967 ( .a(n5755_1), .b(n5754), .o(n5756) );
in01f01 g01968 ( .a(n5756), .o(n5757) );
no03f01 g01969 ( .a(n5296), .b(n5274), .c(n5253), .o(n5758) );
no03f01 g01970 ( .a(n5758), .b(n5309), .c(n5308), .o(n5759) );
no02f01 g01971 ( .a(n5310_1), .b(n5286), .o(n5760_1) );
no02f01 g01972 ( .a(n5760_1), .b(n5759), .o(n5761) );
na02f01 g01973 ( .a(n5760_1), .b(n5759), .o(n5762) );
in01f01 g01974 ( .a(n5762), .o(n5763) );
no02f01 g01975 ( .a(n5763), .b(n5761), .o(n5764) );
no02f01 g01976 ( .a(n5764), .b(n5527), .o(n5765_1) );
no02f01 g01977 ( .a(n5749), .b(n5527), .o(n5766) );
no03f01 g01978 ( .a(n5766), .b(n5765_1), .c(n5757), .o(n5767) );
na02f01 g01979 ( .a(n5764), .b(n5527), .o(n5768) );
in01f01 g01980 ( .a(n5768), .o(n5769_1) );
ao12f01 g01981 ( .a(n5769_1), .b(n5767), .c(n5753), .o(n5770) );
in01f01 g01982 ( .a(n5770), .o(n5771) );
no02f01 g01983 ( .a(n5400_1), .b(n5334), .o(n5772) );
in01f01 g01984 ( .a(n5772), .o(n5773) );
no02f01 g01985 ( .a(n5773), .b(n5312), .o(n5774_1) );
in01f01 g01986 ( .a(n5312), .o(n5775) );
no02f01 g01987 ( .a(n5772), .b(n5775), .o(n5776) );
no02f01 g01988 ( .a(n5776), .b(n5774_1), .o(n5777) );
in01f01 g01989 ( .a(n5777), .o(n5778) );
no02f01 g01990 ( .a(n5778), .b(n5529), .o(n5779_1) );
oa12f01 g01991 ( .a(n5401), .b(n5334), .c(n5775), .o(n5780) );
in01f01 g01992 ( .a(n5780), .o(n5781) );
no02f01 g01993 ( .a(n5403), .b(n5327), .o(n5782) );
no02f01 g01994 ( .a(n5782), .b(n5781), .o(n5783) );
na02f01 g01995 ( .a(n5782), .b(n5781), .o(n5784_1) );
in01f01 g01996 ( .a(n5784_1), .o(n5785) );
no02f01 g01997 ( .a(n5785), .b(n5783), .o(n5786) );
in01f01 g01998 ( .a(n5786), .o(n5787) );
no02f01 g01999 ( .a(n5787), .b(n5529), .o(n5788) );
no02f01 g02000 ( .a(n5403), .b(n5400_1), .o(n5789_1) );
oa12f01 g02001 ( .a(n5789_1), .b(n5336), .c(n5775), .o(n5790) );
in01f01 g02002 ( .a(n5790), .o(n5791) );
no02f01 g02003 ( .a(n5402), .b(n5354), .o(n5792) );
no02f01 g02004 ( .a(n5792), .b(n5791), .o(n5793) );
na02f01 g02005 ( .a(n5792), .b(n5791), .o(n5794_1) );
in01f01 g02006 ( .a(n5794_1), .o(n5795) );
no03f01 g02007 ( .a(n5795), .b(n5793), .c(n5529), .o(n5796) );
no04f01 g02008 ( .a(n5796), .b(n5788), .c(n5779_1), .d(n5771), .o(n5797) );
in01f01 g02009 ( .a(n5354), .o(n5798) );
no02f01 g02010 ( .a(n5336), .b(n5775), .o(n5799_1) );
ao12f01 g02011 ( .a(n5405_1), .b(n5799_1), .c(n5798), .o(n5800) );
in01f01 g02012 ( .a(n5800), .o(n5801) );
no02f01 g02013 ( .a(n5407), .b(n5345_1), .o(n5802) );
in01f01 g02014 ( .a(n5802), .o(n5803) );
no02f01 g02015 ( .a(n5803), .b(n5801), .o(n5804_1) );
no02f01 g02016 ( .a(n5802), .b(n5800), .o(n5805) );
no02f01 g02017 ( .a(n5805), .b(n5804_1), .o(n5806) );
in01f01 g02018 ( .a(n5806), .o(n5807) );
no02f01 g02019 ( .a(n5807), .b(n5527), .o(n5808) );
in01f01 g02020 ( .a(n5808), .o(n5809_1) );
no02f01 g02021 ( .a(n5786), .b(n5527), .o(n5810) );
no02f01 g02022 ( .a(n5777), .b(n5527), .o(n5811) );
no02f01 g02023 ( .a(n5811), .b(n5810), .o(n5812) );
in01f01 g02024 ( .a(n5793), .o(n5813) );
ao12f01 g02025 ( .a(n5527), .b(n5794_1), .c(n5813), .o(n5814_1) );
no02f01 g02026 ( .a(n5806), .b(n5529), .o(n5815) );
no02f01 g02027 ( .a(n5815), .b(n5814_1), .o(n5816) );
ao12f01 g02028 ( .a(n5808), .b(n5816), .c(n5812), .o(n5817) );
ao12f01 g02029 ( .a(n5817), .b(n5809_1), .c(n5797), .o(n5818) );
in01f01 g02030 ( .a(n5387), .o(n5819_1) );
in01f01 g02031 ( .a(n5408), .o(n5820) );
oa12f01 g02032 ( .a(n5376), .b(n5820), .c(n5357), .o(n5821) );
in01f01 g02033 ( .a(n5821), .o(n5822) );
ao12f01 g02034 ( .a(n5417), .b(n5822), .c(n5819_1), .o(n5823) );
in01f01 g02035 ( .a(n5823), .o(n5824_1) );
no02f01 g02036 ( .a(n5419), .b(n5396), .o(n5825) );
in01f01 g02037 ( .a(n5825), .o(n5826) );
no02f01 g02038 ( .a(n5826), .b(n5824_1), .o(n5827) );
no02f01 g02039 ( .a(n5825), .b(n5823), .o(n5828) );
no03f01 g02040 ( .a(n5828), .b(n5827), .c(n5527), .o(n5829_1) );
no02f01 g02041 ( .a(n5820), .b(n5357), .o(n5830) );
no02f01 g02042 ( .a(n5830), .b(n5375_1), .o(n5831) );
no02f01 g02043 ( .a(n5831), .b(n5411), .o(n5832) );
no02f01 g02044 ( .a(n5414), .b(n5367), .o(n5833) );
no02f01 g02045 ( .a(n5833), .b(n5832), .o(n5834_1) );
na02f01 g02046 ( .a(n5833), .b(n5832), .o(n5835) );
in01f01 g02047 ( .a(n5835), .o(n5836) );
no03f01 g02048 ( .a(n5836), .b(n5834_1), .c(n5527), .o(n5837) );
no02f01 g02049 ( .a(n5411), .b(n5375_1), .o(n5838) );
in01f01 g02050 ( .a(n5838), .o(n5839_1) );
no03f01 g02051 ( .a(n5839_1), .b(n5820), .c(n5357), .o(n5840) );
no02f01 g02052 ( .a(n5838), .b(n5830), .o(n5841) );
no03f01 g02053 ( .a(n5841), .b(n5840), .c(n5527), .o(n5842) );
no02f01 g02054 ( .a(n5414), .b(n5411), .o(n5843) );
na02f01 g02055 ( .a(n5843), .b(n5821), .o(n5844_1) );
no02f01 g02056 ( .a(n5415_1), .b(n5387), .o(n5845) );
in01f01 g02057 ( .a(n5845), .o(n5846) );
no02f01 g02058 ( .a(n5846), .b(n5844_1), .o(n5847) );
na02f01 g02059 ( .a(n5846), .b(n5844_1), .o(n5848) );
in01f01 g02060 ( .a(n5848), .o(n5849_1) );
no03f01 g02061 ( .a(n5849_1), .b(n5847), .c(n5527), .o(n5850) );
no04f01 g02062 ( .a(n5850), .b(n5842), .c(n5837), .d(n5829_1), .o(n5851) );
in01f01 g02063 ( .a(n5851), .o(n5852) );
no02f01 g02064 ( .a(n5828), .b(n5827), .o(n5853) );
no02f01 g02065 ( .a(n5853), .b(n5529), .o(n5854_1) );
in01f01 g02066 ( .a(n5834_1), .o(n5855) );
ao12f01 g02067 ( .a(n5529), .b(n5835), .c(n5855), .o(n5856) );
no02f01 g02068 ( .a(n5841), .b(n5840), .o(n5857) );
no02f01 g02069 ( .a(n5857), .b(n5529), .o(n5858) );
no02f01 g02070 ( .a(n5849_1), .b(n5847), .o(n5859_1) );
no02f01 g02071 ( .a(n5859_1), .b(n5529), .o(n5860) );
no04f01 g02072 ( .a(n5860), .b(n5858), .c(n5856), .d(n5854_1), .o(n5861) );
oa12f01 g02073 ( .a(n5861), .b(n5852), .c(n5818), .o(n5862) );
na02f01 g02074 ( .a(n5542), .b(n5529), .o(n5863) );
na02f01 g02075 ( .a(n5553_1), .b(n5529), .o(n5864_1) );
in01f01 g02076 ( .a(n5864_1), .o(n5865) );
na02f01 g02077 ( .a(n5536), .b(n5529), .o(n5866) );
in01f01 g02078 ( .a(n5866), .o(n5867) );
na02f01 g02079 ( .a(n5561), .b(n5529), .o(n5868) );
in01f01 g02080 ( .a(n5868), .o(n5869_1) );
no03f01 g02081 ( .a(n5869_1), .b(n5867), .c(n5865), .o(n5870) );
no02f01 g02082 ( .a(n5580), .b(n5528_1), .o(n5871) );
na04f01 g02083 ( .a(n5871), .b(n5870), .c(n5863), .d(n5862), .o(n5872) );
na02f01 g02084 ( .a(n5872), .b(n5592), .o(n5873) );
in01f01 g02085 ( .a(n5873), .o(n6037) );
no02f01 g02086 ( .a(n5779_1), .b(n5771), .o(n5875) );
in01f01 g02087 ( .a(n5788), .o(n5876) );
in01f01 g02088 ( .a(n5812), .o(n5877) );
ao12f01 g02089 ( .a(n5877), .b(n5876), .c(n5875), .o(n5878_1) );
no02f01 g02090 ( .a(n5814_1), .b(n5796), .o(n5879) );
no02f01 g02091 ( .a(n5879), .b(n5878_1), .o(n5880) );
na02f01 g02092 ( .a(n5879), .b(n5878_1), .o(n5881) );
in01f01 g02093 ( .a(n5881), .o(n5882) );
no02f01 g02094 ( .a(n5882), .b(n5880), .o(n5883_1) );
no02f01 g02095 ( .a(n5883_1), .b(n6037), .o(n5884) );
no02f01 g02096 ( .a(n5811), .b(n5779_1), .o(n5885) );
no02f01 g02097 ( .a(n5885), .b(n5771), .o(n5886) );
na02f01 g02098 ( .a(n5885), .b(n5771), .o(n5887) );
in01f01 g02099 ( .a(n5887), .o(n5888_1) );
no02f01 g02100 ( .a(n5888_1), .b(n5886), .o(n5889) );
no02f01 g02101 ( .a(n5810), .b(n5788), .o(n5890) );
in01f01 g02102 ( .a(n5890), .o(n5891) );
no03f01 g02103 ( .a(n5891), .b(n5811), .c(n5875), .o(n5892) );
no02f01 g02104 ( .a(n5811), .b(n5875), .o(n5893_1) );
no02f01 g02105 ( .a(n5890), .b(n5893_1), .o(n5894) );
no02f01 g02106 ( .a(n5894), .b(n5892), .o(n5895) );
ao12f01 g02107 ( .a(n5873), .b(n5895), .c(n5889), .o(n5896) );
na02f01 g02108 ( .a(n5627), .b(n5626), .o(n5897) );
no02f01 g02109 ( .a(n5897), .b(n5151), .o(n5898_1) );
in01f01 g02110 ( .a(n5898_1), .o(n5899) );
na03f01 g02111 ( .a(n5899), .b(n5872), .c(n5592), .o(n5900) );
no02f01 g02112 ( .a(n5897), .b(cordic_combinational_sub_ln23_0_unr12_z_0_), .o(n5901) );
in01f01 g02113 ( .a(n5901), .o(n5902) );
no02f01 g02114 ( .a(n5631), .b(n5618_1), .o(n5903_1) );
in01f01 g02115 ( .a(n5903_1), .o(n5904) );
no02f01 g02116 ( .a(n5904), .b(n5629), .o(n5905) );
na02f01 g02117 ( .a(n5904), .b(n5629), .o(n5906) );
in01f01 g02118 ( .a(n5906), .o(n5907) );
no02f01 g02119 ( .a(n5907), .b(n5905), .o(n5908_1) );
na02f01 g02120 ( .a(n5908_1), .b(n5873), .o(n5909) );
in01f01 g02121 ( .a(n5909), .o(n5910) );
ao12f01 g02122 ( .a(n5910), .b(n5902), .c(n5900), .o(n5911) );
no02f01 g02123 ( .a(n5908_1), .b(n5873), .o(n5912) );
ao12f01 g02124 ( .a(n5631), .b(n5629), .c(n5619), .o(n5913_1) );
in01f01 g02125 ( .a(n5913_1), .o(n5914) );
no02f01 g02126 ( .a(n5632), .b(n5609), .o(n5915) );
in01f01 g02127 ( .a(n5915), .o(n5916) );
no02f01 g02128 ( .a(n5916), .b(n5914), .o(n5917) );
no02f01 g02129 ( .a(n5915), .b(n5913_1), .o(n5918_1) );
no02f01 g02130 ( .a(n5918_1), .b(n5917), .o(n5919) );
in01f01 g02131 ( .a(n5919), .o(n5920) );
no03f01 g02132 ( .a(n5920), .b(n5912), .c(n5911), .o(n5921) );
na02f01 g02133 ( .a(n5920), .b(n5911), .o(n5922) );
oa12f01 g02134 ( .a(n5922), .b(n5921), .c(n5873), .o(n5923_1) );
no02f01 g02135 ( .a(n5667_1), .b(n5643_1), .o(n5924) );
in01f01 g02136 ( .a(n5924), .o(n5925) );
no02f01 g02137 ( .a(n5925), .b(n5634), .o(n5926) );
no02f01 g02138 ( .a(n5924), .b(n5635), .o(n5927) );
no02f01 g02139 ( .a(n5927), .b(n5926), .o(n5928_1) );
in01f01 g02140 ( .a(n5928_1), .o(n5929) );
no02f01 g02141 ( .a(n5929), .b(n6037), .o(n5930) );
in01f01 g02142 ( .a(n5930), .o(n5931) );
no02f01 g02143 ( .a(n5666), .b(n5663), .o(n5932) );
in01f01 g02144 ( .a(n5932), .o(n5933_1) );
no03f01 g02145 ( .a(n5933_1), .b(n5667_1), .c(n5644), .o(n5934) );
no02f01 g02146 ( .a(n5667_1), .b(n5644), .o(n5935) );
no02f01 g02147 ( .a(n5932), .b(n5935), .o(n5936) );
no02f01 g02148 ( .a(n5936), .b(n5934), .o(n5937) );
na02f01 g02149 ( .a(n5937), .b(n5873), .o(n5938_1) );
no03f01 g02150 ( .a(n5663), .b(n5643_1), .c(n5635), .o(n5939) );
no02f01 g02151 ( .a(n5671), .b(n5655), .o(n5940) );
in01f01 g02152 ( .a(n5940), .o(n5941) );
no03f01 g02153 ( .a(n5941), .b(n5939), .c(n5669), .o(n5942) );
no02f01 g02154 ( .a(n5939), .b(n5669), .o(n5943_1) );
no02f01 g02155 ( .a(n5940), .b(n5943_1), .o(n5944) );
no02f01 g02156 ( .a(n5944), .b(n5942), .o(n5945) );
na02f01 g02157 ( .a(n5945), .b(n5873), .o(n5946) );
na02f01 g02158 ( .a(n5946), .b(n5938_1), .o(n5947) );
in01f01 g02159 ( .a(n5947), .o(n5948_1) );
na03f01 g02160 ( .a(n5948_1), .b(n5931), .c(n5923_1), .o(n5949) );
no02f01 g02161 ( .a(n5945), .b(n5873), .o(n5950) );
in01f01 g02162 ( .a(n5950), .o(n5951) );
no02f01 g02163 ( .a(n5671), .b(n5669), .o(n5952) );
na02f01 g02164 ( .a(n5952), .b(n5665), .o(n5953_1) );
no02f01 g02165 ( .a(n5670), .b(n5600), .o(n5954) );
in01f01 g02166 ( .a(n5954), .o(n5955) );
no02f01 g02167 ( .a(n5955), .b(n5953_1), .o(n5956) );
na02f01 g02168 ( .a(n5955), .b(n5953_1), .o(n5957) );
in01f01 g02169 ( .a(n5957), .o(n5958_1) );
no02f01 g02170 ( .a(n5958_1), .b(n5956), .o(n5959) );
na03f01 g02171 ( .a(n5959), .b(n5951), .c(n5949), .o(n5960) );
ao12f01 g02172 ( .a(n5873), .b(n5937), .c(n5928_1), .o(n5961) );
in01f01 g02173 ( .a(n5961), .o(n5962) );
oa12f01 g02174 ( .a(n5962), .b(n5959), .c(n5949), .o(n5963_1) );
ao12f01 g02175 ( .a(n5963_1), .b(n5960), .c(n6037), .o(n5964) );
in01f01 g02176 ( .a(n5680), .o(n5965) );
ao12f01 g02177 ( .a(n5714), .b(n5965), .c(n5673), .o(n5966) );
no02f01 g02178 ( .a(n5715), .b(n5689), .o(n5967) );
no02f01 g02179 ( .a(n5967), .b(n5966), .o(n5968_1) );
na02f01 g02180 ( .a(n5967), .b(n5966), .o(n5969) );
in01f01 g02181 ( .a(n5969), .o(n5970) );
no02f01 g02182 ( .a(n5970), .b(n5968_1), .o(n5971) );
in01f01 g02183 ( .a(n5971), .o(n5972) );
no02f01 g02184 ( .a(n5972), .b(n6037), .o(n5973_1) );
in01f01 g02185 ( .a(n5673), .o(n5974) );
no02f01 g02186 ( .a(n5714), .b(n5680), .o(n5975) );
no02f01 g02187 ( .a(n5975), .b(n5974), .o(n5976) );
na02f01 g02188 ( .a(n5975), .b(n5974), .o(n5977) );
in01f01 g02189 ( .a(n5977), .o(n5978_1) );
no02f01 g02190 ( .a(n5978_1), .b(n5976), .o(n5979) );
in01f01 g02191 ( .a(n5979), .o(n5980) );
no02f01 g02192 ( .a(n5980), .b(n6037), .o(n5981) );
no02f01 g02193 ( .a(n5981), .b(n5973_1), .o(n5982) );
in01f01 g02194 ( .a(n5982), .o(n5983_1) );
no02f01 g02195 ( .a(n5718), .b(n5717), .o(n5984) );
oa12f01 g02196 ( .a(n5984), .b(n5711_1), .c(n5691), .o(n5985) );
in01f01 g02197 ( .a(n5985), .o(n5986) );
no02f01 g02198 ( .a(n5719), .b(n5703), .o(n5987) );
no02f01 g02199 ( .a(n5987), .b(n5986), .o(n5988_1) );
na02f01 g02200 ( .a(n5987), .b(n5986), .o(n5989) );
in01f01 g02201 ( .a(n5989), .o(n5990) );
no02f01 g02202 ( .a(n5990), .b(n5988_1), .o(n5991) );
in01f01 g02203 ( .a(n5991), .o(n5992) );
no02f01 g02204 ( .a(n5992), .b(n6037), .o(n5993_1) );
na02f01 g02205 ( .a(n5716_1), .b(n5691), .o(n5994) );
in01f01 g02206 ( .a(n5994), .o(n5995) );
no02f01 g02207 ( .a(n5718), .b(n5711_1), .o(n5996) );
no02f01 g02208 ( .a(n5996), .b(n5995), .o(n5997) );
na02f01 g02209 ( .a(n5996), .b(n5995), .o(n5998_1) );
in01f01 g02210 ( .a(n5998_1), .o(n5999) );
no02f01 g02211 ( .a(n5999), .b(n5997), .o(n6000) );
in01f01 g02212 ( .a(n6000), .o(n6001) );
no02f01 g02213 ( .a(n6001), .b(n6037), .o(n6002) );
no03f01 g02214 ( .a(n6002), .b(n5993_1), .c(n5983_1), .o(n6003_1) );
in01f01 g02215 ( .a(n6003_1), .o(n6004) );
ao12f01 g02216 ( .a(n5873), .b(n5979), .c(n5971), .o(n6005) );
ao12f01 g02217 ( .a(n5873), .b(n6000), .c(n5991), .o(n6006) );
no02f01 g02218 ( .a(n6006), .b(n6005), .o(n6007_1) );
oa12f01 g02219 ( .a(n6007_1), .b(n6004), .c(n5964), .o(n6008) );
no02f01 g02220 ( .a(n5755_1), .b(n5732), .o(n6009) );
in01f01 g02221 ( .a(n6009), .o(n6010) );
no02f01 g02222 ( .a(n6010), .b(n5721_1), .o(n6011) );
no02f01 g02223 ( .a(n6009), .b(n5722), .o(n6012_1) );
no02f01 g02224 ( .a(n6012_1), .b(n6011), .o(n6013) );
in01f01 g02225 ( .a(n6013), .o(n6014) );
no02f01 g02226 ( .a(n6014), .b(n6037), .o(n6015) );
no02f01 g02227 ( .a(n5732), .b(n5722), .o(n6016) );
no02f01 g02228 ( .a(n5754), .b(n5742), .o(n6017_1) );
in01f01 g02229 ( .a(n6017_1), .o(n6018) );
no03f01 g02230 ( .a(n6018), .b(n5755_1), .c(n6016), .o(n6019) );
no02f01 g02231 ( .a(n5755_1), .b(n6016), .o(n6020) );
no02f01 g02232 ( .a(n6017_1), .b(n6020), .o(n6021) );
no02f01 g02233 ( .a(n6021), .b(n6019), .o(n6022_1) );
in01f01 g02234 ( .a(n6022_1), .o(n6023) );
no02f01 g02235 ( .a(n6023), .b(n6037), .o(n6024) );
no02f01 g02236 ( .a(n6024), .b(n6015), .o(n6025) );
in01f01 g02237 ( .a(n5766), .o(n6026) );
no02f01 g02238 ( .a(n5757), .b(n5743), .o(n6027_1) );
ao12f01 g02239 ( .a(n5751), .b(n6027_1), .c(n6026), .o(n6028) );
in01f01 g02240 ( .a(n6028), .o(n6029) );
no02f01 g02241 ( .a(n5769_1), .b(n5765_1), .o(n6030) );
no02f01 g02242 ( .a(n6030), .b(n6029), .o(n6031) );
na02f01 g02243 ( .a(n6030), .b(n6029), .o(n6032_1) );
in01f01 g02244 ( .a(n6032_1), .o(n6033) );
no02f01 g02245 ( .a(n6033), .b(n6031), .o(n6034) );
in01f01 g02246 ( .a(n6034), .o(n6035) );
no02f01 g02247 ( .a(n6035), .b(n6037), .o(n6036) );
in01f01 g02248 ( .a(n6036), .o(n6037_1) );
no02f01 g02249 ( .a(n5766), .b(n5751), .o(n6038) );
no02f01 g02250 ( .a(n6038), .b(n6027_1), .o(n6039) );
na02f01 g02251 ( .a(n6038), .b(n6027_1), .o(n6040) );
in01f01 g02252 ( .a(n6040), .o(n6041) );
no02f01 g02253 ( .a(n6041), .b(n6039), .o(n6042_1) );
in01f01 g02254 ( .a(n6042_1), .o(n6043) );
no02f01 g02255 ( .a(n6043), .b(n6037), .o(n6044) );
in01f01 g02256 ( .a(n6044), .o(n6045) );
na04f01 g02257 ( .a(n6045), .b(n6037_1), .c(n6025), .d(n6008), .o(n6046) );
ao12f01 g02258 ( .a(n5873), .b(n6022_1), .c(n6013), .o(n6047_1) );
ao12f01 g02259 ( .a(n5873), .b(n6042_1), .c(n6034), .o(n6048) );
no02f01 g02260 ( .a(n6048), .b(n6047_1), .o(n6049) );
na02f01 g02261 ( .a(n6049), .b(n6046), .o(n6050) );
no02f01 g02262 ( .a(n5895), .b(n5889), .o(n6051_1) );
no02f01 g02263 ( .a(n6051_1), .b(n6037), .o(n6052) );
in01f01 g02264 ( .a(n6052), .o(n6053) );
ao12f01 g02265 ( .a(n5896), .b(n6053), .c(n6050), .o(n6054) );
na02f01 g02266 ( .a(n5883_1), .b(n6037), .o(n6055) );
in01f01 g02267 ( .a(n6055), .o(n6056_1) );
no02f01 g02268 ( .a(n6056_1), .b(n6054), .o(n6057) );
no02f01 g02269 ( .a(n6057), .b(n5884), .o(n6058) );
no02f01 g02270 ( .a(n5814_1), .b(n5877), .o(n6059) );
in01f01 g02271 ( .a(n6059), .o(n6060) );
no02f01 g02272 ( .a(n5815), .b(n5808), .o(n6061_1) );
in01f01 g02273 ( .a(n6061_1), .o(n6062) );
no03f01 g02274 ( .a(n6062), .b(n6060), .c(n5797), .o(n6063) );
no02f01 g02275 ( .a(n6060), .b(n5797), .o(n6064) );
no02f01 g02276 ( .a(n6061_1), .b(n6064), .o(n6065) );
no02f01 g02277 ( .a(n6065), .b(n6063), .o(n6066_1) );
in01f01 g02278 ( .a(n6066_1), .o(n6067) );
no02f01 g02279 ( .a(n6067), .b(n5873), .o(n6068) );
no02f01 g02280 ( .a(n6066_1), .b(n6037), .o(n6069) );
no02f01 g02281 ( .a(n6069), .b(n6068), .o(n6070) );
na02f01 g02282 ( .a(n6070), .b(n6058), .o(n6071_1) );
in01f01 g02283 ( .a(n6070), .o(n6072) );
oa12f01 g02284 ( .a(n6072), .b(n6057), .c(n5884), .o(n6073) );
na02f01 g02285 ( .a(n6073), .b(n6071_1), .o(n208) );
in01f01 g02286 ( .a(n_22641), .o(n6075) );
no02f01 g02287 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_13_), .b(n6075), .o(n6076_1) );
in01f01 g02288 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_7_), .o(n6077) );
in01f01 g02289 ( .a(delay_sub_ln23_unr17_stage6_stallmux_q_1_), .o(n6078) );
in01f01 g02290 ( .a(cordic_combinational_sub_ln23_0_unr20_z_0_), .o(n6079) );
in01f01 g02291 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_1_), .o(n6080) );
ao12f01 g02292 ( .a(delay_sub_ln23_unr17_stage6_stallmux_q_1_), .b(n6080), .c(n6079), .o(n6081_1) );
ao12f01 g02293 ( .a(n6081_1), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_1_), .c(cordic_combinational_sub_ln23_0_unr20_z_0_), .o(n6082) );
no02f01 g02294 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_2_), .b(n6078), .o(n6083) );
no02f01 g02295 ( .a(n6083), .b(n6082), .o(n6084) );
in01f01 g02296 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_3_), .o(n6085) );
in01f01 g02297 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_2_), .o(n6086_1) );
no02f01 g02298 ( .a(n6086_1), .b(delay_sub_ln23_unr17_stage6_stallmux_q_1_), .o(n6087) );
no02f01 g02299 ( .a(n6084), .b(n6087), .o(n6088) );
na02f01 g02300 ( .a(n6088), .b(n6085), .o(n6089) );
ao22f01 g02301 ( .a(n6089), .b(n6078), .c(n6084), .d(delay_sub_ln23_0_unr16_stage6_stallmux_q_3_), .o(n6090) );
no02f01 g02302 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_4_), .b(n6078), .o(n6091_1) );
no02f01 g02303 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_6_), .b(n6078), .o(n6092) );
no02f01 g02304 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_5_), .b(n6078), .o(n6093) );
no04f01 g02305 ( .a(n6093), .b(n6092), .c(n6091_1), .d(n6090), .o(n6094) );
na02f01 g02306 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_6_), .b(n6078), .o(n6095) );
in01f01 g02307 ( .a(n6095), .o(n6096_1) );
no02f01 g02308 ( .a(n6096_1), .b(n6094), .o(n6097) );
ao12f01 g02309 ( .a(delay_sub_ln23_unr17_stage6_stallmux_q_1_), .b(n6097), .c(n6077), .o(n6098) );
in01f01 g02310 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_5_), .o(n6099) );
in01f01 g02311 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_4_), .o(n6100) );
ao12f01 g02312 ( .a(delay_sub_ln23_unr17_stage6_stallmux_q_1_), .b(n6100), .c(n6099), .o(n6101_1) );
ao12f01 g02313 ( .a(n6101_1), .b(n6094), .c(delay_sub_ln23_0_unr16_stage6_stallmux_q_7_), .o(n6102) );
in01f01 g02314 ( .a(n6102), .o(n6103) );
no02f01 g02315 ( .a(n6103), .b(n6098), .o(n6104) );
no02f01 g02316 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_9_), .b(n6078), .o(n6105) );
no02f01 g02317 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_8_), .b(n6078), .o(n6106_1) );
no02f01 g02318 ( .a(n6106_1), .b(n6105), .o(n6107) );
in01f01 g02319 ( .a(n6107), .o(n6108) );
no02f01 g02320 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_11_), .b(n6078), .o(n6109) );
no02f01 g02321 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_10_), .b(n6078), .o(n6110) );
no03f01 g02322 ( .a(n6110), .b(n6109), .c(n6108), .o(n6111_1) );
in01f01 g02323 ( .a(n6111_1), .o(n6112) );
no02f01 g02324 ( .a(n6112), .b(n6104), .o(n6113) );
in01f01 g02325 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_9_), .o(n6114) );
in01f01 g02326 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_8_), .o(n6115) );
ao12f01 g02327 ( .a(delay_sub_ln23_unr17_stage6_stallmux_q_1_), .b(n6115), .c(n6114), .o(n6116_1) );
in01f01 g02328 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_11_), .o(n6117) );
in01f01 g02329 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_10_), .o(n6118) );
ao12f01 g02330 ( .a(delay_sub_ln23_unr17_stage6_stallmux_q_1_), .b(n6118), .c(n6117), .o(n6119) );
no02f01 g02331 ( .a(n6119), .b(n6116_1), .o(n6120) );
in01f01 g02332 ( .a(n6120), .o(n6121_1) );
no02f01 g02333 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_12_), .b(n6078), .o(n6122) );
in01f01 g02334 ( .a(n6122), .o(n6123) );
oa12f01 g02335 ( .a(n6123), .b(n6121_1), .c(n6113), .o(n6124) );
na02f01 g02336 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_12_), .b(n6078), .o(n6125_1) );
in01f01 g02337 ( .a(n6125_1), .o(n6126) );
in01f01 g02338 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_13_), .o(n6127) );
no02f01 g02339 ( .a(n6127), .b(n_22641), .o(n6128) );
no02f01 g02340 ( .a(n6128), .b(n6126), .o(n6129) );
ao12f01 g02341 ( .a(n6076_1), .b(n6129), .c(n6124), .o(n6130_1) );
in01f01 g02342 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_14_), .o(n6131) );
in01f01 g02343 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_15_), .o(n6132) );
ao12f01 g02344 ( .a(n_22641), .b(n6132), .c(n6131), .o(n6133) );
no02f01 g02345 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_14_), .b(n6075), .o(n6134) );
no02f01 g02346 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_15_), .b(n6075), .o(n6135_1) );
no02f01 g02347 ( .a(n6135_1), .b(n6134), .o(n6136) );
oa12f01 g02348 ( .a(n6136), .b(n6133), .c(n6130_1), .o(n6137) );
in01f01 g02349 ( .a(n6137), .o(n6138) );
no02f01 g02350 ( .a(n6075), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_17_), .o(n6139) );
no02f01 g02351 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_16_), .b(n6075), .o(n6140_1) );
no02f01 g02352 ( .a(n6140_1), .b(n6139), .o(n6141) );
no02f01 g02353 ( .a(n6075), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_19_), .o(n6142) );
no02f01 g02354 ( .a(n6075), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_18_), .o(n6143) );
no02f01 g02355 ( .a(n6143), .b(n6142), .o(n6144) );
na02f01 g02356 ( .a(n6144), .b(n6141), .o(n6145_1) );
in01f01 g02357 ( .a(n6145_1), .o(n6146) );
no02f01 g02358 ( .a(n6075), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_20_), .o(n6147) );
no02f01 g02359 ( .a(n6075), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_21_), .o(n6148) );
no02f01 g02360 ( .a(n6148), .b(n6147), .o(n6149_1) );
no02f01 g02361 ( .a(n6075), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_22_), .o(n6150) );
no02f01 g02362 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_23_), .b(n6075), .o(n6151) );
no02f01 g02363 ( .a(n6151), .b(n6150), .o(n6152) );
na03f01 g02364 ( .a(n6152), .b(n6149_1), .c(n6146), .o(n6153) );
in01f01 g02365 ( .a(n6153), .o(n6154_1) );
no02f01 g02366 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_25_), .b(n6075), .o(n6155) );
no02f01 g02367 ( .a(n6075), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_27_), .o(n6156) );
no02f01 g02368 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_24_), .b(n6075), .o(n6157) );
no02f01 g02369 ( .a(n6075), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_26_), .o(n6158) );
no04f01 g02370 ( .a(n6158), .b(n6157), .c(n6156), .d(n6155), .o(n6159_1) );
na02f01 g02371 ( .a(n6159_1), .b(n6154_1), .o(n6160) );
in01f01 g02372 ( .a(n6160), .o(n6161) );
no02f01 g02373 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_28_), .b(n6075), .o(n6162) );
in01f01 g02374 ( .a(n6162), .o(n6163_1) );
na03f01 g02375 ( .a(n6163_1), .b(n6161), .c(n6138), .o(n6164) );
no02f01 g02376 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_30_), .b(n6075), .o(n6165) );
no02f01 g02377 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_29_), .b(n6075), .o(n6166) );
no02f01 g02378 ( .a(n6166), .b(n6165), .o(n6167) );
in01f01 g02379 ( .a(n6167), .o(n6168_1) );
in01f01 g02380 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_17_), .o(n6169) );
in01f01 g02381 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_16_), .o(n6170) );
ao12f01 g02382 ( .a(n_22641), .b(n6170), .c(n6169), .o(n6171) );
in01f01 g02383 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_19_), .o(n6172_1) );
in01f01 g02384 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_18_), .o(n6173) );
ao12f01 g02385 ( .a(n_22641), .b(n6173), .c(n6172_1), .o(n6174) );
no02f01 g02386 ( .a(n6174), .b(n6171), .o(n6175) );
in01f01 g02387 ( .a(n6175), .o(n6176) );
in01f01 g02388 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_21_), .o(n6177_1) );
in01f01 g02389 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_20_), .o(n6178) );
ao12f01 g02390 ( .a(n_22641), .b(n6178), .c(n6177_1), .o(n6179) );
no02f01 g02391 ( .a(n6179), .b(n6176), .o(n6180) );
in01f01 g02392 ( .a(n6180), .o(n6181) );
in01f01 g02393 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_22_), .o(n6182_1) );
in01f01 g02394 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_23_), .o(n6183) );
ao12f01 g02395 ( .a(n_22641), .b(n6183), .c(n6182_1), .o(n6184) );
no02f01 g02396 ( .a(n6184), .b(n6181), .o(n6185) );
in01f01 g02397 ( .a(n6185), .o(n6186) );
in01f01 g02398 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_25_), .o(n6187_1) );
in01f01 g02399 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_24_), .o(n6188) );
ao12f01 g02400 ( .a(n_22641), .b(n6188), .c(n6187_1), .o(n6189) );
no02f01 g02401 ( .a(n6189), .b(n6186), .o(n6190) );
in01f01 g02402 ( .a(n6190), .o(n6191) );
in01f01 g02403 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_26_), .o(n6192_1) );
in01f01 g02404 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_27_), .o(n6193) );
ao12f01 g02405 ( .a(n_22641), .b(n6193), .c(n6192_1), .o(n6194) );
no02f01 g02406 ( .a(n6194), .b(n6191), .o(n6195) );
in01f01 g02407 ( .a(n6195), .o(n6196) );
in01f01 g02408 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_29_), .o(n6197_1) );
in01f01 g02409 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_28_), .o(n6198) );
ao12f01 g02410 ( .a(n_22641), .b(n6198), .c(n6197_1), .o(n6199) );
no02f01 g02411 ( .a(n6199), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_30_), .o(n6200) );
no02f01 g02412 ( .a(n6200), .b(n_22641), .o(n6201) );
no02f01 g02413 ( .a(n6201), .b(n6196), .o(n6202_1) );
oa12f01 g02414 ( .a(n6202_1), .b(n6168_1), .c(n6164), .o(n6203) );
in01f01 g02415 ( .a(n6203), .o(n3633) );
no02f01 g02416 ( .a(n6080), .b(delay_sub_ln23_unr17_stage6_stallmux_q_1_), .o(n6205) );
no02f01 g02417 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_1_), .b(n6078), .o(n6206) );
no03f01 g02418 ( .a(n6206), .b(n6205), .c(cordic_combinational_sub_ln23_0_unr20_z_0_), .o(n6207_1) );
no02f01 g02419 ( .a(n6206), .b(n6205), .o(n6208) );
no02f01 g02420 ( .a(n6208), .b(n6079), .o(n6209) );
no02f01 g02421 ( .a(n6209), .b(n6207_1), .o(n6210) );
ao12f01 g02422 ( .a(n6203), .b(n6210), .c(cordic_combinational_sub_ln23_0_unr20_z_0_), .o(n6211) );
no02f01 g02423 ( .a(n6211), .b(n6207_1), .o(n6212_1) );
in01f01 g02424 ( .a(n6082), .o(n6213) );
no02f01 g02425 ( .a(n6083), .b(n6087), .o(n6214) );
in01f01 g02426 ( .a(n6214), .o(n6215) );
no02f01 g02427 ( .a(n6215), .b(n6213), .o(n6216) );
no02f01 g02428 ( .a(n6214), .b(n6082), .o(n6217_1) );
no02f01 g02429 ( .a(n6217_1), .b(n6216), .o(n6218) );
in01f01 g02430 ( .a(n6218), .o(n6219) );
no02f01 g02431 ( .a(n6219), .b(n3633), .o(n6220) );
no02f01 g02432 ( .a(n6220), .b(n6212_1), .o(n6221) );
no02f01 g02433 ( .a(n6085), .b(delay_sub_ln23_unr17_stage6_stallmux_q_1_), .o(n6222_1) );
no02f01 g02434 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_3_), .b(n6078), .o(n6223) );
no02f01 g02435 ( .a(n6223), .b(n6222_1), .o(n6224) );
no02f01 g02436 ( .a(n6224), .b(n6088), .o(n6225) );
na02f01 g02437 ( .a(n6224), .b(n6088), .o(n6226) );
in01f01 g02438 ( .a(n6226), .o(n6227_1) );
no02f01 g02439 ( .a(n6227_1), .b(n6225), .o(n6228) );
in01f01 g02440 ( .a(n6228), .o(n6229) );
no02f01 g02441 ( .a(n6218), .b(n6203), .o(n6230) );
no02f01 g02442 ( .a(n6230), .b(n6221), .o(n6231_1) );
na02f01 g02443 ( .a(n6228), .b(n6231_1), .o(n6232) );
ao22f01 g02444 ( .a(n6232), .b(n3633), .c(n6229), .d(n6221), .o(n6233) );
in01f01 g02445 ( .a(n6090), .o(n6234) );
no02f01 g02446 ( .a(n6100), .b(delay_sub_ln23_unr17_stage6_stallmux_q_1_), .o(n6235) );
no02f01 g02447 ( .a(n6235), .b(n6091_1), .o(n6236_1) );
in01f01 g02448 ( .a(n6236_1), .o(n6237) );
no02f01 g02449 ( .a(n6237), .b(n6234), .o(n6238) );
no02f01 g02450 ( .a(n6236_1), .b(n6090), .o(n6239) );
no02f01 g02451 ( .a(n6239), .b(n6238), .o(n6240) );
in01f01 g02452 ( .a(n6240), .o(n6241_1) );
no02f01 g02453 ( .a(n6241_1), .b(n3633), .o(n6242) );
in01f01 g02454 ( .a(n6093), .o(n6243) );
no02f01 g02455 ( .a(n6091_1), .b(n6090), .o(n6244) );
ao12f01 g02456 ( .a(n6101_1), .b(n6244), .c(n6243), .o(n6245) );
no02f01 g02457 ( .a(n6096_1), .b(n6092), .o(n6246_1) );
no02f01 g02458 ( .a(n6246_1), .b(n6245), .o(n6247) );
na02f01 g02459 ( .a(n6246_1), .b(n6245), .o(n6248) );
in01f01 g02460 ( .a(n6248), .o(n6249) );
no02f01 g02461 ( .a(n6249), .b(n6247), .o(n6250) );
in01f01 g02462 ( .a(n6250), .o(n6251_1) );
no02f01 g02463 ( .a(n6251_1), .b(n3633), .o(n6252) );
no02f01 g02464 ( .a(n6099), .b(delay_sub_ln23_unr17_stage6_stallmux_q_1_), .o(n6253) );
no02f01 g02465 ( .a(n6253), .b(n6093), .o(n6254) );
in01f01 g02466 ( .a(n6254), .o(n6255) );
no03f01 g02467 ( .a(n6255), .b(n6244), .c(n6235), .o(n6256_1) );
no02f01 g02468 ( .a(n6244), .b(n6235), .o(n6257) );
no02f01 g02469 ( .a(n6254), .b(n6257), .o(n6258) );
no02f01 g02470 ( .a(n6258), .b(n6256_1), .o(n6259) );
in01f01 g02471 ( .a(n6259), .o(n6260_1) );
no02f01 g02472 ( .a(n6260_1), .b(n3633), .o(n6261) );
no04f01 g02473 ( .a(n6261), .b(n6252), .c(n6242), .d(n6233), .o(n6262) );
no02f01 g02474 ( .a(n6250), .b(n6203), .o(n6263) );
in01f01 g02475 ( .a(n6097), .o(n6264) );
no02f01 g02476 ( .a(n6077), .b(delay_sub_ln23_unr17_stage6_stallmux_q_1_), .o(n6265_1) );
no02f01 g02477 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_7_), .b(n6078), .o(n6266) );
no02f01 g02478 ( .a(n6266), .b(n6265_1), .o(n6267) );
in01f01 g02479 ( .a(n6267), .o(n6268) );
no03f01 g02480 ( .a(n6268), .b(n6101_1), .c(n6264), .o(n6269) );
in01f01 g02481 ( .a(n6101_1), .o(n6270) );
ao12f01 g02482 ( .a(n6267), .b(n6270), .c(n6097), .o(n6271) );
no02f01 g02483 ( .a(n6271), .b(n6269), .o(n6272) );
in01f01 g02484 ( .a(n6272), .o(n6273) );
no02f01 g02485 ( .a(n6273), .b(n6263), .o(n6274) );
in01f01 g02486 ( .a(n6274), .o(n6275) );
oa12f01 g02487 ( .a(n3633), .b(n6275), .c(n6262), .o(n6276) );
ao12f01 g02488 ( .a(n6203), .b(n6259), .c(n6240), .o(n6277) );
ao12f01 g02489 ( .a(n6277), .b(n6273), .c(n6262), .o(n6278) );
na02f01 g02490 ( .a(n6278), .b(n6276), .o(n6279) );
no02f01 g02491 ( .a(n6115), .b(delay_sub_ln23_unr17_stage6_stallmux_q_1_), .o(n6280) );
no02f01 g02492 ( .a(n6280), .b(n6106_1), .o(n6281) );
in01f01 g02493 ( .a(n6281), .o(n6282) );
no03f01 g02494 ( .a(n6282), .b(n6103), .c(n6098), .o(n6283) );
no02f01 g02495 ( .a(n6281), .b(n6104), .o(n6284) );
no02f01 g02496 ( .a(n6284), .b(n6283), .o(n6285) );
in01f01 g02497 ( .a(n6285), .o(n6286) );
no02f01 g02498 ( .a(n6106_1), .b(n6104), .o(n6287) );
no02f01 g02499 ( .a(n6114), .b(delay_sub_ln23_unr17_stage6_stallmux_q_1_), .o(n6288) );
no02f01 g02500 ( .a(n6288), .b(n6105), .o(n6289) );
in01f01 g02501 ( .a(n6289), .o(n6290) );
no03f01 g02502 ( .a(n6290), .b(n6287), .c(n6280), .o(n6291) );
no02f01 g02503 ( .a(n6287), .b(n6280), .o(n6292) );
no02f01 g02504 ( .a(n6289), .b(n6292), .o(n6293) );
no02f01 g02505 ( .a(n6293), .b(n6291), .o(n6294) );
in01f01 g02506 ( .a(n6294), .o(n6295) );
ao12f01 g02507 ( .a(n3633), .b(n6295), .c(n6286), .o(n6296) );
in01f01 g02508 ( .a(n6296), .o(n6297) );
no02f01 g02509 ( .a(n6118), .b(delay_sub_ln23_unr17_stage6_stallmux_q_1_), .o(n6298) );
no03f01 g02510 ( .a(n6110), .b(n6108), .c(n6104), .o(n6299) );
no03f01 g02511 ( .a(n6299), .b(n6298), .c(n6116_1), .o(n6300) );
no02f01 g02512 ( .a(n6117), .b(delay_sub_ln23_unr17_stage6_stallmux_q_1_), .o(n6301) );
no02f01 g02513 ( .a(n6301), .b(n6109), .o(n6302) );
no02f01 g02514 ( .a(n6302), .b(n6300), .o(n6303) );
na02f01 g02515 ( .a(n6302), .b(n6300), .o(n6304) );
in01f01 g02516 ( .a(n6304), .o(n6305) );
no02f01 g02517 ( .a(n6305), .b(n6303), .o(n6306) );
in01f01 g02518 ( .a(n6306), .o(n6307) );
no02f01 g02519 ( .a(n6307), .b(n3633), .o(n6308) );
no02f01 g02520 ( .a(n6108), .b(n6104), .o(n6309) );
no02f01 g02521 ( .a(n6309), .b(n6116_1), .o(n6310) );
no02f01 g02522 ( .a(n6298), .b(n6110), .o(n6311) );
no02f01 g02523 ( .a(n6311), .b(n6310), .o(n6312) );
na02f01 g02524 ( .a(n6311), .b(n6310), .o(n6313) );
in01f01 g02525 ( .a(n6313), .o(n6314) );
no02f01 g02526 ( .a(n6314), .b(n6312), .o(n6315) );
in01f01 g02527 ( .a(n6315), .o(n6316) );
no02f01 g02528 ( .a(n6316), .b(n3633), .o(n6317) );
no02f01 g02529 ( .a(n6317), .b(n6308), .o(n6318) );
na03f01 g02530 ( .a(n6318), .b(n6297), .c(n6279), .o(n6319) );
ao12f01 g02531 ( .a(n6203), .b(n6294), .c(n6285), .o(n6320) );
ao12f01 g02532 ( .a(n6203), .b(n6315), .c(n6306), .o(n6321) );
no02f01 g02533 ( .a(n6321), .b(n6320), .o(n6322) );
no02f01 g02534 ( .a(n6121_1), .b(n6113), .o(n6323) );
no02f01 g02535 ( .a(n6126), .b(n6122), .o(n6324) );
no02f01 g02536 ( .a(n6324), .b(n6323), .o(n6325) );
na02f01 g02537 ( .a(n6324), .b(n6323), .o(n6326) );
in01f01 g02538 ( .a(n6326), .o(n6327) );
no02f01 g02539 ( .a(n6327), .b(n6325), .o(n6328) );
na02f01 g02540 ( .a(n6125_1), .b(n6120), .o(n6329) );
ao12f01 g02541 ( .a(n6329), .b(n6123), .c(n6113), .o(n6330) );
no02f01 g02542 ( .a(n6128), .b(n6076_1), .o(n6331) );
no02f01 g02543 ( .a(n6331), .b(n6330), .o(n6332) );
na02f01 g02544 ( .a(n6331), .b(n6330), .o(n6333) );
in01f01 g02545 ( .a(n6333), .o(n6334) );
no02f01 g02546 ( .a(n6334), .b(n6332), .o(n6335) );
no02f01 g02547 ( .a(n6335), .b(n6328), .o(n6336) );
no02f01 g02548 ( .a(n6336), .b(n6203), .o(n6337) );
ao12f01 g02549 ( .a(n6337), .b(n6322), .c(n6319), .o(n6338) );
no02f01 g02550 ( .a(n6131), .b(n_22641), .o(n6339) );
no02f01 g02551 ( .a(n6339), .b(n6130_1), .o(n6340) );
no02f01 g02552 ( .a(n6340), .b(n6134), .o(n6341) );
no02f01 g02553 ( .a(n6132), .b(n_22641), .o(n6342) );
no02f01 g02554 ( .a(n6342), .b(n6135_1), .o(n6343) );
in01f01 g02555 ( .a(n6343), .o(n6344) );
no02f01 g02556 ( .a(n6344), .b(n6341), .o(n6345) );
na02f01 g02557 ( .a(n6344), .b(n6341), .o(n6346) );
in01f01 g02558 ( .a(n6346), .o(n6347) );
no03f01 g02559 ( .a(n6347), .b(n6345), .c(n6203), .o(n6348) );
no02f01 g02560 ( .a(n6134), .b(n6339), .o(n6349) );
in01f01 g02561 ( .a(n6349), .o(n6350) );
no02f01 g02562 ( .a(n6350), .b(n6130_1), .o(n6351) );
in01f01 g02563 ( .a(n6130_1), .o(n6352) );
no02f01 g02564 ( .a(n6349), .b(n6352), .o(n6353) );
no02f01 g02565 ( .a(n6353), .b(n6351), .o(n6354) );
in01f01 g02566 ( .a(n6354), .o(n6355) );
no02f01 g02567 ( .a(n6355), .b(n6203), .o(n6356) );
no02f01 g02568 ( .a(n6356), .b(n6348), .o(n6357) );
ao12f01 g02569 ( .a(n3633), .b(n6335), .c(n6328), .o(n6358) );
no02f01 g02570 ( .a(n6347), .b(n6345), .o(n6359) );
ao12f01 g02571 ( .a(n3633), .b(n6354), .c(n6359), .o(n6360) );
no02f01 g02572 ( .a(n6360), .b(n6358), .o(n6361) );
in01f01 g02573 ( .a(n6361), .o(n6362) );
ao12f01 g02574 ( .a(n6362), .b(n6357), .c(n6338), .o(n6363) );
no02f01 g02575 ( .a(n6145_1), .b(n6137), .o(n6364) );
no02f01 g02576 ( .a(n_22641), .b(n6178), .o(n6365) );
no02f01 g02577 ( .a(n6365), .b(n6147), .o(n6366) );
in01f01 g02578 ( .a(n6366), .o(n6367) );
no03f01 g02579 ( .a(n6367), .b(n6364), .c(n6176), .o(n6368) );
in01f01 g02580 ( .a(n6364), .o(n6369) );
ao12f01 g02581 ( .a(n6366), .b(n6369), .c(n6175), .o(n6370) );
no03f01 g02582 ( .a(n6370), .b(n6368), .c(n6203), .o(n6371) );
no02f01 g02583 ( .a(n6369), .b(n6147), .o(n6372) );
no03f01 g02584 ( .a(n6372), .b(n6365), .c(n6176), .o(n6373) );
in01f01 g02585 ( .a(n6373), .o(n6374) );
no02f01 g02586 ( .a(n_22641), .b(n6177_1), .o(n6375) );
no02f01 g02587 ( .a(n6375), .b(n6148), .o(n6376) );
in01f01 g02588 ( .a(n6376), .o(n6377) );
no02f01 g02589 ( .a(n6377), .b(n6374), .o(n6378) );
no02f01 g02590 ( .a(n6376), .b(n6373), .o(n6379) );
no03f01 g02591 ( .a(n6379), .b(n6378), .c(n6203), .o(n6380) );
na02f01 g02592 ( .a(n6364), .b(n6149_1), .o(n6381) );
in01f01 g02593 ( .a(n6381), .o(n6382) );
no02f01 g02594 ( .a(n_22641), .b(n6182_1), .o(n6383) );
no02f01 g02595 ( .a(n6383), .b(n6150), .o(n6384) );
in01f01 g02596 ( .a(n6384), .o(n6385) );
no03f01 g02597 ( .a(n6385), .b(n6382), .c(n6181), .o(n6386) );
ao12f01 g02598 ( .a(n6384), .b(n6381), .c(n6180), .o(n6387) );
no03f01 g02599 ( .a(n6387), .b(n6386), .c(n6203), .o(n6388) );
no03f01 g02600 ( .a(n6388), .b(n6380), .c(n6371), .o(n6389) );
in01f01 g02601 ( .a(n6389), .o(n6390) );
no02f01 g02602 ( .a(n_22641), .b(n6173), .o(n6391) );
in01f01 g02603 ( .a(n6141), .o(n6392) );
no03f01 g02604 ( .a(n6143), .b(n6392), .c(n6137), .o(n6393) );
no03f01 g02605 ( .a(n6393), .b(n6391), .c(n6171), .o(n6394) );
in01f01 g02606 ( .a(n6394), .o(n6395) );
no02f01 g02607 ( .a(n_22641), .b(n6172_1), .o(n6396) );
no02f01 g02608 ( .a(n6396), .b(n6142), .o(n6397) );
in01f01 g02609 ( .a(n6397), .o(n6398) );
no02f01 g02610 ( .a(n6398), .b(n6395), .o(n6399) );
no02f01 g02611 ( .a(n6397), .b(n6394), .o(n6400) );
no03f01 g02612 ( .a(n6400), .b(n6399), .c(n6203), .o(n6401) );
no02f01 g02613 ( .a(n6170), .b(n_22641), .o(n6402) );
no02f01 g02614 ( .a(n6402), .b(n6140_1), .o(n6403) );
no02f01 g02615 ( .a(n6403), .b(n6137), .o(n6404) );
na02f01 g02616 ( .a(n6403), .b(n6137), .o(n6405) );
in01f01 g02617 ( .a(n6405), .o(n6406) );
no02f01 g02618 ( .a(n6406), .b(n6404), .o(n6407) );
in01f01 g02619 ( .a(n6407), .o(n6408) );
no02f01 g02620 ( .a(n6408), .b(n6203), .o(n6409) );
in01f01 g02621 ( .a(n6140_1), .o(n6410) );
ao12f01 g02622 ( .a(n6402), .b(n6410), .c(n6138), .o(n6411) );
in01f01 g02623 ( .a(n6411), .o(n6412) );
no02f01 g02624 ( .a(n_22641), .b(n6169), .o(n6413) );
no02f01 g02625 ( .a(n6413), .b(n6139), .o(n6414) );
in01f01 g02626 ( .a(n6414), .o(n6415) );
no02f01 g02627 ( .a(n6415), .b(n6412), .o(n6416) );
no02f01 g02628 ( .a(n6414), .b(n6411), .o(n6417) );
no03f01 g02629 ( .a(n6417), .b(n6416), .c(n6203), .o(n6418) );
no02f01 g02630 ( .a(n6418), .b(n6409), .o(n6419) );
in01f01 g02631 ( .a(n6419), .o(n6420) );
ao12f01 g02632 ( .a(n6171), .b(n6141), .c(n6138), .o(n6421) );
in01f01 g02633 ( .a(n6421), .o(n6422) );
no02f01 g02634 ( .a(n6391), .b(n6143), .o(n6423) );
in01f01 g02635 ( .a(n6423), .o(n6424) );
no02f01 g02636 ( .a(n6424), .b(n6422), .o(n6425) );
no02f01 g02637 ( .a(n6423), .b(n6421), .o(n6426) );
no03f01 g02638 ( .a(n6426), .b(n6425), .c(n6203), .o(n6427) );
no03f01 g02639 ( .a(n6427), .b(n6420), .c(n6401), .o(n6428) );
in01f01 g02640 ( .a(n6428), .o(n6429) );
no02f01 g02641 ( .a(n6381), .b(n6150), .o(n6430) );
no03f01 g02642 ( .a(n6430), .b(n6383), .c(n6181), .o(n6431) );
in01f01 g02643 ( .a(n6431), .o(n6432) );
no02f01 g02644 ( .a(n6183), .b(n_22641), .o(n6433) );
no02f01 g02645 ( .a(n6433), .b(n6151), .o(n6434) );
in01f01 g02646 ( .a(n6434), .o(n6435) );
no02f01 g02647 ( .a(n6435), .b(n6432), .o(n6436) );
no02f01 g02648 ( .a(n6434), .b(n6431), .o(n6437) );
no03f01 g02649 ( .a(n6437), .b(n6436), .c(n6203), .o(n6438) );
no03f01 g02650 ( .a(n6438), .b(n6429), .c(n6390), .o(n6439) );
in01f01 g02651 ( .a(n6439), .o(n6440) );
no02f01 g02652 ( .a(n6188), .b(n_22641), .o(n6441) );
no02f01 g02653 ( .a(n6153), .b(n6137), .o(n6442) );
in01f01 g02654 ( .a(n6442), .o(n6443) );
no02f01 g02655 ( .a(n6443), .b(n6157), .o(n6444) );
no03f01 g02656 ( .a(n6444), .b(n6441), .c(n6186), .o(n6445) );
no02f01 g02657 ( .a(n6187_1), .b(n_22641), .o(n6446) );
no02f01 g02658 ( .a(n6446), .b(n6155), .o(n6447) );
no02f01 g02659 ( .a(n6447), .b(n6445), .o(n6448) );
na02f01 g02660 ( .a(n6447), .b(n6445), .o(n6449) );
in01f01 g02661 ( .a(n6449), .o(n6450) );
no03f01 g02662 ( .a(n6450), .b(n6448), .c(n6203), .o(n6451) );
no02f01 g02663 ( .a(n6442), .b(n6186), .o(n6452) );
no02f01 g02664 ( .a(n6441), .b(n6157), .o(n6453) );
no02f01 g02665 ( .a(n6453), .b(n6452), .o(n6454) );
na02f01 g02666 ( .a(n6453), .b(n6452), .o(n6455) );
in01f01 g02667 ( .a(n6455), .o(n6456) );
no03f01 g02668 ( .a(n6456), .b(n6454), .c(n6203), .o(n6457) );
no02f01 g02669 ( .a(n6457), .b(n6451), .o(n6458) );
in01f01 g02670 ( .a(n6458), .o(n6459) );
no03f01 g02671 ( .a(n6443), .b(n6157), .c(n6155), .o(n6460) );
no02f01 g02672 ( .a(n_22641), .b(n6192_1), .o(n6461) );
no02f01 g02673 ( .a(n6461), .b(n6158), .o(n6462) );
in01f01 g02674 ( .a(n6462), .o(n6463) );
no03f01 g02675 ( .a(n6463), .b(n6460), .c(n6191), .o(n6464) );
no02f01 g02676 ( .a(n6460), .b(n6191), .o(n6465) );
no02f01 g02677 ( .a(n6462), .b(n6465), .o(n6466) );
no03f01 g02678 ( .a(n6466), .b(n6464), .c(n6203), .o(n6467) );
no04f01 g02679 ( .a(n6467), .b(n6459), .c(n6440), .d(n6363), .o(n6468) );
in01f01 g02680 ( .a(n6158), .o(n6469) );
na02f01 g02681 ( .a(n6460), .b(n6469), .o(n6470) );
in01f01 g02682 ( .a(n6470), .o(n6471) );
no03f01 g02683 ( .a(n6471), .b(n6461), .c(n6191), .o(n6472) );
in01f01 g02684 ( .a(n6472), .o(n6473) );
no02f01 g02685 ( .a(n_22641), .b(n6193), .o(n6474) );
no02f01 g02686 ( .a(n6474), .b(n6156), .o(n6475) );
in01f01 g02687 ( .a(n6475), .o(n6476) );
no02f01 g02688 ( .a(n6476), .b(n6473), .o(n6477) );
no02f01 g02689 ( .a(n6475), .b(n6472), .o(n6478) );
no02f01 g02690 ( .a(n6478), .b(n6477), .o(n6479) );
in01f01 g02691 ( .a(n6479), .o(n6480) );
no02f01 g02692 ( .a(n6480), .b(n6203), .o(n6481) );
in01f01 g02693 ( .a(n6481), .o(n6482) );
in01f01 g02694 ( .a(n6164), .o(n6483) );
no02f01 g02695 ( .a(n6198), .b(n_22641), .o(n6484) );
no03f01 g02696 ( .a(n6484), .b(n6196), .c(n6483), .o(n6485) );
no02f01 g02697 ( .a(n6197_1), .b(n_22641), .o(n6486) );
no02f01 g02698 ( .a(n6486), .b(n6166), .o(n6487) );
no02f01 g02699 ( .a(n6487), .b(n6485), .o(n6488) );
na02f01 g02700 ( .a(n6487), .b(n6485), .o(n6489) );
in01f01 g02701 ( .a(n6489), .o(n6490) );
no02f01 g02702 ( .a(n6490), .b(n6488), .o(n6491) );
in01f01 g02703 ( .a(n6491), .o(n6492) );
oa12f01 g02704 ( .a(n6195), .b(n6160), .c(n6137), .o(n6493) );
no02f01 g02705 ( .a(n6484), .b(n6162), .o(n6494) );
in01f01 g02706 ( .a(n6494), .o(n6495) );
no02f01 g02707 ( .a(n6495), .b(n6493), .o(n6496) );
na02f01 g02708 ( .a(n6495), .b(n6493), .o(n6497) );
in01f01 g02709 ( .a(n6497), .o(n6498) );
no02f01 g02710 ( .a(n6498), .b(n6496), .o(n6499) );
in01f01 g02711 ( .a(n6499), .o(n6500) );
ao12f01 g02712 ( .a(n6203), .b(n6500), .c(n6492), .o(n6501) );
in01f01 g02713 ( .a(n6501), .o(n6502) );
no02f01 g02714 ( .a(n6199), .b(n6196), .o(n6503) );
oa12f01 g02715 ( .a(n6503), .b(n6166), .c(n6164), .o(n6504) );
in01f01 g02716 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_30_), .o(n6505) );
no02f01 g02717 ( .a(n6505), .b(n_22641), .o(n6506) );
no02f01 g02718 ( .a(n6506), .b(n6165), .o(n6507) );
in01f01 g02719 ( .a(n6507), .o(n6508) );
no02f01 g02720 ( .a(n6508), .b(n6504), .o(n6509) );
na02f01 g02721 ( .a(n6508), .b(n6504), .o(n6510) );
in01f01 g02722 ( .a(n6510), .o(n6511) );
no02f01 g02723 ( .a(n6511), .b(n6509), .o(n6512) );
in01f01 g02724 ( .a(n6512), .o(n6513) );
no02f01 g02725 ( .a(n6513), .b(n6203), .o(n6514) );
in01f01 g02726 ( .a(n6514), .o(n6515) );
na04f01 g02727 ( .a(n6515), .b(n6502), .c(n6482), .d(n6468), .o(n6516) );
no02f01 g02728 ( .a(n6417), .b(n6416), .o(n6517) );
ao12f01 g02729 ( .a(n3633), .b(n6517), .c(n6407), .o(n6518) );
no02f01 g02730 ( .a(n6400), .b(n6399), .o(n6519) );
no02f01 g02731 ( .a(n6426), .b(n6425), .o(n6520) );
ao12f01 g02732 ( .a(n3633), .b(n6520), .c(n6519), .o(n6521) );
no02f01 g02733 ( .a(n6521), .b(n6518), .o(n6522) );
in01f01 g02734 ( .a(n6522), .o(n6523) );
no02f01 g02735 ( .a(n6370), .b(n6368), .o(n6524) );
no02f01 g02736 ( .a(n6379), .b(n6378), .o(n6525) );
ao12f01 g02737 ( .a(n3633), .b(n6525), .c(n6524), .o(n6526) );
no02f01 g02738 ( .a(n6526), .b(n6523), .o(n6527) );
in01f01 g02739 ( .a(n6527), .o(n6528) );
no02f01 g02740 ( .a(n6387), .b(n6386), .o(n6529) );
no02f01 g02741 ( .a(n6437), .b(n6436), .o(n6530) );
ao12f01 g02742 ( .a(n3633), .b(n6530), .c(n6529), .o(n6531) );
no02f01 g02743 ( .a(n6531), .b(n6528), .o(n6532) );
in01f01 g02744 ( .a(n6532), .o(n6533) );
no02f01 g02745 ( .a(n6450), .b(n6448), .o(n6534) );
no02f01 g02746 ( .a(n6456), .b(n6454), .o(n6535) );
ao12f01 g02747 ( .a(n3633), .b(n6535), .c(n6534), .o(n6536) );
no02f01 g02748 ( .a(n6536), .b(n6533), .o(n6537) );
in01f01 g02749 ( .a(n6537), .o(n6538) );
no02f01 g02750 ( .a(n6466), .b(n6464), .o(n6539) );
ao12f01 g02751 ( .a(n3633), .b(n6479), .c(n6539), .o(n6540) );
no02f01 g02752 ( .a(n6540), .b(n6538), .o(n6541) );
in01f01 g02753 ( .a(n6541), .o(n6542) );
ao12f01 g02754 ( .a(n3633), .b(n6499), .c(n6491), .o(n6543) );
no02f01 g02755 ( .a(n6543), .b(n6513), .o(n6544) );
no02f01 g02756 ( .a(n6544), .b(n3633), .o(n6545) );
no02f01 g02757 ( .a(n6545), .b(n6542), .o(n6546) );
na02f01 g02758 ( .a(n6546), .b(n6516), .o(n6547) );
no02f01 g02759 ( .a(n6285), .b(n6203), .o(n6548) );
no02f01 g02760 ( .a(n6286), .b(n3633), .o(n6549) );
no02f01 g02761 ( .a(n6549), .b(n6548), .o(n6550) );
in01f01 g02762 ( .a(n6550), .o(n6551) );
no02f01 g02763 ( .a(n6551), .b(n6279), .o(n6552) );
in01f01 g02764 ( .a(n6279), .o(n6553) );
no02f01 g02765 ( .a(n6550), .b(n6553), .o(n6554) );
no02f01 g02766 ( .a(n6554), .b(n6552), .o(n6555) );
in01f01 g02767 ( .a(n6549), .o(n6556) );
ao12f01 g02768 ( .a(n6548), .b(n6556), .c(n6279), .o(n6557) );
no02f01 g02769 ( .a(n6294), .b(n6203), .o(n6558) );
no02f01 g02770 ( .a(n6295), .b(n3633), .o(n6559) );
no02f01 g02771 ( .a(n6559), .b(n6558), .o(n6560) );
no02f01 g02772 ( .a(n6560), .b(n6557), .o(n6561) );
na02f01 g02773 ( .a(n6560), .b(n6557), .o(n6562) );
in01f01 g02774 ( .a(n6562), .o(n6563) );
no02f01 g02775 ( .a(n6563), .b(n6561), .o(n6564) );
ao12f01 g02776 ( .a(n6547), .b(n6564), .c(n6555), .o(n6565) );
in01f01 g02777 ( .a(n6547), .o(n4043) );
ao12f01 g02778 ( .a(n6320), .b(n6297), .c(n6279), .o(n6567) );
no02f01 g02779 ( .a(n6315), .b(n6203), .o(n6568) );
no02f01 g02780 ( .a(n6568), .b(n6317), .o(n6569) );
no02f01 g02781 ( .a(n6569), .b(n6567), .o(n6570) );
na02f01 g02782 ( .a(n6569), .b(n6567), .o(n6571) );
in01f01 g02783 ( .a(n6571), .o(n6572) );
no02f01 g02784 ( .a(n6572), .b(n6570), .o(n6573) );
no03f01 g02785 ( .a(n6317), .b(n6296), .c(n6553), .o(n6574) );
no03f01 g02786 ( .a(n6574), .b(n6568), .c(n6320), .o(n6575) );
no02f01 g02787 ( .a(n6306), .b(n6203), .o(n6576) );
no02f01 g02788 ( .a(n6576), .b(n6308), .o(n6577) );
no02f01 g02789 ( .a(n6577), .b(n6575), .o(n6578) );
na02f01 g02790 ( .a(n6577), .b(n6575), .o(n6579) );
in01f01 g02791 ( .a(n6579), .o(n6580) );
no02f01 g02792 ( .a(n6580), .b(n6578), .o(n6581) );
ao12f01 g02793 ( .a(n6581), .b(n6573), .c(n4043), .o(n6582) );
in01f01 g02794 ( .a(n6581), .o(n6583) );
no02f01 g02795 ( .a(n6583), .b(n6547), .o(n6584) );
in01f01 g02796 ( .a(n6584), .o(n6585) );
oa12f01 g02797 ( .a(n6585), .b(n6582), .c(n6565), .o(n6586) );
in01f01 g02798 ( .a(n6586), .o(n6587) );
no02f01 g02799 ( .a(n6210), .b(n6203), .o(n6588) );
na02f01 g02800 ( .a(n6210), .b(n6203), .o(n6589) );
in01f01 g02801 ( .a(n6589), .o(n6590) );
no02f01 g02802 ( .a(n6590), .b(n6588), .o(n6591) );
in01f01 g02803 ( .a(n6591), .o(n6592) );
no02f01 g02804 ( .a(n6592), .b(n6079), .o(n6593) );
in01f01 g02805 ( .a(n6593), .o(n6594) );
oa12f01 g02806 ( .a(n4043), .b(n6592), .c(cordic_combinational_sub_ln23_0_unr20_z_0_), .o(n6595) );
no04f01 g02807 ( .a(n6230), .b(n6220), .c(n6211), .d(n6207_1), .o(n6596) );
no02f01 g02808 ( .a(n6230), .b(n6220), .o(n6597) );
no02f01 g02809 ( .a(n6597), .b(n6212_1), .o(n6598) );
no02f01 g02810 ( .a(n6598), .b(n6596), .o(n6599) );
na02f01 g02811 ( .a(n6599), .b(n6547), .o(n6600) );
in01f01 g02812 ( .a(n6600), .o(n6601) );
ao12f01 g02813 ( .a(n6601), .b(n6595), .c(n6594), .o(n6602) );
in01f01 g02814 ( .a(n6602), .o(n6603) );
no02f01 g02815 ( .a(n6228), .b(n6203), .o(n6604) );
no02f01 g02816 ( .a(n6229), .b(n3633), .o(n6605) );
no02f01 g02817 ( .a(n6605), .b(n6604), .o(n6606) );
no02f01 g02818 ( .a(n6606), .b(n6231_1), .o(n6607) );
na02f01 g02819 ( .a(n6606), .b(n6231_1), .o(n6608) );
in01f01 g02820 ( .a(n6608), .o(n6609) );
no02f01 g02821 ( .a(n6609), .b(n6607), .o(n6610) );
in01f01 g02822 ( .a(n6610), .o(n6611) );
no02f01 g02823 ( .a(n6599), .b(n6547), .o(n6612) );
no03f01 g02824 ( .a(n6612), .b(n6611), .c(n6602), .o(n6613) );
oa22f01 g02825 ( .a(n6613), .b(n6547), .c(n6610), .d(n6603), .o(n6614) );
no02f01 g02826 ( .a(n6240), .b(n6203), .o(n6615) );
no02f01 g02827 ( .a(n6615), .b(n6242), .o(n6616) );
no02f01 g02828 ( .a(n6616), .b(n6233), .o(n6617) );
na02f01 g02829 ( .a(n6616), .b(n6233), .o(n6618) );
in01f01 g02830 ( .a(n6618), .o(n6619) );
no02f01 g02831 ( .a(n6619), .b(n6617), .o(n6620) );
in01f01 g02832 ( .a(n6620), .o(n6621) );
no02f01 g02833 ( .a(n6242), .b(n6233), .o(n6622) );
no02f01 g02834 ( .a(n6615), .b(n6622), .o(n6623) );
no02f01 g02835 ( .a(n6259), .b(n6203), .o(n6624) );
no02f01 g02836 ( .a(n6624), .b(n6261), .o(n6625) );
no02f01 g02837 ( .a(n6625), .b(n6623), .o(n6626) );
na02f01 g02838 ( .a(n6625), .b(n6623), .o(n6627) );
in01f01 g02839 ( .a(n6627), .o(n6628) );
no02f01 g02840 ( .a(n6628), .b(n6626), .o(n6629) );
in01f01 g02841 ( .a(n6629), .o(n6630) );
ao12f01 g02842 ( .a(n4043), .b(n6630), .c(n6621), .o(n6631) );
in01f01 g02843 ( .a(n6631), .o(n6632) );
no02f01 g02844 ( .a(n6277), .b(n6263), .o(n6633) );
in01f01 g02845 ( .a(n6633), .o(n6634) );
no02f01 g02846 ( .a(n6273), .b(n3633), .o(n6635) );
no02f01 g02847 ( .a(n6272), .b(n6203), .o(n6636) );
no02f01 g02848 ( .a(n6636), .b(n6635), .o(n6637) );
in01f01 g02849 ( .a(n6637), .o(n6638) );
no03f01 g02850 ( .a(n6638), .b(n6634), .c(n6262), .o(n6639) );
no02f01 g02851 ( .a(n6634), .b(n6262), .o(n6640) );
no02f01 g02852 ( .a(n6637), .b(n6640), .o(n6641) );
no02f01 g02853 ( .a(n6641), .b(n6639), .o(n6642) );
in01f01 g02854 ( .a(n6642), .o(n6643) );
no02f01 g02855 ( .a(n6643), .b(n4043), .o(n6644) );
in01f01 g02856 ( .a(n6644), .o(n6645) );
in01f01 g02857 ( .a(n6261), .o(n6646) );
ao12f01 g02858 ( .a(n6277), .b(n6646), .c(n6622), .o(n6647) );
in01f01 g02859 ( .a(n6647), .o(n6648) );
no02f01 g02860 ( .a(n6263), .b(n6252), .o(n6649) );
in01f01 g02861 ( .a(n6649), .o(n6650) );
no02f01 g02862 ( .a(n6650), .b(n6648), .o(n6651) );
no02f01 g02863 ( .a(n6649), .b(n6647), .o(n6652) );
no02f01 g02864 ( .a(n6652), .b(n6651), .o(n6653) );
in01f01 g02865 ( .a(n6653), .o(n6654) );
no02f01 g02866 ( .a(n6654), .b(n4043), .o(n6655) );
in01f01 g02867 ( .a(n6655), .o(n6656) );
na04f01 g02868 ( .a(n6656), .b(n6645), .c(n6632), .d(n6614), .o(n6657) );
ao12f01 g02869 ( .a(n6547), .b(n6629), .c(n6620), .o(n6658) );
ao12f01 g02870 ( .a(n6547), .b(n6653), .c(n6642), .o(n6659) );
no02f01 g02871 ( .a(n6659), .b(n6658), .o(n6660) );
in01f01 g02872 ( .a(n6555), .o(n6661) );
in01f01 g02873 ( .a(n6564), .o(n6662) );
ao12f01 g02874 ( .a(n4043), .b(n6662), .c(n6661), .o(n6663) );
ao12f01 g02875 ( .a(n6663), .b(n6660), .c(n6657), .o(n6664) );
na02f01 g02876 ( .a(n6573), .b(n6547), .o(n6665) );
in01f01 g02877 ( .a(n6665), .o(n6666) );
no02f01 g02878 ( .a(n6666), .b(n6584), .o(n6667) );
ao12f01 g02879 ( .a(n6587), .b(n6667), .c(n6664), .o(n6668) );
na02f01 g02880 ( .a(n6322), .b(n6319), .o(n6669) );
no02f01 g02881 ( .a(n6328), .b(n3633), .o(n6670) );
na02f01 g02882 ( .a(n6328), .b(n3633), .o(n6671) );
in01f01 g02883 ( .a(n6671), .o(n6672) );
no02f01 g02884 ( .a(n6672), .b(n6670), .o(n6673) );
in01f01 g02885 ( .a(n6673), .o(n6674) );
no02f01 g02886 ( .a(n6674), .b(n6669), .o(n6675) );
ao12f01 g02887 ( .a(n6673), .b(n6322), .c(n6319), .o(n6676) );
no02f01 g02888 ( .a(n6676), .b(n6675), .o(n6677) );
in01f01 g02889 ( .a(n6677), .o(n6678) );
no02f01 g02890 ( .a(n6678), .b(n6547), .o(n6679) );
ao12f01 g02891 ( .a(n6670), .b(n6671), .c(n6669), .o(n6680) );
in01f01 g02892 ( .a(n6335), .o(n6681) );
no02f01 g02893 ( .a(n6681), .b(n6203), .o(n6682) );
no02f01 g02894 ( .a(n6335), .b(n3633), .o(n6683) );
no02f01 g02895 ( .a(n6683), .b(n6682), .o(n6684) );
no02f01 g02896 ( .a(n6684), .b(n6680), .o(n6685) );
na02f01 g02897 ( .a(n6684), .b(n6680), .o(n6686) );
in01f01 g02898 ( .a(n6686), .o(n6687) );
no02f01 g02899 ( .a(n6687), .b(n6685), .o(n6688) );
in01f01 g02900 ( .a(n6688), .o(n6689) );
no02f01 g02901 ( .a(n6689), .b(n6547), .o(n6690) );
no02f01 g02902 ( .a(n6690), .b(n6679), .o(n6691) );
in01f01 g02903 ( .a(n6691), .o(n6692) );
in01f01 g02904 ( .a(n6338), .o(n6693) );
in01f01 g02905 ( .a(n6358), .o(n6694) );
na02f01 g02906 ( .a(n6694), .b(n6693), .o(n6695) );
no02f01 g02907 ( .a(n6354), .b(n3633), .o(n6696) );
no02f01 g02908 ( .a(n6696), .b(n6356), .o(n6697) );
in01f01 g02909 ( .a(n6697), .o(n6698) );
na02f01 g02910 ( .a(n6698), .b(n6695), .o(n6699) );
in01f01 g02911 ( .a(n6699), .o(n6700) );
no02f01 g02912 ( .a(n6698), .b(n6695), .o(n6701) );
no02f01 g02913 ( .a(n6701), .b(n6700), .o(n6702) );
in01f01 g02914 ( .a(n6702), .o(n6703) );
no02f01 g02915 ( .a(n6703), .b(n6547), .o(n6704) );
no02f01 g02916 ( .a(n6696), .b(n6358), .o(n6705) );
oa12f01 g02917 ( .a(n6705), .b(n6356), .c(n6693), .o(n6706) );
no02f01 g02918 ( .a(n6359), .b(n3633), .o(n6707) );
no02f01 g02919 ( .a(n6707), .b(n6348), .o(n6708) );
in01f01 g02920 ( .a(n6708), .o(n6709) );
no02f01 g02921 ( .a(n6709), .b(n6706), .o(n6710) );
na02f01 g02922 ( .a(n6709), .b(n6706), .o(n6711) );
in01f01 g02923 ( .a(n6711), .o(n6712) );
no02f01 g02924 ( .a(n6712), .b(n6710), .o(n6713) );
in01f01 g02925 ( .a(n6713), .o(n6714) );
no02f01 g02926 ( .a(n6714), .b(n6547), .o(n6715) );
no04f01 g02927 ( .a(n6715), .b(n6704), .c(n6692), .d(n6668), .o(n6716) );
ao12f01 g02928 ( .a(n4043), .b(n6713), .c(n6702), .o(n6717) );
ao12f01 g02929 ( .a(n4043), .b(n6688), .c(n6677), .o(n6718) );
no02f01 g02930 ( .a(n6718), .b(n6717), .o(n6719) );
in01f01 g02931 ( .a(n6719), .o(n6720) );
in01f01 g02932 ( .a(n6363), .o(n6721) );
in01f01 g02933 ( .a(n6409), .o(n6722) );
no02f01 g02934 ( .a(n6407), .b(n3633), .o(n6723) );
ao12f01 g02935 ( .a(n6723), .b(n6722), .c(n6721), .o(n6724) );
in01f01 g02936 ( .a(n6724), .o(n6725) );
no02f01 g02937 ( .a(n6517), .b(n3633), .o(n6726) );
no02f01 g02938 ( .a(n6726), .b(n6418), .o(n6727) );
in01f01 g02939 ( .a(n6727), .o(n6728) );
no02f01 g02940 ( .a(n6728), .b(n6725), .o(n6729) );
no02f01 g02941 ( .a(n6727), .b(n6724), .o(n6730) );
no03f01 g02942 ( .a(n6730), .b(n6729), .c(n6547), .o(n6731) );
no02f01 g02943 ( .a(n6723), .b(n6409), .o(n6732) );
no02f01 g02944 ( .a(n6732), .b(n6363), .o(n6733) );
na02f01 g02945 ( .a(n6732), .b(n6363), .o(n6734) );
in01f01 g02946 ( .a(n6734), .o(n6735) );
no02f01 g02947 ( .a(n6735), .b(n6733), .o(n6736) );
in01f01 g02948 ( .a(n6736), .o(n6737) );
no02f01 g02949 ( .a(n6737), .b(n6547), .o(n6738) );
no02f01 g02950 ( .a(n6738), .b(n6731), .o(n6739) );
oa12f01 g02951 ( .a(n6739), .b(n6720), .c(n6716), .o(n6740) );
no02f01 g02952 ( .a(n6420), .b(n6363), .o(n6741) );
in01f01 g02953 ( .a(n6741), .o(n6742) );
no02f01 g02954 ( .a(n6520), .b(n3633), .o(n6743) );
no02f01 g02955 ( .a(n6743), .b(n6518), .o(n6744) );
oa12f01 g02956 ( .a(n6744), .b(n6742), .c(n6427), .o(n6745) );
in01f01 g02957 ( .a(n6745), .o(n6746) );
no02f01 g02958 ( .a(n6519), .b(n3633), .o(n6747) );
no02f01 g02959 ( .a(n6747), .b(n6401), .o(n6748) );
no02f01 g02960 ( .a(n6748), .b(n6746), .o(n6749) );
na02f01 g02961 ( .a(n6748), .b(n6746), .o(n6750) );
in01f01 g02962 ( .a(n6750), .o(n6751) );
no03f01 g02963 ( .a(n6751), .b(n6749), .c(n6547), .o(n6752) );
no02f01 g02964 ( .a(n6741), .b(n6518), .o(n6753) );
no02f01 g02965 ( .a(n6743), .b(n6427), .o(n6754) );
no02f01 g02966 ( .a(n6754), .b(n6753), .o(n6755) );
na02f01 g02967 ( .a(n6754), .b(n6753), .o(n6756) );
in01f01 g02968 ( .a(n6756), .o(n6757) );
no03f01 g02969 ( .a(n6757), .b(n6755), .c(n6547), .o(n6758) );
no02f01 g02970 ( .a(n6758), .b(n6752), .o(n6759) );
in01f01 g02971 ( .a(n6759), .o(n6760) );
no02f01 g02972 ( .a(n6751), .b(n6749), .o(n6761) );
no02f01 g02973 ( .a(n6757), .b(n6755), .o(n6762) );
ao12f01 g02974 ( .a(n4043), .b(n6762), .c(n6761), .o(n6763) );
no02f01 g02975 ( .a(n6730), .b(n6729), .o(n6764) );
ao12f01 g02976 ( .a(n4043), .b(n6736), .c(n6764), .o(n6765) );
no02f01 g02977 ( .a(n6765), .b(n6763), .o(n6766) );
oa12f01 g02978 ( .a(n6766), .b(n6760), .c(n6740), .o(n6767) );
no02f01 g02979 ( .a(n6429), .b(n6363), .o(n6768) );
no02f01 g02980 ( .a(n6524), .b(n3633), .o(n6769) );
no02f01 g02981 ( .a(n6769), .b(n6371), .o(n6770) );
in01f01 g02982 ( .a(n6770), .o(n6771) );
no03f01 g02983 ( .a(n6771), .b(n6768), .c(n6523), .o(n6772) );
in01f01 g02984 ( .a(n6768), .o(n6773) );
ao12f01 g02985 ( .a(n6770), .b(n6773), .c(n6522), .o(n6774) );
no02f01 g02986 ( .a(n6774), .b(n6772), .o(n6775) );
in01f01 g02987 ( .a(n6775), .o(n6776) );
no02f01 g02988 ( .a(n6776), .b(n6547), .o(n6777) );
no02f01 g02989 ( .a(n6769), .b(n6523), .o(n6778) );
oa12f01 g02990 ( .a(n6778), .b(n6773), .c(n6371), .o(n6779) );
in01f01 g02991 ( .a(n6779), .o(n6780) );
no02f01 g02992 ( .a(n6525), .b(n3633), .o(n6781) );
no02f01 g02993 ( .a(n6781), .b(n6380), .o(n6782) );
no02f01 g02994 ( .a(n6782), .b(n6780), .o(n6783) );
na02f01 g02995 ( .a(n6782), .b(n6780), .o(n6784) );
in01f01 g02996 ( .a(n6784), .o(n6785) );
no03f01 g02997 ( .a(n6785), .b(n6783), .c(n6547), .o(n6786) );
no02f01 g02998 ( .a(n6786), .b(n6777), .o(n6787) );
in01f01 g02999 ( .a(n6787), .o(n6788) );
no02f01 g03000 ( .a(n6529), .b(n3633), .o(n6789) );
no02f01 g03001 ( .a(n6789), .b(n6528), .o(n6790) );
oa12f01 g03002 ( .a(n6790), .b(n6773), .c(n6390), .o(n6791) );
no02f01 g03003 ( .a(n6530), .b(n3633), .o(n6792) );
no02f01 g03004 ( .a(n6792), .b(n6438), .o(n6793) );
in01f01 g03005 ( .a(n6793), .o(n6794) );
no02f01 g03006 ( .a(n6794), .b(n6791), .o(n6795) );
na02f01 g03007 ( .a(n6794), .b(n6791), .o(n6796) );
in01f01 g03008 ( .a(n6796), .o(n6797) );
no03f01 g03009 ( .a(n6797), .b(n6795), .c(n6547), .o(n6798) );
no02f01 g03010 ( .a(n6380), .b(n6371), .o(n6799) );
ao12f01 g03011 ( .a(n6528), .b(n6768), .c(n6799), .o(n6800) );
no02f01 g03012 ( .a(n6789), .b(n6388), .o(n6801) );
no02f01 g03013 ( .a(n6801), .b(n6800), .o(n6802) );
na02f01 g03014 ( .a(n6801), .b(n6800), .o(n6803) );
in01f01 g03015 ( .a(n6803), .o(n6804) );
no03f01 g03016 ( .a(n6804), .b(n6802), .c(n6547), .o(n6805) );
no03f01 g03017 ( .a(n6805), .b(n6798), .c(n6788), .o(n6806) );
no02f01 g03018 ( .a(n6797), .b(n6795), .o(n6807) );
no02f01 g03019 ( .a(n6804), .b(n6802), .o(n6808) );
ao12f01 g03020 ( .a(n4043), .b(n6808), .c(n6807), .o(n6809) );
no02f01 g03021 ( .a(n6785), .b(n6783), .o(n6810) );
ao12f01 g03022 ( .a(n4043), .b(n6810), .c(n6775), .o(n6811) );
no02f01 g03023 ( .a(n6811), .b(n6809), .o(n6812) );
in01f01 g03024 ( .a(n6812), .o(n6813) );
ao12f01 g03025 ( .a(n6813), .b(n6806), .c(n6767), .o(n6814) );
no02f01 g03026 ( .a(n6440), .b(n6363), .o(n6815) );
in01f01 g03027 ( .a(n6815), .o(n6816) );
no02f01 g03028 ( .a(n6535), .b(n3633), .o(n6817) );
no02f01 g03029 ( .a(n6817), .b(n6533), .o(n6818) );
oa12f01 g03030 ( .a(n6818), .b(n6457), .c(n6816), .o(n6819) );
no02f01 g03031 ( .a(n6534), .b(n3633), .o(n6820) );
no02f01 g03032 ( .a(n6820), .b(n6451), .o(n6821) );
in01f01 g03033 ( .a(n6821), .o(n6822) );
no02f01 g03034 ( .a(n6822), .b(n6819), .o(n6823) );
na02f01 g03035 ( .a(n6822), .b(n6819), .o(n6824) );
in01f01 g03036 ( .a(n6824), .o(n6825) );
no03f01 g03037 ( .a(n6825), .b(n6823), .c(n6547), .o(n6826) );
no02f01 g03038 ( .a(n6533), .b(n6815), .o(n6827) );
no02f01 g03039 ( .a(n6817), .b(n6457), .o(n6828) );
no02f01 g03040 ( .a(n6828), .b(n6827), .o(n6829) );
na02f01 g03041 ( .a(n6828), .b(n6827), .o(n6830) );
in01f01 g03042 ( .a(n6830), .o(n6831) );
no02f01 g03043 ( .a(n6831), .b(n6829), .o(n6832) );
in01f01 g03044 ( .a(n6832), .o(n6833) );
no02f01 g03045 ( .a(n6833), .b(n6547), .o(n6834) );
no02f01 g03046 ( .a(n6834), .b(n6826), .o(n6835) );
in01f01 g03047 ( .a(n6835), .o(n6836) );
ao12f01 g03048 ( .a(n6538), .b(n6458), .c(n6815), .o(n6837) );
in01f01 g03049 ( .a(n6837), .o(n6838) );
no02f01 g03050 ( .a(n6539), .b(n3633), .o(n6839) );
no02f01 g03051 ( .a(n6839), .b(n6467), .o(n6840) );
in01f01 g03052 ( .a(n6840), .o(n6841) );
no02f01 g03053 ( .a(n6841), .b(n6838), .o(n6842) );
no02f01 g03054 ( .a(n6840), .b(n6837), .o(n6843) );
no03f01 g03055 ( .a(n6843), .b(n6842), .c(n6547), .o(n6844) );
no02f01 g03056 ( .a(n6839), .b(n6538), .o(n6845) );
in01f01 g03057 ( .a(n6845), .o(n6846) );
no02f01 g03058 ( .a(n6479), .b(n3633), .o(n6847) );
no02f01 g03059 ( .a(n6847), .b(n6481), .o(n6848) );
in01f01 g03060 ( .a(n6848), .o(n6849) );
no03f01 g03061 ( .a(n6849), .b(n6846), .c(n6468), .o(n6850) );
no02f01 g03062 ( .a(n6846), .b(n6468), .o(n6851) );
no02f01 g03063 ( .a(n6848), .b(n6851), .o(n6852) );
no03f01 g03064 ( .a(n6852), .b(n6850), .c(n6547), .o(n6853) );
no02f01 g03065 ( .a(n6853), .b(n6844), .o(n6854) );
in01f01 g03066 ( .a(n6854), .o(n6855) );
no02f01 g03067 ( .a(n6500), .b(n6203), .o(n6856) );
no02f01 g03068 ( .a(n6499), .b(n3633), .o(n6857) );
na02f01 g03069 ( .a(n6482), .b(n6468), .o(n6858) );
na02f01 g03070 ( .a(n6541), .b(n6858), .o(n6859) );
no02f01 g03071 ( .a(n6859), .b(n6857), .o(n6860) );
no02f01 g03072 ( .a(n6860), .b(n6856), .o(n6861) );
in01f01 g03073 ( .a(n6861), .o(n6862) );
no02f01 g03074 ( .a(n6492), .b(n6203), .o(n6863) );
no02f01 g03075 ( .a(n6491), .b(n3633), .o(n6864) );
no02f01 g03076 ( .a(n6864), .b(n6863), .o(n6865) );
no02f01 g03077 ( .a(n6865), .b(n6862), .o(n6866) );
na02f01 g03078 ( .a(n6865), .b(n6862), .o(n6867) );
in01f01 g03079 ( .a(n6867), .o(n6868) );
no03f01 g03080 ( .a(n6868), .b(n6866), .c(n6547), .o(n6869) );
no02f01 g03081 ( .a(n6856), .b(n6857), .o(n6870) );
in01f01 g03082 ( .a(n6870), .o(n6871) );
no02f01 g03083 ( .a(n6871), .b(n6859), .o(n6872) );
ao12f01 g03084 ( .a(n6870), .b(n6541), .c(n6858), .o(n6873) );
no03f01 g03085 ( .a(n6873), .b(n6872), .c(n6547), .o(n6874) );
no02f01 g03086 ( .a(n6874), .b(n6869), .o(n6875) );
in01f01 g03087 ( .a(n6875), .o(n6876) );
no02f01 g03088 ( .a(n6543), .b(n6542), .o(n6877) );
oa12f01 g03089 ( .a(n6877), .b(n6501), .c(n6858), .o(n6878) );
no02f01 g03090 ( .a(n6512), .b(n3633), .o(n6879) );
no02f01 g03091 ( .a(n6879), .b(n6514), .o(n6880) );
in01f01 g03092 ( .a(n6880), .o(n6881) );
no02f01 g03093 ( .a(n6881), .b(n6878), .o(n6882) );
na02f01 g03094 ( .a(n6881), .b(n6878), .o(n6883) );
in01f01 g03095 ( .a(n6883), .o(n6884) );
no03f01 g03096 ( .a(n6884), .b(n6882), .c(n6547), .o(n6885) );
no02f01 g03097 ( .a(n6885), .b(n6876), .o(n6886) );
in01f01 g03098 ( .a(n6886), .o(n6887) );
no04f01 g03099 ( .a(n6887), .b(n6855), .c(n6836), .d(n6814), .o(n6888) );
no02f01 g03100 ( .a(n6825), .b(n6823), .o(n6889) );
ao12f01 g03101 ( .a(n4043), .b(n6832), .c(n6889), .o(n6890) );
no02f01 g03102 ( .a(n6843), .b(n6842), .o(n6891) );
no02f01 g03103 ( .a(n6852), .b(n6850), .o(n6892) );
ao12f01 g03104 ( .a(n4043), .b(n6892), .c(n6891), .o(n6893) );
no02f01 g03105 ( .a(n6893), .b(n6890), .o(n6894) );
in01f01 g03106 ( .a(n6894), .o(n6895) );
no02f01 g03107 ( .a(n6884), .b(n6882), .o(n6896) );
no02f01 g03108 ( .a(n6868), .b(n6866), .o(n6897) );
no02f01 g03109 ( .a(n6873), .b(n6872), .o(n6898) );
ao12f01 g03110 ( .a(n4043), .b(n6898), .c(n6897), .o(n6899) );
in01f01 g03111 ( .a(n6899), .o(n6900) );
ao12f01 g03112 ( .a(n4043), .b(n6900), .c(n6896), .o(n6901) );
no02f01 g03113 ( .a(n6901), .b(n6895), .o(n6902) );
in01f01 g03114 ( .a(n6902), .o(n6903) );
no02f01 g03115 ( .a(n6903), .b(n6888), .o(n5001) );
no02f01 g03116 ( .a(n6591), .b(cordic_combinational_sub_ln23_0_unr20_z_0_), .o(n6905) );
no02f01 g03117 ( .a(n6905), .b(n6593), .o(n6906) );
no02f01 g03118 ( .a(n6906), .b(n6547), .o(n6907) );
na02f01 g03119 ( .a(n6906), .b(n6547), .o(n6908) );
in01f01 g03120 ( .a(n6908), .o(n6909) );
no02f01 g03121 ( .a(n6909), .b(n6907), .o(n6910) );
in01f01 g03122 ( .a(n6910), .o(n6911) );
no02f01 g03123 ( .a(n6911), .b(cordic_combinational_sub_ln23_0_unr20_z_0_), .o(n6912) );
no02f01 g03124 ( .a(n6911), .b(n6079), .o(n6913) );
no03f01 g03125 ( .a(n6913), .b(n6903), .c(n6888), .o(n6914) );
na02f01 g03126 ( .a(n6595), .b(n6594), .o(n6915) );
in01f01 g03127 ( .a(n6915), .o(n6916) );
no02f01 g03128 ( .a(n6612), .b(n6601), .o(n6917) );
no02f01 g03129 ( .a(n6917), .b(n6916), .o(n6918) );
na02f01 g03130 ( .a(n6917), .b(n6916), .o(n6919) );
in01f01 g03131 ( .a(n6919), .o(n6920) );
no02f01 g03132 ( .a(n6920), .b(n6918), .o(n6921) );
in01f01 g03133 ( .a(n6921), .o(n6922) );
oa22f01 g03134 ( .a(n6922), .b(n5001), .c(n6914), .d(n6912), .o(n6923) );
in01f01 g03135 ( .a(n6923), .o(n6924) );
no02f01 g03136 ( .a(n6611), .b(n4043), .o(n6925) );
no02f01 g03137 ( .a(n6610), .b(n6547), .o(n6926) );
no02f01 g03138 ( .a(n6926), .b(n6925), .o(n6927) );
in01f01 g03139 ( .a(n6927), .o(n6928) );
no03f01 g03140 ( .a(n6928), .b(n6612), .c(n6602), .o(n6929) );
no02f01 g03141 ( .a(n6612), .b(n6602), .o(n6930) );
no02f01 g03142 ( .a(n6927), .b(n6930), .o(n6931) );
no02f01 g03143 ( .a(n6931), .b(n6929), .o(n6932) );
in01f01 g03144 ( .a(n6932), .o(n6933) );
in01f01 g03145 ( .a(n5001), .o(n6934) );
no02f01 g03146 ( .a(n6921), .b(n6934), .o(n6935) );
in01f01 g03147 ( .a(n6935), .o(n6936) );
na03f01 g03148 ( .a(n6936), .b(n6932), .c(n6923), .o(n6937) );
ao22f01 g03149 ( .a(n6937), .b(n5001), .c(n6933), .d(n6924), .o(n6938) );
in01f01 g03150 ( .a(n6614), .o(n6939) );
no02f01 g03151 ( .a(n6620), .b(n6547), .o(n6940) );
no02f01 g03152 ( .a(n6621), .b(n4043), .o(n6941) );
no02f01 g03153 ( .a(n6941), .b(n6940), .o(n6942) );
no02f01 g03154 ( .a(n6942), .b(n6939), .o(n6943) );
na02f01 g03155 ( .a(n6942), .b(n6939), .o(n6944) );
in01f01 g03156 ( .a(n6944), .o(n6945) );
no02f01 g03157 ( .a(n6945), .b(n6943), .o(n6946) );
in01f01 g03158 ( .a(n6946), .o(n6947) );
no02f01 g03159 ( .a(n6947), .b(n5001), .o(n6948) );
ao12f01 g03160 ( .a(n6658), .b(n6632), .c(n6614), .o(n6949) );
no02f01 g03161 ( .a(n6653), .b(n6547), .o(n6950) );
no02f01 g03162 ( .a(n6950), .b(n6655), .o(n6951) );
no02f01 g03163 ( .a(n6951), .b(n6949), .o(n6952) );
na02f01 g03164 ( .a(n6951), .b(n6949), .o(n6953) );
in01f01 g03165 ( .a(n6953), .o(n6954) );
no02f01 g03166 ( .a(n6954), .b(n6952), .o(n6955) );
na02f01 g03167 ( .a(n6955), .b(n6934), .o(n6956) );
in01f01 g03168 ( .a(n6956), .o(n6957) );
in01f01 g03169 ( .a(n6941), .o(n6958) );
ao12f01 g03170 ( .a(n6940), .b(n6958), .c(n6614), .o(n6959) );
in01f01 g03171 ( .a(n6959), .o(n6960) );
no02f01 g03172 ( .a(n6629), .b(n6547), .o(n6961) );
no02f01 g03173 ( .a(n6630), .b(n4043), .o(n6962) );
no02f01 g03174 ( .a(n6962), .b(n6961), .o(n6963) );
in01f01 g03175 ( .a(n6963), .o(n6964) );
no02f01 g03176 ( .a(n6964), .b(n6960), .o(n6965) );
no02f01 g03177 ( .a(n6963), .b(n6959), .o(n6966) );
no02f01 g03178 ( .a(n6966), .b(n6965), .o(n6967) );
in01f01 g03179 ( .a(n6967), .o(n6968) );
no02f01 g03180 ( .a(n6968), .b(n5001), .o(n6969) );
no02f01 g03181 ( .a(n6969), .b(n6957), .o(n6970) );
in01f01 g03182 ( .a(n6970), .o(n6971) );
na02f01 g03183 ( .a(n6632), .b(n6614), .o(n6972) );
no02f01 g03184 ( .a(n6950), .b(n6658), .o(n6973) );
oa12f01 g03185 ( .a(n6973), .b(n6655), .c(n6972), .o(n6974) );
no02f01 g03186 ( .a(n6642), .b(n6547), .o(n6975) );
no02f01 g03187 ( .a(n6975), .b(n6644), .o(n6976) );
in01f01 g03188 ( .a(n6976), .o(n6977) );
no02f01 g03189 ( .a(n6977), .b(n6974), .o(n6978) );
na02f01 g03190 ( .a(n6977), .b(n6974), .o(n6979) );
in01f01 g03191 ( .a(n6979), .o(n6980) );
no02f01 g03192 ( .a(n6980), .b(n6978), .o(n6981) );
in01f01 g03193 ( .a(n6981), .o(n6982) );
no02f01 g03194 ( .a(n6982), .b(n5001), .o(n6983) );
no04f01 g03195 ( .a(n6983), .b(n6971), .c(n6948), .d(n6938), .o(n6984) );
ao12f01 g03196 ( .a(n6934), .b(n6967), .c(n6946), .o(n6985) );
ao12f01 g03197 ( .a(n6934), .b(n6981), .c(n6955), .o(n6986) );
no02f01 g03198 ( .a(n6986), .b(n6985), .o(n6987) );
in01f01 g03199 ( .a(n6987), .o(n6988) );
no02f01 g03200 ( .a(n6988), .b(n6984), .o(n6989) );
in01f01 g03201 ( .a(n6989), .o(n6990) );
no02f01 g03202 ( .a(n6555), .b(n6547), .o(n6991) );
in01f01 g03203 ( .a(n6657), .o(n6992) );
in01f01 g03204 ( .a(n6660), .o(n6993) );
no02f01 g03205 ( .a(n6993), .b(n6992), .o(n6994) );
no02f01 g03206 ( .a(n6661), .b(n4043), .o(n6995) );
no02f01 g03207 ( .a(n6995), .b(n6994), .o(n6996) );
no02f01 g03208 ( .a(n6996), .b(n6991), .o(n6997) );
no02f01 g03209 ( .a(n6662), .b(n4043), .o(n6998) );
no02f01 g03210 ( .a(n6564), .b(n6547), .o(n6999) );
no02f01 g03211 ( .a(n6999), .b(n6998), .o(n7000) );
no02f01 g03212 ( .a(n7000), .b(n6997), .o(n7001) );
na02f01 g03213 ( .a(n7000), .b(n6997), .o(n7002) );
in01f01 g03214 ( .a(n7002), .o(n7003) );
no02f01 g03215 ( .a(n7003), .b(n7001), .o(n7004) );
in01f01 g03216 ( .a(n7004), .o(n7005) );
no02f01 g03217 ( .a(n7005), .b(n5001), .o(n7006) );
no02f01 g03218 ( .a(n6995), .b(n6991), .o(n7007) );
in01f01 g03219 ( .a(n7007), .o(n7008) );
no03f01 g03220 ( .a(n7008), .b(n6993), .c(n6992), .o(n7009) );
no02f01 g03221 ( .a(n7007), .b(n6994), .o(n7010) );
no02f01 g03222 ( .a(n7010), .b(n7009), .o(n7011) );
in01f01 g03223 ( .a(n7011), .o(n7012) );
no02f01 g03224 ( .a(n7012), .b(n5001), .o(n7013) );
no02f01 g03225 ( .a(n7013), .b(n7006), .o(n7014) );
ao12f01 g03226 ( .a(n6934), .b(n7011), .c(n7004), .o(n7015) );
ao12f01 g03227 ( .a(n7015), .b(n7014), .c(n6990), .o(n7016) );
no02f01 g03228 ( .a(n6573), .b(n6547), .o(n7017) );
no02f01 g03229 ( .a(n6666), .b(n7017), .o(n7018) );
in01f01 g03230 ( .a(n7018), .o(n7019) );
no03f01 g03231 ( .a(n7019), .b(n6664), .c(n6565), .o(n7020) );
no02f01 g03232 ( .a(n6664), .b(n6565), .o(n7021) );
no02f01 g03233 ( .a(n7018), .b(n7021), .o(n7022) );
no02f01 g03234 ( .a(n7022), .b(n7020), .o(n7023) );
in01f01 g03235 ( .a(n7023), .o(n7024) );
no02f01 g03236 ( .a(n7024), .b(n6934), .o(n7025) );
no02f01 g03237 ( .a(n7023), .b(n5001), .o(n7026) );
no02f01 g03238 ( .a(n7026), .b(n7025), .o(n7027) );
na02f01 g03239 ( .a(n7027), .b(n7016), .o(n7028) );
in01f01 g03240 ( .a(n7016), .o(n7029) );
in01f01 g03241 ( .a(n7027), .o(n7030) );
na02f01 g03242 ( .a(n7030), .b(n7029), .o(n7031) );
na02f01 g03243 ( .a(n7031), .b(n7028), .o(n213) );
no02f01 g03244 ( .a(n4792), .b(n4762), .o(n7033) );
na02f01 g03245 ( .a(n7033), .b(n4765), .o(n7034) );
ao12f01 g03246 ( .a(n3821_1), .b(n4793), .c(n4760), .o(n7035) );
no02f01 g03247 ( .a(n7035), .b(n4768), .o(n7036) );
in01f01 g03248 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_28_), .o(n7037) );
no02f01 g03249 ( .a(n3821_1), .b(n7037), .o(n7038) );
in01f01 g03250 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_29_), .o(n7039) );
no02f01 g03251 ( .a(n3821_1), .b(n7039), .o(n7040) );
no02f01 g03252 ( .a(n7040), .b(n7038), .o(n7041) );
na02f01 g03253 ( .a(n7041), .b(n7036), .o(n7042) );
in01f01 g03254 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_30_), .o(n7043) );
no02f01 g03255 ( .a(n3821_1), .b(n7043), .o(n7044) );
no02f01 g03256 ( .a(n7044), .b(n7042), .o(n7045) );
no02f01 g03257 ( .a(n3818), .b(delay_add_ln22_unr20_stage8_stallmux_q_28_), .o(n7046) );
no02f01 g03258 ( .a(n3818), .b(delay_add_ln22_unr20_stage8_stallmux_q_29_), .o(n7047) );
no02f01 g03259 ( .a(n3818), .b(delay_add_ln22_unr20_stage8_stallmux_q_30_), .o(n7048) );
no03f01 g03260 ( .a(n7048), .b(n7047), .c(n7046), .o(n7049) );
in01f01 g03261 ( .a(n7049), .o(n7050) );
ao12f01 g03262 ( .a(n7050), .b(n7045), .c(n7034), .o(n7051) );
in01f01 g03263 ( .a(n7051), .o(n7052) );
no02f01 g03264 ( .a(n3818), .b(delay_add_ln22_unr20_stage8_stallmux_q_31_), .o(n7053) );
na02f01 g03265 ( .a(n3818), .b(delay_add_ln22_unr20_stage8_stallmux_q_31_), .o(n7054) );
in01f01 g03266 ( .a(n7054), .o(n7055) );
no02f01 g03267 ( .a(n7055), .b(n7053), .o(n7056) );
no02f01 g03268 ( .a(n7056), .b(n7052), .o(n7057) );
na02f01 g03269 ( .a(n7056), .b(n7052), .o(n7058) );
in01f01 g03270 ( .a(n7058), .o(n7059) );
no02f01 g03271 ( .a(n7059), .b(n7057), .o(n7060) );
no02f01 g03272 ( .a(n7048), .b(n7044), .o(n7061) );
in01f01 g03273 ( .a(n7034), .o(n7062) );
no02f01 g03274 ( .a(n7047), .b(n7046), .o(n7063) );
ao12f01 g03275 ( .a(n7042), .b(n7063), .c(n7062), .o(n7064) );
no02f01 g03276 ( .a(n7064), .b(n7061), .o(n7065) );
na02f01 g03277 ( .a(n7064), .b(n7061), .o(n7066) );
in01f01 g03278 ( .a(n7066), .o(n7067) );
no02f01 g03279 ( .a(n7067), .b(n7065), .o(n7068) );
in01f01 g03280 ( .a(n7068), .o(n7069) );
ao12f01 g03281 ( .a(n4825_1), .b(n4774), .c(delay_sub_ln23_0_unr21_stage8_stallmux_q), .o(n7070) );
oa12f01 g03282 ( .a(n7070), .b(n4797), .c(n4249), .o(n7071) );
in01f01 g03283 ( .a(n7046), .o(n7072) );
in01f01 g03284 ( .a(n7038), .o(n7073) );
ao22f01 g03285 ( .a(n7072), .b(n7073), .c(n7036), .d(n7034), .o(n7074) );
na02f01 g03286 ( .a(n7073), .b(n7036), .o(n7075) );
no02f01 g03287 ( .a(n7075), .b(n7062), .o(n7076) );
ao12f01 g03288 ( .a(n7074), .b(n7076), .c(n7072), .o(n7077) );
in01f01 g03289 ( .a(n7077), .o(n7078) );
ao12f01 g03290 ( .a(n7071), .b(n7078), .c(delay_sub_ln23_0_unr21_stage8_stallmux_q), .o(n7079) );
no02f01 g03291 ( .a(n7047), .b(n7040), .o(n7080) );
in01f01 g03292 ( .a(n7080), .o(n7081) );
no02f01 g03293 ( .a(n7076), .b(n7046), .o(n7082) );
no02f01 g03294 ( .a(n7082), .b(n7081), .o(n7083) );
na02f01 g03295 ( .a(n7082), .b(n7081), .o(n7084) );
in01f01 g03296 ( .a(n7084), .o(n7085) );
no02f01 g03297 ( .a(n7085), .b(n7083), .o(n7086) );
oa12f01 g03298 ( .a(n7079), .b(n7086), .c(n4249), .o(n7087) );
ao12f01 g03299 ( .a(n7087), .b(n7069), .c(delay_sub_ln23_0_unr21_stage8_stallmux_q), .o(n7088) );
ao12f01 g03300 ( .a(n7088), .b(n7069), .c(n4249), .o(n7089) );
no02f01 g03301 ( .a(n7089), .b(n7060), .o(n7090) );
in01f01 g03302 ( .a(n7060), .o(n7091) );
oa12f01 g03303 ( .a(n4832), .b(n4773), .c(n4249), .o(n7092) );
ao12f01 g03304 ( .a(n7092), .b(n4798), .c(delay_sub_ln23_0_unr21_stage8_stallmux_q), .o(n7093) );
oa12f01 g03305 ( .a(n7093), .b(n7077), .c(n4249), .o(n7094) );
in01f01 g03306 ( .a(n7086), .o(n7095) );
ao12f01 g03307 ( .a(n7094), .b(n7095), .c(delay_sub_ln23_0_unr21_stage8_stallmux_q), .o(n7096) );
oa12f01 g03308 ( .a(n7096), .b(n7068), .c(n4249), .o(n7097) );
oa12f01 g03309 ( .a(n7097), .b(n7068), .c(delay_sub_ln23_0_unr21_stage8_stallmux_q), .o(n7098) );
no02f01 g03310 ( .a(n7098), .b(n7091), .o(n7099) );
no02f01 g03311 ( .a(n4146_1), .b(n4048_1), .o(n7100) );
in01f01 g03312 ( .a(n7100), .o(n7101) );
no02f01 g03313 ( .a(n7101), .b(n4144), .o(n7102) );
no02f01 g03314 ( .a(n7100), .b(n4143), .o(n7103) );
no02f01 g03315 ( .a(n7103), .b(n7102), .o(n7104) );
oa12f01 g03316 ( .a(n7104), .b(n7099), .c(n7090), .o(n7105) );
na02f01 g03317 ( .a(n7069), .b(n7096), .o(n7106) );
na02f01 g03318 ( .a(n7068), .b(n7087), .o(n7107) );
na02f01 g03319 ( .a(n7107), .b(n7106), .o(n7108) );
in01f01 g03320 ( .a(n4140), .o(n7109) );
no02f01 g03321 ( .a(n4141_1), .b(n4055), .o(n7110) );
in01f01 g03322 ( .a(n7110), .o(n7111) );
no02f01 g03323 ( .a(n7111), .b(n7109), .o(n7112) );
no02f01 g03324 ( .a(n7110), .b(n4140), .o(n7113) );
no02f01 g03325 ( .a(n7113), .b(n7112), .o(n7114) );
no02f01 g03326 ( .a(n7114), .b(n7108), .o(n7115) );
in01f01 g03327 ( .a(n7115), .o(n7116) );
na02f01 g03328 ( .a(n7095), .b(n7079), .o(n7117) );
na02f01 g03329 ( .a(n7086), .b(n7094), .o(n7118) );
na02f01 g03330 ( .a(n7118), .b(n7117), .o(n7119) );
in01f01 g03331 ( .a(n4139), .o(n7120) );
no02f01 g03332 ( .a(n7120), .b(n4065), .o(n7121) );
in01f01 g03333 ( .a(n7121), .o(n7122) );
no02f01 g03334 ( .a(n7122), .b(n4138), .o(n7123) );
no02f01 g03335 ( .a(n7121), .b(n4137), .o(n7124) );
no02f01 g03336 ( .a(n7124), .b(n7123), .o(n7125) );
no02f01 g03337 ( .a(n7125), .b(n7119), .o(n7126) );
no02f01 g03338 ( .a(n7078), .b(n7093), .o(n7127) );
no02f01 g03339 ( .a(n7077), .b(n7071), .o(n7128) );
na02f01 g03340 ( .a(n4136_1), .b(n4077), .o(n7129) );
no02f01 g03341 ( .a(n7129), .b(n4135), .o(n7130) );
na02f01 g03342 ( .a(n7129), .b(n4135), .o(n7131) );
in01f01 g03343 ( .a(n7131), .o(n7132) );
no02f01 g03344 ( .a(n7132), .b(n7130), .o(n7133) );
no03f01 g03345 ( .a(n7133), .b(n7128), .c(n7127), .o(n7134) );
in01f01 g03346 ( .a(n7134), .o(n7135) );
no02f01 g03347 ( .a(n7070), .b(n4798), .o(n7136) );
no02f01 g03348 ( .a(n7092), .b(n4797), .o(n7137) );
na02f01 g03349 ( .a(n4132), .b(n4130), .o(n7138) );
in01f01 g03350 ( .a(n7138), .o(n7139) );
in01f01 g03351 ( .a(n4131_1), .o(n7140) );
no02f01 g03352 ( .a(n7140), .b(n4085), .o(n7141) );
no02f01 g03353 ( .a(n7141), .b(n7139), .o(n7142) );
na02f01 g03354 ( .a(n7141), .b(n7139), .o(n7143) );
in01f01 g03355 ( .a(n7143), .o(n7144) );
no02f01 g03356 ( .a(n7144), .b(n7142), .o(n7145) );
no03f01 g03357 ( .a(n7145), .b(n7137), .c(n7136), .o(n7146) );
na03f01 g03358 ( .a(n4839_1), .b(n4833), .c(n4826), .o(n7147) );
oa12f01 g03359 ( .a(n7147), .b(n4886), .c(n4840), .o(n7148) );
oa12f01 g03360 ( .a(n7145), .b(n7137), .c(n7136), .o(n7149) );
ao12f01 g03361 ( .a(n7146), .b(n7149), .c(n7148), .o(n7150) );
no02f01 g03362 ( .a(n7128), .b(n7127), .o(n7151) );
in01f01 g03363 ( .a(n7133), .o(n7152) );
no02f01 g03364 ( .a(n7152), .b(n7151), .o(n7153) );
oa12f01 g03365 ( .a(n7135), .b(n7153), .c(n7150), .o(n7154) );
na02f01 g03366 ( .a(n7125), .b(n7119), .o(n7155) );
ao12f01 g03367 ( .a(n7126), .b(n7155), .c(n7154), .o(n7156) );
in01f01 g03368 ( .a(n7114), .o(n7157) );
ao12f01 g03369 ( .a(n7157), .b(n7107), .c(n7106), .o(n7158) );
oa12f01 g03370 ( .a(n7116), .b(n7158), .c(n7156), .o(n7159) );
no03f01 g03371 ( .a(n7104), .b(n7099), .c(n7090), .o(n7160) );
oa12f01 g03372 ( .a(n7105), .b(n7160), .c(n7159), .o(n7161) );
no02f01 g03373 ( .a(n7091), .b(delay_sub_ln23_0_unr21_stage8_stallmux_q), .o(n7162) );
ao12f01 g03374 ( .a(n4249), .b(n7097), .c(n7060), .o(n7163) );
no02f01 g03375 ( .a(n7163), .b(n7162), .o(n7164) );
in01f01 g03376 ( .a(n4159), .o(n7165) );
no02f01 g03377 ( .a(n4030), .b(n4158), .o(n7166) );
no02f01 g03378 ( .a(n7166), .b(n4032), .o(n7167) );
in01f01 g03379 ( .a(n7167), .o(n7168) );
no03f01 g03380 ( .a(n7168), .b(n7165), .c(n4157), .o(n7169) );
no02f01 g03381 ( .a(n7165), .b(n4157), .o(n7170) );
no02f01 g03382 ( .a(n7167), .b(n7170), .o(n7171) );
no02f01 g03383 ( .a(n7171), .b(n7169), .o(n7172) );
no02f01 g03384 ( .a(n4146_1), .b(n4145), .o(n7173) );
no02f01 g03385 ( .a(n7165), .b(n4154), .o(n7174) );
in01f01 g03386 ( .a(n7174), .o(n7175) );
no02f01 g03387 ( .a(n7175), .b(n7173), .o(n7176) );
na02f01 g03388 ( .a(n7175), .b(n7173), .o(n7177) );
in01f01 g03389 ( .a(n7177), .o(n7178) );
no02f01 g03390 ( .a(n7178), .b(n7176), .o(n7179) );
ao12f01 g03391 ( .a(n7164), .b(n7179), .c(n7172), .o(n7180) );
in01f01 g03392 ( .a(n7180), .o(n7181) );
na02f01 g03393 ( .a(n7172), .b(n7164), .o(n7182) );
na02f01 g03394 ( .a(n7179), .b(n7164), .o(n7183) );
na02f01 g03395 ( .a(n7183), .b(n7182), .o(n7184) );
ao12f01 g03396 ( .a(n7184), .b(n7181), .c(n7161), .o(n7185) );
no02f01 g03397 ( .a(n4030), .b(n4166_1), .o(n7186) );
no02f01 g03398 ( .a(n7186), .b(n4283), .o(n7187) );
no02f01 g03399 ( .a(n7187), .b(n4171_1), .o(n7188) );
in01f01 g03400 ( .a(n7188), .o(n7189) );
no02f01 g03401 ( .a(n4030), .b(n4165), .o(n7190) );
no02f01 g03402 ( .a(n7190), .b(n4170), .o(n7191) );
no02f01 g03403 ( .a(n7191), .b(n7189), .o(n7192) );
na02f01 g03404 ( .a(n7191), .b(n7189), .o(n7193) );
in01f01 g03405 ( .a(n7193), .o(n7194) );
no02f01 g03406 ( .a(n7194), .b(n7192), .o(n7195) );
na02f01 g03407 ( .a(n7195), .b(n7164), .o(n7196) );
in01f01 g03408 ( .a(n4283), .o(n7197) );
no02f01 g03409 ( .a(n7186), .b(n4171_1), .o(n7198) );
no02f01 g03410 ( .a(n7198), .b(n7197), .o(n7199) );
na02f01 g03411 ( .a(n7198), .b(n7197), .o(n7200) );
in01f01 g03412 ( .a(n7200), .o(n7201) );
no02f01 g03413 ( .a(n7201), .b(n7199), .o(n7202) );
na02f01 g03414 ( .a(n7202), .b(n7164), .o(n7203) );
na02f01 g03415 ( .a(n7203), .b(n7196), .o(n7204) );
in01f01 g03416 ( .a(n7164), .o(n7205) );
no02f01 g03417 ( .a(n4030), .b(n4162), .o(n7206) );
no03f01 g03418 ( .a(n4175), .b(n4173), .c(n7197), .o(n7207) );
no03f01 g03419 ( .a(n7207), .b(n4167), .c(n7206), .o(n7208) );
in01f01 g03420 ( .a(n7208), .o(n7209) );
no02f01 g03421 ( .a(n4030), .b(n4163), .o(n7210) );
no02f01 g03422 ( .a(n7210), .b(n4174), .o(n7211) );
in01f01 g03423 ( .a(n7211), .o(n7212) );
no02f01 g03424 ( .a(n7212), .b(n7209), .o(n7213) );
no02f01 g03425 ( .a(n7211), .b(n7208), .o(n7214) );
no02f01 g03426 ( .a(n7214), .b(n7213), .o(n7215) );
in01f01 g03427 ( .a(n7215), .o(n7216) );
no02f01 g03428 ( .a(n7216), .b(n7205), .o(n7217) );
oa12f01 g03429 ( .a(n4172), .b(n4167), .c(n4283), .o(n7218) );
in01f01 g03430 ( .a(n7218), .o(n7219) );
no02f01 g03431 ( .a(n4175), .b(n7206), .o(n7220) );
in01f01 g03432 ( .a(n7220), .o(n7221) );
no02f01 g03433 ( .a(n7221), .b(n7219), .o(n7222) );
no02f01 g03434 ( .a(n7220), .b(n7218), .o(n7223) );
no02f01 g03435 ( .a(n7223), .b(n7222), .o(n7224) );
in01f01 g03436 ( .a(n7224), .o(n7225) );
no02f01 g03437 ( .a(n7225), .b(n7205), .o(n7226) );
no03f01 g03438 ( .a(n7226), .b(n7217), .c(n7204), .o(n7227) );
ao12f01 g03439 ( .a(n7164), .b(n7224), .c(n7215), .o(n7228) );
ao12f01 g03440 ( .a(n7164), .b(n7202), .c(n7195), .o(n7229) );
no02f01 g03441 ( .a(n7229), .b(n7228), .o(n7230) );
in01f01 g03442 ( .a(n7230), .o(n7231) );
ao12f01 g03443 ( .a(n7231), .b(n7227), .c(n7185), .o(n7232) );
no02f01 g03444 ( .a(n4286), .b(n4285_1), .o(n7233) );
in01f01 g03445 ( .a(n7233), .o(n7234) );
no02f01 g03446 ( .a(n4031), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_16_), .o(n7235) );
no02f01 g03447 ( .a(n4030), .b(n4203), .o(n7236) );
no02f01 g03448 ( .a(n7236), .b(n7235), .o(n7237) );
no02f01 g03449 ( .a(n7237), .b(n7234), .o(n7238) );
na02f01 g03450 ( .a(n7237), .b(n7234), .o(n7239) );
in01f01 g03451 ( .a(n7239), .o(n7240) );
no02f01 g03452 ( .a(n7240), .b(n7238), .o(n7241) );
in01f01 g03453 ( .a(n7241), .o(n7242) );
in01f01 g03454 ( .a(n7235), .o(n7243) );
ao12f01 g03455 ( .a(n7236), .b(n7243), .c(n7233), .o(n7244) );
no02f01 g03456 ( .a(n4031), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_17_), .o(n7245) );
no02f01 g03457 ( .a(n4030), .b(n4202), .o(n7246) );
no02f01 g03458 ( .a(n7246), .b(n7245), .o(n7247) );
no02f01 g03459 ( .a(n7247), .b(n7244), .o(n7248) );
na02f01 g03460 ( .a(n7247), .b(n7244), .o(n7249) );
in01f01 g03461 ( .a(n7249), .o(n7250) );
no02f01 g03462 ( .a(n7250), .b(n7248), .o(n7251) );
in01f01 g03463 ( .a(n7251), .o(n7252) );
ao12f01 g03464 ( .a(n7205), .b(n7252), .c(n7242), .o(n7253) );
no02f01 g03465 ( .a(n4030), .b(n4200), .o(n7254) );
no03f01 g03466 ( .a(n4185), .b(n4181_1), .c(n7234), .o(n7255) );
no03f01 g03467 ( .a(n7255), .b(n4204), .c(n7254), .o(n7256) );
no02f01 g03468 ( .a(n4030), .b(n4199), .o(n7257) );
no02f01 g03469 ( .a(n7257), .b(n4182), .o(n7258) );
no02f01 g03470 ( .a(n7258), .b(n7256), .o(n7259) );
na02f01 g03471 ( .a(n7258), .b(n7256), .o(n7260) );
in01f01 g03472 ( .a(n7260), .o(n7261) );
no02f01 g03473 ( .a(n7261), .b(n7259), .o(n7262) );
in01f01 g03474 ( .a(n7262), .o(n7263) );
no02f01 g03475 ( .a(n7263), .b(n7205), .o(n7264) );
no02f01 g03476 ( .a(n4181_1), .b(n7234), .o(n7265) );
no02f01 g03477 ( .a(n7254), .b(n4185), .o(n7266) );
in01f01 g03478 ( .a(n7266), .o(n7267) );
no03f01 g03479 ( .a(n7267), .b(n7265), .c(n4204), .o(n7268) );
no02f01 g03480 ( .a(n7265), .b(n4204), .o(n7269) );
no02f01 g03481 ( .a(n7266), .b(n7269), .o(n7270) );
no02f01 g03482 ( .a(n7270), .b(n7268), .o(n7271) );
in01f01 g03483 ( .a(n7271), .o(n7272) );
no02f01 g03484 ( .a(n7272), .b(n7205), .o(n7273) );
no03f01 g03485 ( .a(n7273), .b(n7264), .c(n7253), .o(n7274) );
in01f01 g03486 ( .a(n7274), .o(n7275) );
no02f01 g03487 ( .a(n4030), .b(n4208), .o(n7276) );
no03f01 g03488 ( .a(n4288), .b(n4177), .c(n7234), .o(n7277) );
no03f01 g03489 ( .a(n7277), .b(n7276), .c(n4206_1), .o(n7278) );
in01f01 g03490 ( .a(n7278), .o(n7279) );
no02f01 g03491 ( .a(n4030), .b(n4207), .o(n7280) );
no02f01 g03492 ( .a(n7280), .b(n4178), .o(n7281) );
in01f01 g03493 ( .a(n7281), .o(n7282) );
no02f01 g03494 ( .a(n7282), .b(n7279), .o(n7283) );
no02f01 g03495 ( .a(n7281), .b(n7278), .o(n7284) );
no02f01 g03496 ( .a(n7284), .b(n7283), .o(n7285) );
na02f01 g03497 ( .a(n7285), .b(n7164), .o(n7286) );
in01f01 g03498 ( .a(n7286), .o(n7287) );
no02f01 g03499 ( .a(n4288), .b(n7234), .o(n7288) );
no02f01 g03500 ( .a(n7276), .b(n4177), .o(n7289) );
in01f01 g03501 ( .a(n7289), .o(n7290) );
no03f01 g03502 ( .a(n7290), .b(n7288), .c(n4206_1), .o(n7291) );
no02f01 g03503 ( .a(n7288), .b(n4206_1), .o(n7292) );
no02f01 g03504 ( .a(n7289), .b(n7292), .o(n7293) );
no02f01 g03505 ( .a(n7293), .b(n7291), .o(n7294) );
na02f01 g03506 ( .a(n7294), .b(n7164), .o(n7295) );
in01f01 g03507 ( .a(n7295), .o(n7296) );
no02f01 g03508 ( .a(n7296), .b(n7287), .o(n7297) );
in01f01 g03509 ( .a(n7297), .o(n7298) );
no02f01 g03510 ( .a(n7205), .b(n4301), .o(n7299) );
no02f01 g03511 ( .a(n7205), .b(n4498_1), .o(n7300) );
no03f01 g03512 ( .a(n7300), .b(n7299), .c(n7298), .o(n7301) );
in01f01 g03513 ( .a(n7301), .o(n7302) );
no02f01 g03514 ( .a(n7205), .b(n4459), .o(n7303) );
no02f01 g03515 ( .a(n7205), .b(n4322), .o(n7304) );
no02f01 g03516 ( .a(n7304), .b(n7303), .o(n7305) );
in01f01 g03517 ( .a(n7305), .o(n7306) );
no04f01 g03518 ( .a(n7306), .b(n7302), .c(n7275), .d(n7232), .o(n7307) );
ao12f01 g03519 ( .a(n7164), .b(n7251), .c(n7241), .o(n7308) );
ao12f01 g03520 ( .a(n7164), .b(n7271), .c(n7262), .o(n7309) );
no02f01 g03521 ( .a(n7309), .b(n7308), .o(n7310) );
in01f01 g03522 ( .a(n7310), .o(n7311) );
ao12f01 g03523 ( .a(n7164), .b(n7294), .c(n7285), .o(n7312) );
ao12f01 g03524 ( .a(n7164), .b(n4454), .c(n4450), .o(n7313) );
no02f01 g03525 ( .a(n7313), .b(n7312), .o(n7314) );
in01f01 g03526 ( .a(n7314), .o(n7315) );
ao12f01 g03527 ( .a(n7315), .b(n7311), .c(n7301), .o(n7316) );
in01f01 g03528 ( .a(n7316), .o(n7317) );
ao12f01 g03529 ( .a(n7164), .b(n4448_1), .c(n4313), .o(n7318) );
no03f01 g03530 ( .a(n7318), .b(n7317), .c(n7307), .o(n7319) );
no02f01 g03531 ( .a(n7164), .b(n4279), .o(n7320) );
no02f01 g03532 ( .a(n7205), .b(n4434_1), .o(n7321) );
no02f01 g03533 ( .a(n7321), .b(n7320), .o(n7322) );
na02f01 g03534 ( .a(n7322), .b(n7319), .o(n7323) );
in01f01 g03535 ( .a(n7323), .o(n7324) );
no02f01 g03536 ( .a(n7322), .b(n7319), .o(n7325) );
no02f01 g03537 ( .a(n7325), .b(n7324), .o(n7326) );
no02f01 g03538 ( .a(n7326), .b(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n7327) );
in01f01 g03539 ( .a(n7300), .o(n7328) );
no02f01 g03540 ( .a(n7164), .b(n4454), .o(n7329) );
no02f01 g03541 ( .a(n7329), .b(n7299), .o(n7330) );
in01f01 g03542 ( .a(n7330), .o(n7331) );
no02f01 g03543 ( .a(n7164), .b(n4450), .o(n7332) );
in01f01 g03544 ( .a(n7332), .o(n7333) );
na02f01 g03545 ( .a(n7098), .b(n7091), .o(n7334) );
na02f01 g03546 ( .a(n7089), .b(n7060), .o(n7335) );
in01f01 g03547 ( .a(n7104), .o(n7336) );
ao12f01 g03548 ( .a(n7336), .b(n7335), .c(n7334), .o(n7337) );
no02f01 g03549 ( .a(n7086), .b(n7094), .o(n7338) );
no02f01 g03550 ( .a(n7095), .b(n7079), .o(n7339) );
no02f01 g03551 ( .a(n7339), .b(n7338), .o(n7340) );
in01f01 g03552 ( .a(n7125), .o(n7341) );
na02f01 g03553 ( .a(n7341), .b(n7340), .o(n7342) );
in01f01 g03554 ( .a(n7146), .o(n7343) );
oa12f01 g03555 ( .a(n4838), .b(n4842), .c(n4841), .o(n7344) );
in01f01 g03556 ( .a(n4852), .o(n7345) );
oa12f01 g03557 ( .a(n7345), .b(n4917_1), .c(n4913), .o(n7346) );
ao12f01 g03558 ( .a(n4843_1), .b(n7346), .c(n7344), .o(n7347) );
na02f01 g03559 ( .a(n7092), .b(n4797), .o(n7348) );
na02f01 g03560 ( .a(n7070), .b(n4798), .o(n7349) );
in01f01 g03561 ( .a(n7145), .o(n7350) );
ao12f01 g03562 ( .a(n7350), .b(n7349), .c(n7348), .o(n7351) );
oa12f01 g03563 ( .a(n7343), .b(n7351), .c(n7347), .o(n7352) );
oa12f01 g03564 ( .a(n7133), .b(n7128), .c(n7127), .o(n7353) );
ao12f01 g03565 ( .a(n7134), .b(n7353), .c(n7352), .o(n7354) );
no02f01 g03566 ( .a(n7341), .b(n7340), .o(n7355) );
oa12f01 g03567 ( .a(n7342), .b(n7355), .c(n7354), .o(n7356) );
in01f01 g03568 ( .a(n7158), .o(n7357) );
ao12f01 g03569 ( .a(n7115), .b(n7357), .c(n7356), .o(n7358) );
na03f01 g03570 ( .a(n7336), .b(n7335), .c(n7334), .o(n7359) );
ao12f01 g03571 ( .a(n7337), .b(n7359), .c(n7358), .o(n7360) );
in01f01 g03572 ( .a(n7184), .o(n7361) );
oa12f01 g03573 ( .a(n7361), .b(n7180), .c(n7360), .o(n7362) );
in01f01 g03574 ( .a(n7227), .o(n7363) );
oa12f01 g03575 ( .a(n7230), .b(n7363), .c(n7362), .o(n7364) );
na03f01 g03576 ( .a(n7297), .b(n7274), .c(n7364), .o(n7365) );
no02f01 g03577 ( .a(n7312), .b(n7311), .o(n7366) );
na03f01 g03578 ( .a(n7366), .b(n7365), .c(n7333), .o(n7367) );
ao12f01 g03579 ( .a(n7331), .b(n7367), .c(n7328), .o(n7368) );
no03f01 g03580 ( .a(n7298), .b(n7275), .c(n7232), .o(n7369) );
in01f01 g03581 ( .a(n7366), .o(n7370) );
no03f01 g03582 ( .a(n7370), .b(n7369), .c(n7332), .o(n7371) );
no03f01 g03583 ( .a(n7371), .b(n7330), .c(n7300), .o(n7372) );
no02f01 g03584 ( .a(n7372), .b(n7368), .o(n7373) );
no02f01 g03585 ( .a(n7164), .b(n4313), .o(n7374) );
no02f01 g03586 ( .a(n7374), .b(n7303), .o(n7375) );
in01f01 g03587 ( .a(n7375), .o(n7376) );
na03f01 g03588 ( .a(n7301), .b(n7274), .c(n7364), .o(n7377) );
na02f01 g03589 ( .a(n7377), .b(n7316), .o(n7378) );
no02f01 g03590 ( .a(n7378), .b(n7376), .o(n7379) );
no03f01 g03591 ( .a(n7302), .b(n7275), .c(n7232), .o(n7380) );
no02f01 g03592 ( .a(n7380), .b(n7317), .o(n7381) );
no02f01 g03593 ( .a(n7381), .b(n7375), .o(n7382) );
no02f01 g03594 ( .a(n7382), .b(n7379), .o(n7383) );
ao12f01 g03595 ( .a(n3789), .b(n7383), .c(n7373), .o(n7384) );
in01f01 g03596 ( .a(n7374), .o(n7385) );
no02f01 g03597 ( .a(n7164), .b(n4448_1), .o(n7386) );
no02f01 g03598 ( .a(n7386), .b(n7304), .o(n7387) );
in01f01 g03599 ( .a(n7303), .o(n7388) );
oa12f01 g03600 ( .a(n7388), .b(n7380), .c(n7317), .o(n7389) );
na03f01 g03601 ( .a(n7389), .b(n7387), .c(n7385), .o(n7390) );
in01f01 g03602 ( .a(n7387), .o(n7391) );
ao12f01 g03603 ( .a(n7303), .b(n7377), .c(n7316), .o(n7392) );
oa12f01 g03604 ( .a(n7391), .b(n7392), .c(n7374), .o(n7393) );
ao12f01 g03605 ( .a(n3789), .b(n7393), .c(n7390), .o(n7394) );
no02f01 g03606 ( .a(n7394), .b(n7384), .o(n7395) );
in01f01 g03607 ( .a(n7325), .o(n7396) );
na02f01 g03608 ( .a(n7396), .b(n7323), .o(n7397) );
na02f01 g03609 ( .a(n7397), .b(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n7398) );
ao12f01 g03610 ( .a(n7327), .b(n7398), .c(n7395), .o(n7399) );
no02f01 g03611 ( .a(n7205), .b(n4373), .o(n7400) );
no02f01 g03612 ( .a(n7164), .b(n4274), .o(n7401) );
no02f01 g03613 ( .a(n7401), .b(n7400), .o(n7402) );
in01f01 g03614 ( .a(n7402), .o(n7403) );
in01f01 g03615 ( .a(n7320), .o(n7404) );
ao12f01 g03616 ( .a(n7321), .b(n7404), .c(n7319), .o(n7405) );
na02f01 g03617 ( .a(n7405), .b(n7403), .o(n7406) );
in01f01 g03618 ( .a(n7406), .o(n7407) );
no02f01 g03619 ( .a(n7405), .b(n7403), .o(n7408) );
no02f01 g03620 ( .a(n7408), .b(n7407), .o(n7409) );
no02f01 g03621 ( .a(n7409), .b(n3789), .o(n7410) );
no02f01 g03622 ( .a(n7410), .b(n7399), .o(n7411) );
no02f01 g03623 ( .a(n7409), .b(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n7412) );
no03f01 g03624 ( .a(n7400), .b(n7321), .c(n7306), .o(n7413) );
ao12f01 g03625 ( .a(n7164), .b(n4279), .c(n4274), .o(n7414) );
no02f01 g03626 ( .a(n7414), .b(n7318), .o(n7415) );
in01f01 g03627 ( .a(n7415), .o(n7416) );
ao12f01 g03628 ( .a(n7416), .b(n7413), .c(n7378), .o(n7417) );
no02f01 g03629 ( .a(n7205), .b(n4412), .o(n7418) );
no02f01 g03630 ( .a(n7164), .b(n4263), .o(n7419) );
no02f01 g03631 ( .a(n7419), .b(n7418), .o(n7420) );
no02f01 g03632 ( .a(n7420), .b(n7417), .o(n7421) );
na02f01 g03633 ( .a(n7420), .b(n7417), .o(n7422) );
in01f01 g03634 ( .a(n7422), .o(n7423) );
no02f01 g03635 ( .a(n7423), .b(n7421), .o(n7424) );
no02f01 g03636 ( .a(n7424), .b(n3789), .o(n7425) );
no02f01 g03637 ( .a(n7424), .b(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n7426) );
no02f01 g03638 ( .a(n7426), .b(n7425), .o(n7427) );
in01f01 g03639 ( .a(n7427), .o(n7428) );
oa12f01 g03640 ( .a(n7428), .b(n7412), .c(n7411), .o(n7429) );
no03f01 g03641 ( .a(n7428), .b(n7412), .c(n7411), .o(n7430) );
in01f01 g03642 ( .a(n7430), .o(n7431) );
no04f01 g03643 ( .a(n4673), .b(n4505), .c(n4441), .d(n4429_1), .o(n7432) );
ao22f01 g03644 ( .a(n4506), .b(n4430), .c(n4669), .d(n4653), .o(n7433) );
no02f01 g03645 ( .a(n7433), .b(n7432), .o(n7434) );
ao12f01 g03646 ( .a(n7434), .b(n7431), .c(n7429), .o(n7435) );
in01f01 g03647 ( .a(n7429), .o(n7436) );
in01f01 g03648 ( .a(n7434), .o(n7437) );
no03f01 g03649 ( .a(n7437), .b(n7430), .c(n7436), .o(n7438) );
no02f01 g03650 ( .a(n7412), .b(n7410), .o(n7439) );
na02f01 g03651 ( .a(n7439), .b(n7399), .o(n7440) );
na02f01 g03652 ( .a(n7397), .b(n3789), .o(n7441) );
oa12f01 g03653 ( .a(n7330), .b(n7371), .c(n7300), .o(n7442) );
na03f01 g03654 ( .a(n7367), .b(n7331), .c(n7328), .o(n7443) );
na02f01 g03655 ( .a(n7443), .b(n7442), .o(n7444) );
in01f01 g03656 ( .a(n7383), .o(n7445) );
oa12f01 g03657 ( .a(delay_sub_ln23_0_unr22_stage8_stallmux_q), .b(n7445), .c(n7444), .o(n7446) );
no03f01 g03658 ( .a(n7392), .b(n7391), .c(n7374), .o(n7447) );
ao12f01 g03659 ( .a(n7387), .b(n7389), .c(n7385), .o(n7448) );
oa12f01 g03660 ( .a(delay_sub_ln23_0_unr22_stage8_stallmux_q), .b(n7448), .c(n7447), .o(n7449) );
na02f01 g03661 ( .a(n7449), .b(n7446), .o(n7450) );
no02f01 g03662 ( .a(n7326), .b(n3789), .o(n7451) );
oa12f01 g03663 ( .a(n7441), .b(n7451), .c(n7450), .o(n7452) );
in01f01 g03664 ( .a(n7408), .o(n7453) );
na02f01 g03665 ( .a(n7453), .b(n7406), .o(n7454) );
na02f01 g03666 ( .a(n7454), .b(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n7455) );
na02f01 g03667 ( .a(n7454), .b(n3789), .o(n7456) );
na02f01 g03668 ( .a(n7456), .b(n7455), .o(n7457) );
na02f01 g03669 ( .a(n7457), .b(n7452), .o(n7458) );
no02f01 g03670 ( .a(n4668), .b(n4467), .o(n7459) );
no02f01 g03671 ( .a(n4445), .b(n4441), .o(n7460) );
no02f01 g03672 ( .a(n7460), .b(n7459), .o(n7461) );
na02f01 g03673 ( .a(n7460), .b(n7459), .o(n7462) );
in01f01 g03674 ( .a(n7462), .o(n7463) );
no02f01 g03675 ( .a(n7463), .b(n7461), .o(n7464) );
ao12f01 g03676 ( .a(n7464), .b(n7458), .c(n7440), .o(n7465) );
in01f01 g03677 ( .a(n7465), .o(n7466) );
no02f01 g03678 ( .a(n7451), .b(n7327), .o(n7467) );
na02f01 g03679 ( .a(n7467), .b(n7450), .o(n7468) );
na02f01 g03680 ( .a(n7398), .b(n7441), .o(n7469) );
na02f01 g03681 ( .a(n7469), .b(n7395), .o(n7470) );
no02f01 g03682 ( .a(n4502), .b(n4479), .o(n7471) );
no02f01 g03683 ( .a(n4667_1), .b(n4467), .o(n7472) );
no02f01 g03684 ( .a(n7472), .b(n7471), .o(n7473) );
na02f01 g03685 ( .a(n7472), .b(n7471), .o(n7474) );
in01f01 g03686 ( .a(n7474), .o(n7475) );
no02f01 g03687 ( .a(n7475), .b(n7473), .o(n7476) );
ao12f01 g03688 ( .a(n7476), .b(n7470), .c(n7468), .o(n7477) );
oa12f01 g03689 ( .a(n3789), .b(n7448), .c(n7447), .o(n7478) );
na02f01 g03690 ( .a(n7478), .b(n7449), .o(n7479) );
no02f01 g03691 ( .a(n7479), .b(n7446), .o(n7480) );
ao12f01 g03692 ( .a(delay_sub_ln23_0_unr22_stage8_stallmux_q), .b(n7393), .c(n7390), .o(n7481) );
no02f01 g03693 ( .a(n7481), .b(n7394), .o(n7482) );
no02f01 g03694 ( .a(n7482), .b(n7384), .o(n7483) );
no02f01 g03695 ( .a(n4658), .b(n4657_1), .o(n7484) );
no04f01 g03696 ( .a(n4662_1), .b(n4493_1), .c(n7484), .d(n4479), .o(n7485) );
in01f01 g03697 ( .a(n7484), .o(n7486) );
ao22f01 g03698 ( .a(n4501), .b(n4494), .c(n7486), .d(n4659), .o(n7487) );
no02f01 g03699 ( .a(n7487), .b(n7485), .o(n7488) );
in01f01 g03700 ( .a(n7488), .o(n7489) );
oa12f01 g03701 ( .a(n7489), .b(n7483), .c(n7480), .o(n7490) );
no03f01 g03702 ( .a(n7489), .b(n7483), .c(n7480), .o(n7491) );
no02f01 g03703 ( .a(n4500), .b(n4499), .o(n7492) );
no02f01 g03704 ( .a(n7492), .b(n4492), .o(n7493) );
na02f01 g03705 ( .a(n7492), .b(n4492), .o(n7494) );
in01f01 g03706 ( .a(n7494), .o(n7495) );
no03f01 g03707 ( .a(n7495), .b(n7493), .c(n4483_1), .o(n7496) );
in01f01 g03708 ( .a(n7493), .o(n7497) );
ao12f01 g03709 ( .a(n4484), .b(n7494), .c(n7497), .o(n7498) );
no02f01 g03710 ( .a(n7498), .b(n7496), .o(n7499) );
na03f01 g03711 ( .a(n7443), .b(n7442), .c(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n7500) );
na03f01 g03712 ( .a(n7443), .b(n7442), .c(n3789), .o(n7501) );
in01f01 g03713 ( .a(n4482), .o(n7502) );
no02f01 g03714 ( .a(n7502), .b(n4450), .o(n7503) );
no02f01 g03715 ( .a(n4482), .b(n4498_1), .o(n7504) );
no02f01 g03716 ( .a(n7504), .b(n7503), .o(n7505) );
in01f01 g03717 ( .a(n7505), .o(n7506) );
na03f01 g03718 ( .a(n7506), .b(n7501), .c(n7500), .o(n7507) );
no02f01 g03719 ( .a(n7507), .b(n7499), .o(n7508) );
na02f01 g03720 ( .a(n7507), .b(n7499), .o(n7509) );
oa12f01 g03721 ( .a(n7445), .b(n7373), .c(n3789), .o(n7510) );
na03f01 g03722 ( .a(n7383), .b(n7444), .c(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n7511) );
na02f01 g03723 ( .a(n7511), .b(n7510), .o(n7512) );
ao12f01 g03724 ( .a(n7508), .b(n7512), .c(n7509), .o(n7513) );
oa12f01 g03725 ( .a(n7490), .b(n7513), .c(n7491), .o(n7514) );
na03f01 g03726 ( .a(n7476), .b(n7470), .c(n7468), .o(n7515) );
ao12f01 g03727 ( .a(n7477), .b(n7515), .c(n7514), .o(n7516) );
no02f01 g03728 ( .a(n7457), .b(n7452), .o(n7517) );
no02f01 g03729 ( .a(n7439), .b(n7399), .o(n7518) );
in01f01 g03730 ( .a(n7464), .o(n7519) );
no03f01 g03731 ( .a(n7519), .b(n7518), .c(n7517), .o(n7520) );
oa12f01 g03732 ( .a(n7466), .b(n7520), .c(n7516), .o(n7521) );
oa12f01 g03733 ( .a(n7521), .b(n7438), .c(n7435), .o(n7522) );
oa12f01 g03734 ( .a(n7437), .b(n7430), .c(n7436), .o(n7523) );
na03f01 g03735 ( .a(n7434), .b(n7431), .c(n7429), .o(n7524) );
in01f01 g03736 ( .a(n7477), .o(n7525) );
na02f01 g03737 ( .a(n7482), .b(n7384), .o(n7526) );
na02f01 g03738 ( .a(n7479), .b(n7446), .o(n7527) );
ao12f01 g03739 ( .a(n7488), .b(n7527), .c(n7526), .o(n7528) );
na03f01 g03740 ( .a(n7488), .b(n7527), .c(n7526), .o(n7529) );
in01f01 g03741 ( .a(n7499), .o(n7530) );
no03f01 g03742 ( .a(n7372), .b(n7368), .c(n3789), .o(n7531) );
no03f01 g03743 ( .a(n7372), .b(n7368), .c(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n7532) );
no03f01 g03744 ( .a(n7505), .b(n7532), .c(n7531), .o(n7533) );
na02f01 g03745 ( .a(n7533), .b(n7530), .o(n7534) );
no02f01 g03746 ( .a(n7533), .b(n7530), .o(n7535) );
ao12f01 g03747 ( .a(n7383), .b(n7444), .c(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n7536) );
no03f01 g03748 ( .a(n7445), .b(n7373), .c(n3789), .o(n7537) );
no02f01 g03749 ( .a(n7537), .b(n7536), .o(n7538) );
oa12f01 g03750 ( .a(n7534), .b(n7538), .c(n7535), .o(n7539) );
ao12f01 g03751 ( .a(n7528), .b(n7539), .c(n7529), .o(n7540) );
no02f01 g03752 ( .a(n7469), .b(n7395), .o(n7541) );
no02f01 g03753 ( .a(n7467), .b(n7450), .o(n7542) );
in01f01 g03754 ( .a(n7476), .o(n7543) );
no03f01 g03755 ( .a(n7543), .b(n7542), .c(n7541), .o(n7544) );
oa12f01 g03756 ( .a(n7525), .b(n7544), .c(n7540), .o(n7545) );
na03f01 g03757 ( .a(n7464), .b(n7458), .c(n7440), .o(n7546) );
ao12f01 g03758 ( .a(n7465), .b(n7546), .c(n7545), .o(n7547) );
na03f01 g03759 ( .a(n7547), .b(n7524), .c(n7523), .o(n7548) );
na02f01 g03760 ( .a(n7548), .b(n7522), .o(n223) );
in01f01 g03761 ( .a(n_17093), .o(n7550) );
no02f01 g03762 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_17_), .b(n7550), .o(n7551) );
in01f01 g03763 ( .a(n7551), .o(n7552) );
in01f01 g03764 ( .a(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .o(n7553) );
in01f01 g03765 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_1_), .o(n7554) );
no02f01 g03766 ( .a(n7554), .b(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .o(n7555) );
na02f01 g03767 ( .a(n7554), .b(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .o(n7556) );
ao12f01 g03768 ( .a(n7555), .b(n7556), .c(cordic_combinational_sub_ln23_0_unr16_z_0_), .o(n7557) );
no02f01 g03769 ( .a(n7553), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_2_), .o(n7558) );
no02f01 g03770 ( .a(n7558), .b(n7557), .o(n7559) );
in01f01 g03771 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_3_), .o(n7560) );
na02f01 g03772 ( .a(n7553), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_2_), .o(n7561) );
in01f01 g03773 ( .a(n7561), .o(n7562) );
no02f01 g03774 ( .a(n7562), .b(n7559), .o(n7563) );
na02f01 g03775 ( .a(n7563), .b(n7560), .o(n7564) );
ao22f01 g03776 ( .a(n7564), .b(n7553), .c(n7559), .d(delay_sub_ln23_0_unr12_stage5_stallmux_q_3_), .o(n7565) );
no02f01 g03777 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_6_), .b(n7553), .o(n7566) );
ao12f01 g03778 ( .a(n7553), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_5_), .c(delay_sub_ln23_0_unr12_stage5_stallmux_q_4_), .o(n7567) );
no02f01 g03779 ( .a(n7567), .b(n7566), .o(n7568) );
in01f01 g03780 ( .a(n7568), .o(n7569) );
no02f01 g03781 ( .a(n7569), .b(n7565), .o(n7570) );
no02f01 g03782 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_7_), .b(n7553), .o(n7571) );
in01f01 g03783 ( .a(n7571), .o(n7572) );
in01f01 g03784 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_4_), .o(n7573) );
in01f01 g03785 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_5_), .o(n7574) );
ao12f01 g03786 ( .a(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .b(n7574), .c(n7573), .o(n7575) );
in01f01 g03787 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_7_), .o(n7576) );
in01f01 g03788 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_6_), .o(n7577) );
ao12f01 g03789 ( .a(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .b(n7577), .c(n7576), .o(n7578) );
no02f01 g03790 ( .a(n7578), .b(n7575), .o(n7579) );
in01f01 g03791 ( .a(n7579), .o(n7580) );
ao12f01 g03792 ( .a(n7580), .b(n7572), .c(n7570), .o(n7581) );
ao12f01 g03793 ( .a(n7553), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_9_), .c(delay_sub_ln23_0_unr12_stage5_stallmux_q_8_), .o(n7582) );
in01f01 g03794 ( .a(n7582), .o(n7583) );
no02f01 g03795 ( .a(n7553), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_11_), .o(n7584) );
no02f01 g03796 ( .a(n7553), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_10_), .o(n7585) );
no02f01 g03797 ( .a(n7585), .b(n7584), .o(n7586) );
na02f01 g03798 ( .a(n7586), .b(n7583), .o(n7587) );
no02f01 g03799 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_12_), .b(n7553), .o(n7588) );
no02f01 g03800 ( .a(n7553), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_13_), .o(n7589) );
no03f01 g03801 ( .a(n7589), .b(n7588), .c(n7587), .o(n7590) );
in01f01 g03802 ( .a(n7590), .o(n7591) );
no02f01 g03803 ( .a(n7591), .b(n7581), .o(n7592) );
no02f01 g03804 ( .a(n7553), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_15_), .o(n7593) );
no02f01 g03805 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_14_), .b(n7553), .o(n7594) );
no02f01 g03806 ( .a(n7594), .b(n7593), .o(n7595) );
in01f01 g03807 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_8_), .o(n7596) );
in01f01 g03808 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_9_), .o(n7597) );
ao12f01 g03809 ( .a(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .b(n7597), .c(n7596), .o(n7598) );
in01f01 g03810 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_10_), .o(n7599) );
in01f01 g03811 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_11_), .o(n7600) );
ao12f01 g03812 ( .a(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .b(n7600), .c(n7599), .o(n7601) );
no02f01 g03813 ( .a(n7601), .b(n7598), .o(n7602) );
in01f01 g03814 ( .a(n7602), .o(n7603) );
in01f01 g03815 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_13_), .o(n7604) );
in01f01 g03816 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_12_), .o(n7605) );
ao12f01 g03817 ( .a(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .b(n7605), .c(n7604), .o(n7606) );
no02f01 g03818 ( .a(n7606), .b(n7603), .o(n7607) );
in01f01 g03819 ( .a(n7607), .o(n7608) );
in01f01 g03820 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_15_), .o(n7609) );
in01f01 g03821 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_14_), .o(n7610) );
ao12f01 g03822 ( .a(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .b(n7610), .c(n7609), .o(n7611) );
no02f01 g03823 ( .a(n7611), .b(n7608), .o(n7612) );
in01f01 g03824 ( .a(n7612), .o(n7613) );
ao12f01 g03825 ( .a(n7613), .b(n7595), .c(n7592), .o(n7614) );
no02f01 g03826 ( .a(n7553), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_16_), .o(n7615) );
no02f01 g03827 ( .a(n7615), .b(n7614), .o(n7616) );
na02f01 g03828 ( .a(n7616), .b(n7552), .o(n7617) );
no02f01 g03829 ( .a(n7550), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_19_), .o(n7618) );
no02f01 g03830 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_18_), .b(n7550), .o(n7619) );
no02f01 g03831 ( .a(n7619), .b(n7618), .o(n7620) );
in01f01 g03832 ( .a(n7620), .o(n7621) );
no02f01 g03833 ( .a(n7621), .b(n7617), .o(n7622) );
na02f01 g03834 ( .a(n7553), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_16_), .o(n7623) );
na02f01 g03835 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_17_), .b(n7550), .o(n7624) );
ao12f01 g03836 ( .a(n7551), .b(n7624), .c(n7623), .o(n7625) );
in01f01 g03837 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_19_), .o(n7626) );
in01f01 g03838 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_18_), .o(n7627) );
ao12f01 g03839 ( .a(n_17093), .b(n7627), .c(n7626), .o(n7628) );
oa12f01 g03840 ( .a(n7620), .b(n7628), .c(n7625), .o(n7629) );
in01f01 g03841 ( .a(n7629), .o(n7630) );
in01f01 g03842 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_21_), .o(n7631) );
in01f01 g03843 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_20_), .o(n7632) );
ao12f01 g03844 ( .a(n_17093), .b(n7632), .c(n7631), .o(n7633) );
in01f01 g03845 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_22_), .o(n7634) );
no02f01 g03846 ( .a(n7634), .b(n_17093), .o(n7635) );
no03f01 g03847 ( .a(n7635), .b(n7633), .c(n7630), .o(n7636) );
in01f01 g03848 ( .a(n7636), .o(n7637) );
in01f01 g03849 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_23_), .o(n7638) );
no02f01 g03850 ( .a(n7638), .b(n_17093), .o(n7639) );
no02f01 g03851 ( .a(n7639), .b(n7637), .o(n7640) );
in01f01 g03852 ( .a(n7640), .o(n7641) );
no02f01 g03853 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_21_), .b(n7550), .o(n7642) );
no02f01 g03854 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_20_), .b(n7550), .o(n7643) );
no02f01 g03855 ( .a(n7643), .b(n7642), .o(n7644) );
in01f01 g03856 ( .a(n7644), .o(n7645) );
no02f01 g03857 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_22_), .b(n7550), .o(n7646) );
no02f01 g03858 ( .a(n7646), .b(n7645), .o(n7647) );
in01f01 g03859 ( .a(n7647), .o(n7648) );
no02f01 g03860 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_23_), .b(n7550), .o(n7649) );
no02f01 g03861 ( .a(n7649), .b(n7648), .o(n7650) );
oa12f01 g03862 ( .a(n7650), .b(n7641), .c(n7622), .o(n7651) );
no02f01 g03863 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_25_), .b(n7550), .o(n7652) );
no02f01 g03864 ( .a(n7550), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_24_), .o(n7653) );
no02f01 g03865 ( .a(n7653), .b(n7652), .o(n7654) );
in01f01 g03866 ( .a(n7654), .o(n7655) );
no02f01 g03867 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_27_), .b(n7550), .o(n7656) );
no02f01 g03868 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_26_), .b(n7550), .o(n7657) );
no03f01 g03869 ( .a(n7657), .b(n7656), .c(n7655), .o(n7658) );
in01f01 g03870 ( .a(n7658), .o(n7659) );
no02f01 g03871 ( .a(n7659), .b(n7651), .o(n7660) );
no02f01 g03872 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_29_), .b(n7550), .o(n7661) );
no02f01 g03873 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_28_), .b(n7550), .o(n7662) );
no02f01 g03874 ( .a(n7662), .b(n7661), .o(n7663) );
in01f01 g03875 ( .a(n7663), .o(n7664) );
no02f01 g03876 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_30_), .b(n7550), .o(n7665) );
no02f01 g03877 ( .a(n7665), .b(n7664), .o(n7666) );
in01f01 g03878 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_29_), .o(n7667) );
in01f01 g03879 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_28_), .o(n7668) );
ao12f01 g03880 ( .a(n_17093), .b(n7668), .c(n7667), .o(n7669) );
oa12f01 g03881 ( .a(n7550), .b(n7669), .c(delay_sub_ln23_0_unr12_stage5_stallmux_q_30_), .o(n7670) );
na02f01 g03882 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_27_), .b(n7550), .o(n7671) );
in01f01 g03883 ( .a(n7671), .o(n7672) );
na02f01 g03884 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_26_), .b(n7550), .o(n7673) );
in01f01 g03885 ( .a(n7673), .o(n7674) );
in01f01 g03886 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_24_), .o(n7675) );
in01f01 g03887 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_25_), .o(n7676) );
ao12f01 g03888 ( .a(n_17093), .b(n7676), .c(n7675), .o(n7677) );
no02f01 g03889 ( .a(n7677), .b(n7674), .o(n7678) );
in01f01 g03890 ( .a(n7678), .o(n7679) );
no02f01 g03891 ( .a(n7679), .b(n7672), .o(n7680) );
na02f01 g03892 ( .a(n7680), .b(n7670), .o(n7681) );
ao12f01 g03893 ( .a(n7681), .b(n7666), .c(n7660), .o(n7682) );
no02f01 g03894 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_3_), .b(n7553), .o(n7683) );
no02f01 g03895 ( .a(n7560), .b(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .o(n7684) );
no02f01 g03896 ( .a(n7684), .b(n7683), .o(n7685) );
in01f01 g03897 ( .a(n7685), .o(n7686) );
no03f01 g03898 ( .a(n7686), .b(n7562), .c(n7559), .o(n7687) );
no02f01 g03899 ( .a(n7685), .b(n7563), .o(n7688) );
no02f01 g03900 ( .a(n7688), .b(n7687), .o(n7689) );
in01f01 g03901 ( .a(n7689), .o(n7690) );
no02f01 g03902 ( .a(n7690), .b(n7682), .o(n7691) );
in01f01 g03903 ( .a(n7557), .o(n7692) );
no02f01 g03904 ( .a(n7562), .b(n7558), .o(n7693) );
in01f01 g03905 ( .a(n7693), .o(n7694) );
no02f01 g03906 ( .a(n7694), .b(n7692), .o(n7695) );
no02f01 g03907 ( .a(n7693), .b(n7557), .o(n7696) );
no02f01 g03908 ( .a(n7696), .b(n7695), .o(n7697) );
in01f01 g03909 ( .a(n7697), .o(n7698) );
no02f01 g03910 ( .a(n7698), .b(n7682), .o(n7699) );
in01f01 g03911 ( .a(n7699), .o(n7700) );
in01f01 g03912 ( .a(n7556), .o(n7701) );
no03f01 g03913 ( .a(n7701), .b(n7555), .c(cordic_combinational_sub_ln23_0_unr16_z_0_), .o(n7702) );
in01f01 g03914 ( .a(cordic_combinational_sub_ln23_0_unr16_z_0_), .o(n7703) );
in01f01 g03915 ( .a(n7555), .o(n7704) );
ao12f01 g03916 ( .a(n7703), .b(n7556), .c(n7704), .o(n7705) );
no02f01 g03917 ( .a(n7705), .b(n7702), .o(n7706) );
in01f01 g03918 ( .a(n7706), .o(n7707) );
no02f01 g03919 ( .a(n7707), .b(n7682), .o(n7708) );
na02f01 g03920 ( .a(n7707), .b(n7682), .o(n7709) );
oa12f01 g03921 ( .a(n7709), .b(n7708), .c(cordic_combinational_sub_ln23_0_unr16_z_0_), .o(n7710) );
na02f01 g03922 ( .a(n7710), .b(n7700), .o(n7711) );
in01f01 g03923 ( .a(n7682), .o(n7712) );
no02f01 g03924 ( .a(n7697), .b(n7712), .o(n7713) );
no02f01 g03925 ( .a(n7689), .b(n7712), .o(n7714) );
no02f01 g03926 ( .a(n7714), .b(n7713), .o(n7715) );
oa12f01 g03927 ( .a(n7715), .b(n7711), .c(n7691), .o(n7716) );
in01f01 g03928 ( .a(n7565), .o(n7717) );
no02f01 g03929 ( .a(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .b(n7573), .o(n7718) );
no02f01 g03930 ( .a(n7553), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_4_), .o(n7719) );
no02f01 g03931 ( .a(n7719), .b(n7718), .o(n7720) );
in01f01 g03932 ( .a(n7720), .o(n7721) );
no02f01 g03933 ( .a(n7721), .b(n7717), .o(n7722) );
no02f01 g03934 ( .a(n7720), .b(n7565), .o(n7723) );
no02f01 g03935 ( .a(n7723), .b(n7722), .o(n7724) );
in01f01 g03936 ( .a(n7724), .o(n7725) );
no02f01 g03937 ( .a(n7725), .b(n7682), .o(n7726) );
in01f01 g03938 ( .a(n7726), .o(n7727) );
na02f01 g03939 ( .a(n7727), .b(n7716), .o(n7728) );
no02f01 g03940 ( .a(n7719), .b(n7565), .o(n7729) );
no02f01 g03941 ( .a(n7729), .b(n7718), .o(n7730) );
no02f01 g03942 ( .a(n7574), .b(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .o(n7731) );
no02f01 g03943 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_5_), .b(n7553), .o(n7732) );
no02f01 g03944 ( .a(n7732), .b(n7731), .o(n7733) );
no02f01 g03945 ( .a(n7733), .b(n7730), .o(n7734) );
na02f01 g03946 ( .a(n7733), .b(n7730), .o(n7735) );
in01f01 g03947 ( .a(n7735), .o(n7736) );
no02f01 g03948 ( .a(n7736), .b(n7734), .o(n7737) );
in01f01 g03949 ( .a(n7737), .o(n7738) );
no02f01 g03950 ( .a(n7738), .b(n7682), .o(n7739) );
in01f01 g03951 ( .a(n7575), .o(n7740) );
oa12f01 g03952 ( .a(n7740), .b(n7567), .c(n7565), .o(n7741) );
no02f01 g03953 ( .a(n7577), .b(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .o(n7742) );
no02f01 g03954 ( .a(n7742), .b(n7566), .o(n7743) );
in01f01 g03955 ( .a(n7743), .o(n7744) );
no02f01 g03956 ( .a(n7744), .b(n7741), .o(n7745) );
na02f01 g03957 ( .a(n7744), .b(n7741), .o(n7746) );
in01f01 g03958 ( .a(n7746), .o(n7747) );
no02f01 g03959 ( .a(n7747), .b(n7745), .o(n7748) );
in01f01 g03960 ( .a(n7748), .o(n7749) );
no02f01 g03961 ( .a(n7749), .b(n7682), .o(n7750) );
no02f01 g03962 ( .a(n7750), .b(n7739), .o(n7751) );
in01f01 g03963 ( .a(n7751), .o(n7752) );
no02f01 g03964 ( .a(n7752), .b(n7728), .o(n7753) );
no03f01 g03965 ( .a(n7742), .b(n7575), .c(n7570), .o(n7754) );
in01f01 g03966 ( .a(n7754), .o(n7755) );
no02f01 g03967 ( .a(n7576), .b(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .o(n7756) );
no02f01 g03968 ( .a(n7756), .b(n7571), .o(n7757) );
in01f01 g03969 ( .a(n7757), .o(n7758) );
no02f01 g03970 ( .a(n7758), .b(n7755), .o(n7759) );
no02f01 g03971 ( .a(n7757), .b(n7754), .o(n7760) );
no02f01 g03972 ( .a(n7760), .b(n7759), .o(n7761) );
in01f01 g03973 ( .a(n7761), .o(n7762) );
no02f01 g03974 ( .a(n7762), .b(n7682), .o(n7763) );
in01f01 g03975 ( .a(n7763), .o(n7764) );
na02f01 g03976 ( .a(n7764), .b(n7753), .o(n7765) );
no02f01 g03977 ( .a(n7737), .b(n7712), .o(n7766) );
no02f01 g03978 ( .a(n7724), .b(n7712), .o(n7767) );
no02f01 g03979 ( .a(n7767), .b(n7766), .o(n7768) );
in01f01 g03980 ( .a(n7768), .o(n7769) );
no02f01 g03981 ( .a(n7761), .b(n7712), .o(n7770) );
no02f01 g03982 ( .a(n7748), .b(n7712), .o(n7771) );
no03f01 g03983 ( .a(n7771), .b(n7770), .c(n7769), .o(n7772) );
na02f01 g03984 ( .a(n7772), .b(n7765), .o(n7773) );
in01f01 g03985 ( .a(n7581), .o(n7774) );
no02f01 g03986 ( .a(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .b(n7596), .o(n7775) );
no02f01 g03987 ( .a(n7553), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_8_), .o(n7776) );
in01f01 g03988 ( .a(n7776), .o(n7777) );
ao12f01 g03989 ( .a(n7775), .b(n7777), .c(n7774), .o(n7778) );
in01f01 g03990 ( .a(n7778), .o(n7779) );
no02f01 g03991 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_9_), .b(n7553), .o(n7780) );
no02f01 g03992 ( .a(n7597), .b(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .o(n7781) );
no02f01 g03993 ( .a(n7781), .b(n7780), .o(n7782) );
in01f01 g03994 ( .a(n7782), .o(n7783) );
no02f01 g03995 ( .a(n7783), .b(n7779), .o(n7784) );
no02f01 g03996 ( .a(n7782), .b(n7778), .o(n7785) );
no02f01 g03997 ( .a(n7785), .b(n7784), .o(n7786) );
in01f01 g03998 ( .a(n7786), .o(n7787) );
no02f01 g03999 ( .a(n7787), .b(n7682), .o(n7788) );
no02f01 g04000 ( .a(n7776), .b(n7775), .o(n7789) );
no02f01 g04001 ( .a(n7789), .b(n7581), .o(n7790) );
na02f01 g04002 ( .a(n7789), .b(n7581), .o(n7791) );
in01f01 g04003 ( .a(n7791), .o(n7792) );
no02f01 g04004 ( .a(n7792), .b(n7790), .o(n7793) );
in01f01 g04005 ( .a(n7793), .o(n7794) );
no02f01 g04006 ( .a(n7794), .b(n7682), .o(n7795) );
no02f01 g04007 ( .a(n7795), .b(n7788), .o(n7796) );
in01f01 g04008 ( .a(n7796), .o(n7797) );
no02f01 g04009 ( .a(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .b(n7599), .o(n7798) );
no03f01 g04010 ( .a(n7585), .b(n7582), .c(n7581), .o(n7799) );
no03f01 g04011 ( .a(n7799), .b(n7798), .c(n7598), .o(n7800) );
in01f01 g04012 ( .a(n7800), .o(n7801) );
no02f01 g04013 ( .a(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .b(n7600), .o(n7802) );
no02f01 g04014 ( .a(n7802), .b(n7584), .o(n7803) );
in01f01 g04015 ( .a(n7803), .o(n7804) );
no02f01 g04016 ( .a(n7804), .b(n7801), .o(n7805) );
no02f01 g04017 ( .a(n7803), .b(n7800), .o(n7806) );
no02f01 g04018 ( .a(n7806), .b(n7805), .o(n7807) );
in01f01 g04019 ( .a(n7807), .o(n7808) );
no02f01 g04020 ( .a(n7808), .b(n7682), .o(n7809) );
ao12f01 g04021 ( .a(n7598), .b(n7583), .c(n7774), .o(n7810) );
no02f01 g04022 ( .a(n7798), .b(n7585), .o(n7811) );
no02f01 g04023 ( .a(n7811), .b(n7810), .o(n7812) );
na02f01 g04024 ( .a(n7811), .b(n7810), .o(n7813) );
in01f01 g04025 ( .a(n7813), .o(n7814) );
no02f01 g04026 ( .a(n7814), .b(n7812), .o(n7815) );
in01f01 g04027 ( .a(n7815), .o(n7816) );
no02f01 g04028 ( .a(n7816), .b(n7682), .o(n7817) );
no03f01 g04029 ( .a(n7817), .b(n7809), .c(n7797), .o(n7818) );
na02f01 g04030 ( .a(n7818), .b(n7773), .o(n7819) );
no02f01 g04031 ( .a(n7605), .b(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .o(n7820) );
no03f01 g04032 ( .a(n7588), .b(n7587), .c(n7581), .o(n7821) );
no03f01 g04033 ( .a(n7821), .b(n7820), .c(n7603), .o(n7822) );
in01f01 g04034 ( .a(n7822), .o(n7823) );
no02f01 g04035 ( .a(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .b(n7604), .o(n7824) );
no02f01 g04036 ( .a(n7824), .b(n7589), .o(n7825) );
in01f01 g04037 ( .a(n7825), .o(n7826) );
no02f01 g04038 ( .a(n7826), .b(n7823), .o(n7827) );
no02f01 g04039 ( .a(n7825), .b(n7822), .o(n7828) );
no02f01 g04040 ( .a(n7828), .b(n7827), .o(n7829) );
in01f01 g04041 ( .a(n7829), .o(n7830) );
no02f01 g04042 ( .a(n7830), .b(n7682), .o(n7831) );
no02f01 g04043 ( .a(n7587), .b(n7581), .o(n7832) );
no02f01 g04044 ( .a(n7832), .b(n7603), .o(n7833) );
no02f01 g04045 ( .a(n7820), .b(n7588), .o(n7834) );
no02f01 g04046 ( .a(n7834), .b(n7833), .o(n7835) );
na02f01 g04047 ( .a(n7834), .b(n7833), .o(n7836) );
in01f01 g04048 ( .a(n7836), .o(n7837) );
no02f01 g04049 ( .a(n7837), .b(n7835), .o(n7838) );
in01f01 g04050 ( .a(n7838), .o(n7839) );
no02f01 g04051 ( .a(n7839), .b(n7682), .o(n7840) );
no02f01 g04052 ( .a(n7840), .b(n7831), .o(n7841) );
in01f01 g04053 ( .a(n7841), .o(n7842) );
no02f01 g04054 ( .a(n7842), .b(n7819), .o(n7843) );
no02f01 g04055 ( .a(n7610), .b(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .o(n7844) );
no03f01 g04056 ( .a(n7594), .b(n7591), .c(n7581), .o(n7845) );
no03f01 g04057 ( .a(n7845), .b(n7844), .c(n7608), .o(n7846) );
in01f01 g04058 ( .a(n7846), .o(n7847) );
no02f01 g04059 ( .a(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .b(n7609), .o(n7848) );
no02f01 g04060 ( .a(n7848), .b(n7593), .o(n7849) );
in01f01 g04061 ( .a(n7849), .o(n7850) );
no02f01 g04062 ( .a(n7850), .b(n7847), .o(n7851) );
no02f01 g04063 ( .a(n7849), .b(n7846), .o(n7852) );
no02f01 g04064 ( .a(n7852), .b(n7851), .o(n7853) );
in01f01 g04065 ( .a(n7853), .o(n7854) );
no02f01 g04066 ( .a(n7854), .b(n7682), .o(n7855) );
no02f01 g04067 ( .a(n7844), .b(n7594), .o(n7856) );
in01f01 g04068 ( .a(n7856), .o(n7857) );
no03f01 g04069 ( .a(n7857), .b(n7608), .c(n7592), .o(n7858) );
no02f01 g04070 ( .a(n7608), .b(n7592), .o(n7859) );
no02f01 g04071 ( .a(n7856), .b(n7859), .o(n7860) );
no02f01 g04072 ( .a(n7860), .b(n7858), .o(n7861) );
in01f01 g04073 ( .a(n7861), .o(n7862) );
no02f01 g04074 ( .a(n7862), .b(n7682), .o(n7863) );
no02f01 g04075 ( .a(n7863), .b(n7855), .o(n7864) );
na02f01 g04076 ( .a(n7864), .b(n7843), .o(n7865) );
no02f01 g04077 ( .a(n7786), .b(n7712), .o(n7866) );
no02f01 g04078 ( .a(n7793), .b(n7712), .o(n7867) );
no02f01 g04079 ( .a(n7867), .b(n7866), .o(n7868) );
no02f01 g04080 ( .a(n7807), .b(n7712), .o(n7869) );
no02f01 g04081 ( .a(n7815), .b(n7712), .o(n7870) );
no02f01 g04082 ( .a(n7870), .b(n7869), .o(n7871) );
na02f01 g04083 ( .a(n7871), .b(n7868), .o(n7872) );
in01f01 g04084 ( .a(n7872), .o(n7873) );
no02f01 g04085 ( .a(n7829), .b(n7712), .o(n7874) );
no02f01 g04086 ( .a(n7838), .b(n7712), .o(n7875) );
no02f01 g04087 ( .a(n7875), .b(n7874), .o(n7876) );
na02f01 g04088 ( .a(n7876), .b(n7873), .o(n7877) );
no02f01 g04089 ( .a(n7853), .b(n7712), .o(n7878) );
no02f01 g04090 ( .a(n7861), .b(n7712), .o(n7879) );
no03f01 g04091 ( .a(n7879), .b(n7878), .c(n7877), .o(n7880) );
na02f01 g04092 ( .a(n7880), .b(n7865), .o(n7881) );
in01f01 g04093 ( .a(n7623), .o(n7882) );
no02f01 g04094 ( .a(n7882), .b(n7616), .o(n7883) );
na02f01 g04095 ( .a(n7624), .b(n7552), .o(n7884) );
in01f01 g04096 ( .a(n7884), .o(n7885) );
no02f01 g04097 ( .a(n7885), .b(n7883), .o(n7886) );
na02f01 g04098 ( .a(n7885), .b(n7883), .o(n7887) );
in01f01 g04099 ( .a(n7887), .o(n7888) );
no02f01 g04100 ( .a(n7888), .b(n7886), .o(n7889) );
in01f01 g04101 ( .a(n7889), .o(n7890) );
no02f01 g04102 ( .a(n7890), .b(n7712), .o(n7891) );
in01f01 g04103 ( .a(n7614), .o(n7892) );
no02f01 g04104 ( .a(n7882), .b(n7615), .o(n7893) );
in01f01 g04105 ( .a(n7893), .o(n7894) );
no02f01 g04106 ( .a(n7894), .b(n7892), .o(n7895) );
no02f01 g04107 ( .a(n7893), .b(n7614), .o(n7896) );
no02f01 g04108 ( .a(n7896), .b(n7895), .o(n7897) );
in01f01 g04109 ( .a(n7897), .o(n7898) );
no02f01 g04110 ( .a(n7898), .b(n7712), .o(n7899) );
no02f01 g04111 ( .a(n7899), .b(n7891), .o(n7900) );
in01f01 g04112 ( .a(n7900), .o(n7901) );
in01f01 g04113 ( .a(n7617), .o(n7902) );
no02f01 g04114 ( .a(n7627), .b(n_17093), .o(n7903) );
no02f01 g04115 ( .a(n7903), .b(n7619), .o(n7904) );
in01f01 g04116 ( .a(n7904), .o(n7905) );
no03f01 g04117 ( .a(n7905), .b(n7625), .c(n7902), .o(n7906) );
no02f01 g04118 ( .a(n7625), .b(n7902), .o(n7907) );
no02f01 g04119 ( .a(n7904), .b(n7907), .o(n7908) );
no02f01 g04120 ( .a(n7908), .b(n7906), .o(n7909) );
in01f01 g04121 ( .a(n7909), .o(n7910) );
no02f01 g04122 ( .a(n7910), .b(n7712), .o(n7911) );
no02f01 g04123 ( .a(n7907), .b(n7619), .o(n7912) );
no02f01 g04124 ( .a(n_17093), .b(n7626), .o(n7913) );
no02f01 g04125 ( .a(n7913), .b(n7618), .o(n7914) );
in01f01 g04126 ( .a(n7914), .o(n7915) );
no03f01 g04127 ( .a(n7915), .b(n7912), .c(n7903), .o(n7916) );
no02f01 g04128 ( .a(n7912), .b(n7903), .o(n7917) );
no02f01 g04129 ( .a(n7914), .b(n7917), .o(n7918) );
no03f01 g04130 ( .a(n7918), .b(n7916), .c(n7712), .o(n7919) );
no03f01 g04131 ( .a(n7919), .b(n7911), .c(n7901), .o(n7920) );
in01f01 g04132 ( .a(n7920), .o(n7921) );
no02f01 g04133 ( .a(n7632), .b(n_17093), .o(n7922) );
no02f01 g04134 ( .a(n7643), .b(n7922), .o(n7923) );
in01f01 g04135 ( .a(n7923), .o(n7924) );
no03f01 g04136 ( .a(n7924), .b(n7630), .c(n7622), .o(n7925) );
no02f01 g04137 ( .a(n7630), .b(n7622), .o(n7926) );
no02f01 g04138 ( .a(n7923), .b(n7926), .o(n7927) );
no02f01 g04139 ( .a(n7927), .b(n7925), .o(n7928) );
in01f01 g04140 ( .a(n7928), .o(n7929) );
no02f01 g04141 ( .a(n7929), .b(n7712), .o(n7930) );
no02f01 g04142 ( .a(n7930), .b(n7921), .o(n7931) );
no02f01 g04143 ( .a(n7926), .b(n7643), .o(n7932) );
no02f01 g04144 ( .a(n7631), .b(n_17093), .o(n7933) );
no02f01 g04145 ( .a(n7933), .b(n7642), .o(n7934) );
in01f01 g04146 ( .a(n7934), .o(n7935) );
no03f01 g04147 ( .a(n7935), .b(n7932), .c(n7922), .o(n7936) );
no02f01 g04148 ( .a(n7932), .b(n7922), .o(n7937) );
no02f01 g04149 ( .a(n7934), .b(n7937), .o(n7938) );
no03f01 g04150 ( .a(n7938), .b(n7936), .c(n7712), .o(n7939) );
no03f01 g04151 ( .a(n7645), .b(n7621), .c(n7617), .o(n7940) );
ao12f01 g04152 ( .a(n7633), .b(n7644), .c(n7630), .o(n7941) );
in01f01 g04153 ( .a(n7941), .o(n7942) );
no02f01 g04154 ( .a(n7646), .b(n7635), .o(n7943) );
in01f01 g04155 ( .a(n7943), .o(n7944) );
no03f01 g04156 ( .a(n7944), .b(n7942), .c(n7940), .o(n7945) );
no02f01 g04157 ( .a(n7942), .b(n7940), .o(n7946) );
no02f01 g04158 ( .a(n7943), .b(n7946), .o(n7947) );
no02f01 g04159 ( .a(n7947), .b(n7945), .o(n7948) );
in01f01 g04160 ( .a(n7948), .o(n7949) );
no02f01 g04161 ( .a(n7949), .b(n7712), .o(n7950) );
in01f01 g04162 ( .a(n7646), .o(n7951) );
no02f01 g04163 ( .a(n7648), .b(n7636), .o(n7952) );
ao12f01 g04164 ( .a(n7952), .b(n7940), .c(n7951), .o(n7953) );
in01f01 g04165 ( .a(n7953), .o(n7954) );
no02f01 g04166 ( .a(n7649), .b(n7639), .o(n7955) );
in01f01 g04167 ( .a(n7955), .o(n7956) );
no02f01 g04168 ( .a(n7956), .b(n7954), .o(n7957) );
no02f01 g04169 ( .a(n7955), .b(n7953), .o(n7958) );
no03f01 g04170 ( .a(n7958), .b(n7957), .c(n7712), .o(n7959) );
no03f01 g04171 ( .a(n7959), .b(n7950), .c(n7939), .o(n7960) );
in01f01 g04172 ( .a(n7657), .o(n7961) );
no02f01 g04173 ( .a(n7655), .b(n7651), .o(n7962) );
ao12f01 g04174 ( .a(n7679), .b(n7962), .c(n7961), .o(n7963) );
in01f01 g04175 ( .a(n7963), .o(n7964) );
no02f01 g04176 ( .a(n7672), .b(n7656), .o(n7965) );
in01f01 g04177 ( .a(n7965), .o(n7966) );
no02f01 g04178 ( .a(n7966), .b(n7964), .o(n7967) );
no02f01 g04179 ( .a(n7965), .b(n7963), .o(n7968) );
no03f01 g04180 ( .a(n7968), .b(n7967), .c(n7712), .o(n7969) );
in01f01 g04181 ( .a(n7651), .o(n7970) );
in01f01 g04182 ( .a(n7653), .o(n7971) );
no02f01 g04183 ( .a(n_17093), .b(n7675), .o(n7972) );
ao12f01 g04184 ( .a(n7972), .b(n7971), .c(n7970), .o(n7973) );
in01f01 g04185 ( .a(n7973), .o(n7974) );
no02f01 g04186 ( .a(n7676), .b(n_17093), .o(n7975) );
no02f01 g04187 ( .a(n7975), .b(n7652), .o(n7976) );
in01f01 g04188 ( .a(n7976), .o(n7977) );
no02f01 g04189 ( .a(n7977), .b(n7974), .o(n7978) );
no02f01 g04190 ( .a(n7976), .b(n7973), .o(n7979) );
no03f01 g04191 ( .a(n7979), .b(n7978), .c(n7712), .o(n7980) );
no02f01 g04192 ( .a(n7674), .b(n7657), .o(n7981) );
in01f01 g04193 ( .a(n7981), .o(n7982) );
no03f01 g04194 ( .a(n7982), .b(n7962), .c(n7677), .o(n7983) );
no02f01 g04195 ( .a(n7962), .b(n7677), .o(n7984) );
no02f01 g04196 ( .a(n7981), .b(n7984), .o(n7985) );
no03f01 g04197 ( .a(n7985), .b(n7983), .c(n7712), .o(n7986) );
no02f01 g04198 ( .a(n7972), .b(n7653), .o(n7987) );
in01f01 g04199 ( .a(n7987), .o(n7988) );
no02f01 g04200 ( .a(n7988), .b(n7970), .o(n7989) );
no02f01 g04201 ( .a(n7987), .b(n7651), .o(n7990) );
no02f01 g04202 ( .a(n7990), .b(n7989), .o(n7991) );
in01f01 g04203 ( .a(n7991), .o(n7992) );
no02f01 g04204 ( .a(n7992), .b(n7712), .o(n7993) );
no04f01 g04205 ( .a(n7993), .b(n7986), .c(n7980), .d(n7969), .o(n7994) );
na03f01 g04206 ( .a(n7994), .b(n7960), .c(n7931), .o(n7995) );
no02f01 g04207 ( .a(n7668), .b(n_17093), .o(n7996) );
in01f01 g04208 ( .a(n7680), .o(n7997) );
in01f01 g04209 ( .a(n7660), .o(n7998) );
no02f01 g04210 ( .a(n7662), .b(n7998), .o(n7999) );
no03f01 g04211 ( .a(n7999), .b(n7997), .c(n7996), .o(n8000) );
in01f01 g04212 ( .a(n8000), .o(n8001) );
no02f01 g04213 ( .a(n7667), .b(n_17093), .o(n8002) );
no02f01 g04214 ( .a(n8002), .b(n7661), .o(n8003) );
in01f01 g04215 ( .a(n8003), .o(n8004) );
no02f01 g04216 ( .a(n8004), .b(n8001), .o(n8005) );
no02f01 g04217 ( .a(n8003), .b(n8000), .o(n8006) );
no03f01 g04218 ( .a(n8006), .b(n8005), .c(n7712), .o(n8007) );
no02f01 g04219 ( .a(n7996), .b(n7662), .o(n8008) );
in01f01 g04220 ( .a(n8008), .o(n8009) );
no03f01 g04221 ( .a(n8009), .b(n7997), .c(n7660), .o(n8010) );
ao12f01 g04222 ( .a(n8008), .b(n7680), .c(n7998), .o(n8011) );
no03f01 g04223 ( .a(n8011), .b(n8010), .c(n7712), .o(n8012) );
no02f01 g04224 ( .a(n8012), .b(n8007), .o(n8013) );
in01f01 g04225 ( .a(n8013), .o(n8014) );
no02f01 g04226 ( .a(n8014), .b(n7995), .o(n8015) );
no02f01 g04227 ( .a(n7968), .b(n7967), .o(n8016) );
no02f01 g04228 ( .a(n8016), .b(n7682), .o(n8017) );
in01f01 g04229 ( .a(n8017), .o(n8018) );
no02f01 g04230 ( .a(n7985), .b(n7983), .o(n8019) );
no02f01 g04231 ( .a(n8019), .b(n7682), .o(n8020) );
no02f01 g04232 ( .a(n7979), .b(n7978), .o(n8021) );
no02f01 g04233 ( .a(n8021), .b(n7682), .o(n8022) );
no02f01 g04234 ( .a(n7991), .b(n7682), .o(n8023) );
no03f01 g04235 ( .a(n8023), .b(n8022), .c(n8020), .o(n8024) );
na02f01 g04236 ( .a(n8024), .b(n8018), .o(n8025) );
no02f01 g04237 ( .a(n7664), .b(n7998), .o(n8026) );
no03f01 g04238 ( .a(n8026), .b(n7997), .c(n7669), .o(n8027) );
na02f01 g04239 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_30_), .b(n7550), .o(n8028) );
in01f01 g04240 ( .a(n8028), .o(n8029) );
no02f01 g04241 ( .a(n8029), .b(n7665), .o(n8030) );
no02f01 g04242 ( .a(n8030), .b(n8027), .o(n8031) );
na02f01 g04243 ( .a(n8030), .b(n8027), .o(n8032) );
in01f01 g04244 ( .a(n8032), .o(n8033) );
no02f01 g04245 ( .a(n8033), .b(n8031), .o(n8034) );
no02f01 g04246 ( .a(n8034), .b(n7682), .o(n8035) );
no02f01 g04247 ( .a(n8006), .b(n8005), .o(n8036) );
no02f01 g04248 ( .a(n8036), .b(n7682), .o(n8037) );
no02f01 g04249 ( .a(n8011), .b(n8010), .o(n8038) );
no02f01 g04250 ( .a(n8038), .b(n7682), .o(n8039) );
no04f01 g04251 ( .a(n8039), .b(n8037), .c(n8035), .d(n8025), .o(n8040) );
in01f01 g04252 ( .a(n8040), .o(n8041) );
ao12f01 g04253 ( .a(n8041), .b(n8015), .c(n7881), .o(n8042) );
na02f01 g04254 ( .a(n8034), .b(n7682), .o(n8043) );
in01f01 g04255 ( .a(n8043), .o(n8044) );
no02f01 g04256 ( .a(n7897), .b(n7682), .o(n8045) );
in01f01 g04257 ( .a(n8045), .o(n8046) );
no02f01 g04258 ( .a(n7909), .b(n7682), .o(n8047) );
no02f01 g04259 ( .a(n7889), .b(n7682), .o(n8048) );
no02f01 g04260 ( .a(n8048), .b(n8047), .o(n8049) );
na02f01 g04261 ( .a(n8049), .b(n8046), .o(n8050) );
no02f01 g04262 ( .a(n7918), .b(n7916), .o(n8051) );
no02f01 g04263 ( .a(n8051), .b(n7682), .o(n8052) );
no02f01 g04264 ( .a(n8052), .b(n8050), .o(n8053) );
no02f01 g04265 ( .a(n7938), .b(n7936), .o(n8054) );
no02f01 g04266 ( .a(n8054), .b(n7682), .o(n8055) );
no02f01 g04267 ( .a(n7928), .b(n7682), .o(n8056) );
no02f01 g04268 ( .a(n8056), .b(n8055), .o(n8057) );
na02f01 g04269 ( .a(n8057), .b(n8053), .o(n8058) );
in01f01 g04270 ( .a(n8058), .o(n8059) );
no02f01 g04271 ( .a(n7958), .b(n7957), .o(n8060) );
no02f01 g04272 ( .a(n8060), .b(n7682), .o(n8061) );
no02f01 g04273 ( .a(n7948), .b(n7682), .o(n8062) );
no02f01 g04274 ( .a(n8062), .b(n8061), .o(n8063) );
na02f01 g04275 ( .a(n8063), .b(n8059), .o(n8064) );
in01f01 g04276 ( .a(n8064), .o(n8065) );
oa12f01 g04277 ( .a(n8065), .b(n8044), .c(n8042), .o(n8066) );
in01f01 g04278 ( .a(n8066), .o(n1821) );
in01f01 g04279 ( .a(n7881), .o(n8068) );
no02f01 g04280 ( .a(n8064), .b(n8025), .o(n8069) );
oa12f01 g04281 ( .a(n8069), .b(n7995), .c(n8068), .o(n8070) );
no02f01 g04282 ( .a(n8070), .b(n8039), .o(n8071) );
no02f01 g04283 ( .a(n8071), .b(n8012), .o(n8072) );
no02f01 g04284 ( .a(n8037), .b(n8007), .o(n8073) );
in01f01 g04285 ( .a(n8073), .o(n8074) );
no02f01 g04286 ( .a(n8074), .b(n8072), .o(n8075) );
na02f01 g04287 ( .a(n8074), .b(n8072), .o(n8076) );
in01f01 g04288 ( .a(n8076), .o(n8077) );
no02f01 g04289 ( .a(n8077), .b(n8075), .o(n8078) );
no02f01 g04290 ( .a(n8039), .b(n8012), .o(n8079) );
in01f01 g04291 ( .a(n8079), .o(n8080) );
no02f01 g04292 ( .a(n8080), .b(n8070), .o(n8081) );
in01f01 g04293 ( .a(n8070), .o(n8082) );
no02f01 g04294 ( .a(n8079), .b(n8082), .o(n8083) );
no02f01 g04295 ( .a(n8083), .b(n8081), .o(n8084) );
ao12f01 g04296 ( .a(n1821), .b(n8084), .c(n8078), .o(n8085) );
in01f01 g04297 ( .a(n8085), .o(n8086) );
no02f01 g04298 ( .a(n8039), .b(n8037), .o(n8087) );
ao12f01 g04299 ( .a(n8014), .b(n8082), .c(n8087), .o(n8088) );
no02f01 g04300 ( .a(n8044), .b(n8035), .o(n8089) );
in01f01 g04301 ( .a(n8089), .o(n8090) );
no02f01 g04302 ( .a(n8090), .b(n8088), .o(n8091) );
na02f01 g04303 ( .a(n8090), .b(n8088), .o(n8092) );
in01f01 g04304 ( .a(n8092), .o(n8093) );
no02f01 g04305 ( .a(n8093), .b(n8091), .o(n8094) );
ao12f01 g04306 ( .a(n1821), .b(n8094), .c(n8086), .o(n8095) );
na02f01 g04307 ( .a(n7960), .b(n7931), .o(n8096) );
no02f01 g04308 ( .a(n8096), .b(n8068), .o(n8097) );
in01f01 g04309 ( .a(n8097), .o(n8098) );
no02f01 g04310 ( .a(n8098), .b(n7993), .o(n8099) );
in01f01 g04311 ( .a(n8099), .o(n8100) );
no02f01 g04312 ( .a(n8064), .b(n8023), .o(n8101) );
in01f01 g04313 ( .a(n8101), .o(n8102) );
no02f01 g04314 ( .a(n8102), .b(n8022), .o(n8103) );
oa12f01 g04315 ( .a(n8103), .b(n8100), .c(n7980), .o(n8104) );
no02f01 g04316 ( .a(n8104), .b(n8020), .o(n8105) );
no02f01 g04317 ( .a(n8105), .b(n7986), .o(n8106) );
in01f01 g04318 ( .a(n8106), .o(n8107) );
no02f01 g04319 ( .a(n8017), .b(n7969), .o(n8108) );
no02f01 g04320 ( .a(n8108), .b(n8107), .o(n8109) );
na02f01 g04321 ( .a(n8108), .b(n8107), .o(n8110) );
in01f01 g04322 ( .a(n8110), .o(n8111) );
no02f01 g04323 ( .a(n8111), .b(n8109), .o(n8112) );
in01f01 g04324 ( .a(n8112), .o(n8113) );
in01f01 g04325 ( .a(n8104), .o(n8114) );
no02f01 g04326 ( .a(n8020), .b(n7986), .o(n8115) );
no02f01 g04327 ( .a(n8115), .b(n8114), .o(n8116) );
na02f01 g04328 ( .a(n8115), .b(n8114), .o(n8117) );
in01f01 g04329 ( .a(n8117), .o(n8118) );
no02f01 g04330 ( .a(n8118), .b(n8116), .o(n8119) );
no02f01 g04331 ( .a(n8119), .b(n1821), .o(n8120) );
oa12f01 g04332 ( .a(n8066), .b(n8120), .c(n8113), .o(n8121) );
no02f01 g04333 ( .a(n8102), .b(n8099), .o(n8122) );
no02f01 g04334 ( .a(n8022), .b(n7980), .o(n8123) );
no02f01 g04335 ( .a(n8123), .b(n8122), .o(n8124) );
na02f01 g04336 ( .a(n8123), .b(n8122), .o(n8125) );
in01f01 g04337 ( .a(n8125), .o(n8126) );
no02f01 g04338 ( .a(n8126), .b(n8124), .o(n8127) );
no02f01 g04339 ( .a(n8097), .b(n8064), .o(n8128) );
no02f01 g04340 ( .a(n8023), .b(n7993), .o(n8129) );
no02f01 g04341 ( .a(n8129), .b(n8128), .o(n8130) );
na02f01 g04342 ( .a(n8129), .b(n8128), .o(n8131) );
in01f01 g04343 ( .a(n8131), .o(n8132) );
no02f01 g04344 ( .a(n8132), .b(n8130), .o(n8133) );
ao12f01 g04345 ( .a(n1821), .b(n8133), .c(n8127), .o(n8134) );
in01f01 g04346 ( .a(n8134), .o(n8135) );
na02f01 g04347 ( .a(n8135), .b(n8121), .o(n8136) );
in01f01 g04348 ( .a(n8136), .o(n8137) );
in01f01 g04349 ( .a(n7843), .o(n8138) );
no02f01 g04350 ( .a(n7879), .b(n7877), .o(n8139) );
oa12f01 g04351 ( .a(n8139), .b(n7863), .c(n8138), .o(n8140) );
no02f01 g04352 ( .a(n7878), .b(n7855), .o(n8141) );
in01f01 g04353 ( .a(n8141), .o(n8142) );
no02f01 g04354 ( .a(n8142), .b(n8140), .o(n8143) );
na02f01 g04355 ( .a(n8142), .b(n8140), .o(n8144) );
in01f01 g04356 ( .a(n8144), .o(n8145) );
no02f01 g04357 ( .a(n8145), .b(n8143), .o(n8146) );
in01f01 g04358 ( .a(n8146), .o(n8147) );
no02f01 g04359 ( .a(n8147), .b(n8066), .o(n8148) );
in01f01 g04360 ( .a(n8148), .o(n8149) );
in01f01 g04361 ( .a(n7709), .o(n8150) );
no02f01 g04362 ( .a(n8150), .b(n7708), .o(n8151) );
no02f01 g04363 ( .a(n8151), .b(cordic_combinational_sub_ln23_0_unr16_z_0_), .o(n8152) );
na02f01 g04364 ( .a(n8151), .b(cordic_combinational_sub_ln23_0_unr16_z_0_), .o(n8153) );
in01f01 g04365 ( .a(n8153), .o(n8154) );
no02f01 g04366 ( .a(n8154), .b(n8152), .o(n8155) );
no02f01 g04367 ( .a(n8155), .b(n8066), .o(n8156) );
na02f01 g04368 ( .a(n8155), .b(n8066), .o(n8157) );
ao12f01 g04369 ( .a(n8156), .b(n8157), .c(cordic_combinational_sub_ln23_0_unr16_z_0_), .o(n8158) );
in01f01 g04370 ( .a(n7710), .o(n8159) );
no02f01 g04371 ( .a(n7713), .b(n7699), .o(n8160) );
no02f01 g04372 ( .a(n8160), .b(n8159), .o(n8161) );
na02f01 g04373 ( .a(n8160), .b(n8159), .o(n8162) );
in01f01 g04374 ( .a(n8162), .o(n8163) );
no02f01 g04375 ( .a(n8163), .b(n8161), .o(n8164) );
in01f01 g04376 ( .a(n8164), .o(n8165) );
no02f01 g04377 ( .a(n8165), .b(n1821), .o(n8166) );
no02f01 g04378 ( .a(n8166), .b(n8158), .o(n8167) );
no02f01 g04379 ( .a(n8164), .b(n8066), .o(n8168) );
no02f01 g04380 ( .a(n8168), .b(n8167), .o(n8169) );
ao12f01 g04381 ( .a(n7713), .b(n7710), .c(n7700), .o(n8170) );
no02f01 g04382 ( .a(n7714), .b(n7691), .o(n8171) );
no02f01 g04383 ( .a(n8171), .b(n8170), .o(n8172) );
na02f01 g04384 ( .a(n8171), .b(n8170), .o(n8173) );
in01f01 g04385 ( .a(n8173), .o(n8174) );
no02f01 g04386 ( .a(n8174), .b(n8172), .o(n8175) );
ao12f01 g04387 ( .a(n8066), .b(n8175), .c(n8169), .o(n8176) );
in01f01 g04388 ( .a(n8175), .o(n8177) );
na02f01 g04389 ( .a(n8177), .b(n8167), .o(n8178) );
in01f01 g04390 ( .a(n8178), .o(n8179) );
no02f01 g04391 ( .a(n8179), .b(n8176), .o(n8180) );
in01f01 g04392 ( .a(n7716), .o(n8181) );
no02f01 g04393 ( .a(n7767), .b(n7726), .o(n8182) );
no02f01 g04394 ( .a(n8182), .b(n8181), .o(n8183) );
na02f01 g04395 ( .a(n8182), .b(n8181), .o(n8184) );
in01f01 g04396 ( .a(n8184), .o(n8185) );
no02f01 g04397 ( .a(n8185), .b(n8183), .o(n8186) );
in01f01 g04398 ( .a(n8186), .o(n8187) );
no02f01 g04399 ( .a(n8187), .b(n1821), .o(n8188) );
no02f01 g04400 ( .a(n8188), .b(n8180), .o(n8189) );
in01f01 g04401 ( .a(n7728), .o(n8190) );
in01f01 g04402 ( .a(n7739), .o(n8191) );
ao12f01 g04403 ( .a(n7769), .b(n8191), .c(n8190), .o(n8192) );
in01f01 g04404 ( .a(n8192), .o(n8193) );
no02f01 g04405 ( .a(n7771), .b(n7750), .o(n8194) );
in01f01 g04406 ( .a(n8194), .o(n8195) );
no02f01 g04407 ( .a(n8195), .b(n8193), .o(n8196) );
no02f01 g04408 ( .a(n8194), .b(n8192), .o(n8197) );
no02f01 g04409 ( .a(n8197), .b(n8196), .o(n8198) );
in01f01 g04410 ( .a(n8198), .o(n8199) );
no02f01 g04411 ( .a(n8199), .b(n1821), .o(n8200) );
no02f01 g04412 ( .a(n7767), .b(n8190), .o(n8201) );
no02f01 g04413 ( .a(n7766), .b(n7739), .o(n8202) );
no02f01 g04414 ( .a(n8202), .b(n8201), .o(n8203) );
na02f01 g04415 ( .a(n8202), .b(n8201), .o(n8204) );
in01f01 g04416 ( .a(n8204), .o(n8205) );
no02f01 g04417 ( .a(n8205), .b(n8203), .o(n8206) );
in01f01 g04418 ( .a(n8206), .o(n8207) );
no02f01 g04419 ( .a(n8207), .b(n1821), .o(n8208) );
no02f01 g04420 ( .a(n8208), .b(n8200), .o(n8209) );
ao12f01 g04421 ( .a(n8066), .b(n8206), .c(n8186), .o(n8210) );
ao12f01 g04422 ( .a(n8210), .b(n8209), .c(n8189), .o(n8211) );
in01f01 g04423 ( .a(n8211), .o(n8212) );
no02f01 g04424 ( .a(n8198), .b(n8066), .o(n8213) );
no02f01 g04425 ( .a(n8213), .b(n8212), .o(n8214) );
in01f01 g04426 ( .a(n8214), .o(n8215) );
no03f01 g04427 ( .a(n7771), .b(n7769), .c(n7753), .o(n8216) );
no02f01 g04428 ( .a(n7770), .b(n7763), .o(n8217) );
no02f01 g04429 ( .a(n8217), .b(n8216), .o(n8218) );
na02f01 g04430 ( .a(n8217), .b(n8216), .o(n8219) );
in01f01 g04431 ( .a(n8219), .o(n8220) );
no02f01 g04432 ( .a(n8220), .b(n8218), .o(n8221) );
in01f01 g04433 ( .a(n8221), .o(n8222) );
no02f01 g04434 ( .a(n8222), .b(n8215), .o(n8223) );
oa12f01 g04435 ( .a(n8066), .b(n8221), .c(n8211), .o(n8224) );
in01f01 g04436 ( .a(n8224), .o(n8225) );
in01f01 g04437 ( .a(n7795), .o(n8226) );
ao12f01 g04438 ( .a(n7867), .b(n8226), .c(n7773), .o(n8227) );
in01f01 g04439 ( .a(n8227), .o(n8228) );
no02f01 g04440 ( .a(n7866), .b(n7788), .o(n8229) );
in01f01 g04441 ( .a(n8229), .o(n8230) );
no02f01 g04442 ( .a(n8230), .b(n8228), .o(n8231) );
no02f01 g04443 ( .a(n8229), .b(n8227), .o(n8232) );
no02f01 g04444 ( .a(n8232), .b(n8231), .o(n8233) );
in01f01 g04445 ( .a(n8233), .o(n8234) );
no02f01 g04446 ( .a(n8234), .b(n1821), .o(n8235) );
in01f01 g04447 ( .a(n7773), .o(n8236) );
no02f01 g04448 ( .a(n7867), .b(n7795), .o(n8237) );
no02f01 g04449 ( .a(n8237), .b(n8236), .o(n8238) );
na02f01 g04450 ( .a(n8237), .b(n8236), .o(n8239) );
in01f01 g04451 ( .a(n8239), .o(n8240) );
no02f01 g04452 ( .a(n8240), .b(n8238), .o(n8241) );
in01f01 g04453 ( .a(n8241), .o(n8242) );
no02f01 g04454 ( .a(n8242), .b(n1821), .o(n8243) );
no02f01 g04455 ( .a(n8243), .b(n8235), .o(n8244) );
in01f01 g04456 ( .a(n8244), .o(n8245) );
no02f01 g04457 ( .a(n7797), .b(n8236), .o(n8246) );
in01f01 g04458 ( .a(n8246), .o(n8247) );
in01f01 g04459 ( .a(n7868), .o(n8248) );
no02f01 g04460 ( .a(n7870), .b(n8248), .o(n8249) );
oa12f01 g04461 ( .a(n8249), .b(n8247), .c(n7817), .o(n8250) );
in01f01 g04462 ( .a(n8250), .o(n8251) );
no02f01 g04463 ( .a(n7869), .b(n7809), .o(n8252) );
no02f01 g04464 ( .a(n8252), .b(n8251), .o(n8253) );
na02f01 g04465 ( .a(n8252), .b(n8251), .o(n8254) );
in01f01 g04466 ( .a(n8254), .o(n8255) );
no03f01 g04467 ( .a(n8255), .b(n8253), .c(n1821), .o(n8256) );
no02f01 g04468 ( .a(n7870), .b(n7817), .o(n8257) );
in01f01 g04469 ( .a(n8257), .o(n8258) );
no03f01 g04470 ( .a(n8258), .b(n8246), .c(n8248), .o(n8259) );
ao12f01 g04471 ( .a(n8257), .b(n8247), .c(n7868), .o(n8260) );
no02f01 g04472 ( .a(n8260), .b(n8259), .o(n8261) );
in01f01 g04473 ( .a(n8261), .o(n8262) );
no02f01 g04474 ( .a(n8262), .b(n1821), .o(n8263) );
no02f01 g04475 ( .a(n8263), .b(n8256), .o(n8264) );
in01f01 g04476 ( .a(n8264), .o(n8265) );
no04f01 g04477 ( .a(n8265), .b(n8245), .c(n8225), .d(n8223), .o(n8266) );
no02f01 g04478 ( .a(n8255), .b(n8253), .o(n8267) );
ao12f01 g04479 ( .a(n8066), .b(n8261), .c(n8267), .o(n8268) );
ao12f01 g04480 ( .a(n8066), .b(n8241), .c(n8233), .o(n8269) );
no02f01 g04481 ( .a(n8269), .b(n8268), .o(n8270) );
in01f01 g04482 ( .a(n8270), .o(n8271) );
no02f01 g04483 ( .a(n8271), .b(n8266), .o(n8272) );
no02f01 g04484 ( .a(n7875), .b(n7872), .o(n8273) );
oa12f01 g04485 ( .a(n8273), .b(n7840), .c(n7819), .o(n8274) );
no02f01 g04486 ( .a(n7874), .b(n7831), .o(n8275) );
in01f01 g04487 ( .a(n8275), .o(n8276) );
no02f01 g04488 ( .a(n8276), .b(n8274), .o(n8277) );
na02f01 g04489 ( .a(n8276), .b(n8274), .o(n8278) );
in01f01 g04490 ( .a(n8278), .o(n8279) );
no02f01 g04491 ( .a(n8279), .b(n8277), .o(n8280) );
in01f01 g04492 ( .a(n8280), .o(n8281) );
no02f01 g04493 ( .a(n8281), .b(n1821), .o(n8282) );
na02f01 g04494 ( .a(n7873), .b(n7819), .o(n8283) );
no02f01 g04495 ( .a(n7875), .b(n7840), .o(n8284) );
in01f01 g04496 ( .a(n8284), .o(n8285) );
no02f01 g04497 ( .a(n8285), .b(n8283), .o(n8286) );
na02f01 g04498 ( .a(n8285), .b(n8283), .o(n8287) );
in01f01 g04499 ( .a(n8287), .o(n8288) );
no02f01 g04500 ( .a(n8288), .b(n8286), .o(n8289) );
in01f01 g04501 ( .a(n8289), .o(n8290) );
no02f01 g04502 ( .a(n8290), .b(n1821), .o(n8291) );
no02f01 g04503 ( .a(n8291), .b(n8282), .o(n8292) );
in01f01 g04504 ( .a(n8292), .o(n8293) );
no02f01 g04505 ( .a(n7879), .b(n7863), .o(n8294) );
in01f01 g04506 ( .a(n8294), .o(n8295) );
no03f01 g04507 ( .a(n8295), .b(n7877), .c(n7843), .o(n8296) );
no02f01 g04508 ( .a(n7877), .b(n7843), .o(n8297) );
no02f01 g04509 ( .a(n8294), .b(n8297), .o(n8298) );
no02f01 g04510 ( .a(n8298), .b(n8296), .o(n8299) );
in01f01 g04511 ( .a(n8299), .o(n8300) );
no02f01 g04512 ( .a(n8300), .b(n1821), .o(n8301) );
no03f01 g04513 ( .a(n8301), .b(n8293), .c(n8272), .o(n8302) );
no02f01 g04514 ( .a(n8299), .b(n8066), .o(n8303) );
ao12f01 g04515 ( .a(n8066), .b(n8289), .c(n8280), .o(n8304) );
no02f01 g04516 ( .a(n8304), .b(n8303), .o(n8305) );
in01f01 g04517 ( .a(n8305), .o(n8306) );
no02f01 g04518 ( .a(n8146), .b(n1821), .o(n8307) );
no02f01 g04519 ( .a(n8307), .b(n8306), .o(n8308) );
in01f01 g04520 ( .a(n8308), .o(n8309) );
oa12f01 g04521 ( .a(n8149), .b(n8309), .c(n8302), .o(n8310) );
in01f01 g04522 ( .a(n7899), .o(n8311) );
ao12f01 g04523 ( .a(n8045), .b(n8311), .c(n7881), .o(n8312) );
in01f01 g04524 ( .a(n8312), .o(n8313) );
no02f01 g04525 ( .a(n8048), .b(n7891), .o(n8314) );
in01f01 g04526 ( .a(n8314), .o(n8315) );
no02f01 g04527 ( .a(n8315), .b(n8313), .o(n8316) );
no02f01 g04528 ( .a(n8314), .b(n8312), .o(n8317) );
no03f01 g04529 ( .a(n8317), .b(n8316), .c(n8066), .o(n8318) );
no02f01 g04530 ( .a(n8045), .b(n7899), .o(n8319) );
no02f01 g04531 ( .a(n8319), .b(n8068), .o(n8320) );
na02f01 g04532 ( .a(n8319), .b(n8068), .o(n8321) );
in01f01 g04533 ( .a(n8321), .o(n8322) );
no02f01 g04534 ( .a(n8322), .b(n8320), .o(n8323) );
in01f01 g04535 ( .a(n8323), .o(n8324) );
no02f01 g04536 ( .a(n8324), .b(n8066), .o(n8325) );
no02f01 g04537 ( .a(n8325), .b(n8318), .o(n8326) );
in01f01 g04538 ( .a(n8326), .o(n8327) );
in01f01 g04539 ( .a(n7911), .o(n8328) );
no02f01 g04540 ( .a(n7901), .b(n8068), .o(n8329) );
ao12f01 g04541 ( .a(n8050), .b(n8329), .c(n8328), .o(n8330) );
no02f01 g04542 ( .a(n8052), .b(n7919), .o(n8331) );
no02f01 g04543 ( .a(n8331), .b(n8330), .o(n8332) );
na02f01 g04544 ( .a(n8331), .b(n8330), .o(n8333) );
in01f01 g04545 ( .a(n8333), .o(n8334) );
no03f01 g04546 ( .a(n8334), .b(n8332), .c(n8066), .o(n8335) );
no03f01 g04547 ( .a(n8329), .b(n8048), .c(n8045), .o(n8336) );
no02f01 g04548 ( .a(n8047), .b(n7911), .o(n8337) );
no02f01 g04549 ( .a(n8337), .b(n8336), .o(n8338) );
na02f01 g04550 ( .a(n8337), .b(n8336), .o(n8339) );
in01f01 g04551 ( .a(n8339), .o(n8340) );
no03f01 g04552 ( .a(n8340), .b(n8338), .c(n8066), .o(n8341) );
no02f01 g04553 ( .a(n8341), .b(n8335), .o(n8342) );
in01f01 g04554 ( .a(n8342), .o(n8343) );
na02f01 g04555 ( .a(n7931), .b(n7881), .o(n8344) );
no02f01 g04556 ( .a(n8344), .b(n7939), .o(n8345) );
in01f01 g04557 ( .a(n8345), .o(n8346) );
no02f01 g04558 ( .a(n8062), .b(n8058), .o(n8347) );
oa12f01 g04559 ( .a(n8347), .b(n8346), .c(n7950), .o(n8348) );
in01f01 g04560 ( .a(n8348), .o(n8349) );
no02f01 g04561 ( .a(n8061), .b(n7959), .o(n8350) );
no02f01 g04562 ( .a(n8350), .b(n8349), .o(n8351) );
na02f01 g04563 ( .a(n8350), .b(n8349), .o(n8352) );
in01f01 g04564 ( .a(n8352), .o(n8353) );
no03f01 g04565 ( .a(n8353), .b(n8351), .c(n8066), .o(n8354) );
no02f01 g04566 ( .a(n8062), .b(n7950), .o(n8355) );
in01f01 g04567 ( .a(n8355), .o(n8356) );
no03f01 g04568 ( .a(n8356), .b(n8345), .c(n8058), .o(n8357) );
ao12f01 g04569 ( .a(n8355), .b(n8346), .c(n8059), .o(n8358) );
no03f01 g04570 ( .a(n8358), .b(n8357), .c(n8066), .o(n8359) );
in01f01 g04571 ( .a(n8053), .o(n8360) );
no02f01 g04572 ( .a(n8056), .b(n8360), .o(n8361) );
na02f01 g04573 ( .a(n8361), .b(n8344), .o(n8362) );
no02f01 g04574 ( .a(n8055), .b(n7939), .o(n8363) );
in01f01 g04575 ( .a(n8363), .o(n8364) );
no02f01 g04576 ( .a(n8364), .b(n8362), .o(n8365) );
na02f01 g04577 ( .a(n8364), .b(n8362), .o(n8366) );
in01f01 g04578 ( .a(n8366), .o(n8367) );
no03f01 g04579 ( .a(n8367), .b(n8365), .c(n8066), .o(n8368) );
ao12f01 g04580 ( .a(n8360), .b(n7920), .c(n7881), .o(n8369) );
in01f01 g04581 ( .a(n8369), .o(n8370) );
no02f01 g04582 ( .a(n8056), .b(n7930), .o(n8371) );
in01f01 g04583 ( .a(n8371), .o(n8372) );
no02f01 g04584 ( .a(n8372), .b(n8370), .o(n8373) );
no02f01 g04585 ( .a(n8371), .b(n8369), .o(n8374) );
no03f01 g04586 ( .a(n8374), .b(n8373), .c(n8066), .o(n8375) );
no02f01 g04587 ( .a(n8375), .b(n8368), .o(n8376) );
in01f01 g04588 ( .a(n8376), .o(n8377) );
no03f01 g04589 ( .a(n8377), .b(n8359), .c(n8354), .o(n8378) );
in01f01 g04590 ( .a(n8378), .o(n8379) );
no04f01 g04591 ( .a(n8379), .b(n8343), .c(n8327), .d(n8310), .o(n8380) );
no02f01 g04592 ( .a(n8317), .b(n8316), .o(n8381) );
ao12f01 g04593 ( .a(n1821), .b(n8323), .c(n8381), .o(n8382) );
no02f01 g04594 ( .a(n8334), .b(n8332), .o(n8383) );
no02f01 g04595 ( .a(n8340), .b(n8338), .o(n8384) );
ao12f01 g04596 ( .a(n1821), .b(n8384), .c(n8383), .o(n8385) );
no02f01 g04597 ( .a(n8385), .b(n8382), .o(n8386) );
in01f01 g04598 ( .a(n8386), .o(n8387) );
no02f01 g04599 ( .a(n8367), .b(n8365), .o(n8388) );
no02f01 g04600 ( .a(n8374), .b(n8373), .o(n8389) );
ao12f01 g04601 ( .a(n1821), .b(n8389), .c(n8388), .o(n8390) );
no02f01 g04602 ( .a(n8353), .b(n8351), .o(n8391) );
no02f01 g04603 ( .a(n8358), .b(n8357), .o(n8392) );
no02f01 g04604 ( .a(n8392), .b(n1821), .o(n8393) );
in01f01 g04605 ( .a(n8393), .o(n8394) );
ao12f01 g04606 ( .a(n1821), .b(n8394), .c(n8391), .o(n8395) );
no03f01 g04607 ( .a(n8395), .b(n8390), .c(n8387), .o(n8396) );
in01f01 g04608 ( .a(n8396), .o(n8397) );
no02f01 g04609 ( .a(n8113), .b(n8066), .o(n8398) );
in01f01 g04610 ( .a(n8398), .o(n8399) );
no03f01 g04611 ( .a(n8126), .b(n8124), .c(n8066), .o(n8400) );
no03f01 g04612 ( .a(n8132), .b(n8130), .c(n8066), .o(n8401) );
no02f01 g04613 ( .a(n8401), .b(n8400), .o(n8402) );
na02f01 g04614 ( .a(n8119), .b(n1821), .o(n8403) );
na03f01 g04615 ( .a(n8403), .b(n8402), .c(n8399), .o(n8404) );
no03f01 g04616 ( .a(n8093), .b(n8091), .c(n8066), .o(n8405) );
no02f01 g04617 ( .a(n8405), .b(n8404), .o(n8406) );
oa12f01 g04618 ( .a(n8406), .b(n8397), .c(n8380), .o(n8407) );
no03f01 g04619 ( .a(n8077), .b(n8075), .c(n8066), .o(n8408) );
no03f01 g04620 ( .a(n8083), .b(n8081), .c(n8066), .o(n8409) );
no02f01 g04621 ( .a(n8409), .b(n8408), .o(n8410) );
in01f01 g04622 ( .a(n8410), .o(n8411) );
ao12f01 g04623 ( .a(n8411), .b(n8407), .c(n8137), .o(n8412) );
no02f01 g04624 ( .a(n8412), .b(n8095), .o(n5973) );
in01f01 g04625 ( .a(n8157), .o(n8414) );
no02f01 g04626 ( .a(n8414), .b(n8156), .o(n8415) );
no02f01 g04627 ( .a(n8415), .b(n7703), .o(n8416) );
na02f01 g04628 ( .a(n8415), .b(n7703), .o(n8417) );
in01f01 g04629 ( .a(n8417), .o(n8418) );
no02f01 g04630 ( .a(n8418), .b(n8416), .o(n8419) );
no03f01 g04631 ( .a(n8419), .b(n8412), .c(n8095), .o(n8420) );
oa12f01 g04632 ( .a(n8419), .b(n8412), .c(n8095), .o(n8421) );
ao12f01 g04633 ( .a(n8420), .b(n8421), .c(n7703), .o(n8422) );
no02f01 g04634 ( .a(n8168), .b(n8166), .o(n8423) );
no02f01 g04635 ( .a(n8423), .b(n8158), .o(n8424) );
na02f01 g04636 ( .a(n8423), .b(n8158), .o(n8425) );
in01f01 g04637 ( .a(n8425), .o(n8426) );
no02f01 g04638 ( .a(n8426), .b(n8424), .o(n8427) );
in01f01 g04639 ( .a(n8427), .o(n8428) );
no02f01 g04640 ( .a(n8428), .b(n5973), .o(n8429) );
na02f01 g04641 ( .a(n8428), .b(n5973), .o(n8430) );
oa12f01 g04642 ( .a(n8430), .b(n8429), .c(n8422), .o(n8431) );
no02f01 g04643 ( .a(n8175), .b(n8066), .o(n8432) );
no02f01 g04644 ( .a(n8177), .b(n1821), .o(n8433) );
no02f01 g04645 ( .a(n8433), .b(n8432), .o(n8434) );
in01f01 g04646 ( .a(n8434), .o(n8435) );
no03f01 g04647 ( .a(n8435), .b(n8168), .c(n8167), .o(n8436) );
no02f01 g04648 ( .a(n8434), .b(n8169), .o(n8437) );
no02f01 g04649 ( .a(n8437), .b(n8436), .o(n8438) );
in01f01 g04650 ( .a(n8438), .o(n8439) );
oa12f01 g04651 ( .a(n5973), .b(n8439), .c(n8431), .o(n8440) );
no03f01 g04652 ( .a(n8438), .b(n8429), .c(n8422), .o(n8441) );
in01f01 g04653 ( .a(n8441), .o(n8442) );
no02f01 g04654 ( .a(n8186), .b(n8066), .o(n8443) );
no02f01 g04655 ( .a(n8443), .b(n8188), .o(n8444) );
in01f01 g04656 ( .a(n8444), .o(n8445) );
no03f01 g04657 ( .a(n8445), .b(n8179), .c(n8176), .o(n8446) );
no02f01 g04658 ( .a(n8444), .b(n8180), .o(n8447) );
no02f01 g04659 ( .a(n8447), .b(n8446), .o(n8448) );
in01f01 g04660 ( .a(n8448), .o(n8449) );
no02f01 g04661 ( .a(n8449), .b(n5973), .o(n8450) );
ao12f01 g04662 ( .a(n8450), .b(n8442), .c(n8440), .o(n8451) );
in01f01 g04663 ( .a(n8208), .o(n8452) );
ao12f01 g04664 ( .a(n8210), .b(n8452), .c(n8189), .o(n8453) );
no02f01 g04665 ( .a(n8213), .b(n8200), .o(n8454) );
no02f01 g04666 ( .a(n8454), .b(n8453), .o(n8455) );
na02f01 g04667 ( .a(n8454), .b(n8453), .o(n8456) );
in01f01 g04668 ( .a(n8456), .o(n8457) );
no02f01 g04669 ( .a(n8457), .b(n8455), .o(n8458) );
in01f01 g04670 ( .a(n8458), .o(n8459) );
no02f01 g04671 ( .a(n8459), .b(n5973), .o(n8460) );
no02f01 g04672 ( .a(n8206), .b(n8066), .o(n8461) );
no02f01 g04673 ( .a(n8461), .b(n8208), .o(n8462) );
in01f01 g04674 ( .a(n8462), .o(n8463) );
no03f01 g04675 ( .a(n8463), .b(n8443), .c(n8189), .o(n8464) );
no02f01 g04676 ( .a(n8443), .b(n8189), .o(n8465) );
no02f01 g04677 ( .a(n8462), .b(n8465), .o(n8466) );
no02f01 g04678 ( .a(n8466), .b(n8464), .o(n8467) );
in01f01 g04679 ( .a(n8467), .o(n8468) );
no02f01 g04680 ( .a(n8468), .b(n5973), .o(n8469) );
no02f01 g04681 ( .a(n8469), .b(n8460), .o(n8470) );
in01f01 g04682 ( .a(n5973), .o(n8471) );
no02f01 g04683 ( .a(n8468), .b(n8449), .o(n8472) );
no02f01 g04684 ( .a(n8472), .b(n8471), .o(n8473) );
ao12f01 g04685 ( .a(n8473), .b(n8470), .c(n8451), .o(n8474) );
no02f01 g04686 ( .a(n8458), .b(n8471), .o(n8475) );
in01f01 g04687 ( .a(n8475), .o(n8476) );
no02f01 g04688 ( .a(n8221), .b(n8066), .o(n8477) );
no02f01 g04689 ( .a(n8222), .b(n1821), .o(n8478) );
no02f01 g04690 ( .a(n8478), .b(n8477), .o(n8479) );
in01f01 g04691 ( .a(n8479), .o(n8480) );
no02f01 g04692 ( .a(n8480), .b(n8215), .o(n8481) );
no02f01 g04693 ( .a(n8479), .b(n8214), .o(n8482) );
no02f01 g04694 ( .a(n8482), .b(n8481), .o(n8483) );
na03f01 g04695 ( .a(n8483), .b(n8476), .c(n8474), .o(n8484) );
oa12f01 g04696 ( .a(n8471), .b(n8483), .c(n8474), .o(n8485) );
no02f01 g04697 ( .a(n8225), .b(n8223), .o(n8486) );
in01f01 g04698 ( .a(n8243), .o(n8487) );
no02f01 g04699 ( .a(n8241), .b(n8066), .o(n8488) );
ao12f01 g04700 ( .a(n8488), .b(n8487), .c(n8486), .o(n8489) );
in01f01 g04701 ( .a(n8489), .o(n8490) );
no02f01 g04702 ( .a(n8233), .b(n8066), .o(n8491) );
no02f01 g04703 ( .a(n8491), .b(n8235), .o(n8492) );
in01f01 g04704 ( .a(n8492), .o(n8493) );
no02f01 g04705 ( .a(n8493), .b(n8490), .o(n8494) );
no02f01 g04706 ( .a(n8492), .b(n8489), .o(n8495) );
no02f01 g04707 ( .a(n8495), .b(n8494), .o(n8496) );
in01f01 g04708 ( .a(n8496), .o(n8497) );
no02f01 g04709 ( .a(n8497), .b(n5973), .o(n8498) );
no02f01 g04710 ( .a(n8488), .b(n8243), .o(n8499) );
in01f01 g04711 ( .a(n8499), .o(n8500) );
no02f01 g04712 ( .a(n8500), .b(n8486), .o(n8501) );
in01f01 g04713 ( .a(n8486), .o(n8502) );
no02f01 g04714 ( .a(n8499), .b(n8502), .o(n8503) );
no02f01 g04715 ( .a(n8503), .b(n8501), .o(n8504) );
in01f01 g04716 ( .a(n8504), .o(n8505) );
no02f01 g04717 ( .a(n8505), .b(n5973), .o(n8506) );
no02f01 g04718 ( .a(n8506), .b(n8498), .o(n8507) );
in01f01 g04719 ( .a(n8507), .o(n8508) );
no02f01 g04720 ( .a(n8245), .b(n8502), .o(n8509) );
no02f01 g04721 ( .a(n8261), .b(n8066), .o(n8510) );
no02f01 g04722 ( .a(n8510), .b(n8263), .o(n8511) );
in01f01 g04723 ( .a(n8511), .o(n8512) );
no03f01 g04724 ( .a(n8512), .b(n8269), .c(n8509), .o(n8513) );
no02f01 g04725 ( .a(n8269), .b(n8509), .o(n8514) );
no02f01 g04726 ( .a(n8511), .b(n8514), .o(n8515) );
no02f01 g04727 ( .a(n8515), .b(n8513), .o(n8516) );
in01f01 g04728 ( .a(n8516), .o(n8517) );
no02f01 g04729 ( .a(n8517), .b(n5973), .o(n8518) );
no03f01 g04730 ( .a(n8263), .b(n8245), .c(n8502), .o(n8519) );
no02f01 g04731 ( .a(n8269), .b(n8510), .o(n8520) );
in01f01 g04732 ( .a(n8520), .o(n8521) );
no02f01 g04733 ( .a(n8267), .b(n8066), .o(n8522) );
no02f01 g04734 ( .a(n8522), .b(n8256), .o(n8523) );
in01f01 g04735 ( .a(n8523), .o(n8524) );
no03f01 g04736 ( .a(n8524), .b(n8521), .c(n8519), .o(n8525) );
no02f01 g04737 ( .a(n8521), .b(n8519), .o(n8526) );
no02f01 g04738 ( .a(n8523), .b(n8526), .o(n8527) );
no02f01 g04739 ( .a(n8527), .b(n8525), .o(n8528) );
in01f01 g04740 ( .a(n8528), .o(n8529) );
no02f01 g04741 ( .a(n8529), .b(n5973), .o(n8530) );
no03f01 g04742 ( .a(n8530), .b(n8518), .c(n8508), .o(n8531) );
na03f01 g04743 ( .a(n8531), .b(n8485), .c(n8484), .o(n8532) );
no02f01 g04744 ( .a(n8505), .b(n8497), .o(n8533) );
no02f01 g04745 ( .a(n8533), .b(n8471), .o(n8534) );
ao12f01 g04746 ( .a(n8471), .b(n8528), .c(n8516), .o(n8535) );
no02f01 g04747 ( .a(n8535), .b(n8534), .o(n8536) );
no02f01 g04748 ( .a(n8289), .b(n8066), .o(n8537) );
no02f01 g04749 ( .a(n8537), .b(n8291), .o(n8538) );
no02f01 g04750 ( .a(n8538), .b(n8272), .o(n8539) );
na02f01 g04751 ( .a(n8538), .b(n8272), .o(n8540) );
in01f01 g04752 ( .a(n8540), .o(n8541) );
no02f01 g04753 ( .a(n8541), .b(n8539), .o(n8542) );
in01f01 g04754 ( .a(n8542), .o(n8543) );
no02f01 g04755 ( .a(n8543), .b(n5973), .o(n8544) );
no02f01 g04756 ( .a(n8291), .b(n8272), .o(n8545) );
no02f01 g04757 ( .a(n8545), .b(n8537), .o(n8546) );
no02f01 g04758 ( .a(n8280), .b(n8066), .o(n8547) );
no02f01 g04759 ( .a(n8547), .b(n8282), .o(n8548) );
no02f01 g04760 ( .a(n8548), .b(n8546), .o(n8549) );
na02f01 g04761 ( .a(n8548), .b(n8546), .o(n8550) );
in01f01 g04762 ( .a(n8550), .o(n8551) );
no02f01 g04763 ( .a(n8551), .b(n8549), .o(n8552) );
in01f01 g04764 ( .a(n8552), .o(n8553) );
no02f01 g04765 ( .a(n8553), .b(n5973), .o(n8554) );
no02f01 g04766 ( .a(n8554), .b(n8544), .o(n8555) );
in01f01 g04767 ( .a(n8555), .o(n8556) );
ao12f01 g04768 ( .a(n8556), .b(n8536), .c(n8532), .o(n8557) );
no02f01 g04769 ( .a(n8542), .b(n8471), .o(n8558) );
no02f01 g04770 ( .a(n8552), .b(n8471), .o(n8559) );
no02f01 g04771 ( .a(n8559), .b(n8558), .o(n8560) );
in01f01 g04772 ( .a(n8560), .o(n8561) );
in01f01 g04773 ( .a(n8301), .o(n8562) );
na02f01 g04774 ( .a(n8292), .b(n8266), .o(n8563) );
na02f01 g04775 ( .a(n8563), .b(n8270), .o(n8564) );
ao12f01 g04776 ( .a(n8306), .b(n8564), .c(n8562), .o(n8565) );
no02f01 g04777 ( .a(n8307), .b(n8148), .o(n8566) );
no02f01 g04778 ( .a(n8566), .b(n8565), .o(n8567) );
na02f01 g04779 ( .a(n8566), .b(n8565), .o(n8568) );
in01f01 g04780 ( .a(n8568), .o(n8569) );
no02f01 g04781 ( .a(n8569), .b(n8567), .o(n8570) );
no02f01 g04782 ( .a(n8303), .b(n8301), .o(n8571) );
in01f01 g04783 ( .a(n8571), .o(n8572) );
no03f01 g04784 ( .a(n8572), .b(n8564), .c(n8304), .o(n8573) );
no02f01 g04785 ( .a(n8564), .b(n8304), .o(n8574) );
no02f01 g04786 ( .a(n8571), .b(n8574), .o(n8575) );
no02f01 g04787 ( .a(n8575), .b(n8573), .o(n8576) );
ao12f01 g04788 ( .a(n5973), .b(n8576), .c(n8570), .o(n8577) );
no03f01 g04789 ( .a(n8577), .b(n8561), .c(n8557), .o(n8578) );
in01f01 g04790 ( .a(n8570), .o(n8579) );
no02f01 g04791 ( .a(n8579), .b(n8471), .o(n8580) );
na02f01 g04792 ( .a(n8576), .b(n5973), .o(n8581) );
in01f01 g04793 ( .a(n8581), .o(n8582) );
no02f01 g04794 ( .a(n8582), .b(n8580), .o(n8583) );
in01f01 g04795 ( .a(n8583), .o(n8584) );
in01f01 g04796 ( .a(n8310), .o(n8585) );
in01f01 g04797 ( .a(n8325), .o(n8586) );
no02f01 g04798 ( .a(n8323), .b(n1821), .o(n8587) );
ao12f01 g04799 ( .a(n8587), .b(n8586), .c(n8585), .o(n8588) );
in01f01 g04800 ( .a(n8588), .o(n8589) );
no02f01 g04801 ( .a(n8381), .b(n1821), .o(n8590) );
no02f01 g04802 ( .a(n8590), .b(n8318), .o(n8591) );
in01f01 g04803 ( .a(n8591), .o(n8592) );
no02f01 g04804 ( .a(n8592), .b(n8589), .o(n8593) );
no02f01 g04805 ( .a(n8591), .b(n8588), .o(n8594) );
no02f01 g04806 ( .a(n8594), .b(n8593), .o(n8595) );
in01f01 g04807 ( .a(n8595), .o(n8596) );
no02f01 g04808 ( .a(n8587), .b(n8325), .o(n8597) );
in01f01 g04809 ( .a(n8597), .o(n8598) );
no02f01 g04810 ( .a(n8598), .b(n8585), .o(n8599) );
no02f01 g04811 ( .a(n8597), .b(n8310), .o(n8600) );
no02f01 g04812 ( .a(n8600), .b(n8599), .o(n8601) );
in01f01 g04813 ( .a(n8601), .o(n8602) );
ao12f01 g04814 ( .a(n8471), .b(n8602), .c(n8596), .o(n8603) );
no03f01 g04815 ( .a(n8603), .b(n8584), .c(n8578), .o(n8604) );
no02f01 g04816 ( .a(n8327), .b(n8310), .o(n8605) );
no02f01 g04817 ( .a(n8382), .b(n8605), .o(n8606) );
no02f01 g04818 ( .a(n8384), .b(n1821), .o(n8607) );
no02f01 g04819 ( .a(n8607), .b(n8341), .o(n8608) );
no02f01 g04820 ( .a(n8608), .b(n8606), .o(n8609) );
na02f01 g04821 ( .a(n8608), .b(n8606), .o(n8610) );
in01f01 g04822 ( .a(n8610), .o(n8611) );
no02f01 g04823 ( .a(n8611), .b(n8609), .o(n8612) );
in01f01 g04824 ( .a(n8612), .o(n8613) );
no02f01 g04825 ( .a(n8613), .b(n8471), .o(n8614) );
in01f01 g04826 ( .a(n8605), .o(n8615) );
no02f01 g04827 ( .a(n8607), .b(n8382), .o(n8616) );
oa12f01 g04828 ( .a(n8616), .b(n8341), .c(n8615), .o(n8617) );
no02f01 g04829 ( .a(n8383), .b(n1821), .o(n8618) );
no02f01 g04830 ( .a(n8618), .b(n8335), .o(n8619) );
in01f01 g04831 ( .a(n8619), .o(n8620) );
no02f01 g04832 ( .a(n8620), .b(n8617), .o(n8621) );
na02f01 g04833 ( .a(n8620), .b(n8617), .o(n8622) );
in01f01 g04834 ( .a(n8622), .o(n8623) );
no03f01 g04835 ( .a(n8623), .b(n8621), .c(n8471), .o(n8624) );
no02f01 g04836 ( .a(n8624), .b(n8614), .o(n8625) );
ao12f01 g04837 ( .a(n8387), .b(n8342), .c(n8605), .o(n8626) );
no02f01 g04838 ( .a(n8626), .b(n8377), .o(n8627) );
no02f01 g04839 ( .a(n8627), .b(n8390), .o(n8628) );
ao12f01 g04840 ( .a(n8359), .b(n8628), .c(n8394), .o(n8629) );
no02f01 g04841 ( .a(n8391), .b(n1821), .o(n8630) );
no02f01 g04842 ( .a(n8630), .b(n8354), .o(n8631) );
in01f01 g04843 ( .a(n8631), .o(n8632) );
no02f01 g04844 ( .a(n8632), .b(n8629), .o(n8633) );
na02f01 g04845 ( .a(n8632), .b(n8629), .o(n8634) );
in01f01 g04846 ( .a(n8634), .o(n8635) );
no03f01 g04847 ( .a(n8635), .b(n8633), .c(n8471), .o(n8636) );
no02f01 g04848 ( .a(n8389), .b(n1821), .o(n8637) );
no02f01 g04849 ( .a(n8637), .b(n8375), .o(n8638) );
no02f01 g04850 ( .a(n8638), .b(n8626), .o(n8639) );
na02f01 g04851 ( .a(n8638), .b(n8626), .o(n8640) );
in01f01 g04852 ( .a(n8640), .o(n8641) );
no02f01 g04853 ( .a(n8641), .b(n8639), .o(n8642) );
in01f01 g04854 ( .a(n8642), .o(n8643) );
no02f01 g04855 ( .a(n8643), .b(n8471), .o(n8644) );
no02f01 g04856 ( .a(n8626), .b(n8375), .o(n8645) );
no02f01 g04857 ( .a(n8645), .b(n8637), .o(n8646) );
no02f01 g04858 ( .a(n8388), .b(n1821), .o(n8647) );
no02f01 g04859 ( .a(n8647), .b(n8368), .o(n8648) );
no02f01 g04860 ( .a(n8648), .b(n8646), .o(n8649) );
na02f01 g04861 ( .a(n8648), .b(n8646), .o(n8650) );
in01f01 g04862 ( .a(n8650), .o(n8651) );
no03f01 g04863 ( .a(n8651), .b(n8649), .c(n8471), .o(n8652) );
no02f01 g04864 ( .a(n8652), .b(n8644), .o(n8653) );
in01f01 g04865 ( .a(n8653), .o(n8654) );
no02f01 g04866 ( .a(n8393), .b(n8359), .o(n8655) );
no02f01 g04867 ( .a(n8655), .b(n8628), .o(n8656) );
na02f01 g04868 ( .a(n8655), .b(n8628), .o(n8657) );
in01f01 g04869 ( .a(n8657), .o(n8658) );
no03f01 g04870 ( .a(n8658), .b(n8656), .c(n8471), .o(n8659) );
no03f01 g04871 ( .a(n8659), .b(n8654), .c(n8636), .o(n8660) );
na03f01 g04872 ( .a(n8660), .b(n8625), .c(n8604), .o(n8661) );
ao12f01 g04873 ( .a(n5973), .b(n8601), .c(n8595), .o(n8662) );
no02f01 g04874 ( .a(n8623), .b(n8621), .o(n8663) );
ao12f01 g04875 ( .a(n5973), .b(n8663), .c(n8612), .o(n8664) );
no02f01 g04876 ( .a(n8664), .b(n8662), .o(n8665) );
in01f01 g04877 ( .a(n8665), .o(n8666) );
no02f01 g04878 ( .a(n8642), .b(n5973), .o(n8667) );
in01f01 g04879 ( .a(n8649), .o(n8668) );
ao12f01 g04880 ( .a(n5973), .b(n8650), .c(n8668), .o(n8669) );
no03f01 g04881 ( .a(n8669), .b(n8667), .c(n8666), .o(n8670) );
in01f01 g04882 ( .a(n8670), .o(n8671) );
no02f01 g04883 ( .a(n8635), .b(n8633), .o(n8672) );
no02f01 g04884 ( .a(n8658), .b(n8656), .o(n8673) );
ao12f01 g04885 ( .a(n5973), .b(n8673), .c(n8672), .o(n8674) );
no02f01 g04886 ( .a(n8674), .b(n8671), .o(n8675) );
no02f01 g04887 ( .a(n8133), .b(n1821), .o(n8676) );
no02f01 g04888 ( .a(n8676), .b(n8401), .o(n8677) );
in01f01 g04889 ( .a(n8677), .o(n8678) );
no03f01 g04890 ( .a(n8678), .b(n8397), .c(n8380), .o(n8679) );
no02f01 g04891 ( .a(n8397), .b(n8380), .o(n8680) );
no02f01 g04892 ( .a(n8677), .b(n8680), .o(n8681) );
no02f01 g04893 ( .a(n8681), .b(n8679), .o(n8682) );
in01f01 g04894 ( .a(n8682), .o(n8683) );
no02f01 g04895 ( .a(n8401), .b(n8680), .o(n8684) );
no02f01 g04896 ( .a(n8684), .b(n8676), .o(n8685) );
no02f01 g04897 ( .a(n8127), .b(n1821), .o(n8686) );
no02f01 g04898 ( .a(n8686), .b(n8400), .o(n8687) );
no02f01 g04899 ( .a(n8687), .b(n8685), .o(n8688) );
na02f01 g04900 ( .a(n8687), .b(n8685), .o(n8689) );
in01f01 g04901 ( .a(n8689), .o(n8690) );
no02f01 g04902 ( .a(n8690), .b(n8688), .o(n8691) );
in01f01 g04903 ( .a(n8691), .o(n8692) );
ao12f01 g04904 ( .a(n8471), .b(n8692), .c(n8683), .o(n8693) );
in01f01 g04905 ( .a(n8403), .o(n8694) );
in01f01 g04906 ( .a(n8402), .o(n8695) );
no02f01 g04907 ( .a(n8695), .b(n8680), .o(n8696) );
in01f01 g04908 ( .a(n8696), .o(n8697) );
no02f01 g04909 ( .a(n8134), .b(n8120), .o(n8698) );
oa12f01 g04910 ( .a(n8698), .b(n8697), .c(n8694), .o(n8699) );
no02f01 g04911 ( .a(n8112), .b(n1821), .o(n8700) );
no02f01 g04912 ( .a(n8700), .b(n8398), .o(n8701) );
in01f01 g04913 ( .a(n8701), .o(n8702) );
no02f01 g04914 ( .a(n8702), .b(n8699), .o(n8703) );
na02f01 g04915 ( .a(n8702), .b(n8699), .o(n8704) );
in01f01 g04916 ( .a(n8704), .o(n8705) );
no02f01 g04917 ( .a(n8705), .b(n8703), .o(n8706) );
in01f01 g04918 ( .a(n8706), .o(n8707) );
no02f01 g04919 ( .a(n8707), .b(n8471), .o(n8708) );
no02f01 g04920 ( .a(n8694), .b(n8120), .o(n8709) );
in01f01 g04921 ( .a(n8709), .o(n8710) );
no03f01 g04922 ( .a(n8710), .b(n8696), .c(n8134), .o(n8711) );
ao12f01 g04923 ( .a(n8709), .b(n8697), .c(n8135), .o(n8712) );
no03f01 g04924 ( .a(n8712), .b(n8711), .c(n8471), .o(n8713) );
no03f01 g04925 ( .a(n8713), .b(n8708), .c(n8693), .o(n8714) );
in01f01 g04926 ( .a(n8714), .o(n8715) );
ao12f01 g04927 ( .a(n8715), .b(n8675), .c(n8661), .o(n8716) );
in01f01 g04928 ( .a(n8716), .o(n8717) );
oa12f01 g04929 ( .a(n8137), .b(n8404), .c(n8680), .o(n8718) );
no02f01 g04930 ( .a(n8084), .b(n1821), .o(n8719) );
no02f01 g04931 ( .a(n8719), .b(n8409), .o(n8720) );
in01f01 g04932 ( .a(n8720), .o(n8721) );
no02f01 g04933 ( .a(n8721), .b(n8718), .o(n8722) );
in01f01 g04934 ( .a(n8718), .o(n8723) );
no02f01 g04935 ( .a(n8720), .b(n8723), .o(n8724) );
no02f01 g04936 ( .a(n8724), .b(n8722), .o(n8725) );
in01f01 g04937 ( .a(n8725), .o(n8726) );
no02f01 g04938 ( .a(n8719), .b(n8718), .o(n8727) );
no02f01 g04939 ( .a(n8727), .b(n8409), .o(n8728) );
no02f01 g04940 ( .a(n8078), .b(n1821), .o(n8729) );
no02f01 g04941 ( .a(n8729), .b(n8408), .o(n8730) );
in01f01 g04942 ( .a(n8730), .o(n8731) );
no02f01 g04943 ( .a(n8731), .b(n8728), .o(n8732) );
na02f01 g04944 ( .a(n8731), .b(n8728), .o(n8733) );
in01f01 g04945 ( .a(n8733), .o(n8734) );
no02f01 g04946 ( .a(n8734), .b(n8732), .o(n8735) );
in01f01 g04947 ( .a(n8735), .o(n8736) );
ao12f01 g04948 ( .a(n8471), .b(n8736), .c(n8726), .o(n8737) );
in01f01 g04949 ( .a(n8737), .o(n8738) );
ao12f01 g04950 ( .a(n8085), .b(n8718), .c(n8410), .o(n8739) );
no02f01 g04951 ( .a(n8094), .b(n1821), .o(n8740) );
no02f01 g04952 ( .a(n8740), .b(n8405), .o(n8741) );
no02f01 g04953 ( .a(n8741), .b(n8739), .o(n8742) );
na02f01 g04954 ( .a(n8741), .b(n8739), .o(n8743) );
in01f01 g04955 ( .a(n8743), .o(n8744) );
no02f01 g04956 ( .a(n8744), .b(n8742), .o(n8745) );
in01f01 g04957 ( .a(n8745), .o(n8746) );
no02f01 g04958 ( .a(n8746), .b(n8471), .o(n8747) );
in01f01 g04959 ( .a(n8747), .o(n8748) );
na02f01 g04960 ( .a(n8748), .b(n8738), .o(n8749) );
no02f01 g04961 ( .a(n8749), .b(n8717), .o(n8750) );
no02f01 g04962 ( .a(n8682), .b(n5973), .o(n8751) );
in01f01 g04963 ( .a(n8751), .o(n8752) );
ao12f01 g04964 ( .a(n5973), .b(n8752), .c(n8691), .o(n8753) );
in01f01 g04965 ( .a(n8753), .o(n8754) );
no02f01 g04966 ( .a(n8712), .b(n8711), .o(n8755) );
no02f01 g04967 ( .a(n8755), .b(n5973), .o(n8756) );
no02f01 g04968 ( .a(n8756), .b(n8707), .o(n8757) );
oa12f01 g04969 ( .a(n8754), .b(n8757), .c(n5973), .o(n8758) );
ao12f01 g04970 ( .a(n5973), .b(n8735), .c(n8725), .o(n8759) );
in01f01 g04971 ( .a(n8759), .o(n8760) );
ao12f01 g04972 ( .a(n5973), .b(n8760), .c(n8745), .o(n8761) );
no03f01 g04973 ( .a(n8761), .b(n8758), .c(n8750), .o(n2131) );
in01f01 g04974 ( .a(n2131), .o(n228) );
in01f01 g04975 ( .a(beta_6), .o(n8764) );
in01f01 g04976 ( .a(beta_31), .o(n8765) );
in01f01 g04977 ( .a(beta_3), .o(n8766) );
na02f01 g04978 ( .a(beta_4), .b(n8765), .o(n8767) );
no02f01 g04979 ( .a(beta_4), .b(n8765), .o(n8768) );
oa12f01 g04980 ( .a(n8767), .b(n8768), .c(n8766), .o(n8769) );
no03f01 g04981 ( .a(n8769), .b(n8765), .c(beta_5), .o(n8770) );
na03f01 g04982 ( .a(n8769), .b(n8765), .c(beta_5), .o(n8771) );
oa12f01 g04983 ( .a(n8771), .b(n8770), .c(n8764), .o(n8772) );
no02f01 g04984 ( .a(n8765), .b(beta_7), .o(n8773) );
in01f01 g04985 ( .a(n8773), .o(n8774) );
oa12f01 g04986 ( .a(beta_8), .b(n8774), .c(n8772), .o(n8775) );
na03f01 g04987 ( .a(n8772), .b(n8765), .c(beta_7), .o(n8776) );
na02f01 g04988 ( .a(n8776), .b(n8775), .o(n8777) );
in01f01 g04989 ( .a(beta_9), .o(n8778) );
in01f01 g04990 ( .a(beta_10), .o(n8779) );
ao12f01 g04991 ( .a(n8765), .b(n8779), .c(n8778), .o(n8780) );
no02f01 g04992 ( .a(beta_31), .b(beta_9), .o(n8781) );
no02f01 g04993 ( .a(beta_31), .b(beta_10), .o(n8782) );
no02f01 g04994 ( .a(n8782), .b(n8781), .o(n8783) );
oa12f01 g04995 ( .a(n8783), .b(n8780), .c(n8777), .o(n8784) );
in01f01 g04996 ( .a(n8784), .o(n8785) );
no02f01 g04997 ( .a(beta_31), .b(beta_11), .o(n8786) );
na02f01 g04998 ( .a(n8786), .b(n8784), .o(n8787) );
in01f01 g04999 ( .a(beta_11), .o(n8788) );
no02f01 g05000 ( .a(n8765), .b(n8788), .o(n8789) );
ao22f01 g05001 ( .a(n8789), .b(n8785), .c(n8787), .d(beta_12), .o(n8790) );
in01f01 g05002 ( .a(beta_13), .o(n8791) );
in01f01 g05003 ( .a(beta_14), .o(n8792) );
ao12f01 g05004 ( .a(n8765), .b(n8792), .c(n8791), .o(n8793) );
in01f01 g05005 ( .a(n8793), .o(n8794) );
no02f01 g05006 ( .a(beta_31), .b(beta_13), .o(n8795) );
no02f01 g05007 ( .a(beta_31), .b(beta_14), .o(n8796) );
no02f01 g05008 ( .a(n8796), .b(n8795), .o(n8797) );
in01f01 g05009 ( .a(n8797), .o(n8798) );
ao12f01 g05010 ( .a(n8798), .b(n8794), .c(n8790), .o(n8799) );
no02f01 g05011 ( .a(beta_31), .b(beta_15), .o(n8800) );
no02f01 g05012 ( .a(beta_31), .b(beta_16), .o(n8801) );
no02f01 g05013 ( .a(n8801), .b(n8800), .o(n8802) );
in01f01 g05014 ( .a(n8802), .o(n8803) );
no02f01 g05015 ( .a(beta_17), .b(beta_31), .o(n8804) );
no02f01 g05016 ( .a(n8804), .b(n8803), .o(n8805) );
in01f01 g05017 ( .a(beta_15), .o(n8806) );
in01f01 g05018 ( .a(beta_16), .o(n8807) );
ao12f01 g05019 ( .a(n8765), .b(n8807), .c(n8806), .o(n8808) );
ao12f01 g05020 ( .a(n8808), .b(n8805), .c(n8799), .o(n8809) );
no02f01 g05021 ( .a(n8765), .b(beta_18), .o(n8810) );
in01f01 g05022 ( .a(beta_18), .o(n8811) );
in01f01 g05023 ( .a(beta_17), .o(n8812) );
ao12f01 g05024 ( .a(n8811), .b(n8812), .c(beta_31), .o(n8813) );
in01f01 g05025 ( .a(n8813), .o(n8814) );
oa12f01 g05026 ( .a(n8814), .b(n8810), .c(n8809), .o(n8815) );
ao12f01 g05027 ( .a(n8765), .b(beta_19), .c(beta_20), .o(n8816) );
no02f01 g05028 ( .a(beta_31), .b(beta_22), .o(n8817) );
no02f01 g05029 ( .a(n8765), .b(beta_21), .o(n8818) );
no03f01 g05030 ( .a(n8818), .b(n8817), .c(n8816), .o(n8819) );
na02f01 g05031 ( .a(n8819), .b(n8815), .o(n8820) );
in01f01 g05032 ( .a(n8820), .o(n8821) );
in01f01 g05033 ( .a(n8817), .o(n8822) );
in01f01 g05034 ( .a(beta_22), .o(n8823) );
in01f01 g05035 ( .a(beta_21), .o(n8824) );
ao12f01 g05036 ( .a(n8823), .b(n8765), .c(n8824), .o(n8825) );
in01f01 g05037 ( .a(beta_20), .o(n8826) );
in01f01 g05038 ( .a(beta_19), .o(n8827) );
ao12f01 g05039 ( .a(beta_31), .b(n8827), .c(n8826), .o(n8828) );
oa12f01 g05040 ( .a(n8822), .b(n8828), .c(n8825), .o(n8829) );
in01f01 g05041 ( .a(n8829), .o(n8830) );
no02f01 g05042 ( .a(n8830), .b(n8821), .o(n8831) );
ao12f01 g05043 ( .a(n8765), .b(beta_23), .c(beta_24), .o(n8832) );
no02f01 g05044 ( .a(beta_31), .b(beta_25), .o(n8833) );
no02f01 g05045 ( .a(beta_26), .b(n8765), .o(n8834) );
no03f01 g05046 ( .a(n8834), .b(n8833), .c(n8832), .o(n8835) );
in01f01 g05047 ( .a(n8835), .o(n8836) );
no02f01 g05048 ( .a(n8836), .b(n8831), .o(n8837) );
in01f01 g05049 ( .a(n8833), .o(n8838) );
in01f01 g05050 ( .a(beta_24), .o(n8839) );
in01f01 g05051 ( .a(beta_23), .o(n8840) );
ao12f01 g05052 ( .a(beta_31), .b(n8840), .c(n8839), .o(n8841) );
in01f01 g05053 ( .a(beta_25), .o(n8842) );
in01f01 g05054 ( .a(beta_26), .o(n8843) );
ao12f01 g05055 ( .a(n8843), .b(beta_31), .c(n8842), .o(n8844) );
ao12f01 g05056 ( .a(n8844), .b(n8841), .c(n8838), .o(n8845) );
in01f01 g05057 ( .a(n8845), .o(n8846) );
no02f01 g05058 ( .a(n8846), .b(n8837), .o(n8847) );
in01f01 g05059 ( .a(n8847), .o(n8848) );
in01f01 g05060 ( .a(beta_27), .o(n8849) );
no02f01 g05061 ( .a(n8765), .b(n8849), .o(n8850) );
na02f01 g05062 ( .a(n8850), .b(n8848), .o(n8851) );
no02f01 g05063 ( .a(beta_31), .b(beta_27), .o(n8852) );
na02f01 g05064 ( .a(n8852), .b(n8847), .o(n8853) );
na02f01 g05065 ( .a(n8853), .b(beta_28), .o(n8854) );
na02f01 g05066 ( .a(n8854), .b(n8851), .o(n8855) );
no02f01 g05067 ( .a(beta_31), .b(beta_29), .o(n8856) );
no02f01 g05068 ( .a(n8765), .b(beta_30), .o(n8857) );
no02f01 g05069 ( .a(n8857), .b(n8856), .o(n8858) );
in01f01 g05070 ( .a(beta_30), .o(n8859) );
in01f01 g05071 ( .a(beta_29), .o(n8860) );
ao12f01 g05072 ( .a(n8859), .b(beta_31), .c(n8860), .o(n8861) );
ao12f01 g05073 ( .a(n8861), .b(n8858), .c(n8855), .o(n8862) );
ao22f01 g05074 ( .a(n8853), .b(beta_28), .c(n8850), .d(n8848), .o(n8863) );
no02f01 g05075 ( .a(n8765), .b(n8860), .o(n8864) );
in01f01 g05076 ( .a(n8864), .o(n8865) );
ao12f01 g05077 ( .a(n8856), .b(n8865), .c(n8863), .o(n8866) );
in01f01 g05078 ( .a(n8866), .o(n8867) );
no02f01 g05079 ( .a(beta_31), .b(n8859), .o(n8868) );
no02f01 g05080 ( .a(n8868), .b(n8857), .o(n8869) );
no02f01 g05081 ( .a(n8869), .b(n8867), .o(n8870) );
na02f01 g05082 ( .a(n8869), .b(n8867), .o(n8871) );
in01f01 g05083 ( .a(n8871), .o(n8872) );
no02f01 g05084 ( .a(n8872), .b(n8870), .o(n8873) );
no02f01 g05085 ( .a(n8873), .b(n8862), .o(n8874) );
no02f01 g05086 ( .a(n8765), .b(n8842), .o(n8875) );
in01f01 g05087 ( .a(n8875), .o(n8876) );
no02f01 g05088 ( .a(n8832), .b(n8831), .o(n8877) );
no02f01 g05089 ( .a(n8877), .b(n8841), .o(n8878) );
ao12f01 g05090 ( .a(n8833), .b(n8878), .c(n8876), .o(n8879) );
in01f01 g05091 ( .a(n8879), .o(n8880) );
no02f01 g05092 ( .a(n8843), .b(beta_31), .o(n8881) );
no02f01 g05093 ( .a(n8881), .b(n8834), .o(n8882) );
no02f01 g05094 ( .a(n8882), .b(n8880), .o(n8883) );
na02f01 g05095 ( .a(n8882), .b(n8880), .o(n8884) );
in01f01 g05096 ( .a(n8884), .o(n8885) );
no03f01 g05097 ( .a(n8885), .b(n8883), .c(n8862), .o(n8886) );
no02f01 g05098 ( .a(beta_31), .b(n8849), .o(n8887) );
no02f01 g05099 ( .a(n8765), .b(beta_27), .o(n8888) );
no02f01 g05100 ( .a(n8888), .b(n8887), .o(n8889) );
in01f01 g05101 ( .a(n8889), .o(n8890) );
no02f01 g05102 ( .a(n8890), .b(n8848), .o(n8891) );
no02f01 g05103 ( .a(n8889), .b(n8847), .o(n8892) );
no02f01 g05104 ( .a(n8892), .b(n8891), .o(n8893) );
in01f01 g05105 ( .a(n8893), .o(n8894) );
no02f01 g05106 ( .a(n8894), .b(n8862), .o(n8895) );
no02f01 g05107 ( .a(n8895), .b(n8886), .o(n8896) );
in01f01 g05108 ( .a(n8858), .o(n8897) );
in01f01 g05109 ( .a(n8861), .o(n8898) );
oa12f01 g05110 ( .a(n8898), .b(n8897), .c(n8863), .o(n8899) );
no02f01 g05111 ( .a(n8885), .b(n8883), .o(n8900) );
ao12f01 g05112 ( .a(n8899), .b(n8893), .c(n8900), .o(n8901) );
no02f01 g05113 ( .a(n8875), .b(n8833), .o(n8902) );
in01f01 g05114 ( .a(n8902), .o(n8903) );
no03f01 g05115 ( .a(n8903), .b(n8877), .c(n8841), .o(n8904) );
no02f01 g05116 ( .a(n8902), .b(n8878), .o(n8905) );
no02f01 g05117 ( .a(n8905), .b(n8904), .o(n8906) );
in01f01 g05118 ( .a(n8831), .o(n8907) );
no02f01 g05119 ( .a(n8840), .b(beta_31), .o(n8908) );
no02f01 g05120 ( .a(beta_23), .b(n8765), .o(n8909) );
in01f01 g05121 ( .a(n8909), .o(n8910) );
ao12f01 g05122 ( .a(n8908), .b(n8910), .c(n8907), .o(n8911) );
in01f01 g05123 ( .a(n8911), .o(n8912) );
no02f01 g05124 ( .a(beta_31), .b(n8839), .o(n8913) );
no02f01 g05125 ( .a(n8765), .b(beta_24), .o(n8914) );
no02f01 g05126 ( .a(n8914), .b(n8913), .o(n8915) );
in01f01 g05127 ( .a(n8915), .o(n8916) );
no02f01 g05128 ( .a(n8916), .b(n8912), .o(n8917) );
no02f01 g05129 ( .a(n8915), .b(n8911), .o(n8918) );
no02f01 g05130 ( .a(n8918), .b(n8917), .o(n8919) );
ao12f01 g05131 ( .a(n8906), .b(n8919), .c(n8862), .o(n8920) );
oa12f01 g05132 ( .a(n8896), .b(n8920), .c(n8901), .o(n8921) );
no02f01 g05133 ( .a(n8808), .b(n8799), .o(n8922) );
no02f01 g05134 ( .a(n8922), .b(n8803), .o(n8923) );
in01f01 g05135 ( .a(n8923), .o(n8924) );
no02f01 g05136 ( .a(n8812), .b(n8765), .o(n8925) );
no02f01 g05137 ( .a(n8925), .b(n8804), .o(n8926) );
no02f01 g05138 ( .a(n8926), .b(n8924), .o(n8927) );
na02f01 g05139 ( .a(n8926), .b(n8924), .o(n8928) );
in01f01 g05140 ( .a(n8928), .o(n8929) );
no02f01 g05141 ( .a(n8929), .b(n8927), .o(n8930) );
in01f01 g05142 ( .a(n8800), .o(n8931) );
no02f01 g05143 ( .a(n8765), .b(n8806), .o(n8932) );
ao12f01 g05144 ( .a(n8932), .b(n8931), .c(n8799), .o(n8933) );
in01f01 g05145 ( .a(n8933), .o(n8934) );
no02f01 g05146 ( .a(n8765), .b(n8807), .o(n8935) );
no02f01 g05147 ( .a(n8935), .b(n8801), .o(n8936) );
in01f01 g05148 ( .a(n8936), .o(n8937) );
no02f01 g05149 ( .a(n8937), .b(n8934), .o(n8938) );
no02f01 g05150 ( .a(n8936), .b(n8933), .o(n8939) );
no02f01 g05151 ( .a(n8939), .b(n8938), .o(n8940) );
ao12f01 g05152 ( .a(n8862), .b(n8940), .c(n8930), .o(n8941) );
in01f01 g05153 ( .a(n8941), .o(n8942) );
in01f01 g05154 ( .a(n8790), .o(n8943) );
no02f01 g05155 ( .a(n8765), .b(n8791), .o(n8944) );
no02f01 g05156 ( .a(n8795), .b(n8944), .o(n8945) );
in01f01 g05157 ( .a(n8945), .o(n8946) );
no02f01 g05158 ( .a(n8946), .b(n8943), .o(n8947) );
no02f01 g05159 ( .a(n8945), .b(n8790), .o(n8948) );
no02f01 g05160 ( .a(n8948), .b(n8947), .o(n8949) );
in01f01 g05161 ( .a(n8949), .o(n8950) );
no02f01 g05162 ( .a(n8950), .b(n8862), .o(n8951) );
in01f01 g05163 ( .a(n8951), .o(n8952) );
no02f01 g05164 ( .a(beta_31), .b(n8788), .o(n8953) );
no02f01 g05165 ( .a(n8765), .b(beta_11), .o(n8954) );
no02f01 g05166 ( .a(n8954), .b(n8784), .o(n8955) );
no02f01 g05167 ( .a(n8955), .b(n8953), .o(n8956) );
no02f01 g05168 ( .a(beta_31), .b(beta_12), .o(n8957) );
na02f01 g05169 ( .a(beta_31), .b(beta_12), .o(n8958) );
in01f01 g05170 ( .a(n8958), .o(n8959) );
no02f01 g05171 ( .a(n8959), .b(n8957), .o(n8960) );
no02f01 g05172 ( .a(n8960), .b(n8956), .o(n8961) );
na02f01 g05173 ( .a(n8960), .b(n8956), .o(n8962) );
in01f01 g05174 ( .a(n8962), .o(n8963) );
no02f01 g05175 ( .a(n8963), .b(n8961), .o(n8964) );
no02f01 g05176 ( .a(n8964), .b(n8862), .o(n8965) );
in01f01 g05177 ( .a(n8965), .o(n8966) );
na02f01 g05178 ( .a(n8899), .b(n8766), .o(n8967) );
in01f01 g05179 ( .a(n8967), .o(n8968) );
in01f01 g05180 ( .a(beta_2), .o(n8969) );
no02f01 g05181 ( .a(n8899), .b(n8969), .o(n8970) );
in01f01 g05182 ( .a(n8970), .o(n8971) );
in01f01 g05183 ( .a(beta_1), .o(n8972) );
in01f01 g05184 ( .a(beta_0), .o(n4932) );
no02f01 g05185 ( .a(n4932), .b(n8972), .o(n8974) );
no02f01 g05186 ( .a(beta_0), .b(beta_1), .o(n8975) );
in01f01 g05187 ( .a(n8975), .o(n8976) );
ao12f01 g05188 ( .a(n8974), .b(n8976), .c(n8899), .o(n8977) );
no02f01 g05189 ( .a(n8862), .b(beta_2), .o(n8978) );
oa12f01 g05190 ( .a(n8971), .b(n8978), .c(n8977), .o(n8979) );
no02f01 g05191 ( .a(n8899), .b(n8766), .o(n8980) );
in01f01 g05192 ( .a(n8980), .o(n8981) );
ao12f01 g05193 ( .a(n8968), .b(n8981), .c(n8979), .o(n8982) );
in01f01 g05194 ( .a(n8767), .o(n8983) );
no02f01 g05195 ( .a(n8768), .b(n8983), .o(n8984) );
no02f01 g05196 ( .a(n8984), .b(n8766), .o(n8985) );
na02f01 g05197 ( .a(n8984), .b(n8766), .o(n8986) );
in01f01 g05198 ( .a(n8986), .o(n8987) );
no02f01 g05199 ( .a(n8987), .b(n8985), .o(n8988) );
in01f01 g05200 ( .a(n8988), .o(n8989) );
no02f01 g05201 ( .a(n8989), .b(n8899), .o(n8990) );
in01f01 g05202 ( .a(beta_5), .o(n8991) );
no02f01 g05203 ( .a(n8765), .b(n8991), .o(n8992) );
no02f01 g05204 ( .a(beta_31), .b(beta_5), .o(n8993) );
no02f01 g05205 ( .a(n8993), .b(n8992), .o(n8994) );
in01f01 g05206 ( .a(n8994), .o(n8995) );
no02f01 g05207 ( .a(n8995), .b(n8769), .o(n8996) );
in01f01 g05208 ( .a(n8769), .o(n8997) );
no02f01 g05209 ( .a(n8994), .b(n8997), .o(n8998) );
no02f01 g05210 ( .a(n8998), .b(n8996), .o(n8999) );
in01f01 g05211 ( .a(n8999), .o(n9000) );
no02f01 g05212 ( .a(n9000), .b(n8899), .o(n9001) );
in01f01 g05213 ( .a(n8993), .o(n9002) );
ao12f01 g05214 ( .a(n8992), .b(n9002), .c(n8769), .o(n9003) );
in01f01 g05215 ( .a(n9003), .o(n9004) );
no02f01 g05216 ( .a(beta_31), .b(n8764), .o(n9005) );
no02f01 g05217 ( .a(n8765), .b(beta_6), .o(n9006) );
no02f01 g05218 ( .a(n9006), .b(n9005), .o(n9007) );
in01f01 g05219 ( .a(n9007), .o(n9008) );
no02f01 g05220 ( .a(n9008), .b(n9004), .o(n9009) );
no02f01 g05221 ( .a(n9007), .b(n9003), .o(n9010) );
no02f01 g05222 ( .a(n9010), .b(n9009), .o(n9011) );
in01f01 g05223 ( .a(n9011), .o(n9012) );
no02f01 g05224 ( .a(n9012), .b(n8899), .o(n9013) );
no02f01 g05225 ( .a(n9013), .b(n9001), .o(n9014) );
in01f01 g05226 ( .a(n9014), .o(n9015) );
no03f01 g05227 ( .a(n9015), .b(n8990), .c(n8982), .o(n9016) );
no02f01 g05228 ( .a(n9011), .b(n8862), .o(n9017) );
no02f01 g05229 ( .a(beta_31), .b(beta_7), .o(n9018) );
in01f01 g05230 ( .a(beta_7), .o(n9019) );
no02f01 g05231 ( .a(n8765), .b(n9019), .o(n9020) );
no02f01 g05232 ( .a(n9020), .b(n9018), .o(n9021) );
in01f01 g05233 ( .a(n9021), .o(n9022) );
no02f01 g05234 ( .a(n9022), .b(n8772), .o(n9023) );
in01f01 g05235 ( .a(n8772), .o(n9024) );
no02f01 g05236 ( .a(n9021), .b(n9024), .o(n9025) );
no02f01 g05237 ( .a(n9025), .b(n9023), .o(n9026) );
in01f01 g05238 ( .a(n9026), .o(n9027) );
no03f01 g05239 ( .a(n9027), .b(n9017), .c(n9016), .o(n9028) );
ao12f01 g05240 ( .a(n8862), .b(n8999), .c(n8988), .o(n9029) );
ao12f01 g05241 ( .a(n9029), .b(n9027), .c(n9016), .o(n9030) );
oa12f01 g05242 ( .a(n9030), .b(n9028), .c(n8862), .o(n9031) );
no02f01 g05243 ( .a(n8765), .b(n8778), .o(n9032) );
no02f01 g05244 ( .a(n8781), .b(n9032), .o(n9033) );
in01f01 g05245 ( .a(n9033), .o(n9034) );
no02f01 g05246 ( .a(n9034), .b(n8777), .o(n9035) );
ao12f01 g05247 ( .a(n9033), .b(n8776), .c(n8775), .o(n9036) );
no02f01 g05248 ( .a(n9036), .b(n9035), .o(n9037) );
in01f01 g05249 ( .a(n9037), .o(n9038) );
in01f01 g05250 ( .a(n9018), .o(n9039) );
ao12f01 g05251 ( .a(n9020), .b(n9039), .c(n8772), .o(n9040) );
in01f01 g05252 ( .a(beta_8), .o(n9041) );
no02f01 g05253 ( .a(beta_31), .b(n9041), .o(n9042) );
no02f01 g05254 ( .a(n8765), .b(beta_8), .o(n9043) );
no02f01 g05255 ( .a(n9043), .b(n9042), .o(n9044) );
no02f01 g05256 ( .a(n9044), .b(n9040), .o(n9045) );
na02f01 g05257 ( .a(n9044), .b(n9040), .o(n9046) );
in01f01 g05258 ( .a(n9046), .o(n9047) );
no02f01 g05259 ( .a(n9047), .b(n9045), .o(n9048) );
in01f01 g05260 ( .a(n9048), .o(n9049) );
ao12f01 g05261 ( .a(n8862), .b(n9049), .c(n9038), .o(n9050) );
in01f01 g05262 ( .a(n9050), .o(n9051) );
no02f01 g05263 ( .a(n9032), .b(n8777), .o(n9052) );
no02f01 g05264 ( .a(n9052), .b(n8781), .o(n9053) );
in01f01 g05265 ( .a(n9053), .o(n9054) );
no02f01 g05266 ( .a(n8765), .b(n8779), .o(n9055) );
no02f01 g05267 ( .a(n9055), .b(n8782), .o(n9056) );
no02f01 g05268 ( .a(n9056), .b(n9054), .o(n9057) );
na02f01 g05269 ( .a(n9056), .b(n9054), .o(n9058) );
in01f01 g05270 ( .a(n9058), .o(n9059) );
no02f01 g05271 ( .a(n9059), .b(n9057), .o(n9060) );
in01f01 g05272 ( .a(n9060), .o(n9061) );
no02f01 g05273 ( .a(n9061), .b(n8862), .o(n9062) );
in01f01 g05274 ( .a(n9062), .o(n9063) );
na03f01 g05275 ( .a(n9063), .b(n9051), .c(n9031), .o(n9064) );
no02f01 g05276 ( .a(n9060), .b(n8899), .o(n9065) );
ao12f01 g05277 ( .a(n8899), .b(n9048), .c(n9037), .o(n9066) );
no02f01 g05278 ( .a(n9066), .b(n9065), .o(n9067) );
no02f01 g05279 ( .a(n8954), .b(n8953), .o(n9068) );
no02f01 g05280 ( .a(n9068), .b(n8784), .o(n9069) );
na02f01 g05281 ( .a(n9068), .b(n8784), .o(n9070) );
in01f01 g05282 ( .a(n9070), .o(n9071) );
no02f01 g05283 ( .a(n9071), .b(n9069), .o(n9072) );
no02f01 g05284 ( .a(n9072), .b(n8862), .o(n9073) );
in01f01 g05285 ( .a(n9073), .o(n9074) );
na03f01 g05286 ( .a(n9074), .b(n9067), .c(n9064), .o(n9075) );
na02f01 g05287 ( .a(n9072), .b(n8862), .o(n9076) );
na02f01 g05288 ( .a(n8964), .b(n8862), .o(n9077) );
na03f01 g05289 ( .a(n9077), .b(n9076), .c(n9075), .o(n9078) );
no02f01 g05290 ( .a(n8949), .b(n8899), .o(n9079) );
in01f01 g05291 ( .a(n9079), .o(n9080) );
na03f01 g05292 ( .a(n9080), .b(n9078), .c(n8966), .o(n9081) );
no02f01 g05293 ( .a(n8795), .b(n8790), .o(n9082) );
no02f01 g05294 ( .a(n8765), .b(n8792), .o(n9083) );
no02f01 g05295 ( .a(n9083), .b(n8796), .o(n9084) );
in01f01 g05296 ( .a(n9084), .o(n9085) );
no03f01 g05297 ( .a(n9085), .b(n9082), .c(n8944), .o(n9086) );
no02f01 g05298 ( .a(n9082), .b(n8944), .o(n9087) );
no02f01 g05299 ( .a(n9084), .b(n9087), .o(n9088) );
no02f01 g05300 ( .a(n9088), .b(n9086), .o(n9089) );
in01f01 g05301 ( .a(n9089), .o(n9090) );
no02f01 g05302 ( .a(n9090), .b(n8862), .o(n9091) );
in01f01 g05303 ( .a(n9091), .o(n9092) );
na03f01 g05304 ( .a(n9092), .b(n9081), .c(n8952), .o(n9093) );
in01f01 g05305 ( .a(n8799), .o(n9094) );
no02f01 g05306 ( .a(n8932), .b(n8800), .o(n9095) );
no02f01 g05307 ( .a(n9095), .b(n9094), .o(n9096) );
na02f01 g05308 ( .a(n9095), .b(n9094), .o(n9097) );
in01f01 g05309 ( .a(n9097), .o(n9098) );
no02f01 g05310 ( .a(n9098), .b(n9096), .o(n9099) );
no02f01 g05311 ( .a(n9099), .b(n8862), .o(n9100) );
no02f01 g05312 ( .a(n9089), .b(n8899), .o(n9101) );
no02f01 g05313 ( .a(n9101), .b(n9100), .o(n9102) );
na02f01 g05314 ( .a(n9102), .b(n9093), .o(n9103) );
na02f01 g05315 ( .a(n9099), .b(n8862), .o(n9104) );
in01f01 g05316 ( .a(n8930), .o(n9105) );
in01f01 g05317 ( .a(n8940), .o(n9106) );
ao12f01 g05318 ( .a(n8899), .b(n9106), .c(n9105), .o(n9107) );
in01f01 g05319 ( .a(n9107), .o(n9108) );
na03f01 g05320 ( .a(n9108), .b(n9104), .c(n9103), .o(n9109) );
no02f01 g05321 ( .a(n8765), .b(beta_19), .o(n9110) );
no02f01 g05322 ( .a(beta_31), .b(n8827), .o(n9111) );
no02f01 g05323 ( .a(n9111), .b(n9110), .o(n9112) );
in01f01 g05324 ( .a(n9112), .o(n9113) );
no02f01 g05325 ( .a(n9113), .b(n8815), .o(n9114) );
in01f01 g05326 ( .a(n8815), .o(n9115) );
no02f01 g05327 ( .a(n9112), .b(n9115), .o(n9116) );
no02f01 g05328 ( .a(n9116), .b(n9114), .o(n9117) );
in01f01 g05329 ( .a(n8805), .o(n9118) );
in01f01 g05330 ( .a(n8925), .o(n9119) );
ao12f01 g05331 ( .a(n9118), .b(n8922), .c(n9119), .o(n9120) );
no02f01 g05332 ( .a(beta_31), .b(n8811), .o(n9121) );
no02f01 g05333 ( .a(n9121), .b(n8810), .o(n9122) );
in01f01 g05334 ( .a(n9122), .o(n9123) );
no02f01 g05335 ( .a(n9123), .b(n9120), .o(n9124) );
na02f01 g05336 ( .a(n9123), .b(n9120), .o(n9125) );
in01f01 g05337 ( .a(n9125), .o(n9126) );
no02f01 g05338 ( .a(n9126), .b(n9124), .o(n9127) );
ao12f01 g05339 ( .a(n8899), .b(n9127), .c(n9117), .o(n9128) );
in01f01 g05340 ( .a(n9128), .o(n9129) );
na03f01 g05341 ( .a(n9129), .b(n9109), .c(n8942), .o(n9130) );
na02f01 g05342 ( .a(n9127), .b(n8899), .o(n9131) );
in01f01 g05343 ( .a(n9131), .o(n9132) );
in01f01 g05344 ( .a(n9117), .o(n9133) );
no02f01 g05345 ( .a(n9133), .b(n8862), .o(n9134) );
no02f01 g05346 ( .a(n9134), .b(n9132), .o(n9135) );
no02f01 g05347 ( .a(n8816), .b(n9115), .o(n9136) );
no02f01 g05348 ( .a(beta_31), .b(n8824), .o(n9137) );
no02f01 g05349 ( .a(n9137), .b(n8818), .o(n9138) );
in01f01 g05350 ( .a(n9138), .o(n9139) );
no03f01 g05351 ( .a(n9139), .b(n9136), .c(n8828), .o(n9140) );
no02f01 g05352 ( .a(n9136), .b(n8828), .o(n9141) );
no02f01 g05353 ( .a(n9138), .b(n9141), .o(n9142) );
no02f01 g05354 ( .a(n9142), .b(n9140), .o(n9143) );
in01f01 g05355 ( .a(n9143), .o(n9144) );
in01f01 g05356 ( .a(n9110), .o(n9145) );
ao12f01 g05357 ( .a(n9111), .b(n9145), .c(n8815), .o(n9146) );
in01f01 g05358 ( .a(n9146), .o(n9147) );
no02f01 g05359 ( .a(beta_31), .b(n8826), .o(n9148) );
no02f01 g05360 ( .a(n8765), .b(beta_20), .o(n9149) );
no02f01 g05361 ( .a(n9149), .b(n9148), .o(n9150) );
in01f01 g05362 ( .a(n9150), .o(n9151) );
no02f01 g05363 ( .a(n9151), .b(n9147), .o(n9152) );
no02f01 g05364 ( .a(n9150), .b(n9146), .o(n9153) );
no02f01 g05365 ( .a(n9153), .b(n9152), .o(n9154) );
no02f01 g05366 ( .a(n9154), .b(n8899), .o(n9155) );
ao12f01 g05367 ( .a(n9155), .b(n9144), .c(n8899), .o(n9156) );
in01f01 g05368 ( .a(n9156), .o(n9157) );
no02f01 g05369 ( .a(n8909), .b(n8908), .o(n9158) );
in01f01 g05370 ( .a(n9158), .o(n9159) );
no02f01 g05371 ( .a(n9159), .b(n8907), .o(n9160) );
no02f01 g05372 ( .a(n9158), .b(n8831), .o(n9161) );
no02f01 g05373 ( .a(n9161), .b(n9160), .o(n9162) );
in01f01 g05374 ( .a(n9162), .o(n9163) );
no02f01 g05375 ( .a(n9163), .b(n8862), .o(n9164) );
no03f01 g05376 ( .a(n8818), .b(n8816), .c(n9115), .o(n9165) );
no03f01 g05377 ( .a(n9165), .b(n8828), .c(n9137), .o(n9166) );
in01f01 g05378 ( .a(n9166), .o(n9167) );
no02f01 g05379 ( .a(n8765), .b(n8823), .o(n9168) );
no02f01 g05380 ( .a(n9168), .b(n8817), .o(n9169) );
in01f01 g05381 ( .a(n9169), .o(n9170) );
no02f01 g05382 ( .a(n9170), .b(n9167), .o(n9171) );
no02f01 g05383 ( .a(n9169), .b(n9166), .o(n9172) );
no02f01 g05384 ( .a(n9172), .b(n9171), .o(n9173) );
in01f01 g05385 ( .a(n9173), .o(n9174) );
no02f01 g05386 ( .a(n9174), .b(n8899), .o(n9175) );
no02f01 g05387 ( .a(n9175), .b(n9164), .o(n9176) );
na04f01 g05388 ( .a(n9176), .b(n9157), .c(n9135), .d(n9130), .o(n9177) );
ao12f01 g05389 ( .a(n9143), .b(n9154), .c(n8899), .o(n9178) );
in01f01 g05390 ( .a(n9178), .o(n9179) );
no02f01 g05391 ( .a(n9179), .b(n9175), .o(n9180) );
in01f01 g05392 ( .a(n9180), .o(n9181) );
no02f01 g05393 ( .a(n9173), .b(n8862), .o(n9182) );
no02f01 g05394 ( .a(n9162), .b(n8899), .o(n9183) );
no02f01 g05395 ( .a(n9183), .b(n9182), .o(n9184) );
ao12f01 g05396 ( .a(n9164), .b(n9184), .c(n9181), .o(n9185) );
in01f01 g05397 ( .a(n9185), .o(n9186) );
na02f01 g05398 ( .a(n9186), .b(n9177), .o(n9187) );
in01f01 g05399 ( .a(n8919), .o(n9188) );
no02f01 g05400 ( .a(n9188), .b(n8862), .o(n9189) );
in01f01 g05401 ( .a(n9189), .o(n9190) );
in01f01 g05402 ( .a(n8906), .o(n9191) );
no02f01 g05403 ( .a(n9191), .b(n8899), .o(n9192) );
in01f01 g05404 ( .a(n9192), .o(n9193) );
na04f01 g05405 ( .a(n9193), .b(n9190), .c(n9187), .d(n8896), .o(n9194) );
na02f01 g05406 ( .a(n9194), .b(n8921), .o(n9195) );
no02f01 g05407 ( .a(n8888), .b(n8847), .o(n9196) );
no02f01 g05408 ( .a(n9196), .b(n8887), .o(n9197) );
no02f01 g05409 ( .a(beta_31), .b(beta_28), .o(n9198) );
na02f01 g05410 ( .a(beta_31), .b(beta_28), .o(n9199) );
in01f01 g05411 ( .a(n9199), .o(n9200) );
no02f01 g05412 ( .a(n9200), .b(n9198), .o(n9201) );
no02f01 g05413 ( .a(n9201), .b(n9197), .o(n9202) );
na02f01 g05414 ( .a(n9201), .b(n9197), .o(n9203) );
in01f01 g05415 ( .a(n9203), .o(n9204) );
no02f01 g05416 ( .a(n9204), .b(n9202), .o(n9205) );
in01f01 g05417 ( .a(n9205), .o(n9206) );
no02f01 g05418 ( .a(n9206), .b(n8862), .o(n9207) );
in01f01 g05419 ( .a(n9207), .o(n9208) );
no02f01 g05420 ( .a(n8864), .b(n8856), .o(n9209) );
in01f01 g05421 ( .a(n9209), .o(n9210) );
no02f01 g05422 ( .a(n9210), .b(n8855), .o(n9211) );
no02f01 g05423 ( .a(n9209), .b(n8863), .o(n9212) );
no02f01 g05424 ( .a(n9212), .b(n9211), .o(n9213) );
no02f01 g05425 ( .a(n9213), .b(n8862), .o(n9214) );
no02f01 g05426 ( .a(n9205), .b(n8899), .o(n9215) );
no02f01 g05427 ( .a(n9215), .b(n9214), .o(n9216) );
in01f01 g05428 ( .a(n9216), .o(n9217) );
ao12f01 g05429 ( .a(n9217), .b(n9208), .c(n9195), .o(n9218) );
na02f01 g05430 ( .a(n9213), .b(n8862), .o(n9219) );
in01f01 g05431 ( .a(n9219), .o(n9220) );
na02f01 g05432 ( .a(n8873), .b(n8862), .o(n9221) );
in01f01 g05433 ( .a(n9221), .o(n9222) );
no03f01 g05434 ( .a(n9222), .b(n9220), .c(n9218), .o(n9223) );
no02f01 g05435 ( .a(n9223), .b(n8874), .o(n9224) );
in01f01 g05436 ( .a(n9224), .o(n9225) );
no02f01 g05437 ( .a(n9225), .b(n8862), .o(n9226) );
no02f01 g05438 ( .a(n9224), .b(n8899), .o(n9227) );
no02f01 g05439 ( .a(n9227), .b(n9226), .o(n9228) );
no02f01 g05440 ( .a(n8862), .b(n8765), .o(n9229) );
no02f01 g05441 ( .a(n8899), .b(beta_31), .o(n9230) );
no02f01 g05442 ( .a(n9230), .b(n9229), .o(n9231) );
in01f01 g05443 ( .a(n9231), .o(n9232) );
no02f01 g05444 ( .a(n9224), .b(n8765), .o(n9233) );
no02f01 g05445 ( .a(n9225), .b(beta_31), .o(n9234) );
no02f01 g05446 ( .a(n9234), .b(n9233), .o(n4201) );
no03f01 g05447 ( .a(n4201), .b(n9232), .c(n9228), .o(n9236) );
in01f01 g05448 ( .a(n9228), .o(n936) );
no02f01 g05449 ( .a(n9232), .b(n936), .o(n9238) );
no02f01 g05450 ( .a(n9231), .b(n9228), .o(n9239) );
no02f01 g05451 ( .a(n9239), .b(n9238), .o(n9240) );
no02f01 g05452 ( .a(n4201), .b(n9232), .o(n9241) );
no02f01 g05453 ( .a(n9241), .b(n9240), .o(n9242) );
no02f01 g05454 ( .a(n9242), .b(n9236), .o(n9243) );
in01f01 g05455 ( .a(n9243), .o(n233) );
in01f01 g05456 ( .a(n9103), .o(n9245) );
in01f01 g05457 ( .a(n9104), .o(n9246) );
no02f01 g05458 ( .a(n9246), .b(n9245), .o(n9247) );
no02f01 g05459 ( .a(n8940), .b(n8862), .o(n9248) );
no02f01 g05460 ( .a(n9106), .b(n8899), .o(n9249) );
in01f01 g05461 ( .a(n9249), .o(n9250) );
ao12f01 g05462 ( .a(n9248), .b(n9250), .c(n9247), .o(n9251) );
in01f01 g05463 ( .a(n9251), .o(n9252) );
no02f01 g05464 ( .a(n9105), .b(n8899), .o(n9253) );
no02f01 g05465 ( .a(n8930), .b(n8862), .o(n9254) );
no02f01 g05466 ( .a(n9254), .b(n9253), .o(n9255) );
in01f01 g05467 ( .a(n9255), .o(n9256) );
no02f01 g05468 ( .a(n9256), .b(n9252), .o(n9257) );
no02f01 g05469 ( .a(n9255), .b(n9251), .o(n9258) );
no02f01 g05470 ( .a(n9258), .b(n9257), .o(n9259) );
no02f01 g05471 ( .a(n9259), .b(n9224), .o(n9260) );
in01f01 g05472 ( .a(n9260), .o(n9261) );
in01f01 g05473 ( .a(n9247), .o(n9262) );
no02f01 g05474 ( .a(n9249), .b(n9248), .o(n9263) );
no02f01 g05475 ( .a(n9263), .b(n9262), .o(n9264) );
na02f01 g05476 ( .a(n9263), .b(n9262), .o(n9265) );
in01f01 g05477 ( .a(n9265), .o(n9266) );
no02f01 g05478 ( .a(n9266), .b(n9264), .o(n9267) );
no02f01 g05479 ( .a(n9267), .b(n9225), .o(n9268) );
in01f01 g05480 ( .a(n9081), .o(n9269) );
no02f01 g05481 ( .a(n9269), .b(n8951), .o(n9270) );
no02f01 g05482 ( .a(n9101), .b(n9270), .o(n9271) );
no02f01 g05483 ( .a(n9271), .b(n9091), .o(n9272) );
in01f01 g05484 ( .a(n9272), .o(n9273) );
no02f01 g05485 ( .a(n9246), .b(n9100), .o(n9274) );
no02f01 g05486 ( .a(n9274), .b(n9273), .o(n9275) );
na02f01 g05487 ( .a(n9274), .b(n9273), .o(n9276) );
in01f01 g05488 ( .a(n9276), .o(n9277) );
no02f01 g05489 ( .a(n9277), .b(n9275), .o(n9278) );
no02f01 g05490 ( .a(n9278), .b(n9225), .o(n9279) );
in01f01 g05491 ( .a(n9279), .o(n9280) );
in01f01 g05492 ( .a(n9270), .o(n9281) );
no02f01 g05493 ( .a(n9101), .b(n9091), .o(n9282) );
no02f01 g05494 ( .a(n9282), .b(n9281), .o(n9283) );
na02f01 g05495 ( .a(n9282), .b(n9281), .o(n9284) );
in01f01 g05496 ( .a(n9284), .o(n9285) );
no02f01 g05497 ( .a(n9285), .b(n9283), .o(n9286) );
no02f01 g05498 ( .a(n9286), .b(n9224), .o(n9287) );
in01f01 g05499 ( .a(n9078), .o(n9288) );
no02f01 g05500 ( .a(n9288), .b(n8965), .o(n9289) );
no02f01 g05501 ( .a(n9079), .b(n8951), .o(n9290) );
no02f01 g05502 ( .a(n9290), .b(n9289), .o(n9291) );
na02f01 g05503 ( .a(n9290), .b(n9289), .o(n9292) );
in01f01 g05504 ( .a(n9292), .o(n9293) );
no02f01 g05505 ( .a(n9293), .b(n9291), .o(n9294) );
no02f01 g05506 ( .a(n9294), .b(n9225), .o(n9295) );
in01f01 g05507 ( .a(n9295), .o(n9296) );
in01f01 g05508 ( .a(n9075), .o(n9297) );
in01f01 g05509 ( .a(n9076), .o(n9298) );
no02f01 g05510 ( .a(n9298), .b(n9297), .o(n9299) );
in01f01 g05511 ( .a(n9299), .o(n9300) );
in01f01 g05512 ( .a(n9077), .o(n9301) );
no02f01 g05513 ( .a(n9301), .b(n8965), .o(n9302) );
no02f01 g05514 ( .a(n9302), .b(n9300), .o(n9303) );
na02f01 g05515 ( .a(n9302), .b(n9300), .o(n9304) );
in01f01 g05516 ( .a(n9304), .o(n9305) );
no02f01 g05517 ( .a(n9305), .b(n9303), .o(n9306) );
no02f01 g05518 ( .a(n9306), .b(n9225), .o(n9307) );
in01f01 g05519 ( .a(n9064), .o(n9308) );
in01f01 g05520 ( .a(n9067), .o(n9309) );
no02f01 g05521 ( .a(n9309), .b(n9308), .o(n9310) );
no02f01 g05522 ( .a(n9298), .b(n9073), .o(n9311) );
no02f01 g05523 ( .a(n9311), .b(n9310), .o(n9312) );
na02f01 g05524 ( .a(n9311), .b(n9310), .o(n9313) );
in01f01 g05525 ( .a(n9313), .o(n9314) );
no02f01 g05526 ( .a(n9314), .b(n9312), .o(n9315) );
in01f01 g05527 ( .a(n9315), .o(n9316) );
no02f01 g05528 ( .a(n9316), .b(n9224), .o(n9317) );
no02f01 g05529 ( .a(n9048), .b(n8899), .o(n9318) );
no02f01 g05530 ( .a(n9049), .b(n8862), .o(n9319) );
in01f01 g05531 ( .a(n9319), .o(n9320) );
ao12f01 g05532 ( .a(n9318), .b(n9320), .c(n9031), .o(n9321) );
no02f01 g05533 ( .a(n9037), .b(n8899), .o(n9322) );
no02f01 g05534 ( .a(n9038), .b(n8862), .o(n9323) );
no02f01 g05535 ( .a(n9323), .b(n9322), .o(n9324) );
no02f01 g05536 ( .a(n9324), .b(n9321), .o(n9325) );
na02f01 g05537 ( .a(n9324), .b(n9321), .o(n9326) );
in01f01 g05538 ( .a(n9326), .o(n9327) );
no02f01 g05539 ( .a(n9327), .b(n9325), .o(n9328) );
no02f01 g05540 ( .a(n9328), .b(n9225), .o(n9329) );
in01f01 g05541 ( .a(n9031), .o(n9330) );
no02f01 g05542 ( .a(n9319), .b(n9318), .o(n9331) );
no02f01 g05543 ( .a(n9331), .b(n9330), .o(n9332) );
na02f01 g05544 ( .a(n9331), .b(n9330), .o(n9333) );
in01f01 g05545 ( .a(n9333), .o(n9334) );
no02f01 g05546 ( .a(n9334), .b(n9332), .o(n9335) );
no02f01 g05547 ( .a(n9335), .b(n9224), .o(n9336) );
in01f01 g05548 ( .a(n9336), .o(n9337) );
in01f01 g05549 ( .a(n8979), .o(n9338) );
no02f01 g05550 ( .a(n8980), .b(n8968), .o(n9339) );
no02f01 g05551 ( .a(n9339), .b(n9338), .o(n9340) );
na02f01 g05552 ( .a(n9339), .b(n9338), .o(n9341) );
in01f01 g05553 ( .a(n9341), .o(n9342) );
no02f01 g05554 ( .a(n9342), .b(n9340), .o(n9343) );
in01f01 g05555 ( .a(n9343), .o(n9344) );
in01f01 g05556 ( .a(n8977), .o(n9345) );
no03f01 g05557 ( .a(n8978), .b(n9345), .c(n8970), .o(n9346) );
no02f01 g05558 ( .a(n8978), .b(n8970), .o(n9347) );
no02f01 g05559 ( .a(n9347), .b(n8977), .o(n9348) );
no02f01 g05560 ( .a(n9348), .b(n9346), .o(n452) );
in01f01 g05561 ( .a(n452), .o(n9350) );
no02f01 g05562 ( .a(n9350), .b(n9344), .o(n9351) );
no03f01 g05563 ( .a(n9351), .b(n9223), .c(n8874), .o(n9352) );
no02f01 g05564 ( .a(n452), .b(n9343), .o(n9353) );
no02f01 g05565 ( .a(n8988), .b(n8862), .o(n9354) );
no02f01 g05566 ( .a(n9354), .b(n8990), .o(n9355) );
no02f01 g05567 ( .a(n9355), .b(n8982), .o(n9356) );
na02f01 g05568 ( .a(n9355), .b(n8982), .o(n9357) );
in01f01 g05569 ( .a(n9357), .o(n9358) );
no02f01 g05570 ( .a(n9358), .b(n9356), .o(n9359) );
no02f01 g05571 ( .a(n8990), .b(n8982), .o(n9360) );
no02f01 g05572 ( .a(n9354), .b(n9360), .o(n9361) );
no02f01 g05573 ( .a(n8999), .b(n8862), .o(n9362) );
no02f01 g05574 ( .a(n9362), .b(n9001), .o(n9363) );
no02f01 g05575 ( .a(n9363), .b(n9361), .o(n9364) );
na02f01 g05576 ( .a(n9363), .b(n9361), .o(n9365) );
in01f01 g05577 ( .a(n9365), .o(n9366) );
no02f01 g05578 ( .a(n9366), .b(n9364), .o(n9367) );
oa22f01 g05579 ( .a(n9367), .b(n9359), .c(n9223), .d(n8874), .o(n9368) );
oa12f01 g05580 ( .a(n9368), .b(n9353), .c(n9352), .o(n9369) );
in01f01 g05581 ( .a(n9359), .o(n9370) );
in01f01 g05582 ( .a(n9367), .o(n9371) );
oa12f01 g05583 ( .a(n9224), .b(n9371), .c(n9370), .o(n9372) );
in01f01 g05584 ( .a(n9001), .o(n9373) );
ao12f01 g05585 ( .a(n9029), .b(n9373), .c(n9360), .o(n9374) );
no02f01 g05586 ( .a(n9017), .b(n9013), .o(n9375) );
no02f01 g05587 ( .a(n9375), .b(n9374), .o(n9376) );
na02f01 g05588 ( .a(n9375), .b(n9374), .o(n9377) );
in01f01 g05589 ( .a(n9377), .o(n9378) );
no02f01 g05590 ( .a(n9378), .b(n9376), .o(n9379) );
in01f01 g05591 ( .a(n9379), .o(n9380) );
no02f01 g05592 ( .a(n9380), .b(n9224), .o(n9381) );
no02f01 g05593 ( .a(n9017), .b(n9016), .o(n9382) );
in01f01 g05594 ( .a(n9029), .o(n9383) );
na02f01 g05595 ( .a(n9383), .b(n9382), .o(n9384) );
in01f01 g05596 ( .a(n9384), .o(n9385) );
no02f01 g05597 ( .a(n9027), .b(n8899), .o(n9386) );
no02f01 g05598 ( .a(n9026), .b(n8862), .o(n9387) );
no02f01 g05599 ( .a(n9387), .b(n9386), .o(n9388) );
no02f01 g05600 ( .a(n9388), .b(n9385), .o(n9389) );
na02f01 g05601 ( .a(n9388), .b(n9385), .o(n9390) );
in01f01 g05602 ( .a(n9390), .o(n9391) );
no02f01 g05603 ( .a(n9391), .b(n9389), .o(n9392) );
in01f01 g05604 ( .a(n9392), .o(n9393) );
no02f01 g05605 ( .a(n9393), .b(n9224), .o(n9394) );
no02f01 g05606 ( .a(n9394), .b(n9381), .o(n9395) );
in01f01 g05607 ( .a(n9395), .o(n9396) );
ao12f01 g05608 ( .a(n9396), .b(n9372), .c(n9369), .o(n9397) );
no02f01 g05609 ( .a(n9379), .b(n9225), .o(n9398) );
no02f01 g05610 ( .a(n9392), .b(n9225), .o(n9399) );
no02f01 g05611 ( .a(n9399), .b(n9398), .o(n9400) );
in01f01 g05612 ( .a(n9400), .o(n9401) );
na02f01 g05613 ( .a(n9335), .b(n9224), .o(n9402) );
oa12f01 g05614 ( .a(n9402), .b(n9401), .c(n9397), .o(n9403) );
na02f01 g05615 ( .a(n9328), .b(n9225), .o(n9404) );
in01f01 g05616 ( .a(n9404), .o(n9405) );
ao12f01 g05617 ( .a(n9405), .b(n9403), .c(n9337), .o(n9406) );
ao12f01 g05618 ( .a(n9066), .b(n9051), .c(n9031), .o(n9407) );
in01f01 g05619 ( .a(n9407), .o(n9408) );
no02f01 g05620 ( .a(n9065), .b(n9062), .o(n9409) );
in01f01 g05621 ( .a(n9409), .o(n9410) );
no02f01 g05622 ( .a(n9410), .b(n9408), .o(n9411) );
no02f01 g05623 ( .a(n9409), .b(n9407), .o(n9412) );
no02f01 g05624 ( .a(n9412), .b(n9411), .o(n9413) );
in01f01 g05625 ( .a(n9413), .o(n9414) );
no02f01 g05626 ( .a(n9414), .b(n9225), .o(n9415) );
in01f01 g05627 ( .a(n9415), .o(n9416) );
oa12f01 g05628 ( .a(n9416), .b(n9406), .c(n9329), .o(n9417) );
no02f01 g05629 ( .a(n9414), .b(n9224), .o(n9418) );
ao12f01 g05630 ( .a(n9418), .b(n9315), .c(n9224), .o(n9419) );
in01f01 g05631 ( .a(n9419), .o(n9420) );
ao12f01 g05632 ( .a(n9317), .b(n9420), .c(n9417), .o(n9421) );
na02f01 g05633 ( .a(n9306), .b(n9225), .o(n9422) );
ao12f01 g05634 ( .a(n9307), .b(n9422), .c(n9421), .o(n9423) );
na02f01 g05635 ( .a(n9294), .b(n9225), .o(n9424) );
in01f01 g05636 ( .a(n9424), .o(n9425) );
oa12f01 g05637 ( .a(n9296), .b(n9425), .c(n9423), .o(n9426) );
na02f01 g05638 ( .a(n9286), .b(n9224), .o(n9427) );
ao12f01 g05639 ( .a(n9287), .b(n9427), .c(n9426), .o(n9428) );
na02f01 g05640 ( .a(n9278), .b(n9225), .o(n9429) );
in01f01 g05641 ( .a(n9429), .o(n9430) );
oa12f01 g05642 ( .a(n9280), .b(n9430), .c(n9428), .o(n9431) );
na02f01 g05643 ( .a(n9267), .b(n9225), .o(n9432) );
ao12f01 g05644 ( .a(n9268), .b(n9432), .c(n9431), .o(n9433) );
na02f01 g05645 ( .a(n9259), .b(n9224), .o(n9434) );
in01f01 g05646 ( .a(n9434), .o(n9435) );
oa12f01 g05647 ( .a(n9261), .b(n9435), .c(n9433), .o(n9436) );
in01f01 g05648 ( .a(n9109), .o(n9437) );
no02f01 g05649 ( .a(n9437), .b(n8941), .o(n9438) );
in01f01 g05650 ( .a(n9438), .o(n9439) );
no02f01 g05651 ( .a(n9127), .b(n8899), .o(n9440) );
ao12f01 g05652 ( .a(n9440), .b(n9131), .c(n9439), .o(n9441) );
no02f01 g05653 ( .a(n9117), .b(n8899), .o(n9442) );
no02f01 g05654 ( .a(n9442), .b(n9134), .o(n9443) );
no02f01 g05655 ( .a(n9443), .b(n9441), .o(n9444) );
na02f01 g05656 ( .a(n9443), .b(n9441), .o(n9445) );
in01f01 g05657 ( .a(n9445), .o(n9446) );
no02f01 g05658 ( .a(n9446), .b(n9444), .o(n9447) );
in01f01 g05659 ( .a(n9447), .o(n9448) );
no02f01 g05660 ( .a(n9132), .b(n9440), .o(n9449) );
in01f01 g05661 ( .a(n9449), .o(n9450) );
no02f01 g05662 ( .a(n9450), .b(n9439), .o(n9451) );
no02f01 g05663 ( .a(n9449), .b(n9438), .o(n9452) );
no02f01 g05664 ( .a(n9452), .b(n9451), .o(n9453) );
in01f01 g05665 ( .a(n9453), .o(n9454) );
ao12f01 g05666 ( .a(n9224), .b(n9454), .c(n9448), .o(n9455) );
in01f01 g05667 ( .a(n9455), .o(n9456) );
in01f01 g05668 ( .a(n9130), .o(n9457) );
in01f01 g05669 ( .a(n9135), .o(n9458) );
no02f01 g05670 ( .a(n9458), .b(n9457), .o(n9459) );
no02f01 g05671 ( .a(n9154), .b(n8862), .o(n9460) );
na02f01 g05672 ( .a(n9154), .b(n8862), .o(n9461) );
in01f01 g05673 ( .a(n9461), .o(n9462) );
no02f01 g05674 ( .a(n9462), .b(n9460), .o(n9463) );
in01f01 g05675 ( .a(n9463), .o(n9464) );
no02f01 g05676 ( .a(n9464), .b(n9459), .o(n9465) );
no03f01 g05677 ( .a(n9463), .b(n9458), .c(n9457), .o(n9466) );
no02f01 g05678 ( .a(n9466), .b(n9465), .o(n9467) );
in01f01 g05679 ( .a(n9467), .o(n9468) );
no02f01 g05680 ( .a(n9468), .b(n9225), .o(n9469) );
ao12f01 g05681 ( .a(n9460), .b(n9461), .c(n9459), .o(n9470) );
no02f01 g05682 ( .a(n9143), .b(n8899), .o(n9471) );
no02f01 g05683 ( .a(n9144), .b(n8862), .o(n9472) );
no02f01 g05684 ( .a(n9472), .b(n9471), .o(n9473) );
no02f01 g05685 ( .a(n9473), .b(n9470), .o(n9474) );
na02f01 g05686 ( .a(n9473), .b(n9470), .o(n9475) );
in01f01 g05687 ( .a(n9475), .o(n9476) );
no02f01 g05688 ( .a(n9476), .b(n9474), .o(n9477) );
in01f01 g05689 ( .a(n9477), .o(n9478) );
no02f01 g05690 ( .a(n9478), .b(n9224), .o(n9479) );
no02f01 g05691 ( .a(n9479), .b(n9469), .o(n9480) );
na03f01 g05692 ( .a(n9480), .b(n9456), .c(n9436), .o(n9481) );
no02f01 g05693 ( .a(n9454), .b(n9448), .o(n9482) );
no03f01 g05694 ( .a(n9482), .b(n9467), .c(n9225), .o(n9483) );
no02f01 g05695 ( .a(n9477), .b(n9225), .o(n9484) );
no02f01 g05696 ( .a(n9467), .b(n9224), .o(n9485) );
no03f01 g05697 ( .a(n9485), .b(n9484), .c(n9483), .o(n9486) );
no02f01 g05698 ( .a(n9486), .b(n9479), .o(n9487) );
in01f01 g05699 ( .a(n9487), .o(n9488) );
in01f01 g05700 ( .a(n9182), .o(n9489) );
ao12f01 g05701 ( .a(n9178), .b(n9157), .c(n9459), .o(n9490) );
ao12f01 g05702 ( .a(n9175), .b(n9490), .c(n9489), .o(n9491) );
no02f01 g05703 ( .a(n9183), .b(n9164), .o(n9492) );
in01f01 g05704 ( .a(n9492), .o(n9493) );
no02f01 g05705 ( .a(n9493), .b(n9491), .o(n9494) );
na02f01 g05706 ( .a(n9493), .b(n9491), .o(n9495) );
in01f01 g05707 ( .a(n9495), .o(n9496) );
no02f01 g05708 ( .a(n9496), .b(n9494), .o(n9497) );
no02f01 g05709 ( .a(n9497), .b(n9224), .o(n9498) );
no02f01 g05710 ( .a(n9182), .b(n9175), .o(n9499) );
no02f01 g05711 ( .a(n9499), .b(n9490), .o(n9500) );
na02f01 g05712 ( .a(n9499), .b(n9490), .o(n9501) );
in01f01 g05713 ( .a(n9501), .o(n9502) );
no02f01 g05714 ( .a(n9502), .b(n9500), .o(n9503) );
no02f01 g05715 ( .a(n9503), .b(n9225), .o(n9504) );
no02f01 g05716 ( .a(n9504), .b(n9498), .o(n9505) );
ao12f01 g05717 ( .a(n9505), .b(n9488), .c(n9481), .o(n9506) );
in01f01 g05718 ( .a(n9187), .o(n9507) );
no02f01 g05719 ( .a(n8919), .b(n8899), .o(n9508) );
no02f01 g05720 ( .a(n9508), .b(n9189), .o(n9509) );
no02f01 g05721 ( .a(n9509), .b(n9507), .o(n9510) );
na02f01 g05722 ( .a(n9509), .b(n9507), .o(n9511) );
in01f01 g05723 ( .a(n9511), .o(n9512) );
no02f01 g05724 ( .a(n9512), .b(n9510), .o(n9513) );
in01f01 g05725 ( .a(n9513), .o(n9514) );
no02f01 g05726 ( .a(n9514), .b(n9224), .o(n9515) );
no02f01 g05727 ( .a(n9189), .b(n9507), .o(n9516) );
no02f01 g05728 ( .a(n9508), .b(n9516), .o(n9517) );
no02f01 g05729 ( .a(n8906), .b(n8862), .o(n9518) );
no02f01 g05730 ( .a(n9518), .b(n9192), .o(n9519) );
no02f01 g05731 ( .a(n9519), .b(n9517), .o(n9520) );
na02f01 g05732 ( .a(n9519), .b(n9517), .o(n9521) );
in01f01 g05733 ( .a(n9521), .o(n9522) );
no02f01 g05734 ( .a(n9522), .b(n9520), .o(n9523) );
in01f01 g05735 ( .a(n9523), .o(n9524) );
no02f01 g05736 ( .a(n9524), .b(n9224), .o(n9525) );
no02f01 g05737 ( .a(n9525), .b(n9515), .o(n9526) );
in01f01 g05738 ( .a(n9525), .o(n9527) );
ao12f01 g05739 ( .a(n9497), .b(n9503), .c(n9225), .o(n9528) );
in01f01 g05740 ( .a(n9528), .o(n9529) );
no02f01 g05741 ( .a(n9513), .b(n9225), .o(n9530) );
no02f01 g05742 ( .a(n9523), .b(n9225), .o(n9531) );
no02f01 g05743 ( .a(n9531), .b(n9530), .o(n9532) );
oa12f01 g05744 ( .a(n9532), .b(n9529), .c(n9515), .o(n9533) );
na02f01 g05745 ( .a(n9533), .b(n9527), .o(n9534) );
in01f01 g05746 ( .a(n9534), .o(n9535) );
ao12f01 g05747 ( .a(n9535), .b(n9526), .c(n9506), .o(n9536) );
ao12f01 g05748 ( .a(n8920), .b(n9193), .c(n9516), .o(n9537) );
in01f01 g05749 ( .a(n9537), .o(n9538) );
no02f01 g05750 ( .a(n8900), .b(n8899), .o(n9539) );
no02f01 g05751 ( .a(n9539), .b(n8886), .o(n9540) );
in01f01 g05752 ( .a(n9540), .o(n9541) );
no02f01 g05753 ( .a(n9541), .b(n9538), .o(n9542) );
no02f01 g05754 ( .a(n9540), .b(n9537), .o(n9543) );
no02f01 g05755 ( .a(n9543), .b(n9542), .o(n9544) );
in01f01 g05756 ( .a(n9544), .o(n9545) );
no02f01 g05757 ( .a(n9545), .b(n9224), .o(n9546) );
in01f01 g05758 ( .a(n9539), .o(n9547) );
ao12f01 g05759 ( .a(n8886), .b(n9537), .c(n9547), .o(n9548) );
in01f01 g05760 ( .a(n9548), .o(n9549) );
no02f01 g05761 ( .a(n8893), .b(n8899), .o(n9550) );
no02f01 g05762 ( .a(n9550), .b(n8895), .o(n9551) );
no02f01 g05763 ( .a(n9551), .b(n9549), .o(n9552) );
na02f01 g05764 ( .a(n9551), .b(n9549), .o(n9553) );
in01f01 g05765 ( .a(n9553), .o(n9554) );
no02f01 g05766 ( .a(n9554), .b(n9552), .o(n9555) );
in01f01 g05767 ( .a(n9555), .o(n9556) );
no02f01 g05768 ( .a(n9556), .b(n9224), .o(n9557) );
no02f01 g05769 ( .a(n9215), .b(n9195), .o(n9558) );
no02f01 g05770 ( .a(n9558), .b(n9207), .o(n9559) );
no02f01 g05771 ( .a(n9220), .b(n9214), .o(n9560) );
in01f01 g05772 ( .a(n9560), .o(n9561) );
no02f01 g05773 ( .a(n9561), .b(n9559), .o(n9562) );
na02f01 g05774 ( .a(n9561), .b(n9559), .o(n9563) );
in01f01 g05775 ( .a(n9563), .o(n9564) );
no03f01 g05776 ( .a(n9564), .b(n9562), .c(n9225), .o(n9565) );
in01f01 g05777 ( .a(n9195), .o(n9566) );
no02f01 g05778 ( .a(n9215), .b(n9207), .o(n9567) );
no02f01 g05779 ( .a(n9567), .b(n9566), .o(n9568) );
na02f01 g05780 ( .a(n9567), .b(n9566), .o(n9569) );
in01f01 g05781 ( .a(n9569), .o(n9570) );
no02f01 g05782 ( .a(n9570), .b(n9568), .o(n9571) );
in01f01 g05783 ( .a(n9571), .o(n9572) );
no02f01 g05784 ( .a(n9572), .b(n9225), .o(n9573) );
no02f01 g05785 ( .a(n9573), .b(n9565), .o(n9574) );
in01f01 g05786 ( .a(n9574), .o(n9575) );
no02f01 g05787 ( .a(n9575), .b(n9557), .o(n9576) );
in01f01 g05788 ( .a(n9576), .o(n9577) );
no03f01 g05789 ( .a(n9577), .b(n9546), .c(n9536), .o(n9578) );
ao12f01 g05790 ( .a(n9225), .b(n9555), .c(n9544), .o(n9579) );
in01f01 g05791 ( .a(n9579), .o(n9580) );
no02f01 g05792 ( .a(n9571), .b(n9224), .o(n9581) );
in01f01 g05793 ( .a(n9562), .o(n9582) );
ao12f01 g05794 ( .a(n9224), .b(n9563), .c(n9582), .o(n9583) );
no02f01 g05795 ( .a(n9583), .b(n9581), .o(n9584) );
oa12f01 g05796 ( .a(n9584), .b(n9580), .c(n9575), .o(n9585) );
no02f01 g05797 ( .a(n9220), .b(n9218), .o(n9586) );
no03f01 g05798 ( .a(n9221), .b(n9586), .c(n8874), .o(n9587) );
in01f01 g05799 ( .a(n9587), .o(n9588) );
oa12f01 g05800 ( .a(n9588), .b(n9585), .c(n9578), .o(n9589) );
na02f01 g05801 ( .a(n9586), .b(n8874), .o(n9590) );
in01f01 g05802 ( .a(n4201), .o(n9591) );
no02f01 g05803 ( .a(n9231), .b(n9224), .o(n9592) );
no02f01 g05804 ( .a(n9232), .b(n9225), .o(n9593) );
no02f01 g05805 ( .a(n9593), .b(n9592), .o(n9594) );
in01f01 g05806 ( .a(n9594), .o(n9595) );
no02f01 g05807 ( .a(n9224), .b(n8862), .o(n9596) );
no03f01 g05808 ( .a(n9596), .b(n9595), .c(n9234), .o(n9597) );
ao12f01 g05809 ( .a(n8899), .b(n9225), .c(n8765), .o(n9598) );
no02f01 g05810 ( .a(n9598), .b(n9597), .o(n9599) );
no02f01 g05811 ( .a(n9594), .b(n8765), .o(n9600) );
no04f01 g05812 ( .a(n9600), .b(n9599), .c(n9591), .d(n9226), .o(n9601) );
ao12f01 g05813 ( .a(n9224), .b(n8862), .c(n8765), .o(n9602) );
no03f01 g05814 ( .a(n9602), .b(n9234), .c(n9227), .o(n9603) );
no02f01 g05815 ( .a(n9603), .b(n9233), .o(n9604) );
no02f01 g05816 ( .a(n9604), .b(n9601), .o(n9605) );
in01f01 g05817 ( .a(n9605), .o(n9606) );
no02f01 g05818 ( .a(n9595), .b(n8765), .o(n9607) );
no02f01 g05819 ( .a(n9594), .b(beta_31), .o(n9608) );
no02f01 g05820 ( .a(n9608), .b(n9607), .o(n9609) );
in01f01 g05821 ( .a(n9609), .o(n9610) );
no02f01 g05822 ( .a(n9610), .b(n9606), .o(n9611) );
no02f01 g05823 ( .a(n9609), .b(n9605), .o(n9612) );
no02f01 g05824 ( .a(n9612), .b(n9611), .o(n9613) );
na03f01 g05825 ( .a(n9613), .b(n9590), .c(n9589), .o(n9614) );
in01f01 g05826 ( .a(n9268), .o(n9615) );
in01f01 g05827 ( .a(n9287), .o(n9616) );
in01f01 g05828 ( .a(n9307), .o(n9617) );
in01f01 g05829 ( .a(n9317), .o(n9618) );
in01f01 g05830 ( .a(n9329), .o(n9619) );
in01f01 g05831 ( .a(n9369), .o(n9620) );
in01f01 g05832 ( .a(n9372), .o(n9621) );
oa12f01 g05833 ( .a(n9395), .b(n9621), .c(n9620), .o(n9622) );
in01f01 g05834 ( .a(n9402), .o(n9623) );
ao12f01 g05835 ( .a(n9623), .b(n9400), .c(n9622), .o(n9624) );
oa12f01 g05836 ( .a(n9404), .b(n9624), .c(n9336), .o(n9625) );
ao12f01 g05837 ( .a(n9415), .b(n9625), .c(n9619), .o(n9626) );
oa12f01 g05838 ( .a(n9618), .b(n9419), .c(n9626), .o(n9627) );
in01f01 g05839 ( .a(n9422), .o(n9628) );
oa12f01 g05840 ( .a(n9617), .b(n9628), .c(n9627), .o(n9629) );
ao12f01 g05841 ( .a(n9295), .b(n9424), .c(n9629), .o(n9630) );
in01f01 g05842 ( .a(n9427), .o(n9631) );
oa12f01 g05843 ( .a(n9616), .b(n9631), .c(n9630), .o(n9632) );
ao12f01 g05844 ( .a(n9279), .b(n9429), .c(n9632), .o(n9633) );
in01f01 g05845 ( .a(n9432), .o(n9634) );
oa12f01 g05846 ( .a(n9615), .b(n9634), .c(n9633), .o(n9635) );
ao12f01 g05847 ( .a(n9260), .b(n9434), .c(n9635), .o(n9636) );
in01f01 g05848 ( .a(n9480), .o(n9637) );
no03f01 g05849 ( .a(n9637), .b(n9455), .c(n9636), .o(n9638) );
oa22f01 g05850 ( .a(n9504), .b(n9498), .c(n9487), .d(n9638), .o(n9639) );
in01f01 g05851 ( .a(n9526), .o(n9640) );
oa12f01 g05852 ( .a(n9534), .b(n9640), .c(n9639), .o(n9641) );
in01f01 g05853 ( .a(n9546), .o(n9642) );
na03f01 g05854 ( .a(n9576), .b(n9642), .c(n9641), .o(n9643) );
in01f01 g05855 ( .a(n9585), .o(n9644) );
ao12f01 g05856 ( .a(n9587), .b(n9644), .c(n9643), .o(n9645) );
in01f01 g05857 ( .a(n9590), .o(n9646) );
in01f01 g05858 ( .a(n9613), .o(n2102) );
oa12f01 g05859 ( .a(n2102), .b(n9646), .c(n9645), .o(n9648) );
na02f01 g05860 ( .a(n9648), .b(n9614), .o(n238) );
no02f01 g05861 ( .a(n6836), .b(n6814), .o(n9650) );
ao12f01 g05862 ( .a(n6895), .b(n6854), .c(n9650), .o(n9651) );
in01f01 g05863 ( .a(n9651), .o(n9652) );
ao12f01 g05864 ( .a(n6899), .b(n9652), .c(n6875), .o(n9653) );
no02f01 g05865 ( .a(n6896), .b(n4043), .o(n9654) );
no02f01 g05866 ( .a(n9654), .b(n6885), .o(n9655) );
no02f01 g05867 ( .a(n9655), .b(n9653), .o(n9656) );
na02f01 g05868 ( .a(n9655), .b(n9653), .o(n9657) );
in01f01 g05869 ( .a(n9657), .o(n9658) );
no02f01 g05870 ( .a(n9658), .b(n9656), .o(n9659) );
in01f01 g05871 ( .a(n6664), .o(n9660) );
no02f01 g05872 ( .a(n7017), .b(n6565), .o(n9661) );
oa12f01 g05873 ( .a(n9661), .b(n6666), .c(n9660), .o(n9662) );
in01f01 g05874 ( .a(n9662), .o(n9663) );
no02f01 g05875 ( .a(n6581), .b(n4043), .o(n9664) );
no02f01 g05876 ( .a(n9664), .b(n6584), .o(n9665) );
no02f01 g05877 ( .a(n9665), .b(n9663), .o(n9666) );
na02f01 g05878 ( .a(n9665), .b(n9663), .o(n9667) );
in01f01 g05879 ( .a(n9667), .o(n9668) );
no02f01 g05880 ( .a(n9668), .b(n9666), .o(n9669) );
in01f01 g05881 ( .a(n9669), .o(n9670) );
ao12f01 g05882 ( .a(n6934), .b(n9670), .c(n7024), .o(n9671) );
in01f01 g05883 ( .a(n9671), .o(n9672) );
na02f01 g05884 ( .a(n9672), .b(n7014), .o(n9673) );
in01f01 g05885 ( .a(n9673), .o(n9674) );
oa12f01 g05886 ( .a(n9674), .b(n6988), .c(n6984), .o(n9675) );
in01f01 g05887 ( .a(n7015), .o(n9676) );
oa12f01 g05888 ( .a(n6934), .b(n9670), .c(n7024), .o(n9677) );
ao12f01 g05889 ( .a(n9671), .b(n9677), .c(n9676), .o(n9678) );
in01f01 g05890 ( .a(n9678), .o(n9679) );
no02f01 g05891 ( .a(n6677), .b(n4043), .o(n9680) );
no02f01 g05892 ( .a(n6679), .b(n6668), .o(n9681) );
no02f01 g05893 ( .a(n9681), .b(n9680), .o(n9682) );
no02f01 g05894 ( .a(n6688), .b(n4043), .o(n9683) );
no02f01 g05895 ( .a(n9683), .b(n6690), .o(n9684) );
no02f01 g05896 ( .a(n9684), .b(n9682), .o(n9685) );
na02f01 g05897 ( .a(n9684), .b(n9682), .o(n9686) );
in01f01 g05898 ( .a(n9686), .o(n9687) );
no02f01 g05899 ( .a(n9687), .b(n9685), .o(n9688) );
in01f01 g05900 ( .a(n6668), .o(n9689) );
no02f01 g05901 ( .a(n9680), .b(n6679), .o(n9690) );
in01f01 g05902 ( .a(n9690), .o(n9691) );
no02f01 g05903 ( .a(n9691), .b(n9689), .o(n9692) );
no02f01 g05904 ( .a(n9690), .b(n6668), .o(n9693) );
no02f01 g05905 ( .a(n9693), .b(n9692), .o(n9694) );
no02f01 g05906 ( .a(n9694), .b(n9688), .o(n9695) );
no02f01 g05907 ( .a(n9695), .b(n6934), .o(n9696) );
ao12f01 g05908 ( .a(n9696), .b(n9679), .c(n9675), .o(n9697) );
ao12f01 g05909 ( .a(n6718), .b(n6691), .c(n9689), .o(n9698) );
in01f01 g05910 ( .a(n9698), .o(n9699) );
no02f01 g05911 ( .a(n6702), .b(n4043), .o(n9700) );
no02f01 g05912 ( .a(n9700), .b(n6704), .o(n9701) );
in01f01 g05913 ( .a(n9701), .o(n9702) );
no02f01 g05914 ( .a(n9702), .b(n9699), .o(n9703) );
no02f01 g05915 ( .a(n9701), .b(n9698), .o(n9704) );
no02f01 g05916 ( .a(n9704), .b(n9703), .o(n9705) );
in01f01 g05917 ( .a(n9705), .o(n9706) );
no02f01 g05918 ( .a(n9706), .b(n6934), .o(n9707) );
in01f01 g05919 ( .a(n9700), .o(n9708) );
ao12f01 g05920 ( .a(n6704), .b(n9698), .c(n9708), .o(n9709) );
no02f01 g05921 ( .a(n6713), .b(n4043), .o(n9710) );
no02f01 g05922 ( .a(n9710), .b(n6715), .o(n9711) );
in01f01 g05923 ( .a(n9711), .o(n9712) );
no02f01 g05924 ( .a(n9712), .b(n9709), .o(n9713) );
na02f01 g05925 ( .a(n9712), .b(n9709), .o(n9714) );
in01f01 g05926 ( .a(n9714), .o(n9715) );
no02f01 g05927 ( .a(n9715), .b(n9713), .o(n9716) );
in01f01 g05928 ( .a(n9716), .o(n9717) );
no02f01 g05929 ( .a(n9717), .b(n6934), .o(n9718) );
no02f01 g05930 ( .a(n9718), .b(n9707), .o(n9719) );
ao12f01 g05931 ( .a(n5001), .b(n9694), .c(n9688), .o(n9720) );
ao12f01 g05932 ( .a(n5001), .b(n9716), .c(n9705), .o(n9721) );
no02f01 g05933 ( .a(n9721), .b(n9720), .o(n9722) );
in01f01 g05934 ( .a(n9722), .o(n9723) );
ao12f01 g05935 ( .a(n9723), .b(n9719), .c(n9697), .o(n9724) );
no02f01 g05936 ( .a(n6720), .b(n6716), .o(n9725) );
in01f01 g05937 ( .a(n9725), .o(n9726) );
in01f01 g05938 ( .a(n6738), .o(n9727) );
no02f01 g05939 ( .a(n6736), .b(n4043), .o(n9728) );
ao12f01 g05940 ( .a(n9728), .b(n9727), .c(n9726), .o(n9729) );
in01f01 g05941 ( .a(n9729), .o(n9730) );
no02f01 g05942 ( .a(n6764), .b(n4043), .o(n9731) );
no02f01 g05943 ( .a(n9731), .b(n6731), .o(n9732) );
in01f01 g05944 ( .a(n9732), .o(n9733) );
no02f01 g05945 ( .a(n9733), .b(n9730), .o(n9734) );
no02f01 g05946 ( .a(n9732), .b(n9729), .o(n9735) );
no02f01 g05947 ( .a(n9735), .b(n9734), .o(n9736) );
in01f01 g05948 ( .a(n9736), .o(n9737) );
no02f01 g05949 ( .a(n9737), .b(n6934), .o(n9738) );
no02f01 g05950 ( .a(n9728), .b(n6738), .o(n9739) );
no02f01 g05951 ( .a(n9739), .b(n9725), .o(n9740) );
na02f01 g05952 ( .a(n9739), .b(n9725), .o(n9741) );
in01f01 g05953 ( .a(n9741), .o(n9742) );
no02f01 g05954 ( .a(n9742), .b(n9740), .o(n9743) );
in01f01 g05955 ( .a(n9743), .o(n9744) );
no02f01 g05956 ( .a(n9744), .b(n6934), .o(n9745) );
no02f01 g05957 ( .a(n9745), .b(n9738), .o(n9746) );
in01f01 g05958 ( .a(n9746), .o(n9747) );
no02f01 g05959 ( .a(n6762), .b(n4043), .o(n9748) );
no02f01 g05960 ( .a(n6765), .b(n9748), .o(n9749) );
oa12f01 g05961 ( .a(n9749), .b(n6758), .c(n6740), .o(n9750) );
no02f01 g05962 ( .a(n6761), .b(n4043), .o(n9751) );
no02f01 g05963 ( .a(n9751), .b(n6752), .o(n9752) );
in01f01 g05964 ( .a(n9752), .o(n9753) );
no02f01 g05965 ( .a(n9753), .b(n9750), .o(n9754) );
na02f01 g05966 ( .a(n9753), .b(n9750), .o(n9755) );
in01f01 g05967 ( .a(n9755), .o(n9756) );
no02f01 g05968 ( .a(n9756), .b(n9754), .o(n9757) );
in01f01 g05969 ( .a(n9757), .o(n9758) );
no02f01 g05970 ( .a(n9758), .b(n6934), .o(n9759) );
in01f01 g05971 ( .a(n6740), .o(n9760) );
no02f01 g05972 ( .a(n9748), .b(n6758), .o(n9761) );
in01f01 g05973 ( .a(n9761), .o(n9762) );
no03f01 g05974 ( .a(n9762), .b(n6765), .c(n9760), .o(n9763) );
in01f01 g05975 ( .a(n6765), .o(n9764) );
ao12f01 g05976 ( .a(n9761), .b(n9764), .c(n6740), .o(n9765) );
no02f01 g05977 ( .a(n9765), .b(n9763), .o(n9766) );
in01f01 g05978 ( .a(n9766), .o(n9767) );
no02f01 g05979 ( .a(n9767), .b(n6934), .o(n9768) );
no02f01 g05980 ( .a(n9768), .b(n9759), .o(n9769) );
in01f01 g05981 ( .a(n9769), .o(n9770) );
no03f01 g05982 ( .a(n9770), .b(n9747), .c(n9724), .o(n9771) );
ao12f01 g05983 ( .a(n5001), .b(n9766), .c(n9757), .o(n9772) );
ao12f01 g05984 ( .a(n5001), .b(n9743), .c(n9736), .o(n9773) );
no02f01 g05985 ( .a(n9773), .b(n9772), .o(n9774) );
in01f01 g05986 ( .a(n9774), .o(n9775) );
no02f01 g05987 ( .a(n6775), .b(n4043), .o(n9776) );
in01f01 g05988 ( .a(n9776), .o(n9777) );
in01f01 g05989 ( .a(n6777), .o(n9778) );
na03f01 g05990 ( .a(n9778), .b(n6759), .c(n9760), .o(n9779) );
na03f01 g05991 ( .a(n9779), .b(n9777), .c(n6766), .o(n9780) );
in01f01 g05992 ( .a(n9780), .o(n9781) );
no02f01 g05993 ( .a(n6810), .b(n4043), .o(n9782) );
no02f01 g05994 ( .a(n9782), .b(n6786), .o(n9783) );
no02f01 g05995 ( .a(n9783), .b(n9781), .o(n9784) );
na02f01 g05996 ( .a(n9783), .b(n9781), .o(n9785) );
in01f01 g05997 ( .a(n9785), .o(n9786) );
no03f01 g05998 ( .a(n9786), .b(n9784), .c(n6934), .o(n9787) );
in01f01 g05999 ( .a(n6767), .o(n9788) );
no02f01 g06000 ( .a(n9776), .b(n6777), .o(n9789) );
no02f01 g06001 ( .a(n9789), .b(n9788), .o(n9790) );
na02f01 g06002 ( .a(n9789), .b(n9788), .o(n9791) );
in01f01 g06003 ( .a(n9791), .o(n9792) );
no02f01 g06004 ( .a(n9792), .b(n9790), .o(n9793) );
in01f01 g06005 ( .a(n9793), .o(n9794) );
no02f01 g06006 ( .a(n9794), .b(n6934), .o(n9795) );
no02f01 g06007 ( .a(n9795), .b(n9787), .o(n9796) );
in01f01 g06008 ( .a(n9796), .o(n9797) );
no02f01 g06009 ( .a(n6808), .b(n4043), .o(n9798) );
in01f01 g06010 ( .a(n9798), .o(n9799) );
ao12f01 g06011 ( .a(n6811), .b(n6787), .c(n6767), .o(n9800) );
ao12f01 g06012 ( .a(n6805), .b(n9800), .c(n9799), .o(n9801) );
no02f01 g06013 ( .a(n6807), .b(n4043), .o(n9802) );
no02f01 g06014 ( .a(n9802), .b(n6798), .o(n9803) );
in01f01 g06015 ( .a(n9803), .o(n9804) );
no02f01 g06016 ( .a(n9804), .b(n9801), .o(n9805) );
na02f01 g06017 ( .a(n9804), .b(n9801), .o(n9806) );
in01f01 g06018 ( .a(n9806), .o(n9807) );
no03f01 g06019 ( .a(n9807), .b(n9805), .c(n6934), .o(n9808) );
in01f01 g06020 ( .a(n9800), .o(n9809) );
no02f01 g06021 ( .a(n9798), .b(n6805), .o(n9810) );
in01f01 g06022 ( .a(n9810), .o(n9811) );
na02f01 g06023 ( .a(n9811), .b(n9809), .o(n9812) );
na02f01 g06024 ( .a(n9810), .b(n9800), .o(n9813) );
na02f01 g06025 ( .a(n9813), .b(n9812), .o(n9814) );
no02f01 g06026 ( .a(n9814), .b(n6934), .o(n9815) );
no03f01 g06027 ( .a(n9815), .b(n9808), .c(n9797), .o(n9816) );
oa12f01 g06028 ( .a(n9816), .b(n9775), .c(n9771), .o(n9817) );
no02f01 g06029 ( .a(n9786), .b(n9784), .o(n9818) );
ao12f01 g06030 ( .a(n5001), .b(n9793), .c(n9818), .o(n9819) );
no02f01 g06031 ( .a(n9807), .b(n9805), .o(n9820) );
na02f01 g06032 ( .a(n9814), .b(n6934), .o(n9821) );
ao12f01 g06033 ( .a(n5001), .b(n9821), .c(n9820), .o(n9822) );
no02f01 g06034 ( .a(n9822), .b(n9819), .o(n9823) );
no02f01 g06035 ( .a(n6832), .b(n4043), .o(n9824) );
no02f01 g06036 ( .a(n9824), .b(n6834), .o(n9825) );
no02f01 g06037 ( .a(n9825), .b(n6814), .o(n9826) );
na02f01 g06038 ( .a(n9825), .b(n6814), .o(n9827) );
in01f01 g06039 ( .a(n9827), .o(n9828) );
no02f01 g06040 ( .a(n9828), .b(n9826), .o(n9829) );
in01f01 g06041 ( .a(n9829), .o(n9830) );
no02f01 g06042 ( .a(n9830), .b(n6934), .o(n9831) );
ao12f01 g06043 ( .a(n9831), .b(n9823), .c(n9817), .o(n9832) );
in01f01 g06044 ( .a(n6814), .o(n9833) );
in01f01 g06045 ( .a(n6834), .o(n9834) );
ao12f01 g06046 ( .a(n9824), .b(n9834), .c(n9833), .o(n9835) );
in01f01 g06047 ( .a(n9835), .o(n9836) );
no02f01 g06048 ( .a(n6889), .b(n4043), .o(n9837) );
no02f01 g06049 ( .a(n9837), .b(n6826), .o(n9838) );
in01f01 g06050 ( .a(n9838), .o(n9839) );
no02f01 g06051 ( .a(n9839), .b(n9836), .o(n9840) );
no02f01 g06052 ( .a(n9838), .b(n9835), .o(n9841) );
no02f01 g06053 ( .a(n9841), .b(n9840), .o(n9842) );
in01f01 g06054 ( .a(n9842), .o(n9843) );
no02f01 g06055 ( .a(n9843), .b(n6934), .o(n9844) );
in01f01 g06056 ( .a(n9844), .o(n9845) );
no02f01 g06057 ( .a(n6891), .b(n4043), .o(n9846) );
no02f01 g06058 ( .a(n9846), .b(n6844), .o(n9847) );
in01f01 g06059 ( .a(n9847), .o(n9848) );
no03f01 g06060 ( .a(n9848), .b(n6890), .c(n9650), .o(n9849) );
no02f01 g06061 ( .a(n6890), .b(n9650), .o(n9850) );
no02f01 g06062 ( .a(n9847), .b(n9850), .o(n9851) );
no02f01 g06063 ( .a(n9851), .b(n9849), .o(n9852) );
in01f01 g06064 ( .a(n9852), .o(n9853) );
no02f01 g06065 ( .a(n9853), .b(n6934), .o(n9854) );
in01f01 g06066 ( .a(n9854), .o(n9855) );
in01f01 g06067 ( .a(n9846), .o(n9856) );
ao12f01 g06068 ( .a(n6844), .b(n9850), .c(n9856), .o(n9857) );
no02f01 g06069 ( .a(n6892), .b(n4043), .o(n9858) );
no02f01 g06070 ( .a(n9858), .b(n6853), .o(n9859) );
in01f01 g06071 ( .a(n9859), .o(n9860) );
no02f01 g06072 ( .a(n9860), .b(n9857), .o(n9861) );
na02f01 g06073 ( .a(n9860), .b(n9857), .o(n9862) );
in01f01 g06074 ( .a(n9862), .o(n9863) );
no02f01 g06075 ( .a(n9863), .b(n9861), .o(n9864) );
in01f01 g06076 ( .a(n9864), .o(n9865) );
no02f01 g06077 ( .a(n9865), .b(n6934), .o(n9866) );
in01f01 g06078 ( .a(n9866), .o(n9867) );
na04f01 g06079 ( .a(n9867), .b(n9855), .c(n9845), .d(n9832), .o(n9868) );
ao12f01 g06080 ( .a(n5001), .b(n9842), .c(n9829), .o(n9869) );
in01f01 g06081 ( .a(n9869), .o(n9870) );
no02f01 g06082 ( .a(n9852), .b(n5001), .o(n9871) );
no02f01 g06083 ( .a(n9871), .b(n9865), .o(n9872) );
oa12f01 g06084 ( .a(n9870), .b(n9872), .c(n5001), .o(n9873) );
in01f01 g06085 ( .a(n9873), .o(n9874) );
no02f01 g06086 ( .a(n6898), .b(n4043), .o(n9875) );
in01f01 g06087 ( .a(n9875), .o(n9876) );
ao12f01 g06088 ( .a(n6874), .b(n9876), .c(n9651), .o(n9877) );
no02f01 g06089 ( .a(n6897), .b(n4043), .o(n9878) );
no02f01 g06090 ( .a(n9878), .b(n6869), .o(n9879) );
in01f01 g06091 ( .a(n9879), .o(n9880) );
no02f01 g06092 ( .a(n9880), .b(n9877), .o(n9881) );
na02f01 g06093 ( .a(n9880), .b(n9877), .o(n9882) );
in01f01 g06094 ( .a(n9882), .o(n9883) );
no03f01 g06095 ( .a(n9883), .b(n9881), .c(n6934), .o(n9884) );
no02f01 g06096 ( .a(n9875), .b(n6874), .o(n9885) );
in01f01 g06097 ( .a(n9885), .o(n9886) );
no02f01 g06098 ( .a(n9886), .b(n9652), .o(n9887) );
no02f01 g06099 ( .a(n9885), .b(n9651), .o(n9888) );
no02f01 g06100 ( .a(n9888), .b(n9887), .o(n9889) );
in01f01 g06101 ( .a(n9889), .o(n9890) );
no02f01 g06102 ( .a(n9890), .b(n6934), .o(n9891) );
no02f01 g06103 ( .a(n9891), .b(n9884), .o(n9892) );
in01f01 g06104 ( .a(n9892), .o(n9893) );
ao12f01 g06105 ( .a(n9893), .b(n9874), .c(n9868), .o(n9894) );
no02f01 g06106 ( .a(n9894), .b(n6934), .o(n9895) );
in01f01 g06107 ( .a(n9881), .o(n9896) );
ao12f01 g06108 ( .a(n5001), .b(n9882), .c(n9896), .o(n9897) );
no02f01 g06109 ( .a(n9889), .b(n5001), .o(n9898) );
no02f01 g06110 ( .a(n9898), .b(n9897), .o(n9899) );
in01f01 g06111 ( .a(n9899), .o(n9900) );
no02f01 g06112 ( .a(n9900), .b(n9894), .o(n9901) );
oa22f01 g06113 ( .a(n9901), .b(n5001), .c(n9895), .d(n9659), .o(n243) );
in01f01 g06114 ( .a(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .o(n9903) );
in01f01 g06115 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_15_), .o(n9904) );
no02f01 g06116 ( .a(n9903), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_7_), .o(n9905) );
in01f01 g06117 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_3_), .o(n9906) );
in01f01 g06118 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_0_), .o(n9907) );
in01f01 g06119 ( .a(delay_sub_ln23_unr25_stage8_stallmux_q_1_), .o(n9908) );
na02f01 g06120 ( .a(n9908), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_1_), .o(n9909) );
no02f01 g06121 ( .a(n9908), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_1_), .o(n9910) );
oa12f01 g06122 ( .a(n9909), .b(n9910), .c(n9907), .o(n9911) );
no02f01 g06123 ( .a(n9908), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_2_), .o(n9912) );
in01f01 g06124 ( .a(n9912), .o(n9913) );
na02f01 g06125 ( .a(n9913), .b(n9911), .o(n9914) );
in01f01 g06126 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_2_), .o(n9915) );
no02f01 g06127 ( .a(delay_sub_ln23_unr25_stage8_stallmux_q_1_), .b(n9915), .o(n9916) );
in01f01 g06128 ( .a(n9916), .o(n9917) );
na02f01 g06129 ( .a(n9914), .b(n9917), .o(n9918) );
no02f01 g06130 ( .a(n9918), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_3_), .o(n9919) );
oa22f01 g06131 ( .a(n9919), .b(delay_sub_ln23_unr25_stage8_stallmux_q_1_), .c(n9914), .d(n9906), .o(n9920) );
no02f01 g06132 ( .a(n9903), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_5_), .o(n9921) );
no02f01 g06133 ( .a(n9908), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_4_), .o(n9922) );
no02f01 g06134 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_6_), .b(n9903), .o(n9923) );
no03f01 g06135 ( .a(n9923), .b(n9922), .c(n9921), .o(n9924) );
na02f01 g06136 ( .a(n9924), .b(n9920), .o(n9925) );
in01f01 g06137 ( .a(n9923), .o(n9926) );
na02f01 g06138 ( .a(n9903), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_5_), .o(n9927) );
na02f01 g06139 ( .a(n9908), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_4_), .o(n9928) );
ao12f01 g06140 ( .a(n9921), .b(n9928), .c(n9927), .o(n9929) );
in01f01 g06141 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_7_), .o(n9930) );
in01f01 g06142 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_6_), .o(n9931) );
ao12f01 g06143 ( .a(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(n9931), .c(n9930), .o(n9932) );
oa12f01 g06144 ( .a(n9926), .b(n9932), .c(n9929), .o(n9933) );
ao12f01 g06145 ( .a(n9905), .b(n9933), .c(n9925), .o(n9934) );
ao12f01 g06146 ( .a(n9903), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_8_), .c(delay_sub_ln23_0_unr24_stage8_stallmux_q_9_), .o(n9935) );
in01f01 g06147 ( .a(n9935), .o(n9936) );
no02f01 g06148 ( .a(n9903), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_11_), .o(n9937) );
no02f01 g06149 ( .a(n9903), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_10_), .o(n9938) );
no02f01 g06150 ( .a(n9938), .b(n9937), .o(n9939) );
na02f01 g06151 ( .a(n9939), .b(n9936), .o(n9940) );
no02f01 g06152 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_12_), .b(n9903), .o(n9941) );
no02f01 g06153 ( .a(n9903), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_13_), .o(n9942) );
no03f01 g06154 ( .a(n9942), .b(n9941), .c(n9940), .o(n9943) );
na02f01 g06155 ( .a(n9943), .b(n9934), .o(n9944) );
no02f01 g06156 ( .a(n9903), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_14_), .o(n9945) );
no02f01 g06157 ( .a(n9945), .b(n9944), .o(n9946) );
na02f01 g06158 ( .a(n9903), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_14_), .o(n9947) );
in01f01 g06159 ( .a(n9947), .o(n9948) );
no02f01 g06160 ( .a(n9948), .b(n9946), .o(n9949) );
na02f01 g06161 ( .a(n9949), .b(n9904), .o(n9950) );
in01f01 g06162 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_9_), .o(n9951) );
in01f01 g06163 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_8_), .o(n9952) );
ao12f01 g06164 ( .a(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(n9952), .c(n9951), .o(n9953) );
in01f01 g06165 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_10_), .o(n9954) );
in01f01 g06166 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_11_), .o(n9955) );
ao12f01 g06167 ( .a(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(n9955), .c(n9954), .o(n9956) );
no02f01 g06168 ( .a(n9956), .b(n9953), .o(n9957) );
in01f01 g06169 ( .a(n9957), .o(n9958) );
in01f01 g06170 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_13_), .o(n9959) );
in01f01 g06171 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_12_), .o(n9960) );
ao12f01 g06172 ( .a(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(n9960), .c(n9959), .o(n9961) );
no02f01 g06173 ( .a(n9961), .b(n9958), .o(n9962) );
in01f01 g06174 ( .a(n9962), .o(n9963) );
ao12f01 g06175 ( .a(n9963), .b(n9946), .c(delay_sub_ln23_0_unr24_stage8_stallmux_q_15_), .o(n9964) );
in01f01 g06176 ( .a(n9964), .o(n9965) );
ao12f01 g06177 ( .a(n9965), .b(n9950), .c(n9903), .o(n9966) );
ao12f01 g06178 ( .a(n9903), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_17_), .c(delay_sub_ln23_0_unr24_stage8_stallmux_q_16_), .o(n9967) );
in01f01 g06179 ( .a(n9967), .o(n9968) );
no02f01 g06180 ( .a(n9903), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_19_), .o(n9969) );
no02f01 g06181 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_18_), .b(n9903), .o(n9970) );
no02f01 g06182 ( .a(n9970), .b(n9969), .o(n9971) );
na02f01 g06183 ( .a(n9971), .b(n9968), .o(n9972) );
no02f01 g06184 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_21_), .b(n9903), .o(n9973) );
no02f01 g06185 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_20_), .b(n9903), .o(n9974) );
no02f01 g06186 ( .a(n9974), .b(n9973), .o(n9975) );
in01f01 g06187 ( .a(n9975), .o(n9976) );
no02f01 g06188 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_22_), .b(n9903), .o(n9977) );
no02f01 g06189 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_23_), .b(n9903), .o(n9978) );
no04f01 g06190 ( .a(n9978), .b(n9977), .c(n9976), .d(n9972), .o(n9979) );
in01f01 g06191 ( .a(n9979), .o(n9980) );
no02f01 g06192 ( .a(n9980), .b(n9966), .o(n9981) );
no02f01 g06193 ( .a(n9903), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_25_), .o(n9982) );
no02f01 g06194 ( .a(n9903), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_24_), .o(n9983) );
no02f01 g06195 ( .a(n9983), .b(n9982), .o(n9984) );
in01f01 g06196 ( .a(n9984), .o(n9985) );
no02f01 g06197 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_27_), .b(n9903), .o(n9986) );
no02f01 g06198 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_26_), .b(n9903), .o(n9987) );
no03f01 g06199 ( .a(n9987), .b(n9986), .c(n9985), .o(n9988) );
na02f01 g06200 ( .a(n9988), .b(n9981), .o(n9989) );
no02f01 g06201 ( .a(n9903), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_28_), .o(n9990) );
no02f01 g06202 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_29_), .b(n9903), .o(n9991) );
no02f01 g06203 ( .a(n9991), .b(n9990), .o(n9992) );
in01f01 g06204 ( .a(n9992), .o(n9993) );
no02f01 g06205 ( .a(n9993), .b(n9989), .o(n9994) );
no02f01 g06206 ( .a(n9903), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_30_), .o(n9995) );
in01f01 g06207 ( .a(n9995), .o(n9996) );
in01f01 g06208 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_19_), .o(n9997) );
no02f01 g06209 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_17_), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_16_), .o(n9998) );
na02f01 g06210 ( .a(n9998), .b(n9997), .o(n9999) );
oa12f01 g06211 ( .a(n9903), .b(n9999), .c(delay_sub_ln23_0_unr24_stage8_stallmux_q_18_), .o(n10000) );
in01f01 g06212 ( .a(n10000), .o(n10001) );
in01f01 g06213 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_21_), .o(n10002) );
in01f01 g06214 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_20_), .o(n10003) );
ao12f01 g06215 ( .a(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(n10003), .c(n10002), .o(n10004) );
no02f01 g06216 ( .a(n10004), .b(n10001), .o(n10005) );
in01f01 g06217 ( .a(n10005), .o(n10006) );
in01f01 g06218 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_23_), .o(n10007) );
in01f01 g06219 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_22_), .o(n10008) );
ao12f01 g06220 ( .a(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(n10008), .c(n10007), .o(n10009) );
no02f01 g06221 ( .a(n10009), .b(n10006), .o(n10010) );
in01f01 g06222 ( .a(n10010), .o(n10011) );
in01f01 g06223 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_24_), .o(n10012) );
in01f01 g06224 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_25_), .o(n10013) );
ao12f01 g06225 ( .a(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(n10013), .c(n10012), .o(n10014) );
no02f01 g06226 ( .a(n10014), .b(n10011), .o(n10015) );
in01f01 g06227 ( .a(n10015), .o(n10016) );
in01f01 g06228 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_27_), .o(n10017) );
in01f01 g06229 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_26_), .o(n10018) );
ao12f01 g06230 ( .a(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(n10018), .c(n10017), .o(n10019) );
no02f01 g06231 ( .a(n10019), .b(n10016), .o(n10020) );
in01f01 g06232 ( .a(n10020), .o(n10021) );
in01f01 g06233 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_28_), .o(n10022) );
in01f01 g06234 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_29_), .o(n10023) );
ao12f01 g06235 ( .a(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(n10023), .c(n10022), .o(n10024) );
no02f01 g06236 ( .a(n10024), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_30_), .o(n10025) );
no02f01 g06237 ( .a(n10025), .b(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .o(n10026) );
no02f01 g06238 ( .a(n10026), .b(n10021), .o(n10027) );
in01f01 g06239 ( .a(n10027), .o(n10028) );
ao12f01 g06240 ( .a(n10028), .b(n9996), .c(n9994), .o(n3055) );
in01f01 g06241 ( .a(n3055), .o(n10030) );
no02f01 g06242 ( .a(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(n10012), .o(n10031) );
in01f01 g06243 ( .a(n9981), .o(n10032) );
no02f01 g06244 ( .a(n9983), .b(n10032), .o(n10033) );
no03f01 g06245 ( .a(n10033), .b(n10031), .c(n10011), .o(n10034) );
no02f01 g06246 ( .a(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(n10013), .o(n10035) );
no02f01 g06247 ( .a(n10035), .b(n9982), .o(n10036) );
no02f01 g06248 ( .a(n10036), .b(n10034), .o(n10037) );
na02f01 g06249 ( .a(n10036), .b(n10034), .o(n10038) );
in01f01 g06250 ( .a(n10038), .o(n10039) );
no02f01 g06251 ( .a(n10039), .b(n10037), .o(n10040) );
in01f01 g06252 ( .a(n10040), .o(n10041) );
no02f01 g06253 ( .a(n10041), .b(n10030), .o(n10042) );
in01f01 g06254 ( .a(n10042), .o(n10043) );
no02f01 g06255 ( .a(n10031), .b(n9983), .o(n10044) );
in01f01 g06256 ( .a(n10044), .o(n10045) );
no03f01 g06257 ( .a(n10045), .b(n10011), .c(n9981), .o(n10046) );
ao12f01 g06258 ( .a(n10044), .b(n10010), .c(n10032), .o(n10047) );
no02f01 g06259 ( .a(n10047), .b(n10046), .o(n10048) );
in01f01 g06260 ( .a(n10048), .o(n10049) );
no02f01 g06261 ( .a(n10049), .b(n10030), .o(n10050) );
in01f01 g06262 ( .a(n9909), .o(n10051) );
no02f01 g06263 ( .a(n9910), .b(n10051), .o(n10052) );
no02f01 g06264 ( .a(n10052), .b(n9907), .o(n10053) );
no03f01 g06265 ( .a(n9910), .b(n10051), .c(delay_sub_ln23_0_unr24_stage8_stallmux_q_0_), .o(n10054) );
no02f01 g06266 ( .a(n10054), .b(n10053), .o(n10055) );
in01f01 g06267 ( .a(n10055), .o(n10056) );
no02f01 g06268 ( .a(n10056), .b(n3055), .o(n10057) );
na02f01 g06269 ( .a(n10056), .b(n3055), .o(n10058) );
oa12f01 g06270 ( .a(n10058), .b(n10057), .c(delay_sub_ln23_0_unr24_stage8_stallmux_q_0_), .o(n10059) );
no02f01 g06271 ( .a(n9912), .b(n9916), .o(n10060) );
in01f01 g06272 ( .a(n10060), .o(n10061) );
no02f01 g06273 ( .a(n10061), .b(n9911), .o(n10062) );
in01f01 g06274 ( .a(n9911), .o(n10063) );
no02f01 g06275 ( .a(n10060), .b(n10063), .o(n10064) );
no02f01 g06276 ( .a(n10064), .b(n10062), .o(n10065) );
na02f01 g06277 ( .a(n10065), .b(n10030), .o(n10066) );
na02f01 g06278 ( .a(n10066), .b(n10059), .o(n10067) );
in01f01 g06279 ( .a(n9918), .o(n10068) );
no02f01 g06280 ( .a(delay_sub_ln23_unr25_stage8_stallmux_q_1_), .b(n9906), .o(n10069) );
no02f01 g06281 ( .a(n9908), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_3_), .o(n10070) );
no02f01 g06282 ( .a(n10070), .b(n10069), .o(n10071) );
no02f01 g06283 ( .a(n10071), .b(n10068), .o(n10072) );
na02f01 g06284 ( .a(n10071), .b(n10068), .o(n10073) );
in01f01 g06285 ( .a(n10073), .o(n10074) );
no02f01 g06286 ( .a(n10074), .b(n10072), .o(n10075) );
no02f01 g06287 ( .a(n10065), .b(n10030), .o(n10076) );
in01f01 g06288 ( .a(n10076), .o(n10077) );
na02f01 g06289 ( .a(n10077), .b(n10067), .o(n10078) );
in01f01 g06290 ( .a(n10075), .o(n10079) );
no02f01 g06291 ( .a(n10079), .b(n10078), .o(n10080) );
oa22f01 g06292 ( .a(n10080), .b(n10030), .c(n10075), .d(n10067), .o(n10081) );
in01f01 g06293 ( .a(n9920), .o(n10082) );
in01f01 g06294 ( .a(n9928), .o(n10083) );
no02f01 g06295 ( .a(n10083), .b(n9922), .o(n10084) );
no02f01 g06296 ( .a(n10084), .b(n10082), .o(n10085) );
na02f01 g06297 ( .a(n10084), .b(n10082), .o(n10086) );
in01f01 g06298 ( .a(n10086), .o(n10087) );
no02f01 g06299 ( .a(n10087), .b(n10085), .o(n10088) );
in01f01 g06300 ( .a(n10088), .o(n10089) );
no02f01 g06301 ( .a(n10089), .b(n10030), .o(n10090) );
no02f01 g06302 ( .a(n9922), .b(n10082), .o(n10091) );
no02f01 g06303 ( .a(n10091), .b(n10083), .o(n10092) );
in01f01 g06304 ( .a(n10092), .o(n10093) );
in01f01 g06305 ( .a(n9921), .o(n10094) );
na02f01 g06306 ( .a(n9927), .b(n10094), .o(n10095) );
no02f01 g06307 ( .a(n10095), .b(n10093), .o(n10096) );
na02f01 g06308 ( .a(n10095), .b(n10093), .o(n10097) );
in01f01 g06309 ( .a(n10097), .o(n10098) );
no02f01 g06310 ( .a(n10098), .b(n10096), .o(n10099) );
in01f01 g06311 ( .a(n10099), .o(n10100) );
no02f01 g06312 ( .a(n10100), .b(n10030), .o(n10101) );
in01f01 g06313 ( .a(n9929), .o(n10102) );
na02f01 g06314 ( .a(n10091), .b(n10094), .o(n10103) );
na02f01 g06315 ( .a(n10103), .b(n10102), .o(n10104) );
no02f01 g06316 ( .a(n9931), .b(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .o(n10105) );
no02f01 g06317 ( .a(n10105), .b(n9923), .o(n10106) );
in01f01 g06318 ( .a(n10106), .o(n10107) );
no02f01 g06319 ( .a(n10107), .b(n10104), .o(n10108) );
na02f01 g06320 ( .a(n10107), .b(n10104), .o(n10109) );
in01f01 g06321 ( .a(n10109), .o(n10110) );
no02f01 g06322 ( .a(n10110), .b(n10108), .o(n10111) );
in01f01 g06323 ( .a(n10111), .o(n10112) );
no02f01 g06324 ( .a(n10112), .b(n10030), .o(n10113) );
no03f01 g06325 ( .a(n10113), .b(n10101), .c(n10090), .o(n10114) );
na02f01 g06326 ( .a(n10114), .b(n10081), .o(n10115) );
no02f01 g06327 ( .a(n10111), .b(n3055), .o(n10116) );
ao12f01 g06328 ( .a(n10105), .b(n9929), .c(n9926), .o(n10117) );
na02f01 g06329 ( .a(n10117), .b(n9925), .o(n10118) );
in01f01 g06330 ( .a(n10118), .o(n10119) );
no02f01 g06331 ( .a(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(n9930), .o(n10120) );
no02f01 g06332 ( .a(n10120), .b(n9905), .o(n10121) );
no02f01 g06333 ( .a(n10121), .b(n10119), .o(n10122) );
na02f01 g06334 ( .a(n10121), .b(n10119), .o(n10123) );
in01f01 g06335 ( .a(n10123), .o(n10124) );
no02f01 g06336 ( .a(n10124), .b(n10122), .o(n10125) );
in01f01 g06337 ( .a(n10125), .o(n10126) );
no02f01 g06338 ( .a(n10126), .b(n10116), .o(n10127) );
na02f01 g06339 ( .a(n10127), .b(n10115), .o(n10128) );
ao12f01 g06340 ( .a(n3055), .b(n10099), .c(n10088), .o(n10129) );
in01f01 g06341 ( .a(n10129), .o(n10130) );
oa12f01 g06342 ( .a(n10130), .b(n10125), .c(n10115), .o(n10131) );
ao12f01 g06343 ( .a(n10131), .b(n10128), .c(n10030), .o(n10132) );
in01f01 g06344 ( .a(n9934), .o(n10133) );
no02f01 g06345 ( .a(n9935), .b(n10133), .o(n10134) );
no02f01 g06346 ( .a(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(n9954), .o(n10135) );
no02f01 g06347 ( .a(n10135), .b(n9938), .o(n10136) );
in01f01 g06348 ( .a(n10136), .o(n10137) );
no03f01 g06349 ( .a(n10137), .b(n10134), .c(n9953), .o(n10138) );
no02f01 g06350 ( .a(n10134), .b(n9953), .o(n10139) );
no02f01 g06351 ( .a(n10136), .b(n10139), .o(n10140) );
no02f01 g06352 ( .a(n10140), .b(n10138), .o(n10141) );
in01f01 g06353 ( .a(n10141), .o(n10142) );
no02f01 g06354 ( .a(n10142), .b(n10030), .o(n10143) );
in01f01 g06355 ( .a(n10143), .o(n10144) );
no03f01 g06356 ( .a(n9938), .b(n9935), .c(n10133), .o(n10145) );
no03f01 g06357 ( .a(n10145), .b(n10135), .c(n9953), .o(n10146) );
no02f01 g06358 ( .a(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(n9955), .o(n10147) );
no02f01 g06359 ( .a(n10147), .b(n9937), .o(n10148) );
no02f01 g06360 ( .a(n10148), .b(n10146), .o(n10149) );
na02f01 g06361 ( .a(n10148), .b(n10146), .o(n10150) );
in01f01 g06362 ( .a(n10150), .o(n10151) );
no02f01 g06363 ( .a(n10151), .b(n10149), .o(n10152) );
in01f01 g06364 ( .a(n10152), .o(n10153) );
no02f01 g06365 ( .a(n10153), .b(n10030), .o(n10154) );
no02f01 g06366 ( .a(n9952), .b(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .o(n10155) );
no02f01 g06367 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_8_), .b(n9903), .o(n10156) );
in01f01 g06368 ( .a(n10156), .o(n10157) );
ao12f01 g06369 ( .a(n10155), .b(n10157), .c(n9934), .o(n10158) );
in01f01 g06370 ( .a(n10158), .o(n10159) );
no02f01 g06371 ( .a(n9903), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_9_), .o(n10160) );
no02f01 g06372 ( .a(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(n9951), .o(n10161) );
no02f01 g06373 ( .a(n10161), .b(n10160), .o(n10162) );
in01f01 g06374 ( .a(n10162), .o(n10163) );
no02f01 g06375 ( .a(n10163), .b(n10159), .o(n10164) );
no02f01 g06376 ( .a(n10162), .b(n10158), .o(n10165) );
no02f01 g06377 ( .a(n10165), .b(n10164), .o(n10166) );
no02f01 g06378 ( .a(n10156), .b(n10155), .o(n10167) );
no02f01 g06379 ( .a(n10167), .b(n10133), .o(n10168) );
na02f01 g06380 ( .a(n10167), .b(n10133), .o(n10169) );
in01f01 g06381 ( .a(n10169), .o(n10170) );
no02f01 g06382 ( .a(n10170), .b(n10168), .o(n10171) );
no02f01 g06383 ( .a(n10171), .b(n10166), .o(n10172) );
no02f01 g06384 ( .a(n10172), .b(n10030), .o(n10173) );
no02f01 g06385 ( .a(n10173), .b(n10154), .o(n10174) );
na02f01 g06386 ( .a(n10174), .b(n10144), .o(n10175) );
no02f01 g06387 ( .a(n9960), .b(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .o(n10176) );
no03f01 g06388 ( .a(n9941), .b(n9940), .c(n10133), .o(n10177) );
no03f01 g06389 ( .a(n10177), .b(n10176), .c(n9958), .o(n10178) );
no02f01 g06390 ( .a(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(n9959), .o(n10179) );
no02f01 g06391 ( .a(n10179), .b(n9942), .o(n10180) );
no02f01 g06392 ( .a(n10180), .b(n10178), .o(n10181) );
na02f01 g06393 ( .a(n10180), .b(n10178), .o(n10182) );
in01f01 g06394 ( .a(n10182), .o(n10183) );
no02f01 g06395 ( .a(n10183), .b(n10181), .o(n10184) );
in01f01 g06396 ( .a(n10184), .o(n10185) );
no02f01 g06397 ( .a(n10185), .b(n10030), .o(n10186) );
no02f01 g06398 ( .a(n9940), .b(n10133), .o(n10187) );
no02f01 g06399 ( .a(n10176), .b(n9941), .o(n10188) );
in01f01 g06400 ( .a(n10188), .o(n10189) );
no03f01 g06401 ( .a(n10189), .b(n10187), .c(n9958), .o(n10190) );
no02f01 g06402 ( .a(n10187), .b(n9958), .o(n10191) );
no02f01 g06403 ( .a(n10188), .b(n10191), .o(n10192) );
no02f01 g06404 ( .a(n10192), .b(n10190), .o(n10193) );
in01f01 g06405 ( .a(n10193), .o(n10194) );
no02f01 g06406 ( .a(n10194), .b(n10030), .o(n10195) );
no03f01 g06407 ( .a(n10195), .b(n10186), .c(n10175), .o(n10196) );
in01f01 g06408 ( .a(n10196), .o(n10197) );
in01f01 g06409 ( .a(n9944), .o(n10198) );
no02f01 g06410 ( .a(n9948), .b(n9945), .o(n10199) );
in01f01 g06411 ( .a(n10199), .o(n10200) );
no03f01 g06412 ( .a(n10200), .b(n9963), .c(n10198), .o(n10201) );
ao12f01 g06413 ( .a(n10199), .b(n9962), .c(n9944), .o(n10202) );
no02f01 g06414 ( .a(n10202), .b(n10201), .o(n10203) );
in01f01 g06415 ( .a(n10203), .o(n10204) );
no02f01 g06416 ( .a(n10204), .b(n10030), .o(n10205) );
no03f01 g06417 ( .a(n10205), .b(n10197), .c(n10132), .o(n10206) );
in01f01 g06418 ( .a(n10206), .o(n10207) );
na02f01 g06419 ( .a(n9962), .b(n9949), .o(n10208) );
no02f01 g06420 ( .a(n9903), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_15_), .o(n10209) );
no02f01 g06421 ( .a(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(n9904), .o(n10210) );
no02f01 g06422 ( .a(n10210), .b(n10209), .o(n10211) );
in01f01 g06423 ( .a(n10211), .o(n10212) );
no02f01 g06424 ( .a(n10212), .b(n10208), .o(n10213) );
na02f01 g06425 ( .a(n10212), .b(n10208), .o(n10214) );
in01f01 g06426 ( .a(n10214), .o(n10215) );
no02f01 g06427 ( .a(n10215), .b(n10213), .o(n10216) );
in01f01 g06428 ( .a(n10216), .o(n10217) );
no02f01 g06429 ( .a(n10217), .b(n10030), .o(n10218) );
ao12f01 g06430 ( .a(n3055), .b(n10171), .c(n10166), .o(n10219) );
ao12f01 g06431 ( .a(n3055), .b(n10152), .c(n10141), .o(n10220) );
no02f01 g06432 ( .a(n10220), .b(n10219), .o(n10221) );
in01f01 g06433 ( .a(n10221), .o(n10222) );
ao12f01 g06434 ( .a(n3055), .b(n10193), .c(n10184), .o(n10223) );
no02f01 g06435 ( .a(n10223), .b(n10222), .o(n10224) );
in01f01 g06436 ( .a(n10224), .o(n10225) );
ao12f01 g06437 ( .a(n3055), .b(n10216), .c(n10203), .o(n10226) );
no02f01 g06438 ( .a(n10226), .b(n10225), .o(n10227) );
oa12f01 g06439 ( .a(n10227), .b(n10218), .c(n10207), .o(n10228) );
in01f01 g06440 ( .a(n9966), .o(n10229) );
in01f01 g06441 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_16_), .o(n10230) );
no02f01 g06442 ( .a(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(n10230), .o(n10231) );
no02f01 g06443 ( .a(n9903), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_16_), .o(n10232) );
in01f01 g06444 ( .a(n10232), .o(n10233) );
ao12f01 g06445 ( .a(n10231), .b(n10233), .c(n10229), .o(n10234) );
in01f01 g06446 ( .a(n10234), .o(n10235) );
no02f01 g06447 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_17_), .b(n9903), .o(n10236) );
na02f01 g06448 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_17_), .b(n9903), .o(n10237) );
in01f01 g06449 ( .a(n10237), .o(n10238) );
no02f01 g06450 ( .a(n10238), .b(n10236), .o(n10239) );
in01f01 g06451 ( .a(n10239), .o(n10240) );
no02f01 g06452 ( .a(n10240), .b(n10235), .o(n10241) );
no02f01 g06453 ( .a(n10239), .b(n10234), .o(n10242) );
no02f01 g06454 ( .a(n10242), .b(n10241), .o(n10243) );
in01f01 g06455 ( .a(n10243), .o(n10244) );
no02f01 g06456 ( .a(n10232), .b(n10231), .o(n10245) );
in01f01 g06457 ( .a(n10245), .o(n10246) );
no02f01 g06458 ( .a(n10246), .b(n10229), .o(n10247) );
no02f01 g06459 ( .a(n10245), .b(n9966), .o(n10248) );
no02f01 g06460 ( .a(n10248), .b(n10247), .o(n10249) );
in01f01 g06461 ( .a(n10249), .o(n10250) );
ao12f01 g06462 ( .a(n10030), .b(n10250), .c(n10244), .o(n10251) );
in01f01 g06463 ( .a(n10251), .o(n10252) );
na02f01 g06464 ( .a(n10252), .b(n10228), .o(n10253) );
no02f01 g06465 ( .a(n9967), .b(n9966), .o(n10254) );
no02f01 g06466 ( .a(n9998), .b(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .o(n10255) );
in01f01 g06467 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_18_), .o(n10256) );
no02f01 g06468 ( .a(n10256), .b(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .o(n10257) );
no02f01 g06469 ( .a(n10257), .b(n9970), .o(n10258) );
in01f01 g06470 ( .a(n10258), .o(n10259) );
no03f01 g06471 ( .a(n10259), .b(n10255), .c(n10254), .o(n10260) );
no02f01 g06472 ( .a(n10255), .b(n10254), .o(n10261) );
no02f01 g06473 ( .a(n10258), .b(n10261), .o(n10262) );
no02f01 g06474 ( .a(n10262), .b(n10260), .o(n10263) );
in01f01 g06475 ( .a(n10263), .o(n10264) );
no02f01 g06476 ( .a(n10264), .b(n10030), .o(n10265) );
no03f01 g06477 ( .a(n9970), .b(n9967), .c(n9966), .o(n10266) );
no03f01 g06478 ( .a(n10266), .b(n10255), .c(n10257), .o(n10267) );
in01f01 g06479 ( .a(n10267), .o(n10268) );
no02f01 g06480 ( .a(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(n9997), .o(n10269) );
no02f01 g06481 ( .a(n10269), .b(n9969), .o(n10270) );
in01f01 g06482 ( .a(n10270), .o(n10271) );
no02f01 g06483 ( .a(n10271), .b(n10268), .o(n10272) );
no02f01 g06484 ( .a(n10270), .b(n10267), .o(n10273) );
no03f01 g06485 ( .a(n10273), .b(n10272), .c(n10030), .o(n10274) );
no02f01 g06486 ( .a(n10274), .b(n10265), .o(n10275) );
in01f01 g06487 ( .a(n10275), .o(n10276) );
no02f01 g06488 ( .a(n10276), .b(n10253), .o(n10277) );
no02f01 g06489 ( .a(n9972), .b(n9966), .o(n10278) );
no02f01 g06490 ( .a(n10003), .b(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .o(n10279) );
no02f01 g06491 ( .a(n10279), .b(n9974), .o(n10280) );
in01f01 g06492 ( .a(n10280), .o(n10281) );
no03f01 g06493 ( .a(n10281), .b(n10278), .c(n10001), .o(n10282) );
in01f01 g06494 ( .a(n10278), .o(n10283) );
ao12f01 g06495 ( .a(n10280), .b(n10283), .c(n10000), .o(n10284) );
no02f01 g06496 ( .a(n10284), .b(n10282), .o(n10285) );
in01f01 g06497 ( .a(n10285), .o(n10286) );
no02f01 g06498 ( .a(n10286), .b(n10030), .o(n10287) );
in01f01 g06499 ( .a(n10287), .o(n10288) );
no02f01 g06500 ( .a(n10283), .b(n9974), .o(n10289) );
no03f01 g06501 ( .a(n10289), .b(n10279), .c(n10001), .o(n10290) );
in01f01 g06502 ( .a(n10290), .o(n10291) );
no02f01 g06503 ( .a(n10002), .b(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .o(n10292) );
no02f01 g06504 ( .a(n10292), .b(n9973), .o(n10293) );
in01f01 g06505 ( .a(n10293), .o(n10294) );
no02f01 g06506 ( .a(n10294), .b(n10291), .o(n10295) );
no02f01 g06507 ( .a(n10293), .b(n10290), .o(n10296) );
no02f01 g06508 ( .a(n10296), .b(n10295), .o(n10297) );
in01f01 g06509 ( .a(n10297), .o(n10298) );
no02f01 g06510 ( .a(n10298), .b(n10030), .o(n10299) );
in01f01 g06511 ( .a(n10299), .o(n10300) );
na03f01 g06512 ( .a(n10300), .b(n10288), .c(n10277), .o(n10301) );
no02f01 g06513 ( .a(n10283), .b(n9976), .o(n10302) );
no02f01 g06514 ( .a(n10008), .b(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .o(n10303) );
no02f01 g06515 ( .a(n10303), .b(n9977), .o(n10304) );
in01f01 g06516 ( .a(n10304), .o(n10305) );
no03f01 g06517 ( .a(n10305), .b(n10302), .c(n10006), .o(n10306) );
no02f01 g06518 ( .a(n10302), .b(n10006), .o(n10307) );
no02f01 g06519 ( .a(n10304), .b(n10307), .o(n10308) );
no03f01 g06520 ( .a(n10308), .b(n10306), .c(n10030), .o(n10309) );
no03f01 g06521 ( .a(n10283), .b(n9977), .c(n9976), .o(n10310) );
no03f01 g06522 ( .a(n10310), .b(n10303), .c(n10006), .o(n10311) );
no02f01 g06523 ( .a(n10007), .b(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .o(n10312) );
no02f01 g06524 ( .a(n10312), .b(n9978), .o(n10313) );
no02f01 g06525 ( .a(n10313), .b(n10311), .o(n10314) );
na02f01 g06526 ( .a(n10313), .b(n10311), .o(n10315) );
in01f01 g06527 ( .a(n10315), .o(n10316) );
no02f01 g06528 ( .a(n10316), .b(n10314), .o(n10317) );
in01f01 g06529 ( .a(n10317), .o(n10318) );
no02f01 g06530 ( .a(n10318), .b(n10030), .o(n10319) );
no04f01 g06531 ( .a(n10319), .b(n10309), .c(n10301), .d(n10050), .o(n10320) );
no02f01 g06532 ( .a(n9985), .b(n10032), .o(n10321) );
no02f01 g06533 ( .a(n10018), .b(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .o(n10322) );
no02f01 g06534 ( .a(n10322), .b(n9987), .o(n10323) );
in01f01 g06535 ( .a(n10323), .o(n10324) );
no03f01 g06536 ( .a(n10324), .b(n10321), .c(n10016), .o(n10325) );
no02f01 g06537 ( .a(n10321), .b(n10016), .o(n10326) );
no02f01 g06538 ( .a(n10323), .b(n10326), .o(n10327) );
no02f01 g06539 ( .a(n10327), .b(n10325), .o(n10328) );
in01f01 g06540 ( .a(n10328), .o(n10329) );
no02f01 g06541 ( .a(n10329), .b(n10030), .o(n10330) );
in01f01 g06542 ( .a(n10330), .o(n10331) );
no03f01 g06543 ( .a(n9987), .b(n9985), .c(n10032), .o(n10332) );
no03f01 g06544 ( .a(n10332), .b(n10322), .c(n10016), .o(n10333) );
in01f01 g06545 ( .a(n10333), .o(n10334) );
no02f01 g06546 ( .a(n10017), .b(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .o(n10335) );
no02f01 g06547 ( .a(n10335), .b(n9986), .o(n10336) );
in01f01 g06548 ( .a(n10336), .o(n10337) );
no02f01 g06549 ( .a(n10337), .b(n10334), .o(n10338) );
no02f01 g06550 ( .a(n10336), .b(n10333), .o(n10339) );
no02f01 g06551 ( .a(n10339), .b(n10338), .o(n10340) );
in01f01 g06552 ( .a(n10340), .o(n10341) );
no02f01 g06553 ( .a(n10341), .b(n10030), .o(n10342) );
in01f01 g06554 ( .a(n10342), .o(n10343) );
na04f01 g06555 ( .a(n10343), .b(n10331), .c(n10320), .d(n10043), .o(n10344) );
ao12f01 g06556 ( .a(n10021), .b(n9988), .c(n9981), .o(n10345) );
no02f01 g06557 ( .a(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(n10022), .o(n10346) );
no02f01 g06558 ( .a(n10346), .b(n9990), .o(n10347) );
no02f01 g06559 ( .a(n10347), .b(n10345), .o(n10348) );
na02f01 g06560 ( .a(n10347), .b(n10345), .o(n10349) );
in01f01 g06561 ( .a(n10349), .o(n10350) );
no03f01 g06562 ( .a(n10350), .b(n10348), .c(n10030), .o(n10351) );
no02f01 g06563 ( .a(n9990), .b(n9989), .o(n10352) );
no03f01 g06564 ( .a(n10352), .b(n10346), .c(n10021), .o(n10353) );
no02f01 g06565 ( .a(n10023), .b(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .o(n10354) );
no02f01 g06566 ( .a(n10354), .b(n9991), .o(n10355) );
no02f01 g06567 ( .a(n10355), .b(n10353), .o(n10356) );
na02f01 g06568 ( .a(n10355), .b(n10353), .o(n10357) );
in01f01 g06569 ( .a(n10357), .o(n10358) );
no03f01 g06570 ( .a(n10358), .b(n10356), .c(n10030), .o(n10359) );
no02f01 g06571 ( .a(n10359), .b(n10351), .o(n10360) );
in01f01 g06572 ( .a(n10360), .o(n10361) );
no03f01 g06573 ( .a(n10024), .b(n10021), .c(n9994), .o(n10362) );
in01f01 g06574 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_30_), .o(n10363) );
no02f01 g06575 ( .a(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(n10363), .o(n10364) );
no02f01 g06576 ( .a(n10364), .b(n9995), .o(n10365) );
no02f01 g06577 ( .a(n10365), .b(n10362), .o(n10366) );
na02f01 g06578 ( .a(n10365), .b(n10362), .o(n10367) );
in01f01 g06579 ( .a(n10367), .o(n10368) );
no03f01 g06580 ( .a(n10368), .b(n10366), .c(n10030), .o(n10369) );
no02f01 g06581 ( .a(n10369), .b(n10361), .o(n10370) );
in01f01 g06582 ( .a(n10370), .o(n10371) );
ao12f01 g06583 ( .a(n3055), .b(n10249), .c(n10243), .o(n10372) );
no02f01 g06584 ( .a(n10273), .b(n10272), .o(n10373) );
ao12f01 g06585 ( .a(n3055), .b(n10373), .c(n10263), .o(n10374) );
no02f01 g06586 ( .a(n10374), .b(n10372), .o(n10375) );
in01f01 g06587 ( .a(n10375), .o(n10376) );
ao12f01 g06588 ( .a(n3055), .b(n10297), .c(n10285), .o(n10377) );
no02f01 g06589 ( .a(n10377), .b(n10376), .o(n10378) );
in01f01 g06590 ( .a(n10378), .o(n10379) );
no02f01 g06591 ( .a(n10308), .b(n10306), .o(n10380) );
ao12f01 g06592 ( .a(n3055), .b(n10317), .c(n10380), .o(n10381) );
no02f01 g06593 ( .a(n10381), .b(n10379), .o(n10382) );
in01f01 g06594 ( .a(n10382), .o(n10383) );
ao12f01 g06595 ( .a(n3055), .b(n10048), .c(n10040), .o(n10384) );
no02f01 g06596 ( .a(n10384), .b(n10383), .o(n10385) );
in01f01 g06597 ( .a(n10385), .o(n10386) );
ao12f01 g06598 ( .a(n3055), .b(n10340), .c(n10328), .o(n10387) );
no02f01 g06599 ( .a(n10387), .b(n10386), .o(n10388) );
in01f01 g06600 ( .a(n10388), .o(n10389) );
no02f01 g06601 ( .a(n10368), .b(n10366), .o(n10390) );
no02f01 g06602 ( .a(n10350), .b(n10348), .o(n10391) );
no02f01 g06603 ( .a(n10358), .b(n10356), .o(n10392) );
ao12f01 g06604 ( .a(n3055), .b(n10392), .c(n10391), .o(n10393) );
in01f01 g06605 ( .a(n10393), .o(n10394) );
ao12f01 g06606 ( .a(n3055), .b(n10394), .c(n10390), .o(n10395) );
no02f01 g06607 ( .a(n10395), .b(n10389), .o(n10396) );
oa12f01 g06608 ( .a(n10396), .b(n10371), .c(n10344), .o(n10397) );
no02f01 g06609 ( .a(n10263), .b(n3055), .o(n10398) );
no02f01 g06610 ( .a(n10398), .b(n10372), .o(n10399) );
oa12f01 g06611 ( .a(n10399), .b(n10265), .c(n10253), .o(n10400) );
in01f01 g06612 ( .a(n10400), .o(n10401) );
no02f01 g06613 ( .a(n10373), .b(n3055), .o(n10402) );
no02f01 g06614 ( .a(n10402), .b(n10274), .o(n10403) );
no02f01 g06615 ( .a(n10403), .b(n10401), .o(n10404) );
na02f01 g06616 ( .a(n10403), .b(n10401), .o(n10405) );
in01f01 g06617 ( .a(n10405), .o(n10406) );
no02f01 g06618 ( .a(n10406), .b(n10404), .o(n10407) );
no02f01 g06619 ( .a(n10376), .b(n10277), .o(n10408) );
no02f01 g06620 ( .a(n10285), .b(n3055), .o(n10409) );
no02f01 g06621 ( .a(n10409), .b(n10287), .o(n10410) );
no02f01 g06622 ( .a(n10410), .b(n10408), .o(n10411) );
na02f01 g06623 ( .a(n10410), .b(n10408), .o(n10412) );
in01f01 g06624 ( .a(n10412), .o(n10413) );
no02f01 g06625 ( .a(n10413), .b(n10411), .o(n10414) );
no02f01 g06626 ( .a(n10414), .b(n10407), .o(n10415) );
no02f01 g06627 ( .a(n10415), .b(n10397), .o(n10416) );
no02f01 g06628 ( .a(n10173), .b(n10132), .o(n10417) );
no02f01 g06629 ( .a(n10417), .b(n10219), .o(n10418) );
no02f01 g06630 ( .a(n10141), .b(n3055), .o(n10419) );
no02f01 g06631 ( .a(n10419), .b(n10143), .o(n10420) );
no02f01 g06632 ( .a(n10420), .b(n10418), .o(n10421) );
na02f01 g06633 ( .a(n10420), .b(n10418), .o(n10422) );
in01f01 g06634 ( .a(n10422), .o(n10423) );
no02f01 g06635 ( .a(n10423), .b(n10421), .o(n10424) );
in01f01 g06636 ( .a(n10424), .o(n10425) );
no02f01 g06637 ( .a(n10425), .b(n10397), .o(n10426) );
in01f01 g06638 ( .a(n10426), .o(n10427) );
in01f01 g06639 ( .a(n10397), .o(n4088) );
in01f01 g06640 ( .a(n10132), .o(n10429) );
no02f01 g06641 ( .a(n10171), .b(n3055), .o(n10430) );
na02f01 g06642 ( .a(n10171), .b(n3055), .o(n10431) );
in01f01 g06643 ( .a(n10431), .o(n10432) );
no02f01 g06644 ( .a(n10432), .b(n10430), .o(n10433) );
in01f01 g06645 ( .a(n10433), .o(n10434) );
no02f01 g06646 ( .a(n10434), .b(n10429), .o(n10435) );
no02f01 g06647 ( .a(n10433), .b(n10132), .o(n10436) );
no02f01 g06648 ( .a(n10436), .b(n10435), .o(n10437) );
no02f01 g06649 ( .a(n10129), .b(n10116), .o(n10438) );
na02f01 g06650 ( .a(n10438), .b(n10115), .o(n10439) );
no02f01 g06651 ( .a(n10126), .b(n10030), .o(n10440) );
no02f01 g06652 ( .a(n10125), .b(n3055), .o(n10441) );
no02f01 g06653 ( .a(n10441), .b(n10440), .o(n10442) );
in01f01 g06654 ( .a(n10442), .o(n10443) );
no02f01 g06655 ( .a(n10443), .b(n10439), .o(n10444) );
na02f01 g06656 ( .a(n10443), .b(n10439), .o(n10445) );
in01f01 g06657 ( .a(n10445), .o(n10446) );
no02f01 g06658 ( .a(n10446), .b(n10444), .o(n10447) );
ao12f01 g06659 ( .a(n4088), .b(n10447), .c(n10437), .o(n10448) );
in01f01 g06660 ( .a(n10448), .o(n10449) );
in01f01 g06661 ( .a(n10081), .o(n10450) );
no02f01 g06662 ( .a(n10088), .b(n3055), .o(n10451) );
no02f01 g06663 ( .a(n10451), .b(n10090), .o(n10452) );
no02f01 g06664 ( .a(n10452), .b(n10450), .o(n10453) );
na02f01 g06665 ( .a(n10452), .b(n10450), .o(n10454) );
in01f01 g06666 ( .a(n10454), .o(n10455) );
no02f01 g06667 ( .a(n10455), .b(n10453), .o(n10456) );
in01f01 g06668 ( .a(n10456), .o(n10457) );
na02f01 g06669 ( .a(n10457), .b(n10397), .o(n10458) );
in01f01 g06670 ( .a(n10078), .o(n10459) );
no02f01 g06671 ( .a(n10079), .b(n3055), .o(n10460) );
no02f01 g06672 ( .a(n10075), .b(n10030), .o(n10461) );
no02f01 g06673 ( .a(n10461), .b(n10460), .o(n10462) );
no02f01 g06674 ( .a(n10462), .b(n10459), .o(n10463) );
na02f01 g06675 ( .a(n10462), .b(n10459), .o(n10464) );
in01f01 g06676 ( .a(n10464), .o(n10465) );
no02f01 g06677 ( .a(n10465), .b(n10463), .o(n10466) );
in01f01 g06678 ( .a(n10466), .o(n10467) );
oa12f01 g06679 ( .a(n10467), .b(n10457), .c(n10397), .o(n10468) );
no02f01 g06680 ( .a(n10090), .b(n10450), .o(n10469) );
no02f01 g06681 ( .a(n10099), .b(n3055), .o(n10470) );
no02f01 g06682 ( .a(n10470), .b(n10101), .o(n10471) );
in01f01 g06683 ( .a(n10471), .o(n10472) );
no03f01 g06684 ( .a(n10472), .b(n10469), .c(n10451), .o(n10473) );
no02f01 g06685 ( .a(n10469), .b(n10451), .o(n10474) );
no02f01 g06686 ( .a(n10471), .b(n10474), .o(n10475) );
no02f01 g06687 ( .a(n10475), .b(n10473), .o(n10476) );
in01f01 g06688 ( .a(n10476), .o(n10477) );
no02f01 g06689 ( .a(n10477), .b(n10397), .o(n10478) );
ao12f01 g06690 ( .a(n10478), .b(n10468), .c(n10458), .o(n10479) );
in01f01 g06691 ( .a(n10101), .o(n10480) );
ao12f01 g06692 ( .a(n10129), .b(n10469), .c(n10480), .o(n10481) );
no02f01 g06693 ( .a(n10116), .b(n10113), .o(n10482) );
no02f01 g06694 ( .a(n10482), .b(n10481), .o(n10483) );
na02f01 g06695 ( .a(n10482), .b(n10481), .o(n10484) );
in01f01 g06696 ( .a(n10484), .o(n10485) );
no02f01 g06697 ( .a(n10485), .b(n10483), .o(n10486) );
in01f01 g06698 ( .a(n10486), .o(n10487) );
na02f01 g06699 ( .a(n10487), .b(n10479), .o(n10488) );
na02f01 g06700 ( .a(n10477), .b(n10397), .o(n10489) );
in01f01 g06701 ( .a(n10489), .o(n10490) );
no03f01 g06702 ( .a(n10490), .b(n10487), .c(n10479), .o(n10491) );
oa12f01 g06703 ( .a(n10488), .b(n10491), .c(n4088), .o(n10492) );
in01f01 g06704 ( .a(n10447), .o(n10493) );
no02f01 g06705 ( .a(n10493), .b(n10397), .o(n10494) );
in01f01 g06706 ( .a(n10494), .o(n10495) );
in01f01 g06707 ( .a(n10437), .o(n10496) );
no02f01 g06708 ( .a(n10496), .b(n10397), .o(n10497) );
in01f01 g06709 ( .a(n10497), .o(n10498) );
ao12f01 g06710 ( .a(n10430), .b(n10431), .c(n10429), .o(n10499) );
in01f01 g06711 ( .a(n10499), .o(n10500) );
in01f01 g06712 ( .a(n10166), .o(n10501) );
no02f01 g06713 ( .a(n10501), .b(n10030), .o(n10502) );
no02f01 g06714 ( .a(n10166), .b(n3055), .o(n10503) );
no02f01 g06715 ( .a(n10503), .b(n10502), .o(n10504) );
in01f01 g06716 ( .a(n10504), .o(n10505) );
no02f01 g06717 ( .a(n10505), .b(n10500), .o(n10506) );
no02f01 g06718 ( .a(n10504), .b(n10499), .o(n10507) );
no02f01 g06719 ( .a(n10507), .b(n10506), .o(n10508) );
in01f01 g06720 ( .a(n10508), .o(n10509) );
no02f01 g06721 ( .a(n10509), .b(n10397), .o(n10510) );
in01f01 g06722 ( .a(n10510), .o(n10511) );
na04f01 g06723 ( .a(n10511), .b(n10498), .c(n10495), .d(n10492), .o(n10512) );
ao12f01 g06724 ( .a(n4088), .b(n10508), .c(n10424), .o(n10513) );
in01f01 g06725 ( .a(n10513), .o(n10514) );
na03f01 g06726 ( .a(n10514), .b(n10512), .c(n10449), .o(n10515) );
na02f01 g06727 ( .a(n10417), .b(n10144), .o(n10516) );
no02f01 g06728 ( .a(n10419), .b(n10219), .o(n10517) );
na02f01 g06729 ( .a(n10517), .b(n10516), .o(n10518) );
no02f01 g06730 ( .a(n10152), .b(n3055), .o(n10519) );
no02f01 g06731 ( .a(n10519), .b(n10154), .o(n10520) );
in01f01 g06732 ( .a(n10520), .o(n10521) );
no02f01 g06733 ( .a(n10521), .b(n10518), .o(n10522) );
na02f01 g06734 ( .a(n10521), .b(n10518), .o(n10523) );
in01f01 g06735 ( .a(n10523), .o(n10524) );
no02f01 g06736 ( .a(n10524), .b(n10522), .o(n10525) );
in01f01 g06737 ( .a(n10525), .o(n10526) );
no02f01 g06738 ( .a(n10175), .b(n10132), .o(n10527) );
no02f01 g06739 ( .a(n10193), .b(n3055), .o(n10528) );
no02f01 g06740 ( .a(n10528), .b(n10195), .o(n10529) );
in01f01 g06741 ( .a(n10529), .o(n10530) );
no03f01 g06742 ( .a(n10530), .b(n10527), .c(n10222), .o(n10531) );
no02f01 g06743 ( .a(n10527), .b(n10222), .o(n10532) );
no02f01 g06744 ( .a(n10529), .b(n10532), .o(n10533) );
no02f01 g06745 ( .a(n10533), .b(n10531), .o(n10534) );
in01f01 g06746 ( .a(n10534), .o(n10535) );
ao12f01 g06747 ( .a(n10397), .b(n10535), .c(n10526), .o(n10536) );
in01f01 g06748 ( .a(n10536), .o(n10537) );
no03f01 g06749 ( .a(n10195), .b(n10175), .c(n10132), .o(n10538) );
no02f01 g06750 ( .a(n10528), .b(n10222), .o(n10539) );
in01f01 g06751 ( .a(n10539), .o(n10540) );
no02f01 g06752 ( .a(n10184), .b(n3055), .o(n10541) );
no02f01 g06753 ( .a(n10541), .b(n10186), .o(n10542) );
in01f01 g06754 ( .a(n10542), .o(n10543) );
no03f01 g06755 ( .a(n10543), .b(n10540), .c(n10538), .o(n10544) );
no02f01 g06756 ( .a(n10540), .b(n10538), .o(n10545) );
no02f01 g06757 ( .a(n10542), .b(n10545), .o(n10546) );
no02f01 g06758 ( .a(n10546), .b(n10544), .o(n10547) );
in01f01 g06759 ( .a(n10547), .o(n10548) );
no02f01 g06760 ( .a(n10548), .b(n10397), .o(n10549) );
ao12f01 g06761 ( .a(n10225), .b(n10196), .c(n10429), .o(n10550) );
no02f01 g06762 ( .a(n10203), .b(n3055), .o(n10551) );
no02f01 g06763 ( .a(n10551), .b(n10205), .o(n10552) );
no02f01 g06764 ( .a(n10552), .b(n10550), .o(n10553) );
na02f01 g06765 ( .a(n10552), .b(n10550), .o(n10554) );
in01f01 g06766 ( .a(n10554), .o(n10555) );
no02f01 g06767 ( .a(n10555), .b(n10553), .o(n10556) );
in01f01 g06768 ( .a(n10556), .o(n10557) );
no02f01 g06769 ( .a(n10557), .b(n10397), .o(n10558) );
no02f01 g06770 ( .a(n10558), .b(n10549), .o(n10559) );
na04f01 g06771 ( .a(n10559), .b(n10537), .c(n10515), .d(n10427), .o(n10560) );
ao12f01 g06772 ( .a(n4088), .b(n10534), .c(n10525), .o(n10561) );
ao12f01 g06773 ( .a(n4088), .b(n10556), .c(n10547), .o(n10562) );
no02f01 g06774 ( .a(n10562), .b(n10561), .o(n10563) );
no02f01 g06775 ( .a(n10551), .b(n10225), .o(n10564) );
na02f01 g06776 ( .a(n10564), .b(n10207), .o(n10565) );
in01f01 g06777 ( .a(n10565), .o(n10566) );
no02f01 g06778 ( .a(n10216), .b(n3055), .o(n10567) );
no02f01 g06779 ( .a(n10567), .b(n10218), .o(n10568) );
no02f01 g06780 ( .a(n10568), .b(n10566), .o(n10569) );
na02f01 g06781 ( .a(n10568), .b(n10566), .o(n10570) );
in01f01 g06782 ( .a(n10570), .o(n10571) );
no02f01 g06783 ( .a(n10571), .b(n10569), .o(n10572) );
in01f01 g06784 ( .a(n10228), .o(n10573) );
no02f01 g06785 ( .a(n10249), .b(n3055), .o(n10574) );
no02f01 g06786 ( .a(n10250), .b(n10030), .o(n10575) );
no02f01 g06787 ( .a(n10575), .b(n10574), .o(n10576) );
no02f01 g06788 ( .a(n10576), .b(n10573), .o(n10577) );
na02f01 g06789 ( .a(n10576), .b(n10573), .o(n10578) );
in01f01 g06790 ( .a(n10578), .o(n10579) );
no02f01 g06791 ( .a(n10579), .b(n10577), .o(n10580) );
no02f01 g06792 ( .a(n10580), .b(n10572), .o(n10581) );
no02f01 g06793 ( .a(n10581), .b(n10397), .o(n10582) );
ao12f01 g06794 ( .a(n10582), .b(n10563), .c(n10560), .o(n10583) );
ao12f01 g06795 ( .a(n10372), .b(n10252), .c(n10228), .o(n10584) );
in01f01 g06796 ( .a(n10584), .o(n10585) );
no02f01 g06797 ( .a(n10398), .b(n10265), .o(n10586) );
in01f01 g06798 ( .a(n10586), .o(n10587) );
no02f01 g06799 ( .a(n10587), .b(n10585), .o(n10588) );
no02f01 g06800 ( .a(n10586), .b(n10584), .o(n10589) );
no02f01 g06801 ( .a(n10589), .b(n10588), .o(n10590) );
in01f01 g06802 ( .a(n10590), .o(n10591) );
no02f01 g06803 ( .a(n10591), .b(n10397), .o(n10592) );
in01f01 g06804 ( .a(n10575), .o(n10593) );
ao12f01 g06805 ( .a(n10574), .b(n10593), .c(n10228), .o(n10594) );
no02f01 g06806 ( .a(n10244), .b(n10030), .o(n10595) );
no02f01 g06807 ( .a(n10243), .b(n3055), .o(n10596) );
no02f01 g06808 ( .a(n10596), .b(n10595), .o(n10597) );
no02f01 g06809 ( .a(n10597), .b(n10594), .o(n10598) );
na02f01 g06810 ( .a(n10597), .b(n10594), .o(n10599) );
in01f01 g06811 ( .a(n10599), .o(n10600) );
no02f01 g06812 ( .a(n10600), .b(n10598), .o(n10601) );
in01f01 g06813 ( .a(n10601), .o(n10602) );
no02f01 g06814 ( .a(n10602), .b(n10397), .o(n10603) );
no02f01 g06815 ( .a(n10603), .b(n10592), .o(n10604) );
ao12f01 g06816 ( .a(n4088), .b(n10580), .c(n10572), .o(n10605) );
ao12f01 g06817 ( .a(n4088), .b(n10601), .c(n10590), .o(n10606) );
no02f01 g06818 ( .a(n10606), .b(n10605), .o(n10607) );
in01f01 g06819 ( .a(n10607), .o(n10608) );
ao12f01 g06820 ( .a(n10608), .b(n10604), .c(n10583), .o(n10609) );
in01f01 g06821 ( .a(n10277), .o(n10610) );
no02f01 g06822 ( .a(n10409), .b(n10376), .o(n10611) );
oa12f01 g06823 ( .a(n10611), .b(n10287), .c(n10610), .o(n10612) );
no02f01 g06824 ( .a(n10297), .b(n3055), .o(n10613) );
no02f01 g06825 ( .a(n10613), .b(n10299), .o(n10614) );
in01f01 g06826 ( .a(n10614), .o(n10615) );
no02f01 g06827 ( .a(n10615), .b(n10612), .o(n10616) );
na02f01 g06828 ( .a(n10615), .b(n10612), .o(n10617) );
in01f01 g06829 ( .a(n10617), .o(n10618) );
no02f01 g06830 ( .a(n10618), .b(n10616), .o(n10619) );
in01f01 g06831 ( .a(n10619), .o(n10620) );
no02f01 g06832 ( .a(n10620), .b(n10397), .o(n10621) );
na02f01 g06833 ( .a(n10378), .b(n10301), .o(n10622) );
in01f01 g06834 ( .a(n10622), .o(n10623) );
no02f01 g06835 ( .a(n10380), .b(n3055), .o(n10624) );
no02f01 g06836 ( .a(n10624), .b(n10309), .o(n10625) );
no02f01 g06837 ( .a(n10625), .b(n10623), .o(n10626) );
na02f01 g06838 ( .a(n10625), .b(n10623), .o(n10627) );
in01f01 g06839 ( .a(n10627), .o(n10628) );
no02f01 g06840 ( .a(n10628), .b(n10626), .o(n10629) );
in01f01 g06841 ( .a(n10629), .o(n10630) );
no02f01 g06842 ( .a(n10630), .b(n10397), .o(n10631) );
no04f01 g06843 ( .a(n10631), .b(n10621), .c(n10609), .d(n10416), .o(n10632) );
ao12f01 g06844 ( .a(n4088), .b(n10414), .c(n10407), .o(n10633) );
ao12f01 g06845 ( .a(n4088), .b(n10629), .c(n10619), .o(n10634) );
no02f01 g06846 ( .a(n10634), .b(n10633), .o(n10635) );
in01f01 g06847 ( .a(n10635), .o(n10636) );
no02f01 g06848 ( .a(n10636), .b(n10632), .o(n10637) );
no02f01 g06849 ( .a(n10309), .b(n10301), .o(n10638) );
in01f01 g06850 ( .a(n10319), .o(n10639) );
ao12f01 g06851 ( .a(n10383), .b(n10639), .c(n10638), .o(n10640) );
no02f01 g06852 ( .a(n10048), .b(n3055), .o(n10641) );
no02f01 g06853 ( .a(n10641), .b(n10050), .o(n10642) );
no02f01 g06854 ( .a(n10642), .b(n10640), .o(n10643) );
na02f01 g06855 ( .a(n10642), .b(n10640), .o(n10644) );
in01f01 g06856 ( .a(n10644), .o(n10645) );
no03f01 g06857 ( .a(n10645), .b(n10643), .c(n10397), .o(n10646) );
no02f01 g06858 ( .a(n10624), .b(n10379), .o(n10647) );
in01f01 g06859 ( .a(n10647), .o(n10648) );
no02f01 g06860 ( .a(n10317), .b(n3055), .o(n10649) );
no02f01 g06861 ( .a(n10649), .b(n10319), .o(n10650) );
in01f01 g06862 ( .a(n10650), .o(n10651) );
no03f01 g06863 ( .a(n10651), .b(n10648), .c(n10638), .o(n10652) );
no02f01 g06864 ( .a(n10648), .b(n10638), .o(n10653) );
no02f01 g06865 ( .a(n10650), .b(n10653), .o(n10654) );
no02f01 g06866 ( .a(n10654), .b(n10652), .o(n10655) );
in01f01 g06867 ( .a(n10655), .o(n10656) );
no02f01 g06868 ( .a(n10656), .b(n10397), .o(n10657) );
no02f01 g06869 ( .a(n10657), .b(n10646), .o(n10658) );
in01f01 g06870 ( .a(n10658), .o(n10659) );
in01f01 g06871 ( .a(n10320), .o(n10660) );
no02f01 g06872 ( .a(n10660), .b(n10042), .o(n10661) );
no02f01 g06873 ( .a(n10386), .b(n10661), .o(n10662) );
no02f01 g06874 ( .a(n10328), .b(n3055), .o(n10663) );
no02f01 g06875 ( .a(n10663), .b(n10330), .o(n10664) );
no02f01 g06876 ( .a(n10664), .b(n10662), .o(n10665) );
na02f01 g06877 ( .a(n10664), .b(n10662), .o(n10666) );
in01f01 g06878 ( .a(n10666), .o(n10667) );
no03f01 g06879 ( .a(n10667), .b(n10665), .c(n10397), .o(n10668) );
no02f01 g06880 ( .a(n10641), .b(n10383), .o(n10669) );
na02f01 g06881 ( .a(n10669), .b(n10660), .o(n10670) );
no02f01 g06882 ( .a(n10040), .b(n3055), .o(n10671) );
no02f01 g06883 ( .a(n10671), .b(n10042), .o(n10672) );
in01f01 g06884 ( .a(n10672), .o(n10673) );
no02f01 g06885 ( .a(n10673), .b(n10670), .o(n10674) );
na02f01 g06886 ( .a(n10673), .b(n10670), .o(n10675) );
in01f01 g06887 ( .a(n10675), .o(n10676) );
no03f01 g06888 ( .a(n10676), .b(n10674), .c(n10397), .o(n10677) );
no03f01 g06889 ( .a(n10677), .b(n10668), .c(n10659), .o(n10678) );
in01f01 g06890 ( .a(n10678), .o(n10679) );
no02f01 g06891 ( .a(n10645), .b(n10643), .o(n10680) );
ao12f01 g06892 ( .a(n4088), .b(n10655), .c(n10680), .o(n10681) );
no02f01 g06893 ( .a(n10667), .b(n10665), .o(n10682) );
no02f01 g06894 ( .a(n10676), .b(n10674), .o(n10683) );
ao12f01 g06895 ( .a(n4088), .b(n10683), .c(n10682), .o(n10684) );
no02f01 g06896 ( .a(n10684), .b(n10681), .o(n10685) );
oa12f01 g06897 ( .a(n10685), .b(n10679), .c(n10637), .o(n10686) );
in01f01 g06898 ( .a(n10661), .o(n10687) );
no02f01 g06899 ( .a(n10663), .b(n10386), .o(n10688) );
oa12f01 g06900 ( .a(n10688), .b(n10330), .c(n10687), .o(n10689) );
no02f01 g06901 ( .a(n10340), .b(n3055), .o(n10690) );
no02f01 g06902 ( .a(n10690), .b(n10342), .o(n10691) );
in01f01 g06903 ( .a(n10691), .o(n10692) );
no02f01 g06904 ( .a(n10692), .b(n10689), .o(n10693) );
na02f01 g06905 ( .a(n10692), .b(n10689), .o(n10694) );
in01f01 g06906 ( .a(n10694), .o(n10695) );
no02f01 g06907 ( .a(n10695), .b(n10693), .o(n10696) );
in01f01 g06908 ( .a(n10696), .o(n10697) );
no02f01 g06909 ( .a(n10697), .b(n10397), .o(n10698) );
in01f01 g06910 ( .a(n10698), .o(n10699) );
in01f01 g06911 ( .a(n10344), .o(n10700) );
no02f01 g06912 ( .a(n10389), .b(n10700), .o(n10701) );
no02f01 g06913 ( .a(n10391), .b(n3055), .o(n10702) );
no02f01 g06914 ( .a(n10702), .b(n10351), .o(n10703) );
no02f01 g06915 ( .a(n10703), .b(n10701), .o(n10704) );
na02f01 g06916 ( .a(n10703), .b(n10701), .o(n10705) );
in01f01 g06917 ( .a(n10705), .o(n10706) );
no02f01 g06918 ( .a(n10706), .b(n10704), .o(n10707) );
in01f01 g06919 ( .a(n10707), .o(n10708) );
no02f01 g06920 ( .a(n10708), .b(n10397), .o(n10709) );
in01f01 g06921 ( .a(n10709), .o(n10710) );
ao12f01 g06922 ( .a(n10361), .b(n10701), .c(n10394), .o(n10711) );
in01f01 g06923 ( .a(n10711), .o(n10712) );
no02f01 g06924 ( .a(n10390), .b(n3055), .o(n10713) );
no02f01 g06925 ( .a(n10713), .b(n10369), .o(n10714) );
no02f01 g06926 ( .a(n10714), .b(n10712), .o(n10715) );
na02f01 g06927 ( .a(n10714), .b(n10712), .o(n10716) );
in01f01 g06928 ( .a(n10716), .o(n10717) );
no03f01 g06929 ( .a(n10717), .b(n10715), .c(n10397), .o(n10718) );
in01f01 g06930 ( .a(n10702), .o(n10719) );
ao12f01 g06931 ( .a(n10351), .b(n10719), .c(n10701), .o(n10720) );
in01f01 g06932 ( .a(n10720), .o(n10721) );
no02f01 g06933 ( .a(n10392), .b(n3055), .o(n10722) );
no02f01 g06934 ( .a(n10722), .b(n10359), .o(n10723) );
no02f01 g06935 ( .a(n10723), .b(n10721), .o(n10724) );
na02f01 g06936 ( .a(n10723), .b(n10721), .o(n10725) );
in01f01 g06937 ( .a(n10725), .o(n10726) );
no03f01 g06938 ( .a(n10726), .b(n10724), .c(n10397), .o(n10727) );
no02f01 g06939 ( .a(n10727), .b(n10718), .o(n10728) );
na04f01 g06940 ( .a(n10728), .b(n10710), .c(n10699), .d(n10686), .o(n10729) );
no02f01 g06941 ( .a(n10717), .b(n10715), .o(n10730) );
no02f01 g06942 ( .a(n10726), .b(n10724), .o(n10731) );
ao12f01 g06943 ( .a(n4088), .b(n10731), .c(n10730), .o(n10732) );
ao12f01 g06944 ( .a(n4088), .b(n10707), .c(n10696), .o(n10733) );
no02f01 g06945 ( .a(n10733), .b(n10732), .o(n10734) );
na02f01 g06946 ( .a(n10734), .b(n10729), .o(n10735) );
in01f01 g06947 ( .a(n10735), .o(n3521) );
in01f01 g06948 ( .a(n10609), .o(n10737) );
no02f01 g06949 ( .a(n10407), .b(n4088), .o(n10738) );
na02f01 g06950 ( .a(n10407), .b(n4088), .o(n10739) );
ao12f01 g06951 ( .a(n10738), .b(n10739), .c(n10737), .o(n10740) );
in01f01 g06952 ( .a(n10414), .o(n10741) );
no02f01 g06953 ( .a(n10741), .b(n10397), .o(n10742) );
no02f01 g06954 ( .a(n10414), .b(n4088), .o(n10743) );
no02f01 g06955 ( .a(n10743), .b(n10742), .o(n10744) );
no02f01 g06956 ( .a(n10744), .b(n10740), .o(n10745) );
na02f01 g06957 ( .a(n10744), .b(n10740), .o(n10746) );
in01f01 g06958 ( .a(n10746), .o(n10747) );
no02f01 g06959 ( .a(n10747), .b(n10745), .o(n10748) );
no02f01 g06960 ( .a(n10609), .b(n10416), .o(n10749) );
no02f01 g06961 ( .a(n10633), .b(n10749), .o(n10750) );
no02f01 g06962 ( .a(n10619), .b(n4088), .o(n10751) );
no02f01 g06963 ( .a(n10751), .b(n10621), .o(n10752) );
no02f01 g06964 ( .a(n10752), .b(n10750), .o(n10753) );
na02f01 g06965 ( .a(n10752), .b(n10750), .o(n10754) );
in01f01 g06966 ( .a(n10754), .o(n10755) );
no02f01 g06967 ( .a(n10755), .b(n10753), .o(n10756) );
ao12f01 g06968 ( .a(n3521), .b(n10756), .c(n10748), .o(n10757) );
no02f01 g06969 ( .a(n10601), .b(n4088), .o(n10758) );
in01f01 g06970 ( .a(n10758), .o(n10759) );
no02f01 g06971 ( .a(n10605), .b(n10583), .o(n10760) );
ao12f01 g06972 ( .a(n10603), .b(n10760), .c(n10759), .o(n10761) );
in01f01 g06973 ( .a(n10761), .o(n10762) );
no02f01 g06974 ( .a(n10590), .b(n4088), .o(n10763) );
no02f01 g06975 ( .a(n10763), .b(n10592), .o(n10764) );
no02f01 g06976 ( .a(n10764), .b(n10762), .o(n10765) );
na02f01 g06977 ( .a(n10764), .b(n10762), .o(n10766) );
in01f01 g06978 ( .a(n10766), .o(n10767) );
no02f01 g06979 ( .a(n10767), .b(n10765), .o(n10768) );
in01f01 g06980 ( .a(n10739), .o(n10769) );
no02f01 g06981 ( .a(n10769), .b(n10738), .o(n10770) );
in01f01 g06982 ( .a(n10770), .o(n10771) );
no02f01 g06983 ( .a(n10771), .b(n10737), .o(n10772) );
no02f01 g06984 ( .a(n10770), .b(n10609), .o(n10773) );
no02f01 g06985 ( .a(n10773), .b(n10772), .o(n10774) );
ao12f01 g06986 ( .a(n3521), .b(n10774), .c(n10768), .o(n10775) );
no02f01 g06987 ( .a(n10775), .b(n10757), .o(n10776) );
in01f01 g06988 ( .a(n10749), .o(n10777) );
no02f01 g06989 ( .a(n10751), .b(n10633), .o(n10778) );
oa12f01 g06990 ( .a(n10778), .b(n10621), .c(n10777), .o(n10779) );
no02f01 g06991 ( .a(n10629), .b(n4088), .o(n10780) );
no02f01 g06992 ( .a(n10780), .b(n10631), .o(n10781) );
in01f01 g06993 ( .a(n10781), .o(n10782) );
no02f01 g06994 ( .a(n10782), .b(n10779), .o(n10783) );
na02f01 g06995 ( .a(n10782), .b(n10779), .o(n10784) );
in01f01 g06996 ( .a(n10784), .o(n10785) );
no02f01 g06997 ( .a(n10785), .b(n10783), .o(n10786) );
no02f01 g06998 ( .a(n10786), .b(n3521), .o(n10787) );
no02f01 g06999 ( .a(n10655), .b(n4088), .o(n10788) );
no02f01 g07000 ( .a(n10788), .b(n10657), .o(n10789) );
no02f01 g07001 ( .a(n10789), .b(n10637), .o(n10790) );
na02f01 g07002 ( .a(n10789), .b(n10637), .o(n10791) );
in01f01 g07003 ( .a(n10791), .o(n10792) );
no02f01 g07004 ( .a(n10792), .b(n10790), .o(n10793) );
no02f01 g07005 ( .a(n10793), .b(n3521), .o(n10794) );
no02f01 g07006 ( .a(n10794), .b(n10787), .o(n10795) );
na02f01 g07007 ( .a(n10795), .b(n10776), .o(n10796) );
in01f01 g07008 ( .a(n10796), .o(n10797) );
in01f01 g07009 ( .a(n10492), .o(n10798) );
no02f01 g07010 ( .a(n10494), .b(n10798), .o(n10799) );
ao12f01 g07011 ( .a(n10448), .b(n10498), .c(n10799), .o(n10800) );
no02f01 g07012 ( .a(n10508), .b(n4088), .o(n10801) );
no02f01 g07013 ( .a(n10801), .b(n10510), .o(n10802) );
no02f01 g07014 ( .a(n10802), .b(n10800), .o(n10803) );
na02f01 g07015 ( .a(n10802), .b(n10800), .o(n10804) );
in01f01 g07016 ( .a(n10804), .o(n10805) );
no02f01 g07017 ( .a(n10805), .b(n10803), .o(n10806) );
in01f01 g07018 ( .a(n10806), .o(n10807) );
no02f01 g07019 ( .a(n10807), .b(n10735), .o(n10808) );
in01f01 g07020 ( .a(n10808), .o(n10809) );
no02f01 g07021 ( .a(n10447), .b(n4088), .o(n10810) );
no02f01 g07022 ( .a(n10810), .b(n10494), .o(n10811) );
no02f01 g07023 ( .a(n10811), .b(n10798), .o(n10812) );
na02f01 g07024 ( .a(n10811), .b(n10798), .o(n10813) );
in01f01 g07025 ( .a(n10813), .o(n10814) );
no02f01 g07026 ( .a(n10814), .b(n10812), .o(n10815) );
no02f01 g07027 ( .a(n10490), .b(n10479), .o(n10816) );
no02f01 g07028 ( .a(n10487), .b(n10397), .o(n10817) );
no02f01 g07029 ( .a(n10486), .b(n4088), .o(n10818) );
no02f01 g07030 ( .a(n10818), .b(n10817), .o(n10819) );
no02f01 g07031 ( .a(n10819), .b(n10816), .o(n10820) );
na02f01 g07032 ( .a(n10819), .b(n10816), .o(n10821) );
in01f01 g07033 ( .a(n10821), .o(n10822) );
no02f01 g07034 ( .a(n10822), .b(n10820), .o(n10823) );
ao12f01 g07035 ( .a(n3521), .b(n10823), .c(n10815), .o(n10824) );
in01f01 g07036 ( .a(n10824), .o(n10825) );
ao12f01 g07037 ( .a(n10467), .b(n10734), .c(n10729), .o(n10826) );
na03f01 g07038 ( .a(n10734), .b(n10729), .c(n10467), .o(n10827) );
in01f01 g07039 ( .a(n10066), .o(n10828) );
no03f01 g07040 ( .a(n10076), .b(n10828), .c(n10059), .o(n10829) );
in01f01 g07041 ( .a(n10059), .o(n10830) );
ao12f01 g07042 ( .a(n10830), .b(n10077), .c(n10066), .o(n10831) );
no02f01 g07043 ( .a(n10831), .b(n10829), .o(n5618) );
in01f01 g07044 ( .a(n5618), .o(n10833) );
ao12f01 g07045 ( .a(n10826), .b(n10833), .c(n10827), .o(n10834) );
in01f01 g07046 ( .a(n10458), .o(n10835) );
no02f01 g07047 ( .a(n10457), .b(n10397), .o(n10836) );
no02f01 g07048 ( .a(n10836), .b(n10835), .o(n10837) );
no02f01 g07049 ( .a(n10837), .b(n10466), .o(n10838) );
na02f01 g07050 ( .a(n10837), .b(n10466), .o(n10839) );
in01f01 g07051 ( .a(n10839), .o(n10840) );
no02f01 g07052 ( .a(n10840), .b(n10838), .o(n10841) );
in01f01 g07053 ( .a(n10841), .o(n10842) );
no02f01 g07054 ( .a(n10842), .b(n10735), .o(n10843) );
no02f01 g07055 ( .a(n10843), .b(n10834), .o(n10844) );
in01f01 g07056 ( .a(n10468), .o(n10845) );
no02f01 g07057 ( .a(n10845), .b(n10835), .o(n10846) );
no02f01 g07058 ( .a(n10490), .b(n10478), .o(n10847) );
no02f01 g07059 ( .a(n10847), .b(n10846), .o(n10848) );
na02f01 g07060 ( .a(n10847), .b(n10846), .o(n10849) );
in01f01 g07061 ( .a(n10849), .o(n10850) );
no02f01 g07062 ( .a(n10850), .b(n10848), .o(n10851) );
in01f01 g07063 ( .a(n10851), .o(n10852) );
na02f01 g07064 ( .a(n10852), .b(n10844), .o(n10853) );
no02f01 g07065 ( .a(n10841), .b(n3521), .o(n10854) );
no03f01 g07066 ( .a(n10854), .b(n10852), .c(n10844), .o(n10855) );
oa12f01 g07067 ( .a(n10853), .b(n10855), .c(n3521), .o(n10856) );
in01f01 g07068 ( .a(n10823), .o(n10857) );
no02f01 g07069 ( .a(n10857), .b(n10735), .o(n10858) );
in01f01 g07070 ( .a(n10858), .o(n10859) );
in01f01 g07071 ( .a(n10815), .o(n10860) );
no02f01 g07072 ( .a(n10860), .b(n10735), .o(n10861) );
in01f01 g07073 ( .a(n10861), .o(n10862) );
no02f01 g07074 ( .a(n10437), .b(n4088), .o(n10863) );
no02f01 g07075 ( .a(n10863), .b(n10497), .o(n10864) );
in01f01 g07076 ( .a(n10864), .o(n10865) );
no03f01 g07077 ( .a(n10865), .b(n10810), .c(n10799), .o(n10866) );
no02f01 g07078 ( .a(n10810), .b(n10799), .o(n10867) );
no02f01 g07079 ( .a(n10864), .b(n10867), .o(n10868) );
no02f01 g07080 ( .a(n10868), .b(n10866), .o(n10869) );
in01f01 g07081 ( .a(n10869), .o(n10870) );
no02f01 g07082 ( .a(n10870), .b(n10735), .o(n10871) );
in01f01 g07083 ( .a(n10871), .o(n10872) );
na04f01 g07084 ( .a(n10872), .b(n10862), .c(n10859), .d(n10856), .o(n10873) );
ao12f01 g07085 ( .a(n3521), .b(n10869), .c(n10806), .o(n10874) );
in01f01 g07086 ( .a(n10874), .o(n10875) );
na03f01 g07087 ( .a(n10875), .b(n10873), .c(n10825), .o(n10876) );
in01f01 g07088 ( .a(n10515), .o(n10877) );
no02f01 g07089 ( .a(n10877), .b(n10426), .o(n10878) );
no02f01 g07090 ( .a(n10525), .b(n4088), .o(n10879) );
no02f01 g07091 ( .a(n10526), .b(n10397), .o(n10880) );
no02f01 g07092 ( .a(n10880), .b(n10879), .o(n10881) );
in01f01 g07093 ( .a(n10881), .o(n10882) );
no02f01 g07094 ( .a(n10882), .b(n10878), .o(n10883) );
in01f01 g07095 ( .a(n10878), .o(n10884) );
no02f01 g07096 ( .a(n10881), .b(n10884), .o(n10885) );
no02f01 g07097 ( .a(n10885), .b(n10883), .o(n10886) );
in01f01 g07098 ( .a(n10886), .o(n10887) );
no02f01 g07099 ( .a(n10887), .b(n10735), .o(n10888) );
in01f01 g07100 ( .a(n10512), .o(n10889) );
no03f01 g07101 ( .a(n10801), .b(n10889), .c(n10448), .o(n10890) );
no02f01 g07102 ( .a(n10424), .b(n4088), .o(n10891) );
no02f01 g07103 ( .a(n10891), .b(n10426), .o(n10892) );
no02f01 g07104 ( .a(n10892), .b(n10890), .o(n10893) );
na02f01 g07105 ( .a(n10892), .b(n10890), .o(n10894) );
in01f01 g07106 ( .a(n10894), .o(n10895) );
no02f01 g07107 ( .a(n10895), .b(n10893), .o(n10896) );
in01f01 g07108 ( .a(n10896), .o(n10897) );
no02f01 g07109 ( .a(n10897), .b(n10735), .o(n10898) );
no02f01 g07110 ( .a(n10898), .b(n10888), .o(n10899) );
in01f01 g07111 ( .a(n10899), .o(n10900) );
in01f01 g07112 ( .a(n10880), .o(n10901) );
ao12f01 g07113 ( .a(n10879), .b(n10901), .c(n10878), .o(n10902) );
in01f01 g07114 ( .a(n10902), .o(n10903) );
no02f01 g07115 ( .a(n10535), .b(n10397), .o(n10904) );
no02f01 g07116 ( .a(n10534), .b(n4088), .o(n10905) );
no02f01 g07117 ( .a(n10905), .b(n10904), .o(n10906) );
in01f01 g07118 ( .a(n10906), .o(n10907) );
no02f01 g07119 ( .a(n10907), .b(n10903), .o(n10908) );
no02f01 g07120 ( .a(n10906), .b(n10902), .o(n10909) );
no02f01 g07121 ( .a(n10909), .b(n10908), .o(n10910) );
in01f01 g07122 ( .a(n10910), .o(n10911) );
no02f01 g07123 ( .a(n10911), .b(n10735), .o(n10912) );
no02f01 g07124 ( .a(n10912), .b(n10900), .o(n10913) );
ao12f01 g07125 ( .a(n10561), .b(n10537), .c(n10878), .o(n10914) );
no02f01 g07126 ( .a(n10547), .b(n4088), .o(n10915) );
no02f01 g07127 ( .a(n10915), .b(n10549), .o(n10916) );
no02f01 g07128 ( .a(n10916), .b(n10914), .o(n10917) );
na02f01 g07129 ( .a(n10916), .b(n10914), .o(n10918) );
in01f01 g07130 ( .a(n10918), .o(n10919) );
no02f01 g07131 ( .a(n10919), .b(n10917), .o(n10920) );
in01f01 g07132 ( .a(n10920), .o(n10921) );
no02f01 g07133 ( .a(n10921), .b(n10735), .o(n10922) );
in01f01 g07134 ( .a(n10922), .o(n10923) );
na04f01 g07135 ( .a(n10923), .b(n10913), .c(n10876), .d(n10809), .o(n10924) );
ao12f01 g07136 ( .a(n3521), .b(n10920), .c(n10910), .o(n10925) );
ao12f01 g07137 ( .a(n3521), .b(n10896), .c(n10886), .o(n10926) );
no02f01 g07138 ( .a(n10926), .b(n10925), .o(n10927) );
na02f01 g07139 ( .a(n10927), .b(n10924), .o(n10928) );
in01f01 g07140 ( .a(n10560), .o(n10929) );
in01f01 g07141 ( .a(n10563), .o(n10930) );
no02f01 g07142 ( .a(n10930), .b(n10929), .o(n10931) );
in01f01 g07143 ( .a(n10931), .o(n10932) );
no02f01 g07144 ( .a(n10572), .b(n4088), .o(n10933) );
na02f01 g07145 ( .a(n10572), .b(n4088), .o(n10934) );
ao12f01 g07146 ( .a(n10933), .b(n10934), .c(n10932), .o(n10935) );
in01f01 g07147 ( .a(n10935), .o(n10936) );
in01f01 g07148 ( .a(n10580), .o(n10937) );
no02f01 g07149 ( .a(n10937), .b(n10397), .o(n10938) );
no02f01 g07150 ( .a(n10580), .b(n4088), .o(n10939) );
no02f01 g07151 ( .a(n10939), .b(n10938), .o(n10940) );
in01f01 g07152 ( .a(n10940), .o(n10941) );
no02f01 g07153 ( .a(n10941), .b(n10936), .o(n10942) );
no02f01 g07154 ( .a(n10940), .b(n10935), .o(n10943) );
no02f01 g07155 ( .a(n10943), .b(n10942), .o(n10944) );
in01f01 g07156 ( .a(n10944), .o(n10945) );
no02f01 g07157 ( .a(n10945), .b(n10735), .o(n10946) );
no02f01 g07158 ( .a(n10758), .b(n10603), .o(n10947) );
no02f01 g07159 ( .a(n10947), .b(n10760), .o(n10948) );
na02f01 g07160 ( .a(n10947), .b(n10760), .o(n10949) );
in01f01 g07161 ( .a(n10949), .o(n10950) );
no02f01 g07162 ( .a(n10950), .b(n10948), .o(n10951) );
in01f01 g07163 ( .a(n10951), .o(n10952) );
no02f01 g07164 ( .a(n10952), .b(n10735), .o(n10953) );
no03f01 g07165 ( .a(n10549), .b(n10536), .c(n10884), .o(n10954) );
no03f01 g07166 ( .a(n10954), .b(n10915), .c(n10561), .o(n10955) );
no02f01 g07167 ( .a(n10556), .b(n4088), .o(n10956) );
no02f01 g07168 ( .a(n10956), .b(n10558), .o(n10957) );
no02f01 g07169 ( .a(n10957), .b(n10955), .o(n10958) );
na02f01 g07170 ( .a(n10957), .b(n10955), .o(n10959) );
in01f01 g07171 ( .a(n10959), .o(n10960) );
no02f01 g07172 ( .a(n10960), .b(n10958), .o(n10961) );
in01f01 g07173 ( .a(n10961), .o(n10962) );
in01f01 g07174 ( .a(n10934), .o(n10963) );
no02f01 g07175 ( .a(n10963), .b(n10933), .o(n10964) );
no02f01 g07176 ( .a(n10964), .b(n10931), .o(n10965) );
na02f01 g07177 ( .a(n10964), .b(n10931), .o(n10966) );
in01f01 g07178 ( .a(n10966), .o(n10967) );
no02f01 g07179 ( .a(n10967), .b(n10965), .o(n10968) );
in01f01 g07180 ( .a(n10968), .o(n10969) );
ao12f01 g07181 ( .a(n10735), .b(n10969), .c(n10962), .o(n10970) );
no03f01 g07182 ( .a(n10970), .b(n10953), .c(n10946), .o(n10971) );
ao12f01 g07183 ( .a(n3521), .b(n10968), .c(n10961), .o(n10972) );
ao12f01 g07184 ( .a(n3521), .b(n10951), .c(n10944), .o(n10973) );
no02f01 g07185 ( .a(n10973), .b(n10972), .o(n10974) );
in01f01 g07186 ( .a(n10974), .o(n10975) );
ao12f01 g07187 ( .a(n10975), .b(n10971), .c(n10928), .o(n10976) );
in01f01 g07188 ( .a(n10774), .o(n10977) );
no02f01 g07189 ( .a(n10977), .b(n10735), .o(n10978) );
in01f01 g07190 ( .a(n10768), .o(n10979) );
no02f01 g07191 ( .a(n10979), .b(n10735), .o(n10980) );
no02f01 g07192 ( .a(n10980), .b(n10978), .o(n10981) );
in01f01 g07193 ( .a(n10981), .o(n10982) );
in01f01 g07194 ( .a(n10756), .o(n10983) );
no02f01 g07195 ( .a(n10983), .b(n10735), .o(n10984) );
na02f01 g07196 ( .a(n10748), .b(n3521), .o(n10985) );
in01f01 g07197 ( .a(n10985), .o(n10986) );
no03f01 g07198 ( .a(n10986), .b(n10984), .c(n10982), .o(n10987) );
in01f01 g07199 ( .a(n10987), .o(n10988) );
no02f01 g07200 ( .a(n10988), .b(n10976), .o(n10989) );
na02f01 g07201 ( .a(n10786), .b(n3521), .o(n10990) );
in01f01 g07202 ( .a(n10990), .o(n10991) );
na02f01 g07203 ( .a(n10793), .b(n3521), .o(n10992) );
in01f01 g07204 ( .a(n10992), .o(n10993) );
no02f01 g07205 ( .a(n10993), .b(n10991), .o(n10994) );
na02f01 g07206 ( .a(n10994), .b(n10989), .o(n10995) );
in01f01 g07207 ( .a(n10632), .o(n10996) );
no02f01 g07208 ( .a(n10788), .b(n10636), .o(n10997) );
oa12f01 g07209 ( .a(n10997), .b(n10657), .c(n10996), .o(n10998) );
no02f01 g07210 ( .a(n10680), .b(n4088), .o(n10999) );
no02f01 g07211 ( .a(n10999), .b(n10646), .o(n11000) );
in01f01 g07212 ( .a(n11000), .o(n11001) );
no02f01 g07213 ( .a(n11001), .b(n10998), .o(n11002) );
na02f01 g07214 ( .a(n11001), .b(n10998), .o(n11003) );
in01f01 g07215 ( .a(n11003), .o(n11004) );
no02f01 g07216 ( .a(n11004), .b(n11002), .o(n11005) );
in01f01 g07217 ( .a(n11005), .o(n11006) );
no02f01 g07218 ( .a(n11006), .b(n10735), .o(n11007) );
no02f01 g07219 ( .a(n11005), .b(n3521), .o(n11008) );
no02f01 g07220 ( .a(n11008), .b(n11007), .o(n11009) );
na03f01 g07221 ( .a(n11009), .b(n10995), .c(n10797), .o(n11010) );
na02f01 g07222 ( .a(n10995), .b(n10797), .o(n11011) );
in01f01 g07223 ( .a(n11009), .o(n11012) );
na02f01 g07224 ( .a(n11012), .b(n11011), .o(n11013) );
na02f01 g07225 ( .a(n11013), .b(n11010), .o(n248) );
in01f01 g07226 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_22_), .o(n11015) );
in01f01 g07227 ( .a(delay_xor_ln23_unr3_stage2_stallmux_q), .o(n11016) );
no02f01 g07228 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(n11016), .o(n11017) );
in01f01 g07229 ( .a(n11017), .o(n11018) );
no02f01 g07230 ( .a(n11018), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_18_), .o(n11019) );
in01f01 g07231 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_17_), .o(n11020) );
in01f01 g07232 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(n11021) );
no02f01 g07233 ( .a(n11021), .b(delay_xor_ln23_unr3_stage2_stallmux_q), .o(n11022) );
no02f01 g07234 ( .a(n11022), .b(n11020), .o(n11023) );
no02f01 g07235 ( .a(n11018), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_16_), .o(n11024) );
in01f01 g07236 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_15_), .o(n11025) );
no02f01 g07237 ( .a(n11022), .b(n11025), .o(n11026) );
in01f01 g07238 ( .a(n11026), .o(n11027) );
na02f01 g07239 ( .a(n11018), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_16_), .o(n11028) );
ao12f01 g07240 ( .a(n11024), .b(n11028), .c(n11027), .o(n11029) );
in01f01 g07241 ( .a(n11022), .o(n11030) );
no02f01 g07242 ( .a(n11030), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_17_), .o(n11031) );
in01f01 g07243 ( .a(n11031), .o(n11032) );
ao12f01 g07244 ( .a(n11023), .b(n11032), .c(n11029), .o(n11033) );
na02f01 g07245 ( .a(n11018), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_18_), .o(n11034) );
ao12f01 g07246 ( .a(n11019), .b(n11034), .c(n11033), .o(n11035) );
in01f01 g07247 ( .a(n11035), .o(n11036) );
in01f01 g07248 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_20_), .o(n11037) );
in01f01 g07249 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_19_), .o(n11038) );
ao12f01 g07250 ( .a(n11017), .b(n11038), .c(n11037), .o(n11039) );
in01f01 g07251 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_21_), .o(n11040) );
no02f01 g07252 ( .a(n11017), .b(n11040), .o(n11041) );
no02f01 g07253 ( .a(n11041), .b(n11039), .o(n11042) );
na02f01 g07254 ( .a(n11042), .b(n11036), .o(n11043) );
in01f01 g07255 ( .a(n11043), .o(n11044) );
ao22f01 g07256 ( .a(n11044), .b(n11015), .c(n11036), .d(n11017), .o(n11045) );
in01f01 g07257 ( .a(n11045), .o(n11046) );
in01f01 g07258 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_12_), .o(n11047) );
in01f01 g07259 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_11_), .o(n11048) );
ao12f01 g07260 ( .a(n11017), .b(n11048), .c(n11047), .o(n11049) );
in01f01 g07261 ( .a(n11049), .o(n11050) );
no02f01 g07262 ( .a(n11030), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_13_), .o(n11051) );
no02f01 g07263 ( .a(n11051), .b(n11050), .o(n11052) );
no02f01 g07264 ( .a(n11018), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_14_), .o(n11053) );
in01f01 g07265 ( .a(n11053), .o(n11054) );
no02f01 g07266 ( .a(n11030), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_6_), .o(n11055) );
in01f01 g07267 ( .a(n11055), .o(n11056) );
in01f01 g07268 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_2_), .o(n11057) );
in01f01 g07269 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_0_), .o(n11058) );
no02f01 g07270 ( .a(n11017), .b(n11058), .o(n11059) );
in01f01 g07271 ( .a(n11059), .o(n11060) );
no02f01 g07272 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln23_unr3_stage2_stallmux_q), .o(n11061) );
in01f01 g07273 ( .a(n11061), .o(n11062) );
na02f01 g07274 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln23_unr3_stage2_stallmux_q), .o(n11063) );
na02f01 g07275 ( .a(n11063), .b(n11062), .o(n11064) );
no02f01 g07276 ( .a(n11064), .b(delay_sub_ln23_0_unr1_stage2_stallmux_q_1_), .o(n11065) );
no02f01 g07277 ( .a(n11018), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_0_), .o(n11066) );
oa12f01 g07278 ( .a(n11060), .b(n11066), .c(n11065), .o(n11067) );
no02f01 g07279 ( .a(n11030), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_1_), .o(n11068) );
in01f01 g07280 ( .a(n11068), .o(n11069) );
in01f01 g07281 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_1_), .o(n11070) );
no02f01 g07282 ( .a(n11022), .b(n11070), .o(n11071) );
ao12f01 g07283 ( .a(n11071), .b(n11069), .c(n11067), .o(n11072) );
ao12f01 g07284 ( .a(n11022), .b(n11072), .c(n11057), .o(n11073) );
in01f01 g07285 ( .a(n11067), .o(n11074) );
no03f01 g07286 ( .a(n11068), .b(n11074), .c(n11057), .o(n11075) );
no02f01 g07287 ( .a(n11075), .b(n11073), .o(n11076) );
no02f01 g07288 ( .a(n11030), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_4_), .o(n11077) );
no02f01 g07289 ( .a(n11018), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_3_), .o(n11078) );
no02f01 g07290 ( .a(n11018), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_5_), .o(n11079) );
no04f01 g07291 ( .a(n11079), .b(n11078), .c(n11077), .d(n11076), .o(n11080) );
in01f01 g07292 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_6_), .o(n11081) );
na02f01 g07293 ( .a(n11018), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_5_), .o(n11082) );
in01f01 g07294 ( .a(n11082), .o(n11083) );
no02f01 g07295 ( .a(n11083), .b(n11030), .o(n11084) );
na02f01 g07296 ( .a(n11030), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_4_), .o(n11085) );
na02f01 g07297 ( .a(n11018), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_3_), .o(n11086) );
ao12f01 g07298 ( .a(n11077), .b(n11086), .c(n11085), .o(n11087) );
in01f01 g07299 ( .a(n11087), .o(n11088) );
no02f01 g07300 ( .a(n11088), .b(n11079), .o(n11089) );
in01f01 g07301 ( .a(n11089), .o(n11090) );
oa12f01 g07302 ( .a(n11090), .b(n11084), .c(n11081), .o(n11091) );
oa12f01 g07303 ( .a(n11056), .b(n11091), .c(n11080), .o(n11092) );
no02f01 g07304 ( .a(n11018), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_8_), .o(n11093) );
no02f01 g07305 ( .a(n11018), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_7_), .o(n11094) );
no02f01 g07306 ( .a(n11094), .b(n11093), .o(n11095) );
in01f01 g07307 ( .a(n11095), .o(n11096) );
no02f01 g07308 ( .a(n11018), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_9_), .o(n11097) );
no03f01 g07309 ( .a(n11097), .b(n11096), .c(n11092), .o(n11098) );
in01f01 g07310 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_8_), .o(n11099) );
in01f01 g07311 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_7_), .o(n11100) );
ao12f01 g07312 ( .a(n11017), .b(n11100), .c(n11099), .o(n11101) );
na02f01 g07313 ( .a(n11018), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_9_), .o(n11102) );
in01f01 g07314 ( .a(n11102), .o(n11103) );
in01f01 g07315 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_10_), .o(n11104) );
no02f01 g07316 ( .a(n11022), .b(n11104), .o(n11105) );
no03f01 g07317 ( .a(n11105), .b(n11103), .c(n11101), .o(n11106) );
in01f01 g07318 ( .a(n11106), .o(n11107) );
no02f01 g07319 ( .a(n11030), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_10_), .o(n11108) );
in01f01 g07320 ( .a(n11108), .o(n11109) );
oa12f01 g07321 ( .a(n11109), .b(n11107), .c(n11098), .o(n11110) );
no02f01 g07322 ( .a(n11018), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_12_), .o(n11111) );
no02f01 g07323 ( .a(n11018), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_11_), .o(n11112) );
no03f01 g07324 ( .a(n11112), .b(n11111), .c(n11051), .o(n11113) );
in01f01 g07325 ( .a(n11113), .o(n11114) );
na02f01 g07326 ( .a(n11030), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_13_), .o(n11115) );
in01f01 g07327 ( .a(n11115), .o(n11116) );
in01f01 g07328 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_14_), .o(n11117) );
no02f01 g07329 ( .a(n11017), .b(n11117), .o(n11118) );
no02f01 g07330 ( .a(n11118), .b(n11116), .o(n11119) );
oa12f01 g07331 ( .a(n11119), .b(n11114), .c(n11110), .o(n11120) );
ao12f01 g07332 ( .a(n11052), .b(n11120), .c(n11054), .o(n11121) );
no02f01 g07333 ( .a(n11030), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_15_), .o(n11122) );
no03f01 g07334 ( .a(n11122), .b(n11031), .c(n11024), .o(n11123) );
in01f01 g07335 ( .a(n11123), .o(n11124) );
no02f01 g07336 ( .a(n11124), .b(n11019), .o(n11125) );
in01f01 g07337 ( .a(n11125), .o(n11126) );
oa12f01 g07338 ( .a(n11046), .b(n11126), .c(n11121), .o(n11127) );
no02f01 g07339 ( .a(n11018), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_20_), .o(n11128) );
no02f01 g07340 ( .a(n11018), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_19_), .o(n11129) );
no02f01 g07341 ( .a(n11129), .b(n11128), .o(n11130) );
in01f01 g07342 ( .a(n11130), .o(n11131) );
no02f01 g07343 ( .a(n11018), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_21_), .o(n11132) );
no02f01 g07344 ( .a(n11018), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_22_), .o(n11133) );
no03f01 g07345 ( .a(n11133), .b(n11132), .c(n11131), .o(n11134) );
no02f01 g07346 ( .a(n11030), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_26_), .o(n11135) );
no02f01 g07347 ( .a(n11030), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_25_), .o(n11136) );
no02f01 g07348 ( .a(n11136), .b(n11135), .o(n11137) );
ao12f01 g07349 ( .a(n11018), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_23_), .c(delay_sub_ln23_0_unr2_stage2_stallmux_q_24_), .o(n11138) );
in01f01 g07350 ( .a(n11138), .o(n11139) );
na04f01 g07351 ( .a(n11139), .b(n11137), .c(n11134), .d(n11127), .o(n11140) );
in01f01 g07352 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_24_), .o(n11141) );
in01f01 g07353 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_23_), .o(n11142) );
ao12f01 g07354 ( .a(n11017), .b(n11142), .c(n11141), .o(n11143) );
in01f01 g07355 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_26_), .o(n11144) );
in01f01 g07356 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_25_), .o(n11145) );
ao12f01 g07357 ( .a(n11022), .b(n11145), .c(n11144), .o(n11146) );
oa12f01 g07358 ( .a(n11137), .b(n11146), .c(n11143), .o(n11147) );
in01f01 g07359 ( .a(n11147), .o(n11148) );
in01f01 g07360 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_28_), .o(n11149) );
in01f01 g07361 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_27_), .o(n11150) );
ao12f01 g07362 ( .a(n11022), .b(n11150), .c(n11149), .o(n11151) );
no02f01 g07363 ( .a(n11151), .b(n11148), .o(n11152) );
na02f01 g07364 ( .a(n11152), .b(n11140), .o(n11153) );
in01f01 g07365 ( .a(n11063), .o(n11154) );
no02f01 g07366 ( .a(n11030), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_28_), .o(n11155) );
no02f01 g07367 ( .a(n11030), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_27_), .o(n11156) );
no03f01 g07368 ( .a(n11156), .b(n11155), .c(n11154), .o(n11157) );
na02f01 g07369 ( .a(n11157), .b(n11153), .o(n11158) );
no02f01 g07370 ( .a(n11022), .b(n11150), .o(n11159) );
na02f01 g07371 ( .a(n11147), .b(n11140), .o(n11160) );
no02f01 g07372 ( .a(n11160), .b(n11159), .o(n11161) );
no02f01 g07373 ( .a(n11161), .b(n11156), .o(n11162) );
in01f01 g07374 ( .a(n11162), .o(n11163) );
no02f01 g07375 ( .a(n11022), .b(n11149), .o(n11164) );
no02f01 g07376 ( .a(n11164), .b(n11155), .o(n11165) );
no02f01 g07377 ( .a(n11165), .b(n11163), .o(n11166) );
na02f01 g07378 ( .a(n11165), .b(n11163), .o(n11167) );
in01f01 g07379 ( .a(n11167), .o(n11168) );
no02f01 g07380 ( .a(n11168), .b(n11166), .o(n11169) );
no02f01 g07381 ( .a(n11156), .b(n11159), .o(n11170) );
in01f01 g07382 ( .a(n11170), .o(n11171) );
no02f01 g07383 ( .a(n11171), .b(n11160), .o(n11172) );
ao12f01 g07384 ( .a(n11170), .b(n11147), .c(n11140), .o(n11173) );
no02f01 g07385 ( .a(n11173), .b(n11172), .o(n11174) );
no02f01 g07386 ( .a(n11174), .b(n11158), .o(n11175) );
in01f01 g07387 ( .a(n11175), .o(n11176) );
ao12f01 g07388 ( .a(n11158), .b(n11176), .c(n11169), .o(n11177) );
in01f01 g07389 ( .a(n11157), .o(n11178) );
ao12f01 g07390 ( .a(n11178), .b(n11152), .c(n11140), .o(n11179) );
in01f01 g07391 ( .a(n11110), .o(n11180) );
in01f01 g07392 ( .a(n11112), .o(n11181) );
no02f01 g07393 ( .a(n11017), .b(n11048), .o(n11182) );
ao12f01 g07394 ( .a(n11182), .b(n11181), .c(n11180), .o(n11183) );
in01f01 g07395 ( .a(n11183), .o(n11184) );
no02f01 g07396 ( .a(n11017), .b(n11047), .o(n11185) );
no02f01 g07397 ( .a(n11185), .b(n11111), .o(n11186) );
in01f01 g07398 ( .a(n11186), .o(n11187) );
no02f01 g07399 ( .a(n11187), .b(n11184), .o(n11188) );
no02f01 g07400 ( .a(n11186), .b(n11183), .o(n11189) );
no02f01 g07401 ( .a(n11189), .b(n11188), .o(n11190) );
in01f01 g07402 ( .a(n11190), .o(n11191) );
no02f01 g07403 ( .a(n11191), .b(n11179), .o(n11192) );
in01f01 g07404 ( .a(n11092), .o(n11193) );
in01f01 g07405 ( .a(n11094), .o(n11194) );
no02f01 g07406 ( .a(n11017), .b(n11100), .o(n11195) );
ao12f01 g07407 ( .a(n11195), .b(n11194), .c(n11193), .o(n11196) );
in01f01 g07408 ( .a(n11196), .o(n11197) );
no02f01 g07409 ( .a(n11017), .b(n11099), .o(n11198) );
no02f01 g07410 ( .a(n11198), .b(n11093), .o(n11199) );
in01f01 g07411 ( .a(n11199), .o(n11200) );
no02f01 g07412 ( .a(n11200), .b(n11197), .o(n11201) );
no02f01 g07413 ( .a(n11199), .b(n11196), .o(n11202) );
no02f01 g07414 ( .a(n11202), .b(n11201), .o(n11203) );
no02f01 g07415 ( .a(n11195), .b(n11094), .o(n11204) );
no02f01 g07416 ( .a(n11204), .b(n11092), .o(n11205) );
na02f01 g07417 ( .a(n11204), .b(n11092), .o(n11206) );
in01f01 g07418 ( .a(n11206), .o(n11207) );
no02f01 g07419 ( .a(n11207), .b(n11205), .o(n11208) );
ao12f01 g07420 ( .a(n11203), .b(n11208), .c(n11158), .o(n11209) );
ao12f01 g07421 ( .a(n11101), .b(n11095), .c(n11193), .o(n11210) );
in01f01 g07422 ( .a(n11210), .o(n11211) );
no02f01 g07423 ( .a(n11103), .b(n11097), .o(n11212) );
in01f01 g07424 ( .a(n11212), .o(n11213) );
no02f01 g07425 ( .a(n11213), .b(n11211), .o(n11214) );
no02f01 g07426 ( .a(n11212), .b(n11210), .o(n11215) );
no02f01 g07427 ( .a(n11215), .b(n11214), .o(n11216) );
in01f01 g07428 ( .a(n11216), .o(n11217) );
no02f01 g07429 ( .a(n11217), .b(n11158), .o(n11218) );
in01f01 g07430 ( .a(n11218), .o(n11219) );
na02f01 g07431 ( .a(n11219), .b(n11209), .o(n11220) );
no03f01 g07432 ( .a(n11103), .b(n11101), .c(n11098), .o(n11221) );
in01f01 g07433 ( .a(n11221), .o(n11222) );
no02f01 g07434 ( .a(n11108), .b(n11105), .o(n11223) );
in01f01 g07435 ( .a(n11223), .o(n11224) );
no02f01 g07436 ( .a(n11224), .b(n11222), .o(n11225) );
no02f01 g07437 ( .a(n11223), .b(n11221), .o(n11226) );
no02f01 g07438 ( .a(n11226), .b(n11225), .o(n11227) );
no02f01 g07439 ( .a(n11227), .b(n11158), .o(n11228) );
no02f01 g07440 ( .a(n11216), .b(n11179), .o(n11229) );
no02f01 g07441 ( .a(n11229), .b(n11228), .o(n11230) );
na02f01 g07442 ( .a(n11227), .b(n11158), .o(n11231) );
in01f01 g07443 ( .a(n11231), .o(n11232) );
ao12f01 g07444 ( .a(n11232), .b(n11230), .c(n11220), .o(n11233) );
no02f01 g07445 ( .a(n11030), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_2_), .o(n11234) );
no02f01 g07446 ( .a(n11022), .b(n11057), .o(n11235) );
no02f01 g07447 ( .a(n11235), .b(n11234), .o(n11236) );
no02f01 g07448 ( .a(n11236), .b(n11072), .o(n11237) );
na02f01 g07449 ( .a(n11236), .b(n11072), .o(n11238) );
in01f01 g07450 ( .a(n11238), .o(n11239) );
no02f01 g07451 ( .a(n11239), .b(n11237), .o(n11240) );
in01f01 g07452 ( .a(n11240), .o(n11241) );
no02f01 g07453 ( .a(n11241), .b(n11158), .o(n11242) );
in01f01 g07454 ( .a(n11242), .o(n11243) );
no02f01 g07455 ( .a(n11240), .b(n11179), .o(n11244) );
no02f01 g07456 ( .a(n11071), .b(n11068), .o(n11245) );
in01f01 g07457 ( .a(n11245), .o(n11246) );
no02f01 g07458 ( .a(n11246), .b(n11067), .o(n11247) );
no02f01 g07459 ( .a(n11245), .b(n11074), .o(n11248) );
no02f01 g07460 ( .a(n11248), .b(n11247), .o(n11249) );
no02f01 g07461 ( .a(n11249), .b(n11158), .o(n11250) );
in01f01 g07462 ( .a(n11250), .o(n11251) );
no02f01 g07463 ( .a(n11066), .b(n11059), .o(n11252) );
no02f01 g07464 ( .a(n11252), .b(n11065), .o(n11253) );
na02f01 g07465 ( .a(n11252), .b(n11065), .o(n11254) );
in01f01 g07466 ( .a(n11254), .o(n11255) );
no02f01 g07467 ( .a(n11255), .b(n11253), .o(n11256) );
no02f01 g07468 ( .a(n11256), .b(n11179), .o(n11257) );
na02f01 g07469 ( .a(n11256), .b(n11179), .o(n11258) );
in01f01 g07470 ( .a(delay_sub_ln23_0_unr1_stage2_stallmux_q_1_), .o(n11259) );
no02f01 g07471 ( .a(n11064), .b(n11259), .o(n11260) );
ao12f01 g07472 ( .a(delay_sub_ln23_0_unr1_stage2_stallmux_q_1_), .b(n11063), .c(n11062), .o(n11261) );
no02f01 g07473 ( .a(n11261), .b(n11260), .o(n11262) );
ao12f01 g07474 ( .a(n11257), .b(n11262), .c(n11258), .o(n11263) );
na02f01 g07475 ( .a(n11249), .b(n11158), .o(n11264) );
in01f01 g07476 ( .a(n11264), .o(n11265) );
oa12f01 g07477 ( .a(n11251), .b(n11265), .c(n11263), .o(n11266) );
oa12f01 g07478 ( .a(n11243), .b(n11266), .c(n11244), .o(n11267) );
in01f01 g07479 ( .a(n11077), .o(n11268) );
no02f01 g07480 ( .a(n11078), .b(n11076), .o(n11269) );
ao12f01 g07481 ( .a(n11087), .b(n11269), .c(n11268), .o(n11270) );
in01f01 g07482 ( .a(n11270), .o(n11271) );
no02f01 g07483 ( .a(n11083), .b(n11079), .o(n11272) );
in01f01 g07484 ( .a(n11272), .o(n11273) );
no02f01 g07485 ( .a(n11273), .b(n11271), .o(n11274) );
no02f01 g07486 ( .a(n11272), .b(n11270), .o(n11275) );
no02f01 g07487 ( .a(n11275), .b(n11274), .o(n11276) );
in01f01 g07488 ( .a(n11276), .o(n11277) );
no02f01 g07489 ( .a(n11277), .b(n11179), .o(n11278) );
in01f01 g07490 ( .a(n11086), .o(n11279) );
no02f01 g07491 ( .a(n11279), .b(n11078), .o(n11280) );
in01f01 g07492 ( .a(n11280), .o(n11281) );
no03f01 g07493 ( .a(n11281), .b(n11075), .c(n11073), .o(n11282) );
no02f01 g07494 ( .a(n11280), .b(n11076), .o(n11283) );
no02f01 g07495 ( .a(n11283), .b(n11282), .o(n11284) );
in01f01 g07496 ( .a(n11284), .o(n11285) );
no02f01 g07497 ( .a(n11285), .b(n11158), .o(n11286) );
no02f01 g07498 ( .a(n11269), .b(n11279), .o(n11287) );
in01f01 g07499 ( .a(n11287), .o(n11288) );
na02f01 g07500 ( .a(n11085), .b(n11268), .o(n11289) );
no02f01 g07501 ( .a(n11289), .b(n11288), .o(n11290) );
na02f01 g07502 ( .a(n11289), .b(n11288), .o(n11291) );
in01f01 g07503 ( .a(n11291), .o(n11292) );
no02f01 g07504 ( .a(n11292), .b(n11290), .o(n11293) );
in01f01 g07505 ( .a(n11293), .o(n11294) );
no02f01 g07506 ( .a(n11294), .b(n11158), .o(n11295) );
no03f01 g07507 ( .a(n11295), .b(n11286), .c(n11278), .o(n11296) );
in01f01 g07508 ( .a(n11296), .o(n11297) );
no02f01 g07509 ( .a(n11297), .b(n11267), .o(n11298) );
in01f01 g07510 ( .a(n11298), .o(n11299) );
in01f01 g07511 ( .a(n11080), .o(n11300) );
na03f01 g07512 ( .a(n11090), .b(n11082), .c(n11300), .o(n11301) );
no02f01 g07513 ( .a(n11022), .b(n11081), .o(n11302) );
no02f01 g07514 ( .a(n11302), .b(n11055), .o(n11303) );
in01f01 g07515 ( .a(n11303), .o(n11304) );
no02f01 g07516 ( .a(n11304), .b(n11301), .o(n11305) );
na02f01 g07517 ( .a(n11304), .b(n11301), .o(n11306) );
in01f01 g07518 ( .a(n11306), .o(n11307) );
no02f01 g07519 ( .a(n11307), .b(n11305), .o(n11308) );
no02f01 g07520 ( .a(n11308), .b(n11179), .o(n11309) );
no02f01 g07521 ( .a(n11276), .b(n11158), .o(n11310) );
no02f01 g07522 ( .a(n11310), .b(n11309), .o(n11311) );
na02f01 g07523 ( .a(n11311), .b(n11299), .o(n11312) );
na02f01 g07524 ( .a(n11308), .b(n11179), .o(n11313) );
ao12f01 g07525 ( .a(n11179), .b(n11293), .c(n11284), .o(n11314) );
in01f01 g07526 ( .a(n11314), .o(n11315) );
no02f01 g07527 ( .a(n11315), .b(n11278), .o(n11316) );
ao12f01 g07528 ( .a(n11316), .b(n11313), .c(n11312), .o(n11317) );
na02f01 g07529 ( .a(n11208), .b(n11179), .o(n11318) );
in01f01 g07530 ( .a(n11318), .o(n11319) );
in01f01 g07531 ( .a(n11203), .o(n11320) );
no02f01 g07532 ( .a(n11320), .b(n11179), .o(n11321) );
no03f01 g07533 ( .a(n11232), .b(n11218), .c(n11321), .o(n11322) );
in01f01 g07534 ( .a(n11322), .o(n11323) );
no03f01 g07535 ( .a(n11323), .b(n11319), .c(n11317), .o(n11324) );
no02f01 g07536 ( .a(n11182), .b(n11112), .o(n11325) );
no02f01 g07537 ( .a(n11325), .b(n11110), .o(n11326) );
na02f01 g07538 ( .a(n11325), .b(n11110), .o(n11327) );
in01f01 g07539 ( .a(n11327), .o(n11328) );
no02f01 g07540 ( .a(n11328), .b(n11326), .o(n11329) );
in01f01 g07541 ( .a(n11329), .o(n11330) );
no02f01 g07542 ( .a(n11330), .b(n11158), .o(n11331) );
in01f01 g07543 ( .a(n11331), .o(n11332) );
oa12f01 g07544 ( .a(n11332), .b(n11324), .c(n11233), .o(n11333) );
no02f01 g07545 ( .a(n11190), .b(n11158), .o(n11334) );
no02f01 g07546 ( .a(n11329), .b(n11179), .o(n11335) );
no02f01 g07547 ( .a(n11335), .b(n11334), .o(n11336) );
ao12f01 g07548 ( .a(n11192), .b(n11336), .c(n11333), .o(n11337) );
no02f01 g07549 ( .a(n11112), .b(n11111), .o(n11338) );
ao12f01 g07550 ( .a(n11049), .b(n11338), .c(n11180), .o(n11339) );
no02f01 g07551 ( .a(n11116), .b(n11051), .o(n11340) );
no02f01 g07552 ( .a(n11340), .b(n11339), .o(n11341) );
na02f01 g07553 ( .a(n11340), .b(n11339), .o(n11342) );
in01f01 g07554 ( .a(n11342), .o(n11343) );
no02f01 g07555 ( .a(n11343), .b(n11341), .o(n11344) );
in01f01 g07556 ( .a(n11344), .o(n11345) );
no02f01 g07557 ( .a(n11345), .b(n11158), .o(n11346) );
in01f01 g07558 ( .a(n11346), .o(n11347) );
no02f01 g07559 ( .a(n11344), .b(n11179), .o(n11348) );
ao12f01 g07560 ( .a(n11051), .b(n11339), .c(n11115), .o(n11349) );
no02f01 g07561 ( .a(n11118), .b(n11053), .o(n11350) );
in01f01 g07562 ( .a(n11350), .o(n11351) );
no02f01 g07563 ( .a(n11351), .b(n11349), .o(n11352) );
na02f01 g07564 ( .a(n11351), .b(n11349), .o(n11353) );
in01f01 g07565 ( .a(n11353), .o(n11354) );
no02f01 g07566 ( .a(n11354), .b(n11352), .o(n11355) );
no02f01 g07567 ( .a(n11355), .b(n11158), .o(n11356) );
no02f01 g07568 ( .a(n11356), .b(n11348), .o(n11357) );
in01f01 g07569 ( .a(n11357), .o(n11358) );
ao12f01 g07570 ( .a(n11358), .b(n11347), .c(n11337), .o(n11359) );
na02f01 g07571 ( .a(n11355), .b(n11158), .o(n11360) );
in01f01 g07572 ( .a(n11360), .o(n11361) );
no02f01 g07573 ( .a(n11122), .b(n11121), .o(n11362) );
no02f01 g07574 ( .a(n11362), .b(n11026), .o(n11363) );
in01f01 g07575 ( .a(n11363), .o(n11364) );
in01f01 g07576 ( .a(n11024), .o(n11365) );
na02f01 g07577 ( .a(n11028), .b(n11365), .o(n11366) );
no02f01 g07578 ( .a(n11366), .b(n11364), .o(n11367) );
na02f01 g07579 ( .a(n11366), .b(n11364), .o(n11368) );
in01f01 g07580 ( .a(n11368), .o(n11369) );
no03f01 g07581 ( .a(n11369), .b(n11367), .c(n11158), .o(n11370) );
in01f01 g07582 ( .a(n11121), .o(n11371) );
no02f01 g07583 ( .a(n11122), .b(n11026), .o(n11372) );
in01f01 g07584 ( .a(n11372), .o(n11373) );
no02f01 g07585 ( .a(n11373), .b(n11371), .o(n11374) );
no02f01 g07586 ( .a(n11372), .b(n11121), .o(n11375) );
no02f01 g07587 ( .a(n11375), .b(n11374), .o(n11376) );
in01f01 g07588 ( .a(n11376), .o(n11377) );
no02f01 g07589 ( .a(n11377), .b(n11158), .o(n11378) );
no02f01 g07590 ( .a(n11378), .b(n11370), .o(n11379) );
in01f01 g07591 ( .a(n11379), .o(n11380) );
ao12f01 g07592 ( .a(n11029), .b(n11362), .c(n11365), .o(n11381) );
in01f01 g07593 ( .a(n11381), .o(n11382) );
no02f01 g07594 ( .a(n11031), .b(n11023), .o(n11383) );
in01f01 g07595 ( .a(n11383), .o(n11384) );
no02f01 g07596 ( .a(n11384), .b(n11382), .o(n11385) );
no02f01 g07597 ( .a(n11383), .b(n11381), .o(n11386) );
no03f01 g07598 ( .a(n11386), .b(n11385), .c(n11158), .o(n11387) );
no02f01 g07599 ( .a(n11124), .b(n11121), .o(n11388) );
in01f01 g07600 ( .a(n11388), .o(n11389) );
na02f01 g07601 ( .a(n11389), .b(n11033), .o(n11390) );
in01f01 g07602 ( .a(n11019), .o(n11391) );
na02f01 g07603 ( .a(n11034), .b(n11391), .o(n11392) );
no02f01 g07604 ( .a(n11392), .b(n11390), .o(n11393) );
na02f01 g07605 ( .a(n11392), .b(n11390), .o(n11394) );
in01f01 g07606 ( .a(n11394), .o(n11395) );
no03f01 g07607 ( .a(n11395), .b(n11393), .c(n11158), .o(n11396) );
no03f01 g07608 ( .a(n11396), .b(n11387), .c(n11380), .o(n11397) );
in01f01 g07609 ( .a(n11397), .o(n11398) );
in01f01 g07610 ( .a(n11129), .o(n11399) );
no02f01 g07611 ( .a(n11017), .b(n11038), .o(n11400) );
no02f01 g07612 ( .a(n11389), .b(n11019), .o(n11401) );
no02f01 g07613 ( .a(n11401), .b(n11035), .o(n11402) );
in01f01 g07614 ( .a(n11402), .o(n11403) );
ao12f01 g07615 ( .a(n11400), .b(n11403), .c(n11399), .o(n11404) );
in01f01 g07616 ( .a(n11404), .o(n11405) );
no02f01 g07617 ( .a(n11017), .b(n11037), .o(n11406) );
no02f01 g07618 ( .a(n11406), .b(n11128), .o(n11407) );
in01f01 g07619 ( .a(n11407), .o(n11408) );
no02f01 g07620 ( .a(n11408), .b(n11405), .o(n11409) );
no02f01 g07621 ( .a(n11407), .b(n11404), .o(n11410) );
no03f01 g07622 ( .a(n11410), .b(n11409), .c(n11158), .o(n11411) );
no02f01 g07623 ( .a(n11400), .b(n11129), .o(n11412) );
no02f01 g07624 ( .a(n11412), .b(n11402), .o(n11413) );
na02f01 g07625 ( .a(n11412), .b(n11402), .o(n11414) );
in01f01 g07626 ( .a(n11414), .o(n11415) );
no03f01 g07627 ( .a(n11415), .b(n11413), .c(n11158), .o(n11416) );
na02f01 g07628 ( .a(n11401), .b(n11130), .o(n11417) );
ao12f01 g07629 ( .a(n11039), .b(n11130), .c(n11035), .o(n11418) );
na02f01 g07630 ( .a(n11418), .b(n11417), .o(n11419) );
in01f01 g07631 ( .a(n11419), .o(n11420) );
no02f01 g07632 ( .a(n11132), .b(n11041), .o(n11421) );
no02f01 g07633 ( .a(n11421), .b(n11420), .o(n11422) );
na02f01 g07634 ( .a(n11421), .b(n11420), .o(n11423) );
in01f01 g07635 ( .a(n11423), .o(n11424) );
no03f01 g07636 ( .a(n11424), .b(n11422), .c(n11158), .o(n11425) );
oa12f01 g07637 ( .a(n11130), .b(n11401), .c(n11043), .o(n11426) );
no02f01 g07638 ( .a(n11426), .b(n11132), .o(n11427) );
no02f01 g07639 ( .a(n11017), .b(n11015), .o(n11428) );
no02f01 g07640 ( .a(n11428), .b(n11133), .o(n11429) );
in01f01 g07641 ( .a(n11429), .o(n11430) );
no02f01 g07642 ( .a(n11430), .b(n11427), .o(n11431) );
na02f01 g07643 ( .a(n11430), .b(n11427), .o(n11432) );
in01f01 g07644 ( .a(n11432), .o(n11433) );
no03f01 g07645 ( .a(n11433), .b(n11431), .c(n11158), .o(n11434) );
no04f01 g07646 ( .a(n11434), .b(n11425), .c(n11416), .d(n11411), .o(n11435) );
in01f01 g07647 ( .a(n11435), .o(n11436) );
no04f01 g07648 ( .a(n11436), .b(n11398), .c(n11361), .d(n11359), .o(n11437) );
no02f01 g07649 ( .a(n11424), .b(n11422), .o(n11438) );
no02f01 g07650 ( .a(n11433), .b(n11431), .o(n11439) );
ao12f01 g07651 ( .a(n11179), .b(n11439), .c(n11438), .o(n11440) );
no02f01 g07652 ( .a(n11410), .b(n11409), .o(n11441) );
no02f01 g07653 ( .a(n11415), .b(n11413), .o(n11442) );
ao12f01 g07654 ( .a(n11179), .b(n11442), .c(n11441), .o(n11443) );
no02f01 g07655 ( .a(n11369), .b(n11367), .o(n11444) );
ao12f01 g07656 ( .a(n11179), .b(n11376), .c(n11444), .o(n11445) );
no02f01 g07657 ( .a(n11386), .b(n11385), .o(n11446) );
no02f01 g07658 ( .a(n11395), .b(n11393), .o(n11447) );
ao12f01 g07659 ( .a(n11179), .b(n11447), .c(n11446), .o(n11448) );
no02f01 g07660 ( .a(n11448), .b(n11445), .o(n11449) );
in01f01 g07661 ( .a(n11449), .o(n11450) );
no02f01 g07662 ( .a(n11450), .b(n11443), .o(n11451) );
in01f01 g07663 ( .a(n11451), .o(n11452) );
no02f01 g07664 ( .a(n11452), .b(n11440), .o(n11453) );
in01f01 g07665 ( .a(n11453), .o(n11454) );
in01f01 g07666 ( .a(n11127), .o(n11455) );
in01f01 g07667 ( .a(n11134), .o(n11456) );
no02f01 g07668 ( .a(n11456), .b(n11455), .o(n11457) );
no02f01 g07669 ( .a(n11017), .b(n11142), .o(n11458) );
no02f01 g07670 ( .a(n11018), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_23_), .o(n11459) );
in01f01 g07671 ( .a(n11459), .o(n11460) );
ao12f01 g07672 ( .a(n11458), .b(n11460), .c(n11457), .o(n11461) );
in01f01 g07673 ( .a(n11461), .o(n11462) );
no02f01 g07674 ( .a(n11017), .b(n11141), .o(n11463) );
no02f01 g07675 ( .a(n11018), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_24_), .o(n11464) );
no02f01 g07676 ( .a(n11464), .b(n11463), .o(n11465) );
in01f01 g07677 ( .a(n11465), .o(n11466) );
no02f01 g07678 ( .a(n11466), .b(n11462), .o(n11467) );
no02f01 g07679 ( .a(n11465), .b(n11461), .o(n11468) );
no03f01 g07680 ( .a(n11468), .b(n11467), .c(n11179), .o(n11469) );
no02f01 g07681 ( .a(n11459), .b(n11458), .o(n11470) );
in01f01 g07682 ( .a(n11470), .o(n11471) );
no02f01 g07683 ( .a(n11471), .b(n11457), .o(n11472) );
no03f01 g07684 ( .a(n11470), .b(n11456), .c(n11455), .o(n11473) );
no02f01 g07685 ( .a(n11473), .b(n11472), .o(n11474) );
in01f01 g07686 ( .a(n11474), .o(n11475) );
no02f01 g07687 ( .a(n11475), .b(n11158), .o(n11476) );
no02f01 g07688 ( .a(n11476), .b(n11469), .o(n11477) );
oa12f01 g07689 ( .a(n11477), .b(n11454), .c(n11437), .o(n11478) );
no02f01 g07690 ( .a(n11022), .b(n11145), .o(n11479) );
in01f01 g07691 ( .a(n11479), .o(n11480) );
ao12f01 g07692 ( .a(n11143), .b(n11139), .c(n11457), .o(n11481) );
ao12f01 g07693 ( .a(n11136), .b(n11481), .c(n11480), .o(n11482) );
no02f01 g07694 ( .a(n11022), .b(n11144), .o(n11483) );
no02f01 g07695 ( .a(n11483), .b(n11135), .o(n11484) );
in01f01 g07696 ( .a(n11484), .o(n11485) );
no02f01 g07697 ( .a(n11485), .b(n11482), .o(n11486) );
na02f01 g07698 ( .a(n11485), .b(n11482), .o(n11487) );
in01f01 g07699 ( .a(n11487), .o(n11488) );
no02f01 g07700 ( .a(n11488), .b(n11486), .o(n11489) );
in01f01 g07701 ( .a(n11489), .o(n11490) );
in01f01 g07702 ( .a(n11481), .o(n11491) );
no02f01 g07703 ( .a(n11479), .b(n11136), .o(n11492) );
in01f01 g07704 ( .a(n11492), .o(n11493) );
no02f01 g07705 ( .a(n11493), .b(n11491), .o(n11494) );
no02f01 g07706 ( .a(n11492), .b(n11481), .o(n11495) );
no02f01 g07707 ( .a(n11495), .b(n11494), .o(n11496) );
no02f01 g07708 ( .a(n11496), .b(n11158), .o(n11497) );
no02f01 g07709 ( .a(n11497), .b(n11490), .o(n11498) );
no02f01 g07710 ( .a(n11468), .b(n11467), .o(n11499) );
ao12f01 g07711 ( .a(n11499), .b(n11474), .c(n11158), .o(n11500) );
in01f01 g07712 ( .a(n11500), .o(n11501) );
oa12f01 g07713 ( .a(n11501), .b(n11498), .c(n11158), .o(n11502) );
in01f01 g07714 ( .a(n11502), .o(n11503) );
no02f01 g07715 ( .a(n11490), .b(n11179), .o(n11504) );
na02f01 g07716 ( .a(n11496), .b(n11158), .o(n11505) );
in01f01 g07717 ( .a(n11505), .o(n11506) );
no02f01 g07718 ( .a(n11506), .b(n11504), .o(n11507) );
in01f01 g07719 ( .a(n11507), .o(n11508) );
ao12f01 g07720 ( .a(n11508), .b(n11503), .c(n11478), .o(n11509) );
no03f01 g07721 ( .a(n11168), .b(n11166), .c(n11179), .o(n11510) );
na02f01 g07722 ( .a(n11174), .b(n11158), .o(n11511) );
in01f01 g07723 ( .a(n11511), .o(n11512) );
no02f01 g07724 ( .a(n11512), .b(n11510), .o(n11513) );
oa12f01 g07725 ( .a(n11513), .b(n11509), .c(n11177), .o(n11514) );
in01f01 g07726 ( .a(n11514), .o(n11515) );
in01f01 g07727 ( .a(n11509), .o(n11516) );
ao12f01 g07728 ( .a(n11512), .b(n11516), .c(n11176), .o(n11517) );
in01f01 g07729 ( .a(n11517), .o(n11518) );
no02f01 g07730 ( .a(n11169), .b(n11158), .o(n11519) );
no02f01 g07731 ( .a(n11519), .b(n11510), .o(n11520) );
no02f01 g07732 ( .a(n11520), .b(n11518), .o(n11521) );
na02f01 g07733 ( .a(n11520), .b(n11518), .o(n11522) );
in01f01 g07734 ( .a(n11522), .o(n11523) );
no02f01 g07735 ( .a(n11523), .b(n11521), .o(n11524) );
in01f01 g07736 ( .a(n11524), .o(n11525) );
no02f01 g07737 ( .a(n11525), .b(n11515), .o(n11526) );
no02f01 g07738 ( .a(n11474), .b(n11179), .o(n11527) );
no02f01 g07739 ( .a(n11527), .b(n11476), .o(n11528) );
in01f01 g07740 ( .a(n11528), .o(n11529) );
no03f01 g07741 ( .a(n11529), .b(n11454), .c(n11437), .o(n11530) );
no02f01 g07742 ( .a(n11454), .b(n11437), .o(n11531) );
no02f01 g07743 ( .a(n11528), .b(n11531), .o(n11532) );
no02f01 g07744 ( .a(n11532), .b(n11530), .o(n11533) );
in01f01 g07745 ( .a(n11533), .o(n11534) );
no02f01 g07746 ( .a(n11534), .b(n11515), .o(n11535) );
no02f01 g07747 ( .a(n11438), .b(n11179), .o(n11536) );
in01f01 g07748 ( .a(n11536), .o(n11537) );
no02f01 g07749 ( .a(n11361), .b(n11359), .o(n11538) );
in01f01 g07750 ( .a(n11538), .o(n11539) );
no02f01 g07751 ( .a(n11398), .b(n11539), .o(n11540) );
no02f01 g07752 ( .a(n11416), .b(n11411), .o(n11541) );
ao12f01 g07753 ( .a(n11452), .b(n11541), .c(n11540), .o(n11542) );
ao12f01 g07754 ( .a(n11425), .b(n11542), .c(n11537), .o(n11543) );
in01f01 g07755 ( .a(n11543), .o(n11544) );
no02f01 g07756 ( .a(n11439), .b(n11179), .o(n11545) );
no02f01 g07757 ( .a(n11545), .b(n11434), .o(n11546) );
no02f01 g07758 ( .a(n11546), .b(n11544), .o(n11547) );
na02f01 g07759 ( .a(n11546), .b(n11544), .o(n11548) );
in01f01 g07760 ( .a(n11548), .o(n11549) );
no02f01 g07761 ( .a(n11549), .b(n11547), .o(n11550) );
no02f01 g07762 ( .a(n11550), .b(n11515), .o(n11551) );
no02f01 g07763 ( .a(n11324), .b(n11233), .o(n11552) );
no02f01 g07764 ( .a(n11335), .b(n11331), .o(n11553) );
no02f01 g07765 ( .a(n11553), .b(n11552), .o(n11554) );
na02f01 g07766 ( .a(n11553), .b(n11552), .o(n11555) );
in01f01 g07767 ( .a(n11555), .o(n11556) );
no02f01 g07768 ( .a(n11556), .b(n11554), .o(n11557) );
in01f01 g07769 ( .a(n11557), .o(n11558) );
no02f01 g07770 ( .a(n11558), .b(n11515), .o(n11559) );
in01f01 g07771 ( .a(n11559), .o(n11560) );
in01f01 g07772 ( .a(n11321), .o(n11561) );
no02f01 g07773 ( .a(n11319), .b(n11317), .o(n11562) );
ao12f01 g07774 ( .a(n11209), .b(n11562), .c(n11561), .o(n11563) );
in01f01 g07775 ( .a(n11563), .o(n11564) );
ao12f01 g07776 ( .a(n11229), .b(n11564), .c(n11219), .o(n11565) );
no02f01 g07777 ( .a(n11232), .b(n11228), .o(n11566) );
no02f01 g07778 ( .a(n11566), .b(n11565), .o(n11567) );
na02f01 g07779 ( .a(n11566), .b(n11565), .o(n11568) );
in01f01 g07780 ( .a(n11568), .o(n11569) );
no02f01 g07781 ( .a(n11569), .b(n11567), .o(n11570) );
no02f01 g07782 ( .a(n11570), .b(n11515), .o(n11571) );
in01f01 g07783 ( .a(n11571), .o(n11572) );
no02f01 g07784 ( .a(n11229), .b(n11218), .o(n11573) );
in01f01 g07785 ( .a(n11573), .o(n11574) );
no02f01 g07786 ( .a(n11574), .b(n11564), .o(n11575) );
no02f01 g07787 ( .a(n11573), .b(n11563), .o(n11576) );
no02f01 g07788 ( .a(n11576), .b(n11575), .o(n11577) );
in01f01 g07789 ( .a(n11577), .o(n11578) );
no02f01 g07790 ( .a(n11578), .b(n11515), .o(n11579) );
in01f01 g07791 ( .a(n11579), .o(n11580) );
no02f01 g07792 ( .a(n11284), .b(n11179), .o(n11581) );
no02f01 g07793 ( .a(n11286), .b(n11267), .o(n11582) );
no02f01 g07794 ( .a(n11582), .b(n11581), .o(n11583) );
no02f01 g07795 ( .a(n11293), .b(n11179), .o(n11584) );
no02f01 g07796 ( .a(n11584), .b(n11295), .o(n11585) );
no02f01 g07797 ( .a(n11585), .b(n11583), .o(n11586) );
na02f01 g07798 ( .a(n11585), .b(n11583), .o(n11587) );
in01f01 g07799 ( .a(n11587), .o(n11588) );
no02f01 g07800 ( .a(n11588), .b(n11586), .o(n11589) );
no02f01 g07801 ( .a(n11589), .b(n11515), .o(n11590) );
in01f01 g07802 ( .a(n11267), .o(n11591) );
no02f01 g07803 ( .a(n11581), .b(n11286), .o(n11592) );
in01f01 g07804 ( .a(n11592), .o(n11593) );
no02f01 g07805 ( .a(n11593), .b(n11591), .o(n11594) );
no02f01 g07806 ( .a(n11592), .b(n11267), .o(n11595) );
no02f01 g07807 ( .a(n11595), .b(n11594), .o(n11596) );
in01f01 g07808 ( .a(n11596), .o(n11597) );
no02f01 g07809 ( .a(n11597), .b(n11515), .o(n11598) );
in01f01 g07810 ( .a(n11598), .o(n11599) );
no02f01 g07811 ( .a(n11244), .b(n11242), .o(n11600) );
in01f01 g07812 ( .a(n11600), .o(n11601) );
no02f01 g07813 ( .a(n11601), .b(n11266), .o(n11602) );
in01f01 g07814 ( .a(n11266), .o(n11603) );
no02f01 g07815 ( .a(n11600), .b(n11603), .o(n11604) );
no02f01 g07816 ( .a(n11604), .b(n11602), .o(n11605) );
no02f01 g07817 ( .a(n11605), .b(n11515), .o(n11606) );
in01f01 g07818 ( .a(n11263), .o(n11607) );
no03f01 g07819 ( .a(n11265), .b(n11607), .c(n11250), .o(n11608) );
ao12f01 g07820 ( .a(n11263), .b(n11264), .c(n11251), .o(n11609) );
no02f01 g07821 ( .a(n11609), .b(n11608), .o(n11610) );
no02f01 g07822 ( .a(n11610), .b(n11515), .o(n11611) );
in01f01 g07823 ( .a(n11258), .o(n11612) );
no03f01 g07824 ( .a(n11262), .b(n11612), .c(n11257), .o(n11613) );
in01f01 g07825 ( .a(n11257), .o(n11614) );
in01f01 g07826 ( .a(n11262), .o(n11615) );
ao12f01 g07827 ( .a(n11615), .b(n11258), .c(n11614), .o(n11616) );
no02f01 g07828 ( .a(n11616), .b(n11613), .o(n11617) );
no02f01 g07829 ( .a(n11617), .b(n11514), .o(n11618) );
na02f01 g07830 ( .a(n11515), .b(n11262), .o(n11619) );
no02f01 g07831 ( .a(n11515), .b(n11262), .o(n11620) );
ao12f01 g07832 ( .a(n11620), .b(n11619), .c(delay_sub_ln23_0_unr1_stage2_stallmux_q_0_), .o(n11621) );
in01f01 g07833 ( .a(n11621), .o(n11622) );
in01f01 g07834 ( .a(n11617), .o(n11623) );
no02f01 g07835 ( .a(n11623), .b(n11515), .o(n11624) );
in01f01 g07836 ( .a(n11624), .o(n11625) );
ao12f01 g07837 ( .a(n11618), .b(n11625), .c(n11622), .o(n11626) );
in01f01 g07838 ( .a(n11626), .o(n11627) );
na02f01 g07839 ( .a(n11610), .b(n11515), .o(n11628) );
ao12f01 g07840 ( .a(n11611), .b(n11628), .c(n11627), .o(n11629) );
in01f01 g07841 ( .a(n11629), .o(n11630) );
na02f01 g07842 ( .a(n11605), .b(n11515), .o(n11631) );
ao12f01 g07843 ( .a(n11606), .b(n11631), .c(n11630), .o(n11632) );
no02f01 g07844 ( .a(n11596), .b(n11514), .o(n11633) );
in01f01 g07845 ( .a(n11633), .o(n11634) );
na02f01 g07846 ( .a(n11634), .b(n11632), .o(n11635) );
na02f01 g07847 ( .a(n11635), .b(n11599), .o(n11636) );
na02f01 g07848 ( .a(n11589), .b(n11515), .o(n11637) );
in01f01 g07849 ( .a(n11637), .o(n11638) );
no02f01 g07850 ( .a(n11638), .b(n11636), .o(n11639) );
no02f01 g07851 ( .a(n11639), .b(n11590), .o(n11640) );
no03f01 g07852 ( .a(n11295), .b(n11286), .c(n11267), .o(n11641) );
no02f01 g07853 ( .a(n11310), .b(n11278), .o(n11642) );
in01f01 g07854 ( .a(n11642), .o(n11643) );
no03f01 g07855 ( .a(n11643), .b(n11641), .c(n11314), .o(n11644) );
no02f01 g07856 ( .a(n11641), .b(n11314), .o(n11645) );
no02f01 g07857 ( .a(n11642), .b(n11645), .o(n11646) );
no02f01 g07858 ( .a(n11646), .b(n11644), .o(n11647) );
no02f01 g07859 ( .a(n11647), .b(n11514), .o(n11648) );
in01f01 g07860 ( .a(n11648), .o(n11649) );
na02f01 g07861 ( .a(n11649), .b(n11640), .o(n11650) );
na02f01 g07862 ( .a(n11647), .b(n11514), .o(n11651) );
no02f01 g07863 ( .a(n11316), .b(n11310), .o(n11652) );
na02f01 g07864 ( .a(n11652), .b(n11299), .o(n11653) );
in01f01 g07865 ( .a(n11653), .o(n11654) );
in01f01 g07866 ( .a(n11313), .o(n11655) );
no02f01 g07867 ( .a(n11655), .b(n11309), .o(n11656) );
no02f01 g07868 ( .a(n11656), .b(n11654), .o(n11657) );
na02f01 g07869 ( .a(n11656), .b(n11654), .o(n11658) );
in01f01 g07870 ( .a(n11658), .o(n11659) );
no02f01 g07871 ( .a(n11659), .b(n11657), .o(n11660) );
in01f01 g07872 ( .a(n11660), .o(n11661) );
no02f01 g07873 ( .a(n11661), .b(n11514), .o(n11662) );
in01f01 g07874 ( .a(n11662), .o(n11663) );
in01f01 g07875 ( .a(n11317), .o(n11664) );
no02f01 g07876 ( .a(n11208), .b(n11179), .o(n11665) );
no02f01 g07877 ( .a(n11319), .b(n11665), .o(n11666) );
in01f01 g07878 ( .a(n11666), .o(n11667) );
no02f01 g07879 ( .a(n11667), .b(n11664), .o(n11668) );
no02f01 g07880 ( .a(n11666), .b(n11317), .o(n11669) );
no02f01 g07881 ( .a(n11669), .b(n11668), .o(n11670) );
in01f01 g07882 ( .a(n11670), .o(n11671) );
no02f01 g07883 ( .a(n11671), .b(n11515), .o(n11672) );
in01f01 g07884 ( .a(n11672), .o(n11673) );
na04f01 g07885 ( .a(n11673), .b(n11663), .c(n11651), .d(n11650), .o(n11674) );
ao12f01 g07886 ( .a(n11670), .b(n11660), .c(n11514), .o(n11675) );
in01f01 g07887 ( .a(n11675), .o(n11676) );
no02f01 g07888 ( .a(n11203), .b(n11158), .o(n11677) );
no02f01 g07889 ( .a(n11677), .b(n11321), .o(n11678) );
in01f01 g07890 ( .a(n11678), .o(n11679) );
no03f01 g07891 ( .a(n11679), .b(n11562), .c(n11665), .o(n11680) );
no02f01 g07892 ( .a(n11562), .b(n11665), .o(n11681) );
no02f01 g07893 ( .a(n11678), .b(n11681), .o(n11682) );
no02f01 g07894 ( .a(n11682), .b(n11680), .o(n11683) );
in01f01 g07895 ( .a(n11683), .o(n11684) );
no02f01 g07896 ( .a(n11684), .b(n11514), .o(n11685) );
ao12f01 g07897 ( .a(n11685), .b(n11676), .c(n11674), .o(n11686) );
no02f01 g07898 ( .a(n11577), .b(n11514), .o(n11687) );
no02f01 g07899 ( .a(n11683), .b(n11515), .o(n11688) );
no02f01 g07900 ( .a(n11688), .b(n11687), .o(n11689) );
in01f01 g07901 ( .a(n11689), .o(n11690) );
oa12f01 g07902 ( .a(n11580), .b(n11690), .c(n11686), .o(n11691) );
na02f01 g07903 ( .a(n11570), .b(n11515), .o(n11692) );
in01f01 g07904 ( .a(n11692), .o(n11693) );
oa12f01 g07905 ( .a(n11572), .b(n11693), .c(n11691), .o(n11694) );
no02f01 g07906 ( .a(n11557), .b(n11514), .o(n11695) );
oa12f01 g07907 ( .a(n11560), .b(n11695), .c(n11694), .o(n11696) );
in01f01 g07908 ( .a(n11335), .o(n11697) );
na02f01 g07909 ( .a(n11697), .b(n11333), .o(n11698) );
no02f01 g07910 ( .a(n11334), .b(n11192), .o(n11699) );
in01f01 g07911 ( .a(n11699), .o(n11700) );
no02f01 g07912 ( .a(n11700), .b(n11698), .o(n11701) );
na02f01 g07913 ( .a(n11700), .b(n11698), .o(n11702) );
in01f01 g07914 ( .a(n11702), .o(n11703) );
no02f01 g07915 ( .a(n11703), .b(n11701), .o(n11704) );
in01f01 g07916 ( .a(n11704), .o(n11705) );
no02f01 g07917 ( .a(n11705), .b(n11514), .o(n11706) );
no02f01 g07918 ( .a(n11704), .b(n11515), .o(n11707) );
in01f01 g07919 ( .a(n11337), .o(n11708) );
no02f01 g07920 ( .a(n11348), .b(n11346), .o(n11709) );
no02f01 g07921 ( .a(n11709), .b(n11708), .o(n11710) );
na02f01 g07922 ( .a(n11709), .b(n11708), .o(n11711) );
in01f01 g07923 ( .a(n11711), .o(n11712) );
no02f01 g07924 ( .a(n11712), .b(n11710), .o(n11713) );
no02f01 g07925 ( .a(n11713), .b(n11515), .o(n11714) );
no02f01 g07926 ( .a(n11714), .b(n11707), .o(n11715) );
oa12f01 g07927 ( .a(n11715), .b(n11706), .c(n11696), .o(n11716) );
na02f01 g07928 ( .a(n11713), .b(n11515), .o(n11717) );
no02f01 g07929 ( .a(n11376), .b(n11179), .o(n11718) );
no02f01 g07930 ( .a(n11718), .b(n11378), .o(n11719) );
no02f01 g07931 ( .a(n11719), .b(n11539), .o(n11720) );
na02f01 g07932 ( .a(n11719), .b(n11539), .o(n11721) );
in01f01 g07933 ( .a(n11721), .o(n11722) );
no02f01 g07934 ( .a(n11722), .b(n11720), .o(n11723) );
in01f01 g07935 ( .a(n11723), .o(n11724) );
no02f01 g07936 ( .a(n11724), .b(n11514), .o(n11725) );
oa12f01 g07937 ( .a(n11347), .b(n11348), .c(n11337), .o(n11726) );
in01f01 g07938 ( .a(n11726), .o(n11727) );
no02f01 g07939 ( .a(n11361), .b(n11356), .o(n11728) );
in01f01 g07940 ( .a(n11728), .o(n11729) );
no02f01 g07941 ( .a(n11729), .b(n11727), .o(n11730) );
no02f01 g07942 ( .a(n11728), .b(n11726), .o(n11731) );
no02f01 g07943 ( .a(n11731), .b(n11730), .o(n11732) );
in01f01 g07944 ( .a(n11732), .o(n11733) );
no02f01 g07945 ( .a(n11733), .b(n11514), .o(n11734) );
no02f01 g07946 ( .a(n11734), .b(n11725), .o(n11735) );
in01f01 g07947 ( .a(n11378), .o(n11736) );
ao12f01 g07948 ( .a(n11718), .b(n11736), .c(n11538), .o(n11737) );
in01f01 g07949 ( .a(n11737), .o(n11738) );
no02f01 g07950 ( .a(n11444), .b(n11179), .o(n11739) );
no02f01 g07951 ( .a(n11739), .b(n11370), .o(n11740) );
in01f01 g07952 ( .a(n11740), .o(n11741) );
no02f01 g07953 ( .a(n11741), .b(n11738), .o(n11742) );
no02f01 g07954 ( .a(n11740), .b(n11737), .o(n11743) );
no02f01 g07955 ( .a(n11743), .b(n11742), .o(n11744) );
in01f01 g07956 ( .a(n11744), .o(n11745) );
no02f01 g07957 ( .a(n11745), .b(n11514), .o(n11746) );
ao12f01 g07958 ( .a(n11445), .b(n11379), .c(n11538), .o(n11747) );
no02f01 g07959 ( .a(n11446), .b(n11179), .o(n11748) );
no02f01 g07960 ( .a(n11748), .b(n11387), .o(n11749) );
no02f01 g07961 ( .a(n11749), .b(n11747), .o(n11750) );
na02f01 g07962 ( .a(n11749), .b(n11747), .o(n11751) );
in01f01 g07963 ( .a(n11751), .o(n11752) );
no02f01 g07964 ( .a(n11752), .b(n11750), .o(n11753) );
in01f01 g07965 ( .a(n11753), .o(n11754) );
no02f01 g07966 ( .a(n11754), .b(n11514), .o(n11755) );
no02f01 g07967 ( .a(n11755), .b(n11746), .o(n11756) );
na04f01 g07968 ( .a(n11756), .b(n11735), .c(n11717), .d(n11716), .o(n11757) );
no02f01 g07969 ( .a(n11732), .b(n11515), .o(n11758) );
no02f01 g07970 ( .a(n11723), .b(n11515), .o(n11759) );
no02f01 g07971 ( .a(n11759), .b(n11758), .o(n11760) );
in01f01 g07972 ( .a(n11760), .o(n11761) );
no02f01 g07973 ( .a(n11744), .b(n11515), .o(n11762) );
no02f01 g07974 ( .a(n11753), .b(n11515), .o(n11763) );
no03f01 g07975 ( .a(n11763), .b(n11762), .c(n11761), .o(n11764) );
na02f01 g07976 ( .a(n11764), .b(n11757), .o(n11765) );
no03f01 g07977 ( .a(n11387), .b(n11380), .c(n11539), .o(n11766) );
no03f01 g07978 ( .a(n11766), .b(n11748), .c(n11445), .o(n11767) );
no02f01 g07979 ( .a(n11447), .b(n11179), .o(n11768) );
no02f01 g07980 ( .a(n11768), .b(n11396), .o(n11769) );
no02f01 g07981 ( .a(n11769), .b(n11767), .o(n11770) );
na02f01 g07982 ( .a(n11769), .b(n11767), .o(n11771) );
in01f01 g07983 ( .a(n11771), .o(n11772) );
no02f01 g07984 ( .a(n11772), .b(n11770), .o(n11773) );
in01f01 g07985 ( .a(n11773), .o(n11774) );
no02f01 g07986 ( .a(n11774), .b(n11514), .o(n11775) );
in01f01 g07987 ( .a(n11775), .o(n11776) );
no02f01 g07988 ( .a(n11442), .b(n11179), .o(n11777) );
no02f01 g07989 ( .a(n11777), .b(n11416), .o(n11778) );
in01f01 g07990 ( .a(n11778), .o(n11779) );
no03f01 g07991 ( .a(n11779), .b(n11450), .c(n11540), .o(n11780) );
no02f01 g07992 ( .a(n11450), .b(n11540), .o(n11781) );
no02f01 g07993 ( .a(n11778), .b(n11781), .o(n11782) );
no02f01 g07994 ( .a(n11782), .b(n11780), .o(n11783) );
in01f01 g07995 ( .a(n11783), .o(n11784) );
no02f01 g07996 ( .a(n11784), .b(n11514), .o(n11785) );
in01f01 g07997 ( .a(n11785), .o(n11786) );
no03f01 g07998 ( .a(n11416), .b(n11398), .c(n11539), .o(n11787) );
no03f01 g07999 ( .a(n11787), .b(n11450), .c(n11777), .o(n11788) );
no02f01 g08000 ( .a(n11441), .b(n11179), .o(n11789) );
no02f01 g08001 ( .a(n11789), .b(n11411), .o(n11790) );
no02f01 g08002 ( .a(n11790), .b(n11788), .o(n11791) );
na02f01 g08003 ( .a(n11790), .b(n11788), .o(n11792) );
in01f01 g08004 ( .a(n11792), .o(n11793) );
no03f01 g08005 ( .a(n11793), .b(n11791), .c(n11514), .o(n11794) );
no02f01 g08006 ( .a(n11536), .b(n11425), .o(n11795) );
no02f01 g08007 ( .a(n11795), .b(n11542), .o(n11796) );
na02f01 g08008 ( .a(n11795), .b(n11542), .o(n11797) );
in01f01 g08009 ( .a(n11797), .o(n11798) );
no03f01 g08010 ( .a(n11798), .b(n11796), .c(n11514), .o(n11799) );
no02f01 g08011 ( .a(n11799), .b(n11794), .o(n11800) );
na04f01 g08012 ( .a(n11800), .b(n11786), .c(n11776), .d(n11765), .o(n11801) );
no02f01 g08013 ( .a(n11773), .b(n11515), .o(n11802) );
no02f01 g08014 ( .a(n11783), .b(n11515), .o(n11803) );
no02f01 g08015 ( .a(n11803), .b(n11802), .o(n11804) );
no02f01 g08016 ( .a(n11804), .b(n11794), .o(n11805) );
in01f01 g08017 ( .a(n11796), .o(n11806) );
ao12f01 g08018 ( .a(n11515), .b(n11797), .c(n11806), .o(n11807) );
in01f01 g08019 ( .a(n11791), .o(n11808) );
ao12f01 g08020 ( .a(n11515), .b(n11792), .c(n11808), .o(n11809) );
no03f01 g08021 ( .a(n11809), .b(n11807), .c(n11805), .o(n11810) );
no02f01 g08022 ( .a(n11810), .b(n11799), .o(n11811) );
in01f01 g08023 ( .a(n11811), .o(n11812) );
na02f01 g08024 ( .a(n11550), .b(n11515), .o(n11813) );
in01f01 g08025 ( .a(n11813), .o(n11814) );
ao12f01 g08026 ( .a(n11814), .b(n11812), .c(n11801), .o(n11815) );
no02f01 g08027 ( .a(n11533), .b(n11514), .o(n11816) );
no03f01 g08028 ( .a(n11816), .b(n11815), .c(n11551), .o(n11817) );
in01f01 g08029 ( .a(n11476), .o(n11818) );
na02f01 g08030 ( .a(n11818), .b(n11437), .o(n11819) );
no02f01 g08031 ( .a(n11527), .b(n11454), .o(n11820) );
na02f01 g08032 ( .a(n11820), .b(n11819), .o(n11821) );
in01f01 g08033 ( .a(n11821), .o(n11822) );
no02f01 g08034 ( .a(n11499), .b(n11158), .o(n11823) );
no02f01 g08035 ( .a(n11823), .b(n11469), .o(n11824) );
no02f01 g08036 ( .a(n11824), .b(n11822), .o(n11825) );
na02f01 g08037 ( .a(n11824), .b(n11822), .o(n11826) );
in01f01 g08038 ( .a(n11826), .o(n11827) );
no03f01 g08039 ( .a(n11827), .b(n11825), .c(n11515), .o(n11828) );
in01f01 g08040 ( .a(n11478), .o(n11829) );
no02f01 g08041 ( .a(n11500), .b(n11829), .o(n11830) );
in01f01 g08042 ( .a(n11830), .o(n11831) );
no02f01 g08043 ( .a(n11506), .b(n11497), .o(n11832) );
in01f01 g08044 ( .a(n11832), .o(n11833) );
no02f01 g08045 ( .a(n11833), .b(n11831), .o(n11834) );
no02f01 g08046 ( .a(n11832), .b(n11830), .o(n11835) );
no03f01 g08047 ( .a(n11835), .b(n11834), .c(n11515), .o(n11836) );
no02f01 g08048 ( .a(n11836), .b(n11828), .o(n11837) );
in01f01 g08049 ( .a(n11837), .o(n11838) );
no03f01 g08050 ( .a(n11838), .b(n11817), .c(n11535), .o(n11839) );
in01f01 g08051 ( .a(n11825), .o(n11840) );
ao12f01 g08052 ( .a(n11514), .b(n11826), .c(n11840), .o(n11841) );
no02f01 g08053 ( .a(n11835), .b(n11834), .o(n11842) );
no02f01 g08054 ( .a(n11842), .b(n11514), .o(n11843) );
no02f01 g08055 ( .a(n11843), .b(n11841), .o(n11844) );
in01f01 g08056 ( .a(n11844), .o(n11845) );
oa12f01 g08057 ( .a(n11505), .b(n11831), .c(n11497), .o(n11846) );
no02f01 g08058 ( .a(n11489), .b(n11158), .o(n11847) );
no02f01 g08059 ( .a(n11847), .b(n11504), .o(n11848) );
no02f01 g08060 ( .a(n11848), .b(n11846), .o(n11849) );
na02f01 g08061 ( .a(n11848), .b(n11846), .o(n11850) );
in01f01 g08062 ( .a(n11850), .o(n11851) );
no02f01 g08063 ( .a(n11851), .b(n11849), .o(n11852) );
in01f01 g08064 ( .a(n11852), .o(n11853) );
no02f01 g08065 ( .a(n11853), .b(n11515), .o(n11854) );
no02f01 g08066 ( .a(n11512), .b(n11175), .o(n11855) );
no02f01 g08067 ( .a(n11855), .b(n11516), .o(n11856) );
na02f01 g08068 ( .a(n11855), .b(n11516), .o(n11857) );
in01f01 g08069 ( .a(n11857), .o(n11858) );
no03f01 g08070 ( .a(n11858), .b(n11856), .c(n11515), .o(n11859) );
no02f01 g08071 ( .a(n11859), .b(n11854), .o(n11860) );
oa12f01 g08072 ( .a(n11860), .b(n11845), .c(n11839), .o(n11861) );
no02f01 g08073 ( .a(n11852), .b(n11514), .o(n11862) );
in01f01 g08074 ( .a(n11856), .o(n11863) );
ao12f01 g08075 ( .a(n11514), .b(n11857), .c(n11863), .o(n11864) );
no02f01 g08076 ( .a(n11864), .b(n11862), .o(n11865) );
in01f01 g08077 ( .a(n11865), .o(n11866) );
no02f01 g08078 ( .a(n11524), .b(n11514), .o(n11867) );
no02f01 g08079 ( .a(n11867), .b(n11866), .o(n11868) );
ao12f01 g08080 ( .a(n11526), .b(n11868), .c(n11861), .o(n4116) );
in01f01 g08081 ( .a(delay_add_ln22_unr2_stage2_stallmux_q_23_), .o(n11870) );
no02f01 g08082 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_4_), .b(n11021), .o(n11871) );
no02f01 g08083 ( .a(n11021), .b(delay_xor_ln22_unr3_stage2_stallmux_q_3_), .o(n11872) );
in01f01 g08084 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_0_), .o(n11873) );
na02f01 g08085 ( .a(n11873), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(n11874) );
in01f01 g08086 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_1_), .o(n11875) );
na02f01 g08087 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(n11875), .o(n11876) );
in01f01 g08088 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_2_), .o(n11877) );
na02f01 g08089 ( .a(n11877), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(n11878) );
na03f01 g08090 ( .a(n11878), .b(n11876), .c(n11874), .o(n11879) );
no03f01 g08091 ( .a(n11879), .b(n11872), .c(n11871), .o(n11880) );
in01f01 g08092 ( .a(n11880), .o(n11881) );
no02f01 g08093 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_5_), .b(n11021), .o(n11882) );
no02f01 g08094 ( .a(n11882), .b(n11881), .o(n11883) );
no02f01 g08095 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_6_), .b(n11021), .o(n11884) );
no02f01 g08096 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_8_), .b(n11021), .o(n11885) );
no02f01 g08097 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_7_), .b(n11021), .o(n11886) );
no03f01 g08098 ( .a(n11886), .b(n11885), .c(n11884), .o(n11887) );
na02f01 g08099 ( .a(n11887), .b(n11883), .o(n11888) );
no02f01 g08100 ( .a(n11021), .b(delay_xor_ln22_unr3_stage2_stallmux_q_9_), .o(n11889) );
no02f01 g08101 ( .a(n11889), .b(n11888), .o(n11890) );
in01f01 g08102 ( .a(n11890), .o(n11891) );
no02f01 g08103 ( .a(n11021), .b(delay_xor_ln22_unr3_stage2_stallmux_q_10_), .o(n11892) );
no02f01 g08104 ( .a(n11892), .b(n11891), .o(n11893) );
in01f01 g08105 ( .a(n11893), .o(n11894) );
no02f01 g08106 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_11_), .b(n11021), .o(n11895) );
no02f01 g08107 ( .a(n11895), .b(n11894), .o(n11896) );
in01f01 g08108 ( .a(n11896), .o(n11897) );
no02f01 g08109 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_12_), .b(n11021), .o(n11898) );
no02f01 g08110 ( .a(n11898), .b(n11897), .o(n11899) );
in01f01 g08111 ( .a(n11899), .o(n11900) );
no02f01 g08112 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_13_), .b(n11021), .o(n11901) );
no02f01 g08113 ( .a(n11901), .b(n11900), .o(n11902) );
in01f01 g08114 ( .a(n11902), .o(n11903) );
no02f01 g08115 ( .a(n11021), .b(delay_xor_ln22_unr3_stage2_stallmux_q_14_), .o(n11904) );
no02f01 g08116 ( .a(n11904), .b(n11903), .o(n11905) );
in01f01 g08117 ( .a(n11905), .o(n11906) );
no02f01 g08118 ( .a(n11021), .b(delay_xor_ln22_unr3_stage2_stallmux_q_15_), .o(n11907) );
no02f01 g08119 ( .a(n11907), .b(n11906), .o(n11908) );
in01f01 g08120 ( .a(n11908), .o(n11909) );
no02f01 g08121 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_16_), .b(n11021), .o(n11910) );
no02f01 g08122 ( .a(n11910), .b(n11909), .o(n11911) );
in01f01 g08123 ( .a(n11911), .o(n11912) );
no02f01 g08124 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_17_), .b(n11021), .o(n11913) );
no02f01 g08125 ( .a(n11913), .b(n11912), .o(n11914) );
in01f01 g08126 ( .a(n11914), .o(n11915) );
no02f01 g08127 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_18_), .b(n11021), .o(n11916) );
no02f01 g08128 ( .a(n11916), .b(n11915), .o(n11917) );
in01f01 g08129 ( .a(n11917), .o(n11918) );
no02f01 g08130 ( .a(n11021), .b(delay_xor_ln22_unr3_stage2_stallmux_q_19_), .o(n11919) );
no02f01 g08131 ( .a(n11919), .b(n11918), .o(n11920) );
in01f01 g08132 ( .a(n11920), .o(n11921) );
no02f01 g08133 ( .a(n11021), .b(delay_xor_ln22_unr3_stage2_stallmux_q_20_), .o(n11922) );
no02f01 g08134 ( .a(n11922), .b(n11921), .o(n11923) );
in01f01 g08135 ( .a(n11923), .o(n11924) );
no02f01 g08136 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_21_), .b(n11021), .o(n11925) );
no02f01 g08137 ( .a(n11925), .b(n11924), .o(n11926) );
in01f01 g08138 ( .a(n11926), .o(n11927) );
no02f01 g08139 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_22_), .b(n11021), .o(n11928) );
no02f01 g08140 ( .a(n11928), .b(n11927), .o(n11929) );
no02f01 g08141 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_23_), .b(n11021), .o(n11930) );
in01f01 g08142 ( .a(n11930), .o(n11931) );
na02f01 g08143 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_23_), .b(n11021), .o(n11932) );
na02f01 g08144 ( .a(n11932), .b(n11931), .o(n11933) );
no02f01 g08145 ( .a(n11933), .b(n11929), .o(n11934) );
na02f01 g08146 ( .a(n11933), .b(n11929), .o(n11935) );
in01f01 g08147 ( .a(n11935), .o(n11936) );
no02f01 g08148 ( .a(n11936), .b(n11934), .o(n11937) );
no02f01 g08149 ( .a(n11937), .b(n11870), .o(n11938) );
na02f01 g08150 ( .a(n11937), .b(n11870), .o(n11939) );
in01f01 g08151 ( .a(n11939), .o(n11940) );
no02f01 g08152 ( .a(n11940), .b(n11938), .o(n11941) );
in01f01 g08153 ( .a(n11941), .o(n11942) );
na02f01 g08154 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_22_), .b(n11021), .o(n11943) );
in01f01 g08155 ( .a(n11943), .o(n11944) );
no02f01 g08156 ( .a(n11944), .b(n11928), .o(n11945) );
in01f01 g08157 ( .a(n11945), .o(n11946) );
no02f01 g08158 ( .a(n11946), .b(n11926), .o(n11947) );
no02f01 g08159 ( .a(n11945), .b(n11927), .o(n11948) );
no02f01 g08160 ( .a(n11948), .b(n11947), .o(n11949) );
in01f01 g08161 ( .a(n11949), .o(n11950) );
no02f01 g08162 ( .a(n11950), .b(delay_add_ln22_unr2_stage2_stallmux_q_22_), .o(n11951) );
in01f01 g08163 ( .a(n11951), .o(n11952) );
in01f01 g08164 ( .a(delay_add_ln22_unr2_stage2_stallmux_q_20_), .o(n11953) );
na02f01 g08165 ( .a(n11021), .b(delay_xor_ln22_unr3_stage2_stallmux_q_20_), .o(n11954) );
in01f01 g08166 ( .a(n11954), .o(n11955) );
no02f01 g08167 ( .a(n11955), .b(n11922), .o(n11956) );
in01f01 g08168 ( .a(n11956), .o(n11957) );
no02f01 g08169 ( .a(n11957), .b(n11920), .o(n11958) );
no02f01 g08170 ( .a(n11956), .b(n11921), .o(n11959) );
no02f01 g08171 ( .a(n11959), .b(n11958), .o(n11960) );
no02f01 g08172 ( .a(n11960), .b(n11953), .o(n11961) );
in01f01 g08173 ( .a(n11961), .o(n11962) );
na02f01 g08174 ( .a(n11021), .b(delay_xor_ln22_unr3_stage2_stallmux_q_19_), .o(n11963) );
in01f01 g08175 ( .a(n11963), .o(n11964) );
no02f01 g08176 ( .a(n11964), .b(n11919), .o(n11965) );
no02f01 g08177 ( .a(n11965), .b(n11918), .o(n11966) );
na02f01 g08178 ( .a(n11965), .b(n11918), .o(n11967) );
in01f01 g08179 ( .a(n11967), .o(n11968) );
no02f01 g08180 ( .a(n11968), .b(n11966), .o(n11969) );
in01f01 g08181 ( .a(n11969), .o(n11970) );
no02f01 g08182 ( .a(n11970), .b(delay_add_ln22_unr2_stage2_stallmux_q_19_), .o(n11971) );
in01f01 g08183 ( .a(delay_add_ln22_unr2_stage2_stallmux_q_17_), .o(n11972) );
na02f01 g08184 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_17_), .b(n11021), .o(n11973) );
in01f01 g08185 ( .a(n11973), .o(n11974) );
no02f01 g08186 ( .a(n11974), .b(n11913), .o(n11975) );
in01f01 g08187 ( .a(n11975), .o(n11976) );
no02f01 g08188 ( .a(n11976), .b(n11911), .o(n11977) );
no02f01 g08189 ( .a(n11975), .b(n11912), .o(n11978) );
no02f01 g08190 ( .a(n11978), .b(n11977), .o(n11979) );
no02f01 g08191 ( .a(n11979), .b(n11972), .o(n11980) );
in01f01 g08192 ( .a(n11980), .o(n11981) );
in01f01 g08193 ( .a(delay_add_ln22_unr2_stage2_stallmux_q_16_), .o(n11982) );
na02f01 g08194 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_16_), .b(n11021), .o(n11983) );
in01f01 g08195 ( .a(n11983), .o(n11984) );
no02f01 g08196 ( .a(n11984), .b(n11910), .o(n11985) );
in01f01 g08197 ( .a(n11985), .o(n11986) );
no02f01 g08198 ( .a(n11986), .b(n11908), .o(n11987) );
no02f01 g08199 ( .a(n11985), .b(n11909), .o(n11988) );
no02f01 g08200 ( .a(n11988), .b(n11987), .o(n11989) );
no02f01 g08201 ( .a(n11989), .b(n11982), .o(n11990) );
in01f01 g08202 ( .a(n11990), .o(n11991) );
in01f01 g08203 ( .a(delay_add_ln22_unr2_stage2_stallmux_q_15_), .o(n11992) );
na02f01 g08204 ( .a(n11021), .b(delay_xor_ln22_unr3_stage2_stallmux_q_15_), .o(n11993) );
in01f01 g08205 ( .a(n11993), .o(n11994) );
no02f01 g08206 ( .a(n11994), .b(n11907), .o(n11995) );
no02f01 g08207 ( .a(n11995), .b(n11906), .o(n11996) );
na02f01 g08208 ( .a(n11995), .b(n11906), .o(n11997) );
in01f01 g08209 ( .a(n11997), .o(n11998) );
no02f01 g08210 ( .a(n11998), .b(n11996), .o(n11999) );
no02f01 g08211 ( .a(n11999), .b(n11992), .o(n12000) );
in01f01 g08212 ( .a(n12000), .o(n12001) );
in01f01 g08213 ( .a(delay_add_ln22_unr2_stage2_stallmux_q_13_), .o(n12002) );
na02f01 g08214 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_13_), .b(n11021), .o(n12003) );
in01f01 g08215 ( .a(n12003), .o(n12004) );
no02f01 g08216 ( .a(n12004), .b(n11901), .o(n12005) );
in01f01 g08217 ( .a(n12005), .o(n12006) );
no02f01 g08218 ( .a(n12006), .b(n11899), .o(n12007) );
no02f01 g08219 ( .a(n12005), .b(n11900), .o(n12008) );
no02f01 g08220 ( .a(n12008), .b(n12007), .o(n12009) );
no02f01 g08221 ( .a(n12009), .b(n12002), .o(n12010) );
in01f01 g08222 ( .a(n12010), .o(n12011) );
na02f01 g08223 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_12_), .b(n11021), .o(n12012) );
in01f01 g08224 ( .a(n12012), .o(n12013) );
no02f01 g08225 ( .a(n12013), .b(n11898), .o(n12014) );
in01f01 g08226 ( .a(n12014), .o(n12015) );
no02f01 g08227 ( .a(n12015), .b(n11896), .o(n12016) );
no02f01 g08228 ( .a(n12014), .b(n11897), .o(n12017) );
no02f01 g08229 ( .a(n12017), .b(n12016), .o(n12018) );
in01f01 g08230 ( .a(n12018), .o(n12019) );
no02f01 g08231 ( .a(n12019), .b(delay_add_ln22_unr2_stage2_stallmux_q_12_), .o(n12020) );
na02f01 g08232 ( .a(n12019), .b(delay_add_ln22_unr2_stage2_stallmux_q_12_), .o(n12021) );
na02f01 g08233 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_11_), .b(n11021), .o(n12022) );
in01f01 g08234 ( .a(n12022), .o(n12023) );
no02f01 g08235 ( .a(n12023), .b(n11895), .o(n12024) );
in01f01 g08236 ( .a(n12024), .o(n12025) );
no02f01 g08237 ( .a(n12025), .b(n11893), .o(n12026) );
no02f01 g08238 ( .a(n12024), .b(n11894), .o(n12027) );
no02f01 g08239 ( .a(n12027), .b(n12026), .o(n12028) );
in01f01 g08240 ( .a(n12028), .o(n12029) );
no02f01 g08241 ( .a(n12029), .b(delay_add_ln22_unr2_stage2_stallmux_q_11_), .o(n12030) );
in01f01 g08242 ( .a(n12030), .o(n12031) );
in01f01 g08243 ( .a(delay_add_ln22_unr2_stage2_stallmux_q_10_), .o(n12032) );
na02f01 g08244 ( .a(n11021), .b(delay_xor_ln22_unr3_stage2_stallmux_q_10_), .o(n12033) );
in01f01 g08245 ( .a(n12033), .o(n12034) );
no02f01 g08246 ( .a(n12034), .b(n11892), .o(n12035) );
in01f01 g08247 ( .a(n12035), .o(n12036) );
no02f01 g08248 ( .a(n12036), .b(n11890), .o(n12037) );
no02f01 g08249 ( .a(n12035), .b(n11891), .o(n12038) );
no02f01 g08250 ( .a(n12038), .b(n12037), .o(n12039) );
no02f01 g08251 ( .a(n12039), .b(n12032), .o(n12040) );
in01f01 g08252 ( .a(n12040), .o(n12041) );
in01f01 g08253 ( .a(delay_add_ln22_unr2_stage2_stallmux_q_9_), .o(n12042) );
na02f01 g08254 ( .a(n11021), .b(delay_xor_ln22_unr3_stage2_stallmux_q_9_), .o(n12043) );
in01f01 g08255 ( .a(n12043), .o(n12044) );
no02f01 g08256 ( .a(n12044), .b(n11889), .o(n12045) );
in01f01 g08257 ( .a(n12045), .o(n12046) );
ao12f01 g08258 ( .a(n12046), .b(n11887), .c(n11883), .o(n12047) );
no02f01 g08259 ( .a(n12045), .b(n11888), .o(n12048) );
no02f01 g08260 ( .a(n12048), .b(n12047), .o(n12049) );
no02f01 g08261 ( .a(n12049), .b(n12042), .o(n12050) );
in01f01 g08262 ( .a(delay_add_ln22_unr2_stage2_stallmux_q_4_), .o(n12051) );
no02f01 g08263 ( .a(n11879), .b(n11872), .o(n12052) );
na02f01 g08264 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_4_), .b(n11021), .o(n12053) );
in01f01 g08265 ( .a(n12053), .o(n12054) );
no02f01 g08266 ( .a(n12054), .b(n11871), .o(n12055) );
in01f01 g08267 ( .a(n12055), .o(n12056) );
na02f01 g08268 ( .a(n12056), .b(n12052), .o(n12057) );
in01f01 g08269 ( .a(n12057), .o(n12058) );
no02f01 g08270 ( .a(n12056), .b(n12052), .o(n12059) );
no02f01 g08271 ( .a(n12059), .b(n12058), .o(n12060) );
no02f01 g08272 ( .a(n12060), .b(n12051), .o(n12061) );
in01f01 g08273 ( .a(n12061), .o(n12062) );
in01f01 g08274 ( .a(delay_add_ln22_unr2_stage2_stallmux_q_3_), .o(n12063) );
in01f01 g08275 ( .a(n11879), .o(n12064) );
na02f01 g08276 ( .a(n11021), .b(delay_xor_ln22_unr3_stage2_stallmux_q_3_), .o(n12065) );
in01f01 g08277 ( .a(n12065), .o(n12066) );
no03f01 g08278 ( .a(n12066), .b(n12064), .c(n11872), .o(n12067) );
in01f01 g08279 ( .a(n11872), .o(n12068) );
ao12f01 g08280 ( .a(n11879), .b(n12065), .c(n12068), .o(n12069) );
no02f01 g08281 ( .a(n12069), .b(n12067), .o(n12070) );
no02f01 g08282 ( .a(n12070), .b(n12063), .o(n12071) );
in01f01 g08283 ( .a(delay_add_ln22_unr2_stage2_stallmux_q_1_), .o(n12072) );
na02f01 g08284 ( .a(n11021), .b(delay_xor_ln22_unr3_stage2_stallmux_q_1_), .o(n12073) );
na02f01 g08285 ( .a(n12073), .b(n11876), .o(n12074) );
no02f01 g08286 ( .a(n12074), .b(n11874), .o(n12075) );
in01f01 g08287 ( .a(n11874), .o(n12076) );
ao12f01 g08288 ( .a(n12076), .b(n12073), .c(n11876), .o(n12077) );
no02f01 g08289 ( .a(n12077), .b(n12075), .o(n12078) );
no02f01 g08290 ( .a(n12078), .b(n12072), .o(n12079) );
na02f01 g08291 ( .a(n11876), .b(n11874), .o(n12080) );
in01f01 g08292 ( .a(n12080), .o(n12081) );
no02f01 g08293 ( .a(n11877), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(n12082) );
in01f01 g08294 ( .a(n12082), .o(n12083) );
na02f01 g08295 ( .a(n12083), .b(n11878), .o(n12084) );
na02f01 g08296 ( .a(n12084), .b(n12081), .o(n12085) );
na03f01 g08297 ( .a(n12083), .b(n12080), .c(n11878), .o(n12086) );
na02f01 g08298 ( .a(n12086), .b(n12085), .o(n12087) );
oa12f01 g08299 ( .a(n12087), .b(n12079), .c(delay_add_ln22_unr2_stage2_stallmux_q_2_), .o(n12088) );
na02f01 g08300 ( .a(n12079), .b(delay_add_ln22_unr2_stage2_stallmux_q_2_), .o(n12089) );
na02f01 g08301 ( .a(n12089), .b(n12088), .o(n12090) );
no03f01 g08302 ( .a(n12069), .b(n12067), .c(delay_add_ln22_unr2_stage2_stallmux_q_3_), .o(n12091) );
in01f01 g08303 ( .a(n12091), .o(n12092) );
ao12f01 g08304 ( .a(n12071), .b(n12092), .c(n12090), .o(n12093) );
no03f01 g08305 ( .a(n12059), .b(n12058), .c(delay_add_ln22_unr2_stage2_stallmux_q_4_), .o(n12094) );
oa12f01 g08306 ( .a(n12062), .b(n12094), .c(n12093), .o(n12095) );
in01f01 g08307 ( .a(delay_add_ln22_unr2_stage2_stallmux_q_5_), .o(n12096) );
na02f01 g08308 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_5_), .b(n11021), .o(n12097) );
in01f01 g08309 ( .a(n12097), .o(n12098) );
no02f01 g08310 ( .a(n12098), .b(n11882), .o(n12099) );
no02f01 g08311 ( .a(n12099), .b(n11881), .o(n12100) );
na02f01 g08312 ( .a(n12099), .b(n11881), .o(n12101) );
in01f01 g08313 ( .a(n12101), .o(n12102) );
no02f01 g08314 ( .a(n12102), .b(n12100), .o(n12103) );
na02f01 g08315 ( .a(n12103), .b(n12096), .o(n12104) );
no02f01 g08316 ( .a(n12103), .b(n12096), .o(n12105) );
ao12f01 g08317 ( .a(n12105), .b(n12104), .c(n12095), .o(n12106) );
in01f01 g08318 ( .a(delay_add_ln22_unr2_stage2_stallmux_q_6_), .o(n12107) );
in01f01 g08319 ( .a(n11884), .o(n12108) );
na02f01 g08320 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_6_), .b(n11021), .o(n12109) );
na02f01 g08321 ( .a(n12109), .b(n12108), .o(n12110) );
no02f01 g08322 ( .a(n12110), .b(n11883), .o(n12111) );
na02f01 g08323 ( .a(n12110), .b(n11883), .o(n12112) );
in01f01 g08324 ( .a(n12112), .o(n12113) );
no02f01 g08325 ( .a(n12113), .b(n12111), .o(n12114) );
na02f01 g08326 ( .a(n12114), .b(n12107), .o(n12115) );
in01f01 g08327 ( .a(n12115), .o(n12116) );
no02f01 g08328 ( .a(n12114), .b(n12107), .o(n12117) );
in01f01 g08329 ( .a(n12117), .o(n12118) );
oa12f01 g08330 ( .a(n12118), .b(n12116), .c(n12106), .o(n12119) );
na02f01 g08331 ( .a(n12108), .b(n11883), .o(n12120) );
in01f01 g08332 ( .a(n11886), .o(n12121) );
na02f01 g08333 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_7_), .b(n11021), .o(n12122) );
na02f01 g08334 ( .a(n12122), .b(n12121), .o(n12123) );
in01f01 g08335 ( .a(n12123), .o(n12124) );
no02f01 g08336 ( .a(n12124), .b(n12120), .o(n12125) );
ao12f01 g08337 ( .a(n12123), .b(n12108), .c(n11883), .o(n12126) );
no02f01 g08338 ( .a(n12126), .b(n12125), .o(n12127) );
in01f01 g08339 ( .a(n12127), .o(n12128) );
no02f01 g08340 ( .a(n12128), .b(delay_add_ln22_unr2_stage2_stallmux_q_7_), .o(n12129) );
in01f01 g08341 ( .a(n12129), .o(n12130) );
na02f01 g08342 ( .a(n12128), .b(delay_add_ln22_unr2_stage2_stallmux_q_7_), .o(n12131) );
in01f01 g08343 ( .a(n12131), .o(n12132) );
ao12f01 g08344 ( .a(n12132), .b(n12130), .c(n12119), .o(n12133) );
in01f01 g08345 ( .a(n12133), .o(n12134) );
no02f01 g08346 ( .a(n12120), .b(n11886), .o(n12135) );
na02f01 g08347 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_8_), .b(n11021), .o(n12136) );
in01f01 g08348 ( .a(n12136), .o(n12137) );
no02f01 g08349 ( .a(n12137), .b(n11885), .o(n12138) );
in01f01 g08350 ( .a(n12138), .o(n12139) );
no02f01 g08351 ( .a(n12139), .b(n12135), .o(n12140) );
na02f01 g08352 ( .a(n12139), .b(n12135), .o(n12141) );
in01f01 g08353 ( .a(n12141), .o(n12142) );
no02f01 g08354 ( .a(n12142), .b(n12140), .o(n12143) );
in01f01 g08355 ( .a(n12143), .o(n12144) );
no02f01 g08356 ( .a(n12144), .b(delay_add_ln22_unr2_stage2_stallmux_q_8_), .o(n12145) );
in01f01 g08357 ( .a(n12145), .o(n12146) );
na02f01 g08358 ( .a(n12144), .b(delay_add_ln22_unr2_stage2_stallmux_q_8_), .o(n12147) );
in01f01 g08359 ( .a(n12147), .o(n12148) );
ao12f01 g08360 ( .a(n12148), .b(n12146), .c(n12134), .o(n12149) );
in01f01 g08361 ( .a(n12149), .o(n12150) );
na02f01 g08362 ( .a(n12049), .b(n12042), .o(n12151) );
ao12f01 g08363 ( .a(n12050), .b(n12151), .c(n12150), .o(n12152) );
na02f01 g08364 ( .a(n12039), .b(n12032), .o(n12153) );
in01f01 g08365 ( .a(n12153), .o(n12154) );
oa12f01 g08366 ( .a(n12041), .b(n12154), .c(n12152), .o(n12155) );
na02f01 g08367 ( .a(n12155), .b(n12031), .o(n12156) );
na02f01 g08368 ( .a(n12029), .b(delay_add_ln22_unr2_stage2_stallmux_q_11_), .o(n12157) );
na02f01 g08369 ( .a(n12157), .b(n12156), .o(n12158) );
in01f01 g08370 ( .a(n12158), .o(n12159) );
ao12f01 g08371 ( .a(n12020), .b(n12159), .c(n12021), .o(n12160) );
na02f01 g08372 ( .a(n12009), .b(n12002), .o(n12161) );
na02f01 g08373 ( .a(n12161), .b(n12160), .o(n12162) );
na02f01 g08374 ( .a(n12162), .b(n12011), .o(n12163) );
na02f01 g08375 ( .a(n11021), .b(delay_xor_ln22_unr3_stage2_stallmux_q_14_), .o(n12164) );
in01f01 g08376 ( .a(n12164), .o(n12165) );
no02f01 g08377 ( .a(n12165), .b(n11904), .o(n12166) );
no02f01 g08378 ( .a(n12166), .b(n11903), .o(n12167) );
na02f01 g08379 ( .a(n12166), .b(n11903), .o(n12168) );
in01f01 g08380 ( .a(n12168), .o(n12169) );
no02f01 g08381 ( .a(n12169), .b(n12167), .o(n12170) );
in01f01 g08382 ( .a(n12170), .o(n12171) );
no02f01 g08383 ( .a(n12171), .b(delay_add_ln22_unr2_stage2_stallmux_q_14_), .o(n12172) );
in01f01 g08384 ( .a(n12172), .o(n12173) );
na02f01 g08385 ( .a(n12173), .b(n12163), .o(n12174) );
na02f01 g08386 ( .a(n12171), .b(delay_add_ln22_unr2_stage2_stallmux_q_14_), .o(n12175) );
na02f01 g08387 ( .a(n12175), .b(n12174), .o(n12176) );
na02f01 g08388 ( .a(n11999), .b(n11992), .o(n12177) );
na02f01 g08389 ( .a(n12177), .b(n12176), .o(n12178) );
na02f01 g08390 ( .a(n12178), .b(n12001), .o(n12179) );
na02f01 g08391 ( .a(n11989), .b(n11982), .o(n12180) );
na02f01 g08392 ( .a(n12180), .b(n12179), .o(n12181) );
na02f01 g08393 ( .a(n12181), .b(n11991), .o(n12182) );
na02f01 g08394 ( .a(n11979), .b(n11972), .o(n12183) );
na02f01 g08395 ( .a(n12183), .b(n12182), .o(n12184) );
na02f01 g08396 ( .a(n12184), .b(n11981), .o(n12185) );
na02f01 g08397 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_18_), .b(n11021), .o(n12186) );
in01f01 g08398 ( .a(n12186), .o(n12187) );
no02f01 g08399 ( .a(n12187), .b(n11916), .o(n12188) );
no02f01 g08400 ( .a(n12188), .b(n11915), .o(n12189) );
na02f01 g08401 ( .a(n12188), .b(n11915), .o(n12190) );
in01f01 g08402 ( .a(n12190), .o(n12191) );
no02f01 g08403 ( .a(n12191), .b(n12189), .o(n12192) );
in01f01 g08404 ( .a(n12192), .o(n12193) );
no02f01 g08405 ( .a(n12193), .b(delay_add_ln22_unr2_stage2_stallmux_q_18_), .o(n12194) );
in01f01 g08406 ( .a(n12194), .o(n12195) );
na02f01 g08407 ( .a(n12195), .b(n12185), .o(n12196) );
na02f01 g08408 ( .a(n12193), .b(delay_add_ln22_unr2_stage2_stallmux_q_18_), .o(n12197) );
na02f01 g08409 ( .a(n12197), .b(n12196), .o(n12198) );
na02f01 g08410 ( .a(n11970), .b(delay_add_ln22_unr2_stage2_stallmux_q_19_), .o(n12199) );
in01f01 g08411 ( .a(n12199), .o(n12200) );
no02f01 g08412 ( .a(n12200), .b(n12198), .o(n12201) );
no02f01 g08413 ( .a(n12201), .b(n11971), .o(n12202) );
na02f01 g08414 ( .a(n11960), .b(n11953), .o(n12203) );
na02f01 g08415 ( .a(n12203), .b(n12202), .o(n12204) );
na02f01 g08416 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_21_), .b(n11021), .o(n12205) );
in01f01 g08417 ( .a(n12205), .o(n12206) );
no02f01 g08418 ( .a(n12206), .b(n11925), .o(n12207) );
in01f01 g08419 ( .a(n12207), .o(n12208) );
no02f01 g08420 ( .a(n12208), .b(n11923), .o(n12209) );
no02f01 g08421 ( .a(n12207), .b(n11924), .o(n12210) );
no02f01 g08422 ( .a(n12210), .b(n12209), .o(n12211) );
in01f01 g08423 ( .a(n12211), .o(n12212) );
no02f01 g08424 ( .a(n12212), .b(delay_add_ln22_unr2_stage2_stallmux_q_21_), .o(n12213) );
ao12f01 g08425 ( .a(n12213), .b(n12204), .c(n11962), .o(n12214) );
na02f01 g08426 ( .a(n12212), .b(delay_add_ln22_unr2_stage2_stallmux_q_21_), .o(n12215) );
in01f01 g08427 ( .a(n12215), .o(n12216) );
no02f01 g08428 ( .a(n12216), .b(n12214), .o(n12217) );
na02f01 g08429 ( .a(n11950), .b(delay_add_ln22_unr2_stage2_stallmux_q_22_), .o(n12218) );
na02f01 g08430 ( .a(n12218), .b(n12217), .o(n12219) );
na03f01 g08431 ( .a(n12219), .b(n11952), .c(n11942), .o(n12220) );
na02f01 g08432 ( .a(n12204), .b(n11962), .o(n12221) );
in01f01 g08433 ( .a(n12213), .o(n12222) );
na02f01 g08434 ( .a(n12222), .b(n12221), .o(n12223) );
na02f01 g08435 ( .a(n12215), .b(n12223), .o(n12224) );
in01f01 g08436 ( .a(n12218), .o(n12225) );
no02f01 g08437 ( .a(n12225), .b(n12224), .o(n12226) );
oa12f01 g08438 ( .a(n11941), .b(n12226), .c(n11951), .o(n12227) );
ao12f01 g08439 ( .a(n11158), .b(n12227), .c(n12220), .o(n12228) );
in01f01 g08440 ( .a(n12203), .o(n12229) );
no02f01 g08441 ( .a(n12229), .b(n11961), .o(n12230) );
in01f01 g08442 ( .a(n12230), .o(n12231) );
na02f01 g08443 ( .a(n12231), .b(n12202), .o(n12232) );
in01f01 g08444 ( .a(n12232), .o(n12233) );
no02f01 g08445 ( .a(n12231), .b(n12202), .o(n12234) );
no02f01 g08446 ( .a(n12234), .b(n12233), .o(n12235) );
no02f01 g08447 ( .a(n12235), .b(n11158), .o(n12236) );
in01f01 g08448 ( .a(n12221), .o(n12237) );
no02f01 g08449 ( .a(n12216), .b(n12213), .o(n12238) );
no02f01 g08450 ( .a(n12238), .b(n12237), .o(n12239) );
in01f01 g08451 ( .a(n12239), .o(n12240) );
na02f01 g08452 ( .a(n12238), .b(n12237), .o(n12241) );
na02f01 g08453 ( .a(n12241), .b(n12240), .o(n12242) );
ao12f01 g08454 ( .a(n12236), .b(n12242), .c(n11179), .o(n12243) );
no02f01 g08455 ( .a(n12225), .b(n11951), .o(n12244) );
no02f01 g08456 ( .a(n12244), .b(n12217), .o(n12245) );
in01f01 g08457 ( .a(n12244), .o(n12246) );
no02f01 g08458 ( .a(n12246), .b(n12224), .o(n12247) );
oa12f01 g08459 ( .a(n11179), .b(n12247), .c(n12245), .o(n12248) );
na02f01 g08460 ( .a(n12248), .b(n12243), .o(n12249) );
na02f01 g08461 ( .a(n12227), .b(n12220), .o(n12250) );
na02f01 g08462 ( .a(n12250), .b(n11158), .o(n12251) );
oa12f01 g08463 ( .a(n12251), .b(n12249), .c(n12228), .o(n12252) );
in01f01 g08464 ( .a(n12241), .o(n12253) );
no02f01 g08465 ( .a(n12253), .b(n12239), .o(n12254) );
in01f01 g08466 ( .a(n12235), .o(n12255) );
no02f01 g08467 ( .a(n12200), .b(n11971), .o(n12256) );
in01f01 g08468 ( .a(n12256), .o(n12257) );
no02f01 g08469 ( .a(n12257), .b(n12198), .o(n12258) );
na02f01 g08470 ( .a(n12257), .b(n12198), .o(n12259) );
in01f01 g08471 ( .a(n12259), .o(n12260) );
no02f01 g08472 ( .a(n12260), .b(n12258), .o(n12261) );
no02f01 g08473 ( .a(n12261), .b(n11179), .o(n12262) );
in01f01 g08474 ( .a(n12183), .o(n12263) );
no02f01 g08475 ( .a(n12263), .b(n11980), .o(n12264) );
in01f01 g08476 ( .a(n12264), .o(n12265) );
no02f01 g08477 ( .a(n12265), .b(n12182), .o(n12266) );
ao12f01 g08478 ( .a(n12264), .b(n12181), .c(n11991), .o(n12267) );
no02f01 g08479 ( .a(n12267), .b(n12266), .o(n12268) );
no02f01 g08480 ( .a(n12268), .b(n11179), .o(n12269) );
in01f01 g08481 ( .a(n12155), .o(n12270) );
na02f01 g08482 ( .a(n12157), .b(n12031), .o(n12271) );
in01f01 g08483 ( .a(n12271), .o(n12272) );
no02f01 g08484 ( .a(n12272), .b(n12270), .o(n12273) );
no02f01 g08485 ( .a(n12271), .b(n12155), .o(n12274) );
no02f01 g08486 ( .a(n12274), .b(n12273), .o(n12275) );
in01f01 g08487 ( .a(n12151), .o(n12276) );
no02f01 g08488 ( .a(n12276), .b(n12050), .o(n12277) );
in01f01 g08489 ( .a(n12277), .o(n12278) );
no02f01 g08490 ( .a(n12278), .b(n12150), .o(n12279) );
no02f01 g08491 ( .a(n12277), .b(n12149), .o(n12280) );
no02f01 g08492 ( .a(n12280), .b(n12279), .o(n12281) );
no02f01 g08493 ( .a(n12132), .b(n12129), .o(n12282) );
in01f01 g08494 ( .a(n12282), .o(n12283) );
no02f01 g08495 ( .a(n12283), .b(n12119), .o(n12284) );
na02f01 g08496 ( .a(n12283), .b(n12119), .o(n12285) );
in01f01 g08497 ( .a(n12285), .o(n12286) );
no02f01 g08498 ( .a(n12286), .b(n12284), .o(n12287) );
no02f01 g08499 ( .a(n12287), .b(n11179), .o(n12288) );
in01f01 g08500 ( .a(n12288), .o(n12289) );
in01f01 g08501 ( .a(n12093), .o(n12290) );
no02f01 g08502 ( .a(n12094), .b(n12061), .o(n12291) );
in01f01 g08503 ( .a(n12291), .o(n12292) );
no02f01 g08504 ( .a(n12292), .b(n12290), .o(n12293) );
no02f01 g08505 ( .a(n12291), .b(n12093), .o(n12294) );
no02f01 g08506 ( .a(n12294), .b(n12293), .o(n12295) );
in01f01 g08507 ( .a(n12295), .o(n12296) );
in01f01 g08508 ( .a(n12104), .o(n12297) );
no02f01 g08509 ( .a(n12105), .b(n12297), .o(n12298) );
in01f01 g08510 ( .a(n12298), .o(n12299) );
no02f01 g08511 ( .a(n12299), .b(n12095), .o(n12300) );
in01f01 g08512 ( .a(n12095), .o(n12301) );
no02f01 g08513 ( .a(n12298), .b(n12301), .o(n12302) );
no02f01 g08514 ( .a(n12302), .b(n12300), .o(n12303) );
in01f01 g08515 ( .a(n12303), .o(n12304) );
oa12f01 g08516 ( .a(n11158), .b(n12304), .c(n12296), .o(n12305) );
in01f01 g08517 ( .a(n12305), .o(n12306) );
no02f01 g08518 ( .a(n12117), .b(n12116), .o(n12307) );
no02f01 g08519 ( .a(n12307), .b(n12106), .o(n12308) );
na02f01 g08520 ( .a(n12307), .b(n12106), .o(n12309) );
in01f01 g08521 ( .a(n12309), .o(n12310) );
no02f01 g08522 ( .a(n12310), .b(n12308), .o(n12311) );
in01f01 g08523 ( .a(n12311), .o(n12312) );
ao12f01 g08524 ( .a(n12306), .b(n12312), .c(n11158), .o(n12313) );
na02f01 g08525 ( .a(n12313), .b(n12289), .o(n12314) );
no02f01 g08526 ( .a(n12148), .b(n12145), .o(n12315) );
in01f01 g08527 ( .a(n12315), .o(n12316) );
no02f01 g08528 ( .a(n12316), .b(n12134), .o(n12317) );
no02f01 g08529 ( .a(n12315), .b(n12133), .o(n12318) );
no02f01 g08530 ( .a(n12318), .b(n12317), .o(n12319) );
no02f01 g08531 ( .a(n12319), .b(n11179), .o(n12320) );
no02f01 g08532 ( .a(n12320), .b(n12314), .o(n12321) );
oa12f01 g08533 ( .a(n12321), .b(n12281), .c(n11179), .o(n12322) );
no02f01 g08534 ( .a(n12154), .b(n12040), .o(n12323) );
no02f01 g08535 ( .a(n12323), .b(n12152), .o(n12324) );
na02f01 g08536 ( .a(n12323), .b(n12152), .o(n12325) );
in01f01 g08537 ( .a(n12325), .o(n12326) );
no02f01 g08538 ( .a(n12326), .b(n12324), .o(n12327) );
no02f01 g08539 ( .a(n12327), .b(n11179), .o(n12328) );
no02f01 g08540 ( .a(n12328), .b(n12322), .o(n12329) );
oa12f01 g08541 ( .a(n12329), .b(n12275), .c(n11179), .o(n12330) );
in01f01 g08542 ( .a(n12021), .o(n12331) );
no02f01 g08543 ( .a(n12331), .b(n12020), .o(n12332) );
in01f01 g08544 ( .a(n12332), .o(n12333) );
no02f01 g08545 ( .a(n12333), .b(n12158), .o(n12334) );
no02f01 g08546 ( .a(n12332), .b(n12159), .o(n12335) );
no02f01 g08547 ( .a(n12335), .b(n12334), .o(n12336) );
in01f01 g08548 ( .a(n12336), .o(n12337) );
ao12f01 g08549 ( .a(n12330), .b(n12337), .c(n11158), .o(n12338) );
na02f01 g08550 ( .a(n12161), .b(n12011), .o(n12339) );
no02f01 g08551 ( .a(n12339), .b(n12160), .o(n12340) );
na02f01 g08552 ( .a(n12339), .b(n12160), .o(n12341) );
in01f01 g08553 ( .a(n12341), .o(n12342) );
no02f01 g08554 ( .a(n12342), .b(n12340), .o(n12343) );
oa12f01 g08555 ( .a(n12338), .b(n12343), .c(n11179), .o(n12344) );
na02f01 g08556 ( .a(n12175), .b(n12173), .o(n12345) );
in01f01 g08557 ( .a(n12345), .o(n12346) );
ao12f01 g08558 ( .a(n12346), .b(n12162), .c(n12011), .o(n12347) );
no02f01 g08559 ( .a(n12345), .b(n12163), .o(n12348) );
no02f01 g08560 ( .a(n12348), .b(n12347), .o(n12349) );
in01f01 g08561 ( .a(n12349), .o(n12350) );
ao12f01 g08562 ( .a(n12344), .b(n12350), .c(n11158), .o(n12351) );
na02f01 g08563 ( .a(n12177), .b(n12001), .o(n12352) );
no02f01 g08564 ( .a(n12352), .b(n12176), .o(n12353) );
na02f01 g08565 ( .a(n12352), .b(n12176), .o(n12354) );
in01f01 g08566 ( .a(n12354), .o(n12355) );
no02f01 g08567 ( .a(n12355), .b(n12353), .o(n12356) );
oa12f01 g08568 ( .a(n12351), .b(n12356), .c(n11179), .o(n12357) );
in01f01 g08569 ( .a(n12356), .o(n12358) );
ao12f01 g08570 ( .a(n11158), .b(n12343), .c(n12336), .o(n12359) );
ao12f01 g08571 ( .a(n12359), .b(n12350), .c(n11179), .o(n12360) );
in01f01 g08572 ( .a(n12360), .o(n12361) );
ao12f01 g08573 ( .a(n12361), .b(n12358), .c(n11179), .o(n12362) );
na02f01 g08574 ( .a(n12362), .b(n12357), .o(n12363) );
na02f01 g08575 ( .a(n12180), .b(n11991), .o(n12364) );
no02f01 g08576 ( .a(n12364), .b(n12179), .o(n12365) );
na02f01 g08577 ( .a(n12364), .b(n12179), .o(n12366) );
in01f01 g08578 ( .a(n12366), .o(n12367) );
no02f01 g08579 ( .a(n12367), .b(n12365), .o(n12368) );
no02f01 g08580 ( .a(n12368), .b(n11179), .o(n12369) );
in01f01 g08581 ( .a(n12369), .o(n12370) );
na02f01 g08582 ( .a(n12370), .b(n12363), .o(n12371) );
no02f01 g08583 ( .a(n12371), .b(n12269), .o(n12372) );
in01f01 g08584 ( .a(n12197), .o(n12373) );
no02f01 g08585 ( .a(n12373), .b(n12194), .o(n12374) );
in01f01 g08586 ( .a(n12374), .o(n12375) );
no02f01 g08587 ( .a(n12375), .b(n12185), .o(n12376) );
na02f01 g08588 ( .a(n12375), .b(n12185), .o(n12377) );
in01f01 g08589 ( .a(n12377), .o(n12378) );
no02f01 g08590 ( .a(n12378), .b(n12376), .o(n12379) );
no02f01 g08591 ( .a(n12379), .b(n11179), .o(n12380) );
in01f01 g08592 ( .a(n12380), .o(n12381) );
na02f01 g08593 ( .a(n12381), .b(n12372), .o(n12382) );
no02f01 g08594 ( .a(n12382), .b(n12262), .o(n12383) );
no02f01 g08595 ( .a(n12261), .b(n11158), .o(n12384) );
in01f01 g08596 ( .a(n12379), .o(n12385) );
na02f01 g08597 ( .a(n12385), .b(n11179), .o(n12386) );
ao12f01 g08598 ( .a(n11158), .b(n12368), .c(n12268), .o(n12387) );
in01f01 g08599 ( .a(n12387), .o(n12388) );
na02f01 g08600 ( .a(n12388), .b(n12386), .o(n12389) );
no03f01 g08601 ( .a(n12389), .b(n12384), .c(n12383), .o(n12390) );
ao12f01 g08602 ( .a(n12390), .b(n12255), .c(n11158), .o(n12391) );
oa12f01 g08603 ( .a(n12391), .b(n12254), .c(n11179), .o(n12392) );
oa12f01 g08604 ( .a(n11158), .b(n12247), .c(n12245), .o(n12393) );
in01f01 g08605 ( .a(n12393), .o(n12394) );
no02f01 g08606 ( .a(n12394), .b(n12392), .o(n12395) );
na02f01 g08607 ( .a(n12395), .b(n12251), .o(n12396) );
na02f01 g08608 ( .a(n12396), .b(n12252), .o(n12397) );
oa12f01 g08609 ( .a(n11952), .b(n12216), .c(n12214), .o(n12398) );
ao12f01 g08610 ( .a(n11940), .b(n12398), .c(n12218), .o(n12399) );
no02f01 g08611 ( .a(n12399), .b(n11938), .o(n12400) );
in01f01 g08612 ( .a(n12400), .o(n12401) );
in01f01 g08613 ( .a(delay_add_ln22_unr2_stage2_stallmux_q_24_), .o(n12402) );
na02f01 g08614 ( .a(n11931), .b(n11929), .o(n12403) );
no02f01 g08615 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_24_), .b(n11021), .o(n12404) );
in01f01 g08616 ( .a(n12404), .o(n12405) );
na02f01 g08617 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_24_), .b(n11021), .o(n12406) );
na02f01 g08618 ( .a(n12406), .b(n12405), .o(n12407) );
in01f01 g08619 ( .a(n12407), .o(n12408) );
no02f01 g08620 ( .a(n12408), .b(n12403), .o(n12409) );
ao12f01 g08621 ( .a(n12407), .b(n11931), .c(n11929), .o(n12410) );
no02f01 g08622 ( .a(n12410), .b(n12409), .o(n12411) );
no02f01 g08623 ( .a(n12411), .b(n12402), .o(n12412) );
na02f01 g08624 ( .a(n12411), .b(n12402), .o(n12413) );
in01f01 g08625 ( .a(n12413), .o(n12414) );
no02f01 g08626 ( .a(n12414), .b(n12412), .o(n12415) );
in01f01 g08627 ( .a(n12415), .o(n12416) );
no02f01 g08628 ( .a(n12416), .b(n12401), .o(n12417) );
no02f01 g08629 ( .a(n12415), .b(n12400), .o(n12418) );
no02f01 g08630 ( .a(n12418), .b(n12417), .o(n12419) );
in01f01 g08631 ( .a(n12419), .o(n12420) );
na02f01 g08632 ( .a(n12420), .b(n12397), .o(n12421) );
na02f01 g08633 ( .a(n12250), .b(n11179), .o(n12422) );
in01f01 g08634 ( .a(n12236), .o(n12423) );
oa12f01 g08635 ( .a(n12423), .b(n12254), .c(n11158), .o(n12424) );
in01f01 g08636 ( .a(n12248), .o(n12425) );
no02f01 g08637 ( .a(n12425), .b(n12424), .o(n12426) );
ao12f01 g08638 ( .a(n11179), .b(n12227), .c(n12220), .o(n12427) );
ao12f01 g08639 ( .a(n12427), .b(n12426), .c(n12422), .o(n12428) );
in01f01 g08640 ( .a(n12395), .o(n12429) );
no02f01 g08641 ( .a(n12429), .b(n12427), .o(n12430) );
no02f01 g08642 ( .a(n12430), .b(n12428), .o(n12431) );
na02f01 g08643 ( .a(n12419), .b(n12431), .o(n12432) );
no02f01 g08644 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_3_), .b(n11021), .o(n12433) );
no02f01 g08645 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_2_), .b(n11021), .o(n12434) );
in01f01 g08646 ( .a(n12434), .o(n12435) );
no02f01 g08647 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_1_), .b(n11021), .o(n12436) );
no02f01 g08648 ( .a(n11021), .b(delay_xor_ln21_unr3_stage2_stallmux_q_0_), .o(n12437) );
no02f01 g08649 ( .a(n12437), .b(n12436), .o(n12438) );
na02f01 g08650 ( .a(n12438), .b(n12435), .o(n12439) );
no02f01 g08651 ( .a(n12439), .b(n12433), .o(n12440) );
no02f01 g08652 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_4_), .b(n11021), .o(n12441) );
in01f01 g08653 ( .a(n12441), .o(n12442) );
na02f01 g08654 ( .a(n12442), .b(n12440), .o(n12443) );
no02f01 g08655 ( .a(n11021), .b(delay_xor_ln21_unr3_stage2_stallmux_q_5_), .o(n12444) );
no02f01 g08656 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_6_), .b(n11021), .o(n12445) );
no03f01 g08657 ( .a(n12445), .b(n12444), .c(n12443), .o(n12446) );
no02f01 g08658 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_7_), .b(n11021), .o(n12447) );
in01f01 g08659 ( .a(n12447), .o(n12448) );
na02f01 g08660 ( .a(n12448), .b(n12446), .o(n12449) );
no02f01 g08661 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_8_), .b(n11021), .o(n12450) );
no02f01 g08662 ( .a(n12450), .b(n12449), .o(n12451) );
in01f01 g08663 ( .a(n12451), .o(n12452) );
no02f01 g08664 ( .a(n11021), .b(delay_xor_ln21_unr3_stage2_stallmux_q_9_), .o(n12453) );
no02f01 g08665 ( .a(n12453), .b(n12452), .o(n12454) );
in01f01 g08666 ( .a(n12454), .o(n12455) );
no02f01 g08667 ( .a(n11021), .b(delay_xor_ln21_unr3_stage2_stallmux_q_10_), .o(n12456) );
no02f01 g08668 ( .a(n12456), .b(n12455), .o(n12457) );
no02f01 g08669 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_11_), .b(n11021), .o(n12458) );
in01f01 g08670 ( .a(n12458), .o(n12459) );
na02f01 g08671 ( .a(n12459), .b(n12457), .o(n12460) );
no02f01 g08672 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_12_), .b(n11021), .o(n12461) );
no02f01 g08673 ( .a(n12461), .b(n12460), .o(n12462) );
in01f01 g08674 ( .a(n12462), .o(n12463) );
no02f01 g08675 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_13_), .b(n11021), .o(n12464) );
no02f01 g08676 ( .a(n12464), .b(n12463), .o(n12465) );
in01f01 g08677 ( .a(n12465), .o(n12466) );
no02f01 g08678 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_14_), .b(n11021), .o(n12467) );
no02f01 g08679 ( .a(n12467), .b(n12466), .o(n12468) );
in01f01 g08680 ( .a(n12468), .o(n12469) );
no02f01 g08681 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_15_), .b(n11021), .o(n12470) );
no02f01 g08682 ( .a(n12470), .b(n12469), .o(n12471) );
in01f01 g08683 ( .a(n12471), .o(n12472) );
no02f01 g08684 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_16_), .b(n11021), .o(n12473) );
no02f01 g08685 ( .a(n12473), .b(n12472), .o(n12474) );
in01f01 g08686 ( .a(n12474), .o(n12475) );
no02f01 g08687 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_17_), .b(n11021), .o(n12476) );
no02f01 g08688 ( .a(n12476), .b(n12475), .o(n12477) );
in01f01 g08689 ( .a(n12477), .o(n12478) );
no02f01 g08690 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_18_), .b(n11021), .o(n12479) );
no02f01 g08691 ( .a(n12479), .b(n12478), .o(n12480) );
no02f01 g08692 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_19_), .b(n11021), .o(n12481) );
in01f01 g08693 ( .a(n12481), .o(n12482) );
na02f01 g08694 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_19_), .b(n11021), .o(n12483) );
na02f01 g08695 ( .a(n12483), .b(n12482), .o(n12484) );
no02f01 g08696 ( .a(n12484), .b(n12480), .o(n12485) );
na02f01 g08697 ( .a(n12484), .b(n12480), .o(n12486) );
in01f01 g08698 ( .a(n12486), .o(n12487) );
no02f01 g08699 ( .a(n12487), .b(n12485), .o(n12488) );
no02f01 g08700 ( .a(n12488), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_19_), .o(n12489) );
in01f01 g08701 ( .a(n12489), .o(n12490) );
in01f01 g08702 ( .a(delay_sub_ln21_0_unr2_stage2_stallmux_q_16_), .o(n12491) );
na02f01 g08703 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_16_), .b(n11021), .o(n12492) );
in01f01 g08704 ( .a(n12492), .o(n12493) );
no02f01 g08705 ( .a(n12493), .b(n12473), .o(n12494) );
in01f01 g08706 ( .a(n12494), .o(n12495) );
no02f01 g08707 ( .a(n12495), .b(n12471), .o(n12496) );
no02f01 g08708 ( .a(n12494), .b(n12472), .o(n12497) );
no03f01 g08709 ( .a(n12497), .b(n12496), .c(n12491), .o(n12498) );
in01f01 g08710 ( .a(delay_sub_ln21_0_unr2_stage2_stallmux_q_15_), .o(n12499) );
na02f01 g08711 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_15_), .b(n11021), .o(n12500) );
in01f01 g08712 ( .a(n12500), .o(n12501) );
no02f01 g08713 ( .a(n12501), .b(n12470), .o(n12502) );
no02f01 g08714 ( .a(n12502), .b(n12469), .o(n12503) );
in01f01 g08715 ( .a(n12503), .o(n12504) );
na02f01 g08716 ( .a(n12502), .b(n12469), .o(n12505) );
na02f01 g08717 ( .a(n12505), .b(n12504), .o(n12506) );
no02f01 g08718 ( .a(n12506), .b(n12499), .o(n12507) );
in01f01 g08719 ( .a(n12507), .o(n12508) );
in01f01 g08720 ( .a(delay_sub_ln21_0_unr2_stage2_stallmux_q_13_), .o(n12509) );
na02f01 g08721 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_13_), .b(n11021), .o(n12510) );
in01f01 g08722 ( .a(n12510), .o(n12511) );
no02f01 g08723 ( .a(n12511), .b(n12464), .o(n12512) );
no02f01 g08724 ( .a(n12512), .b(n12463), .o(n12513) );
na02f01 g08725 ( .a(n12512), .b(n12463), .o(n12514) );
in01f01 g08726 ( .a(n12514), .o(n12515) );
no02f01 g08727 ( .a(n12515), .b(n12513), .o(n12516) );
in01f01 g08728 ( .a(n12516), .o(n12517) );
no02f01 g08729 ( .a(n12517), .b(n12509), .o(n12518) );
in01f01 g08730 ( .a(n12518), .o(n12519) );
na02f01 g08731 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_12_), .b(n11021), .o(n12520) );
in01f01 g08732 ( .a(n12520), .o(n12521) );
no02f01 g08733 ( .a(n12521), .b(n12461), .o(n12522) );
na02f01 g08734 ( .a(n12522), .b(n12460), .o(n12523) );
in01f01 g08735 ( .a(n12523), .o(n12524) );
no02f01 g08736 ( .a(n12522), .b(n12460), .o(n12525) );
no02f01 g08737 ( .a(n12525), .b(n12524), .o(n12526) );
no02f01 g08738 ( .a(n12526), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_12_), .o(n12527) );
in01f01 g08739 ( .a(n12527), .o(n12528) );
in01f01 g08740 ( .a(n12437), .o(n12529) );
in01f01 g08741 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_1_), .o(n12530) );
na02f01 g08742 ( .a(n12530), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(n12531) );
na02f01 g08743 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_1_), .b(n11021), .o(n12532) );
na02f01 g08744 ( .a(n12532), .b(n12531), .o(n12533) );
no02f01 g08745 ( .a(n12533), .b(n12529), .o(n12534) );
ao12f01 g08746 ( .a(n12437), .b(n12532), .c(n12531), .o(n12535) );
no02f01 g08747 ( .a(n12535), .b(n12534), .o(n12536) );
na02f01 g08748 ( .a(n12536), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_1_), .o(n12537) );
no02f01 g08749 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln21_unr3_stage2_stallmux_q_0_), .o(n12538) );
na02f01 g08750 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln21_unr3_stage2_stallmux_q_0_), .o(n12539) );
in01f01 g08751 ( .a(n12539), .o(n12540) );
no02f01 g08752 ( .a(n12540), .b(n12538), .o(n12541) );
in01f01 g08753 ( .a(n12541), .o(n12542) );
no02f01 g08754 ( .a(n12542), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_0_), .o(n12543) );
no02f01 g08755 ( .a(n12536), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_1_), .o(n12544) );
oa12f01 g08756 ( .a(n12537), .b(n12544), .c(n12543), .o(n12545) );
in01f01 g08757 ( .a(delay_sub_ln21_0_unr2_stage2_stallmux_q_2_), .o(n12546) );
na02f01 g08758 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_2_), .b(n11021), .o(n12547) );
na02f01 g08759 ( .a(n12547), .b(n12435), .o(n12548) );
no02f01 g08760 ( .a(n12548), .b(n12438), .o(n12549) );
in01f01 g08761 ( .a(n12549), .o(n12550) );
na02f01 g08762 ( .a(n12548), .b(n12438), .o(n12551) );
na02f01 g08763 ( .a(n12551), .b(n12550), .o(n12552) );
na02f01 g08764 ( .a(n12552), .b(n12546), .o(n12553) );
no02f01 g08765 ( .a(n12552), .b(n12546), .o(n12554) );
ao12f01 g08766 ( .a(n12554), .b(n12553), .c(n12545), .o(n12555) );
in01f01 g08767 ( .a(n12439), .o(n12556) );
na02f01 g08768 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_3_), .b(n11021), .o(n12557) );
in01f01 g08769 ( .a(n12557), .o(n12558) );
no02f01 g08770 ( .a(n12558), .b(n12433), .o(n12559) );
in01f01 g08771 ( .a(n12559), .o(n12560) );
no02f01 g08772 ( .a(n12560), .b(n12556), .o(n12561) );
no02f01 g08773 ( .a(n12559), .b(n12439), .o(n12562) );
no02f01 g08774 ( .a(n12562), .b(n12561), .o(n12563) );
no02f01 g08775 ( .a(n12563), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_3_), .o(n12564) );
na02f01 g08776 ( .a(n12563), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_3_), .o(n12565) );
oa12f01 g08777 ( .a(n12565), .b(n12564), .c(n12555), .o(n12566) );
na02f01 g08778 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_4_), .b(n11021), .o(n12567) );
na02f01 g08779 ( .a(n12567), .b(n12442), .o(n12568) );
no02f01 g08780 ( .a(n12568), .b(n12440), .o(n12569) );
na02f01 g08781 ( .a(n12568), .b(n12440), .o(n12570) );
in01f01 g08782 ( .a(n12570), .o(n12571) );
no02f01 g08783 ( .a(n12571), .b(n12569), .o(n12572) );
no02f01 g08784 ( .a(n12572), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_4_), .o(n12573) );
in01f01 g08785 ( .a(n12573), .o(n12574) );
na02f01 g08786 ( .a(n12572), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_4_), .o(n12575) );
in01f01 g08787 ( .a(n12575), .o(n12576) );
ao12f01 g08788 ( .a(n12576), .b(n12574), .c(n12566), .o(n12577) );
na02f01 g08789 ( .a(n11021), .b(delay_xor_ln21_unr3_stage2_stallmux_q_5_), .o(n12578) );
in01f01 g08790 ( .a(n12578), .o(n12579) );
no02f01 g08791 ( .a(n12579), .b(n12444), .o(n12580) );
no02f01 g08792 ( .a(n12580), .b(n12443), .o(n12581) );
na02f01 g08793 ( .a(n12580), .b(n12443), .o(n12582) );
in01f01 g08794 ( .a(n12582), .o(n12583) );
no02f01 g08795 ( .a(n12583), .b(n12581), .o(n12584) );
no02f01 g08796 ( .a(n12584), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_5_), .o(n12585) );
in01f01 g08797 ( .a(delay_sub_ln21_0_unr2_stage2_stallmux_q_5_), .o(n12586) );
in01f01 g08798 ( .a(n12584), .o(n12587) );
no02f01 g08799 ( .a(n12587), .b(n12586), .o(n12588) );
in01f01 g08800 ( .a(n12588), .o(n12589) );
oa12f01 g08801 ( .a(n12589), .b(n12585), .c(n12577), .o(n12590) );
no02f01 g08802 ( .a(n12444), .b(n12443), .o(n12591) );
na02f01 g08803 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_6_), .b(n11021), .o(n12592) );
in01f01 g08804 ( .a(n12592), .o(n12593) );
no02f01 g08805 ( .a(n12593), .b(n12445), .o(n12594) );
in01f01 g08806 ( .a(n12594), .o(n12595) );
na02f01 g08807 ( .a(n12595), .b(n12591), .o(n12596) );
in01f01 g08808 ( .a(n12596), .o(n12597) );
no02f01 g08809 ( .a(n12595), .b(n12591), .o(n12598) );
no02f01 g08810 ( .a(n12598), .b(n12597), .o(n12599) );
no02f01 g08811 ( .a(n12599), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_6_), .o(n12600) );
in01f01 g08812 ( .a(n12600), .o(n12601) );
na02f01 g08813 ( .a(n12599), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_6_), .o(n12602) );
in01f01 g08814 ( .a(n12602), .o(n12603) );
ao12f01 g08815 ( .a(n12603), .b(n12601), .c(n12590), .o(n12604) );
na02f01 g08816 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_7_), .b(n11021), .o(n12605) );
na02f01 g08817 ( .a(n12605), .b(n12448), .o(n12606) );
na02f01 g08818 ( .a(n12606), .b(n12446), .o(n12607) );
in01f01 g08819 ( .a(n12607), .o(n12608) );
no02f01 g08820 ( .a(n12606), .b(n12446), .o(n12609) );
no02f01 g08821 ( .a(n12609), .b(n12608), .o(n12610) );
no02f01 g08822 ( .a(n12610), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_7_), .o(n12611) );
na02f01 g08823 ( .a(n12610), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_7_), .o(n12612) );
oa12f01 g08824 ( .a(n12612), .b(n12611), .c(n12604), .o(n12613) );
na02f01 g08825 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_8_), .b(n11021), .o(n12614) );
in01f01 g08826 ( .a(n12614), .o(n12615) );
no02f01 g08827 ( .a(n12615), .b(n12450), .o(n12616) );
no02f01 g08828 ( .a(n12616), .b(n12449), .o(n12617) );
na02f01 g08829 ( .a(n12616), .b(n12449), .o(n12618) );
in01f01 g08830 ( .a(n12618), .o(n12619) );
no02f01 g08831 ( .a(n12619), .b(n12617), .o(n12620) );
no02f01 g08832 ( .a(n12620), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_8_), .o(n12621) );
in01f01 g08833 ( .a(n12621), .o(n12622) );
in01f01 g08834 ( .a(delay_sub_ln21_0_unr2_stage2_stallmux_q_8_), .o(n12623) );
in01f01 g08835 ( .a(n12620), .o(n12624) );
no02f01 g08836 ( .a(n12624), .b(n12623), .o(n12625) );
ao12f01 g08837 ( .a(n12625), .b(n12622), .c(n12613), .o(n12626) );
na02f01 g08838 ( .a(n11021), .b(delay_xor_ln21_unr3_stage2_stallmux_q_9_), .o(n12627) );
in01f01 g08839 ( .a(n12627), .o(n12628) );
no02f01 g08840 ( .a(n12628), .b(n12453), .o(n12629) );
in01f01 g08841 ( .a(n12629), .o(n12630) );
no02f01 g08842 ( .a(n12630), .b(n12451), .o(n12631) );
no02f01 g08843 ( .a(n12629), .b(n12452), .o(n12632) );
no02f01 g08844 ( .a(n12632), .b(n12631), .o(n12633) );
no02f01 g08845 ( .a(n12633), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_9_), .o(n12634) );
na02f01 g08846 ( .a(n12633), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_9_), .o(n12635) );
oa12f01 g08847 ( .a(n12635), .b(n12634), .c(n12626), .o(n12636) );
na02f01 g08848 ( .a(n11021), .b(delay_xor_ln21_unr3_stage2_stallmux_q_10_), .o(n12637) );
in01f01 g08849 ( .a(n12637), .o(n12638) );
no02f01 g08850 ( .a(n12638), .b(n12456), .o(n12639) );
in01f01 g08851 ( .a(n12639), .o(n12640) );
no02f01 g08852 ( .a(n12640), .b(n12454), .o(n12641) );
na02f01 g08853 ( .a(n12640), .b(n12454), .o(n12642) );
in01f01 g08854 ( .a(n12642), .o(n12643) );
no02f01 g08855 ( .a(n12643), .b(n12641), .o(n12644) );
no02f01 g08856 ( .a(n12644), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_10_), .o(n12645) );
in01f01 g08857 ( .a(n12645), .o(n12646) );
in01f01 g08858 ( .a(delay_sub_ln21_0_unr2_stage2_stallmux_q_10_), .o(n12647) );
in01f01 g08859 ( .a(n12644), .o(n12648) );
no02f01 g08860 ( .a(n12648), .b(n12647), .o(n12649) );
ao12f01 g08861 ( .a(n12649), .b(n12646), .c(n12636), .o(n12650) );
na02f01 g08862 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_11_), .b(n11021), .o(n12651) );
na02f01 g08863 ( .a(n12651), .b(n12459), .o(n12652) );
in01f01 g08864 ( .a(n12652), .o(n12653) );
no03f01 g08865 ( .a(n12653), .b(n12456), .c(n12455), .o(n12654) );
no02f01 g08866 ( .a(n12652), .b(n12457), .o(n12655) );
no02f01 g08867 ( .a(n12655), .b(n12654), .o(n12656) );
in01f01 g08868 ( .a(n12656), .o(n12657) );
no02f01 g08869 ( .a(n12657), .b(n12650), .o(n12658) );
in01f01 g08870 ( .a(delay_sub_ln21_0_unr2_stage2_stallmux_q_12_), .o(n12659) );
no03f01 g08871 ( .a(n12525), .b(n12524), .c(n12659), .o(n12660) );
oa12f01 g08872 ( .a(n12528), .b(n12660), .c(n12658), .o(n12661) );
no02f01 g08873 ( .a(n12516), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_13_), .o(n12662) );
oa12f01 g08874 ( .a(n12519), .b(n12662), .c(n12661), .o(n12663) );
na02f01 g08875 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_14_), .b(n11021), .o(n12664) );
in01f01 g08876 ( .a(n12664), .o(n12665) );
no02f01 g08877 ( .a(n12665), .b(n12467), .o(n12666) );
in01f01 g08878 ( .a(n12666), .o(n12667) );
no02f01 g08879 ( .a(n12667), .b(n12465), .o(n12668) );
no02f01 g08880 ( .a(n12666), .b(n12466), .o(n12669) );
no02f01 g08881 ( .a(n12669), .b(n12668), .o(n12670) );
na02f01 g08882 ( .a(n12670), .b(n12663), .o(n12671) );
ao12f01 g08883 ( .a(delay_sub_ln21_0_unr2_stage2_stallmux_q_15_), .b(n12505), .c(n12504), .o(n12672) );
oa12f01 g08884 ( .a(n12508), .b(n12672), .c(n12671), .o(n12673) );
no02f01 g08885 ( .a(n12497), .b(n12496), .o(n12674) );
no02f01 g08886 ( .a(n12674), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_16_), .o(n12675) );
in01f01 g08887 ( .a(n12675), .o(n12676) );
ao12f01 g08888 ( .a(n12498), .b(n12676), .c(n12673), .o(n12677) );
na02f01 g08889 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_17_), .b(n11021), .o(n12678) );
in01f01 g08890 ( .a(n12678), .o(n12679) );
no02f01 g08891 ( .a(n12679), .b(n12476), .o(n12680) );
no02f01 g08892 ( .a(n12680), .b(n12475), .o(n12681) );
na02f01 g08893 ( .a(n12680), .b(n12475), .o(n12682) );
in01f01 g08894 ( .a(n12682), .o(n12683) );
no02f01 g08895 ( .a(n12683), .b(n12681), .o(n12684) );
na02f01 g08896 ( .a(n12684), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_17_), .o(n12685) );
no02f01 g08897 ( .a(n12684), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_17_), .o(n12686) );
ao12f01 g08898 ( .a(n12686), .b(n12685), .c(n12677), .o(n12687) );
na02f01 g08899 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_18_), .b(n11021), .o(n12688) );
in01f01 g08900 ( .a(n12688), .o(n12689) );
no02f01 g08901 ( .a(n12689), .b(n12479), .o(n12690) );
no02f01 g08902 ( .a(n12690), .b(n12478), .o(n12691) );
na02f01 g08903 ( .a(n12690), .b(n12478), .o(n12692) );
in01f01 g08904 ( .a(n12692), .o(n12693) );
no02f01 g08905 ( .a(n12693), .b(n12691), .o(n12694) );
no02f01 g08906 ( .a(n12694), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_18_), .o(n12695) );
in01f01 g08907 ( .a(n12695), .o(n12696) );
na02f01 g08908 ( .a(n12694), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_18_), .o(n12697) );
in01f01 g08909 ( .a(n12697), .o(n12698) );
ao12f01 g08910 ( .a(n12698), .b(n12696), .c(n12687), .o(n12699) );
na02f01 g08911 ( .a(n12488), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_19_), .o(n12700) );
na02f01 g08912 ( .a(n12700), .b(n12699), .o(n12701) );
na02f01 g08913 ( .a(n12482), .b(n12480), .o(n12702) );
in01f01 g08914 ( .a(n12702), .o(n12703) );
no02f01 g08915 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_20_), .b(n11021), .o(n12704) );
in01f01 g08916 ( .a(n12704), .o(n12705) );
na02f01 g08917 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_20_), .b(n11021), .o(n12706) );
na02f01 g08918 ( .a(n12706), .b(n12705), .o(n12707) );
no02f01 g08919 ( .a(n12707), .b(n12703), .o(n12708) );
na02f01 g08920 ( .a(n12707), .b(n12703), .o(n12709) );
in01f01 g08921 ( .a(n12709), .o(n12710) );
no02f01 g08922 ( .a(n12710), .b(n12708), .o(n12711) );
no02f01 g08923 ( .a(n12711), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_20_), .o(n12712) );
na02f01 g08924 ( .a(n12711), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_20_), .o(n12713) );
in01f01 g08925 ( .a(n12713), .o(n12714) );
no02f01 g08926 ( .a(n12714), .b(n12712), .o(n12715) );
in01f01 g08927 ( .a(n12715), .o(n12716) );
ao12f01 g08928 ( .a(n12716), .b(n12701), .c(n12490), .o(n12717) );
na02f01 g08929 ( .a(n12701), .b(n12490), .o(n12718) );
no02f01 g08930 ( .a(n12715), .b(n12718), .o(n12719) );
no02f01 g08931 ( .a(n12719), .b(n12717), .o(n12720) );
in01f01 g08932 ( .a(n12720), .o(n12721) );
ao12f01 g08933 ( .a(n12721), .b(n12432), .c(n12421), .o(n12722) );
no02f01 g08934 ( .a(n12419), .b(n12431), .o(n12723) );
no02f01 g08935 ( .a(n12420), .b(n12397), .o(n12724) );
no03f01 g08936 ( .a(n12720), .b(n12724), .c(n12723), .o(n12725) );
no02f01 g08937 ( .a(n12725), .b(n12722), .o(n12726) );
oa22f01 g08938 ( .a(n12395), .b(n12249), .c(n12427), .d(n12228), .o(n12727) );
in01f01 g08939 ( .a(n12727), .o(n12728) );
no04f01 g08940 ( .a(n12395), .b(n12427), .c(n12249), .d(n12228), .o(n12729) );
na02f01 g08941 ( .a(n12700), .b(n12490), .o(n12730) );
in01f01 g08942 ( .a(n12730), .o(n12731) );
no02f01 g08943 ( .a(n12731), .b(n12699), .o(n12732) );
na02f01 g08944 ( .a(n12731), .b(n12699), .o(n12733) );
in01f01 g08945 ( .a(n12733), .o(n12734) );
no02f01 g08946 ( .a(n12734), .b(n12732), .o(n12735) );
no03f01 g08947 ( .a(n12735), .b(n12729), .c(n12728), .o(n12736) );
ao22f01 g08948 ( .a(n12393), .b(n12248), .c(n12392), .d(n12243), .o(n12737) );
na02f01 g08949 ( .a(n12392), .b(n12243), .o(n12738) );
na02f01 g08950 ( .a(n12393), .b(n12248), .o(n12739) );
no02f01 g08951 ( .a(n12739), .b(n12738), .o(n12740) );
no02f01 g08952 ( .a(n12698), .b(n12695), .o(n12741) );
in01f01 g08953 ( .a(n12741), .o(n12742) );
no02f01 g08954 ( .a(n12742), .b(n12687), .o(n12743) );
na02f01 g08955 ( .a(n12742), .b(n12687), .o(n12744) );
in01f01 g08956 ( .a(n12744), .o(n12745) );
no02f01 g08957 ( .a(n12745), .b(n12743), .o(n12746) );
no03f01 g08958 ( .a(n12746), .b(n12740), .c(n12737), .o(n12747) );
in01f01 g08959 ( .a(n12747), .o(n12748) );
oa12f01 g08960 ( .a(n12242), .b(n12391), .c(n12236), .o(n12749) );
no02f01 g08961 ( .a(n12389), .b(n12384), .o(n12750) );
oa12f01 g08962 ( .a(n12750), .b(n12382), .c(n12262), .o(n12751) );
oa12f01 g08963 ( .a(n12751), .b(n12235), .c(n11179), .o(n12752) );
na03f01 g08964 ( .a(n12752), .b(n12254), .c(n12423), .o(n12753) );
in01f01 g08965 ( .a(n12685), .o(n12754) );
no02f01 g08966 ( .a(n12686), .b(n12754), .o(n12755) );
no02f01 g08967 ( .a(n12755), .b(n12677), .o(n12756) );
na02f01 g08968 ( .a(n12755), .b(n12677), .o(n12757) );
in01f01 g08969 ( .a(n12757), .o(n12758) );
no02f01 g08970 ( .a(n12758), .b(n12756), .o(n12759) );
in01f01 g08971 ( .a(n12759), .o(n12760) );
ao12f01 g08972 ( .a(n12760), .b(n12753), .c(n12749), .o(n12761) );
in01f01 g08973 ( .a(n12761), .o(n12762) );
na02f01 g08974 ( .a(n12390), .b(n12235), .o(n12763) );
na02f01 g08975 ( .a(n12751), .b(n12255), .o(n12764) );
in01f01 g08976 ( .a(n12673), .o(n12765) );
no02f01 g08977 ( .a(n12675), .b(n12498), .o(n12766) );
no02f01 g08978 ( .a(n12766), .b(n12765), .o(n12767) );
na02f01 g08979 ( .a(n12766), .b(n12765), .o(n12768) );
in01f01 g08980 ( .a(n12768), .o(n12769) );
no02f01 g08981 ( .a(n12769), .b(n12767), .o(n12770) );
in01f01 g08982 ( .a(n12770), .o(n12771) );
na03f01 g08983 ( .a(n12771), .b(n12764), .c(n12763), .o(n12772) );
in01f01 g08984 ( .a(n12261), .o(n12773) );
no02f01 g08985 ( .a(n12387), .b(n12372), .o(n12774) );
na02f01 g08986 ( .a(n12774), .b(n12386), .o(n12775) );
ao12f01 g08987 ( .a(n12773), .b(n12775), .c(n12381), .o(n12776) );
in01f01 g08988 ( .a(n12776), .o(n12777) );
na03f01 g08989 ( .a(n12775), .b(n12381), .c(n12773), .o(n12778) );
no02f01 g08990 ( .a(n12672), .b(n12507), .o(n12779) );
in01f01 g08991 ( .a(n12779), .o(n12780) );
ao12f01 g08992 ( .a(n12780), .b(n12670), .c(n12663), .o(n12781) );
no02f01 g08993 ( .a(n12779), .b(n12671), .o(n12782) );
no02f01 g08994 ( .a(n12782), .b(n12781), .o(n12783) );
in01f01 g08995 ( .a(n12783), .o(n12784) );
ao12f01 g08996 ( .a(n12784), .b(n12778), .c(n12777), .o(n12785) );
in01f01 g08997 ( .a(n12785), .o(n12786) );
in01f01 g08998 ( .a(n12268), .o(n12787) );
in01f01 g08999 ( .a(n12362), .o(n12788) );
no02f01 g09000 ( .a(n12368), .b(n11158), .o(n12789) );
no02f01 g09001 ( .a(n12369), .b(n12357), .o(n12790) );
no03f01 g09002 ( .a(n12790), .b(n12789), .c(n12788), .o(n12791) );
in01f01 g09003 ( .a(n12791), .o(n12792) );
no02f01 g09004 ( .a(n12792), .b(n12787), .o(n12793) );
no02f01 g09005 ( .a(n12791), .b(n12268), .o(n12794) );
no02f01 g09006 ( .a(n12794), .b(n12793), .o(n12795) );
no02f01 g09007 ( .a(n12662), .b(n12518), .o(n12796) );
no02f01 g09008 ( .a(n12796), .b(n12661), .o(n12797) );
na02f01 g09009 ( .a(n12796), .b(n12661), .o(n12798) );
in01f01 g09010 ( .a(n12798), .o(n12799) );
no02f01 g09011 ( .a(n12799), .b(n12797), .o(n12800) );
in01f01 g09012 ( .a(n12800), .o(n12801) );
no02f01 g09013 ( .a(n12801), .b(n12795), .o(n12802) );
in01f01 g09014 ( .a(n12802), .o(n12803) );
in01f01 g09015 ( .a(n12368), .o(n12804) );
no02f01 g09016 ( .a(n12804), .b(n12363), .o(n12805) );
na02f01 g09017 ( .a(n12804), .b(n12363), .o(n12806) );
in01f01 g09018 ( .a(n12806), .o(n12807) );
no02f01 g09019 ( .a(n12807), .b(n12805), .o(n12808) );
in01f01 g09020 ( .a(n12808), .o(n12809) );
no02f01 g09021 ( .a(n12660), .b(n12527), .o(n12810) );
in01f01 g09022 ( .a(n12810), .o(n12811) );
no02f01 g09023 ( .a(n12811), .b(n12658), .o(n12812) );
no03f01 g09024 ( .a(n12810), .b(n12657), .c(n12650), .o(n12813) );
no02f01 g09025 ( .a(n12813), .b(n12812), .o(n12814) );
no02f01 g09026 ( .a(n12814), .b(n12809), .o(n12815) );
no02f01 g09027 ( .a(n12656), .b(n12650), .o(n12816) );
in01f01 g09028 ( .a(n12650), .o(n12817) );
no02f01 g09029 ( .a(n12657), .b(n12817), .o(n12818) );
no02f01 g09030 ( .a(n12818), .b(n12816), .o(n12819) );
in01f01 g09031 ( .a(n12819), .o(n12820) );
in01f01 g09032 ( .a(n12343), .o(n12821) );
no02f01 g09033 ( .a(n12821), .b(n12338), .o(n12822) );
na02f01 g09034 ( .a(n12821), .b(n12338), .o(n12823) );
in01f01 g09035 ( .a(n12823), .o(n12824) );
no02f01 g09036 ( .a(n12824), .b(n12822), .o(n12825) );
in01f01 g09037 ( .a(n12635), .o(n12826) );
no02f01 g09038 ( .a(n12826), .b(n12634), .o(n12827) );
no02f01 g09039 ( .a(n12827), .b(n12626), .o(n12828) );
na02f01 g09040 ( .a(n12827), .b(n12626), .o(n12829) );
in01f01 g09041 ( .a(n12829), .o(n12830) );
no02f01 g09042 ( .a(n12830), .b(n12828), .o(n12831) );
in01f01 g09043 ( .a(n12831), .o(n12832) );
no02f01 g09044 ( .a(n12832), .b(n12825), .o(n12833) );
no02f01 g09045 ( .a(n12336), .b(n12330), .o(n12834) );
na02f01 g09046 ( .a(n12336), .b(n12330), .o(n12835) );
in01f01 g09047 ( .a(n12835), .o(n12836) );
no02f01 g09048 ( .a(n12836), .b(n12834), .o(n12837) );
in01f01 g09049 ( .a(n12837), .o(n12838) );
in01f01 g09050 ( .a(n12613), .o(n12839) );
no02f01 g09051 ( .a(n12625), .b(n12621), .o(n12840) );
no02f01 g09052 ( .a(n12840), .b(n12839), .o(n12841) );
na02f01 g09053 ( .a(n12840), .b(n12839), .o(n12842) );
in01f01 g09054 ( .a(n12842), .o(n12843) );
no02f01 g09055 ( .a(n12843), .b(n12841), .o(n12844) );
no02f01 g09056 ( .a(n12844), .b(n12838), .o(n12845) );
in01f01 g09057 ( .a(n12604), .o(n12846) );
in01f01 g09058 ( .a(n12612), .o(n12847) );
no02f01 g09059 ( .a(n12847), .b(n12611), .o(n12848) );
in01f01 g09060 ( .a(n12848), .o(n12849) );
no02f01 g09061 ( .a(n12849), .b(n12846), .o(n12850) );
no02f01 g09062 ( .a(n12848), .b(n12604), .o(n12851) );
no02f01 g09063 ( .a(n12851), .b(n12850), .o(n12852) );
in01f01 g09064 ( .a(n12852), .o(n12853) );
in01f01 g09065 ( .a(n12281), .o(n12854) );
na02f01 g09066 ( .a(n12321), .b(n12854), .o(n12855) );
oa12f01 g09067 ( .a(n12281), .b(n12320), .c(n12314), .o(n12856) );
na02f01 g09068 ( .a(n12856), .b(n12855), .o(n12857) );
in01f01 g09069 ( .a(n12857), .o(n12858) );
in01f01 g09070 ( .a(n12577), .o(n12859) );
no02f01 g09071 ( .a(n12588), .b(n12585), .o(n12860) );
in01f01 g09072 ( .a(n12860), .o(n12861) );
no02f01 g09073 ( .a(n12861), .b(n12859), .o(n12862) );
no02f01 g09074 ( .a(n12860), .b(n12577), .o(n12863) );
no02f01 g09075 ( .a(n12863), .b(n12862), .o(n12864) );
in01f01 g09076 ( .a(n12864), .o(n12865) );
no02f01 g09077 ( .a(n12865), .b(n12858), .o(n12866) );
na02f01 g09078 ( .a(n12319), .b(n12314), .o(n12867) );
in01f01 g09079 ( .a(n12867), .o(n12868) );
no02f01 g09080 ( .a(n12319), .b(n12314), .o(n12869) );
no02f01 g09081 ( .a(n12869), .b(n12868), .o(n12870) );
in01f01 g09082 ( .a(n12566), .o(n12871) );
no02f01 g09083 ( .a(n12576), .b(n12573), .o(n12872) );
no02f01 g09084 ( .a(n12872), .b(n12871), .o(n12873) );
na02f01 g09085 ( .a(n12872), .b(n12871), .o(n12874) );
in01f01 g09086 ( .a(n12874), .o(n12875) );
no02f01 g09087 ( .a(n12875), .b(n12873), .o(n12876) );
in01f01 g09088 ( .a(n12876), .o(n12877) );
no02f01 g09089 ( .a(n12877), .b(n12870), .o(n12878) );
in01f01 g09090 ( .a(n12287), .o(n12879) );
no02f01 g09091 ( .a(n12313), .b(n12879), .o(n12880) );
in01f01 g09092 ( .a(n12880), .o(n12881) );
na02f01 g09093 ( .a(n12313), .b(n12879), .o(n12882) );
na02f01 g09094 ( .a(n12882), .b(n12881), .o(n12883) );
in01f01 g09095 ( .a(n12565), .o(n12884) );
no02f01 g09096 ( .a(n12884), .b(n12564), .o(n12885) );
no02f01 g09097 ( .a(n12885), .b(n12555), .o(n12886) );
na02f01 g09098 ( .a(n12885), .b(n12555), .o(n12887) );
in01f01 g09099 ( .a(n12887), .o(n12888) );
no02f01 g09100 ( .a(n12888), .b(n12886), .o(n12889) );
no02f01 g09101 ( .a(n12889), .b(n12883), .o(n12890) );
na02f01 g09102 ( .a(n12889), .b(n12883), .o(n12891) );
no02f01 g09103 ( .a(n12295), .b(n11179), .o(n12892) );
na02f01 g09104 ( .a(n12303), .b(n12892), .o(n12893) );
oa12f01 g09105 ( .a(n12304), .b(n12295), .c(n11179), .o(n12894) );
na02f01 g09106 ( .a(n12894), .b(n12893), .o(n12895) );
no02f01 g09107 ( .a(n12541), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_0_), .o(n12896) );
in01f01 g09108 ( .a(delay_sub_ln21_0_unr2_stage2_stallmux_q_0_), .o(n12897) );
no02f01 g09109 ( .a(n12542), .b(n12897), .o(n12898) );
no02f01 g09110 ( .a(n12898), .b(n12896), .o(n12899) );
no02f01 g09111 ( .a(n12899), .b(n12295), .o(n12900) );
in01f01 g09112 ( .a(n12537), .o(n12901) );
no02f01 g09113 ( .a(n12544), .b(n12901), .o(n12902) );
no02f01 g09114 ( .a(n12902), .b(n12543), .o(n12903) );
na02f01 g09115 ( .a(n12902), .b(n12543), .o(n12904) );
in01f01 g09116 ( .a(n12904), .o(n12905) );
no02f01 g09117 ( .a(n12905), .b(n12903), .o(n12906) );
ao12f01 g09118 ( .a(n12895), .b(n12906), .c(n12900), .o(n12907) );
no02f01 g09119 ( .a(n12906), .b(n12900), .o(n12908) );
in01f01 g09120 ( .a(n12545), .o(n12909) );
in01f01 g09121 ( .a(n12553), .o(n12910) );
no02f01 g09122 ( .a(n12554), .b(n12910), .o(n12911) );
no02f01 g09123 ( .a(n12911), .b(n12909), .o(n12912) );
na02f01 g09124 ( .a(n12911), .b(n12909), .o(n12913) );
in01f01 g09125 ( .a(n12913), .o(n12914) );
no02f01 g09126 ( .a(n12914), .b(n12912), .o(n12915) );
in01f01 g09127 ( .a(n12915), .o(n12916) );
no03f01 g09128 ( .a(n12916), .b(n12908), .c(n12907), .o(n12917) );
na02f01 g09129 ( .a(n12311), .b(n12306), .o(n12918) );
in01f01 g09130 ( .a(n12918), .o(n12919) );
no02f01 g09131 ( .a(n12311), .b(n12306), .o(n12920) );
no02f01 g09132 ( .a(n12920), .b(n12919), .o(n12921) );
in01f01 g09133 ( .a(n12921), .o(n12922) );
oa12f01 g09134 ( .a(n12916), .b(n12908), .c(n12907), .o(n12923) );
oa12f01 g09135 ( .a(n12923), .b(n12922), .c(n12917), .o(n12924) );
ao12f01 g09136 ( .a(n12890), .b(n12924), .c(n12891), .o(n12925) );
no02f01 g09137 ( .a(n12925), .b(n12878), .o(n12926) );
in01f01 g09138 ( .a(n12870), .o(n12927) );
no02f01 g09139 ( .a(n12876), .b(n12927), .o(n12928) );
no02f01 g09140 ( .a(n12864), .b(n12857), .o(n12929) );
no03f01 g09141 ( .a(n12929), .b(n12928), .c(n12926), .o(n12930) );
no02f01 g09142 ( .a(n12327), .b(n12322), .o(n12931) );
na02f01 g09143 ( .a(n12327), .b(n12322), .o(n12932) );
in01f01 g09144 ( .a(n12932), .o(n12933) );
no02f01 g09145 ( .a(n12933), .b(n12931), .o(n12934) );
in01f01 g09146 ( .a(n12590), .o(n12935) );
no02f01 g09147 ( .a(n12603), .b(n12600), .o(n12936) );
no02f01 g09148 ( .a(n12936), .b(n12935), .o(n12937) );
na02f01 g09149 ( .a(n12936), .b(n12935), .o(n12938) );
in01f01 g09150 ( .a(n12938), .o(n12939) );
no02f01 g09151 ( .a(n12939), .b(n12937), .o(n12940) );
in01f01 g09152 ( .a(n12940), .o(n12941) );
no02f01 g09153 ( .a(n12941), .b(n12934), .o(n12942) );
no03f01 g09154 ( .a(n12942), .b(n12930), .c(n12866), .o(n12943) );
na02f01 g09155 ( .a(n12941), .b(n12934), .o(n12944) );
in01f01 g09156 ( .a(n12944), .o(n12945) );
oa12f01 g09157 ( .a(n12853), .b(n12945), .c(n12943), .o(n12946) );
no03f01 g09158 ( .a(n12328), .b(n12322), .c(n12275), .o(n12947) );
in01f01 g09159 ( .a(n12275), .o(n12948) );
no02f01 g09160 ( .a(n12329), .b(n12948), .o(n12949) );
no02f01 g09161 ( .a(n12949), .b(n12947), .o(n12950) );
na02f01 g09162 ( .a(n12944), .b(n12852), .o(n12951) );
oa12f01 g09163 ( .a(n12950), .b(n12951), .c(n12943), .o(n12952) );
in01f01 g09164 ( .a(n12844), .o(n12953) );
no02f01 g09165 ( .a(n12953), .b(n12837), .o(n12954) );
ao12f01 g09166 ( .a(n12954), .b(n12952), .c(n12946), .o(n12955) );
na02f01 g09167 ( .a(n12832), .b(n12825), .o(n12956) );
in01f01 g09168 ( .a(n12956), .o(n12957) );
no03f01 g09169 ( .a(n12957), .b(n12955), .c(n12845), .o(n12958) );
in01f01 g09170 ( .a(n12359), .o(n12959) );
na02f01 g09171 ( .a(n12959), .b(n12344), .o(n12960) );
no02f01 g09172 ( .a(n12960), .b(n12350), .o(n12961) );
na02f01 g09173 ( .a(n12960), .b(n12350), .o(n12962) );
in01f01 g09174 ( .a(n12962), .o(n12963) );
no02f01 g09175 ( .a(n12963), .b(n12961), .o(n12964) );
in01f01 g09176 ( .a(n12636), .o(n12965) );
no02f01 g09177 ( .a(n12649), .b(n12645), .o(n12966) );
no02f01 g09178 ( .a(n12966), .b(n12965), .o(n12967) );
na02f01 g09179 ( .a(n12966), .b(n12965), .o(n12968) );
in01f01 g09180 ( .a(n12968), .o(n12969) );
no02f01 g09181 ( .a(n12969), .b(n12967), .o(n12970) );
in01f01 g09182 ( .a(n12970), .o(n12971) );
no02f01 g09183 ( .a(n12971), .b(n12964), .o(n12972) );
no03f01 g09184 ( .a(n12972), .b(n12958), .c(n12833), .o(n12973) );
na02f01 g09185 ( .a(n12971), .b(n12964), .o(n12974) );
in01f01 g09186 ( .a(n12974), .o(n12975) );
oa12f01 g09187 ( .a(n12820), .b(n12975), .c(n12973), .o(n12976) );
no02f01 g09188 ( .a(n12361), .b(n12351), .o(n12977) );
no02f01 g09189 ( .a(n12977), .b(n12356), .o(n12978) );
na02f01 g09190 ( .a(n12977), .b(n12356), .o(n12979) );
in01f01 g09191 ( .a(n12979), .o(n12980) );
no02f01 g09192 ( .a(n12980), .b(n12978), .o(n12981) );
na02f01 g09193 ( .a(n12974), .b(n12819), .o(n12982) );
oa12f01 g09194 ( .a(n12981), .b(n12982), .c(n12973), .o(n12983) );
na02f01 g09195 ( .a(n12983), .b(n12976), .o(n12984) );
in01f01 g09196 ( .a(n12814), .o(n12985) );
no02f01 g09197 ( .a(n12985), .b(n12808), .o(n12986) );
in01f01 g09198 ( .a(n12986), .o(n12987) );
ao12f01 g09199 ( .a(n12815), .b(n12987), .c(n12984), .o(n12988) );
na02f01 g09200 ( .a(n12801), .b(n12795), .o(n12989) );
na02f01 g09201 ( .a(n12989), .b(n12988), .o(n12990) );
na02f01 g09202 ( .a(n12774), .b(n12379), .o(n12991) );
oa12f01 g09203 ( .a(n12385), .b(n12387), .c(n12372), .o(n12992) );
na02f01 g09204 ( .a(n12992), .b(n12991), .o(n12993) );
in01f01 g09205 ( .a(n12670), .o(n12994) );
no02f01 g09206 ( .a(n12994), .b(n12663), .o(n12995) );
in01f01 g09207 ( .a(n12663), .o(n12996) );
no02f01 g09208 ( .a(n12670), .b(n12996), .o(n12997) );
no02f01 g09209 ( .a(n12997), .b(n12995), .o(n12998) );
na02f01 g09210 ( .a(n12998), .b(n12993), .o(n12999) );
na03f01 g09211 ( .a(n12999), .b(n12990), .c(n12803), .o(n13000) );
na03f01 g09212 ( .a(n12784), .b(n12778), .c(n12777), .o(n13001) );
in01f01 g09213 ( .a(n12998), .o(n13002) );
na03f01 g09214 ( .a(n13002), .b(n12992), .c(n12991), .o(n13003) );
na02f01 g09215 ( .a(n13003), .b(n13001), .o(n13004) );
in01f01 g09216 ( .a(n13004), .o(n13005) );
na02f01 g09217 ( .a(n13005), .b(n13000), .o(n13006) );
ao12f01 g09218 ( .a(n12771), .b(n12764), .c(n12763), .o(n13007) );
in01f01 g09219 ( .a(n13007), .o(n13008) );
na03f01 g09220 ( .a(n13008), .b(n13006), .c(n12786), .o(n13009) );
na03f01 g09221 ( .a(n12760), .b(n12753), .c(n12749), .o(n13010) );
na03f01 g09222 ( .a(n13010), .b(n13009), .c(n12772), .o(n13011) );
oa12f01 g09223 ( .a(n12746), .b(n12740), .c(n12737), .o(n13012) );
na03f01 g09224 ( .a(n13012), .b(n13011), .c(n12762), .o(n13013) );
in01f01 g09225 ( .a(n12729), .o(n13014) );
in01f01 g09226 ( .a(n12735), .o(n13015) );
ao12f01 g09227 ( .a(n13015), .b(n13014), .c(n12727), .o(n13016) );
ao12f01 g09228 ( .a(n13016), .b(n13013), .c(n12748), .o(n13017) );
no02f01 g09229 ( .a(n13017), .b(n12736), .o(n13018) );
no02f01 g09230 ( .a(n13018), .b(n12726), .o(n13019) );
oa12f01 g09231 ( .a(n12720), .b(n12724), .c(n12723), .o(n13020) );
na03f01 g09232 ( .a(n12721), .b(n12432), .c(n12421), .o(n13021) );
na02f01 g09233 ( .a(n13021), .b(n13020), .o(n13022) );
in01f01 g09234 ( .a(n12736), .o(n13023) );
in01f01 g09235 ( .a(n12772), .o(n13024) );
ao12f01 g09236 ( .a(n12802), .b(n12989), .c(n12988), .o(n13025) );
ao12f01 g09237 ( .a(n13004), .b(n12999), .c(n13025), .o(n13026) );
no03f01 g09238 ( .a(n13007), .b(n13026), .c(n12785), .o(n13027) );
in01f01 g09239 ( .a(n13010), .o(n13028) );
no03f01 g09240 ( .a(n13028), .b(n13027), .c(n13024), .o(n13029) );
in01f01 g09241 ( .a(n12737), .o(n13030) );
na04f01 g09242 ( .a(n12393), .b(n12392), .c(n12248), .d(n12243), .o(n13031) );
in01f01 g09243 ( .a(n12746), .o(n13032) );
ao12f01 g09244 ( .a(n13032), .b(n13031), .c(n13030), .o(n13033) );
no03f01 g09245 ( .a(n13033), .b(n13029), .c(n12761), .o(n13034) );
oa12f01 g09246 ( .a(n12735), .b(n12729), .c(n12728), .o(n13035) );
oa12f01 g09247 ( .a(n13035), .b(n13034), .c(n12747), .o(n13036) );
na02f01 g09248 ( .a(n13036), .b(n13023), .o(n13037) );
no02f01 g09249 ( .a(n13037), .b(n13022), .o(n13038) );
no02f01 g09250 ( .a(n13038), .b(n13019), .o(n13039) );
no02f01 g09251 ( .a(n13039), .b(n11515), .o(n13040) );
no02f01 g09252 ( .a(n12928), .b(n12926), .o(n13041) );
no02f01 g09253 ( .a(n12929), .b(n12866), .o(n13042) );
no02f01 g09254 ( .a(n13042), .b(n13041), .o(n13043) );
na02f01 g09255 ( .a(n13042), .b(n13041), .o(n13044) );
in01f01 g09256 ( .a(n13044), .o(n13045) );
no02f01 g09257 ( .a(n13045), .b(n13043), .o(n13046) );
in01f01 g09258 ( .a(n13046), .o(n13047) );
no02f01 g09259 ( .a(n12930), .b(n12866), .o(n13048) );
no03f01 g09260 ( .a(n12945), .b(n12942), .c(n13048), .o(n13049) );
in01f01 g09261 ( .a(n13048), .o(n13050) );
no02f01 g09262 ( .a(n12945), .b(n12942), .o(n13051) );
no02f01 g09263 ( .a(n13051), .b(n13050), .o(n13052) );
no02f01 g09264 ( .a(n13052), .b(n13049), .o(n13053) );
in01f01 g09265 ( .a(n13053), .o(n13054) );
oa12f01 g09266 ( .a(n11514), .b(n13054), .c(n13047), .o(n13055) );
ao12f01 g09267 ( .a(n12942), .b(n12944), .c(n13050), .o(n13056) );
in01f01 g09268 ( .a(n13056), .o(n13057) );
no02f01 g09269 ( .a(n12950), .b(n12853), .o(n13058) );
no03f01 g09270 ( .a(n12949), .b(n12947), .c(n12852), .o(n13059) );
no02f01 g09271 ( .a(n13059), .b(n13058), .o(n13060) );
no02f01 g09272 ( .a(n13060), .b(n13057), .o(n13061) );
na02f01 g09273 ( .a(n13060), .b(n13057), .o(n13062) );
in01f01 g09274 ( .a(n13062), .o(n13063) );
no02f01 g09275 ( .a(n13063), .b(n13061), .o(n13064) );
in01f01 g09276 ( .a(n13064), .o(n13065) );
na02f01 g09277 ( .a(n13065), .b(n11514), .o(n13066) );
na02f01 g09278 ( .a(n13066), .b(n13055), .o(n13067) );
in01f01 g09279 ( .a(n12946), .o(n13068) );
in01f01 g09280 ( .a(n12952), .o(n13069) );
no04f01 g09281 ( .a(n12954), .b(n13069), .c(n13068), .d(n12845), .o(n13070) );
no02f01 g09282 ( .a(n12954), .b(n12845), .o(n13071) );
ao12f01 g09283 ( .a(n13071), .b(n12952), .c(n12946), .o(n13072) );
no02f01 g09284 ( .a(n13072), .b(n13070), .o(n13073) );
in01f01 g09285 ( .a(n13073), .o(n13074) );
na02f01 g09286 ( .a(n13074), .b(n11514), .o(n13075) );
in01f01 g09287 ( .a(n13075), .o(n13076) );
no02f01 g09288 ( .a(n13073), .b(n11514), .o(n13077) );
no02f01 g09289 ( .a(n13064), .b(n11514), .o(n13078) );
no02f01 g09290 ( .a(n13078), .b(n13077), .o(n13079) );
oa12f01 g09291 ( .a(n13079), .b(n13076), .c(n13067), .o(n13080) );
no04f01 g09292 ( .a(n12957), .b(n12955), .c(n12845), .d(n12833), .o(n13081) );
no02f01 g09293 ( .a(n12955), .b(n12845), .o(n13082) );
no02f01 g09294 ( .a(n12957), .b(n12833), .o(n13083) );
no02f01 g09295 ( .a(n13083), .b(n13082), .o(n13084) );
no02f01 g09296 ( .a(n13084), .b(n13081), .o(n13085) );
no02f01 g09297 ( .a(n13085), .b(n11515), .o(n13086) );
no02f01 g09298 ( .a(n12958), .b(n12833), .o(n13087) );
no03f01 g09299 ( .a(n12975), .b(n12972), .c(n13087), .o(n13088) );
in01f01 g09300 ( .a(n13087), .o(n13089) );
no02f01 g09301 ( .a(n12975), .b(n12972), .o(n13090) );
no02f01 g09302 ( .a(n13090), .b(n13089), .o(n13091) );
no02f01 g09303 ( .a(n13091), .b(n13088), .o(n13092) );
no02f01 g09304 ( .a(n13092), .b(n11515), .o(n13093) );
no02f01 g09305 ( .a(n13093), .b(n13086), .o(n13094) );
na02f01 g09306 ( .a(n13094), .b(n13080), .o(n13095) );
in01f01 g09307 ( .a(n13095), .o(n13096) );
ao12f01 g09308 ( .a(n12972), .b(n12974), .c(n13089), .o(n13097) );
no02f01 g09309 ( .a(n12981), .b(n12820), .o(n13098) );
no03f01 g09310 ( .a(n12980), .b(n12978), .c(n12819), .o(n13099) );
no02f01 g09311 ( .a(n13099), .b(n13098), .o(n13100) );
in01f01 g09312 ( .a(n13100), .o(n13101) );
no02f01 g09313 ( .a(n13101), .b(n13097), .o(n13102) );
na02f01 g09314 ( .a(n13101), .b(n13097), .o(n13103) );
in01f01 g09315 ( .a(n13103), .o(n13104) );
no02f01 g09316 ( .a(n13104), .b(n13102), .o(n13105) );
no02f01 g09317 ( .a(n13105), .b(n11515), .o(n13106) );
in01f01 g09318 ( .a(n13106), .o(n13107) );
no02f01 g09319 ( .a(n13085), .b(n11514), .o(n13108) );
no02f01 g09320 ( .a(n13092), .b(n11514), .o(n13109) );
no02f01 g09321 ( .a(n13109), .b(n13108), .o(n13110) );
no02f01 g09322 ( .a(n13105), .b(n11514), .o(n13111) );
in01f01 g09323 ( .a(n13111), .o(n13112) );
no02f01 g09324 ( .a(n12986), .b(n12815), .o(n13113) );
in01f01 g09325 ( .a(n13113), .o(n13114) );
no02f01 g09326 ( .a(n13114), .b(n12984), .o(n13115) );
in01f01 g09327 ( .a(n13115), .o(n13116) );
na02f01 g09328 ( .a(n13114), .b(n12984), .o(n13117) );
na02f01 g09329 ( .a(n13117), .b(n13116), .o(n13118) );
na02f01 g09330 ( .a(n13118), .b(n11515), .o(n13119) );
na03f01 g09331 ( .a(n13119), .b(n13112), .c(n13110), .o(n13120) );
oa12f01 g09332 ( .a(n13107), .b(n13120), .c(n13096), .o(n13121) );
in01f01 g09333 ( .a(n13118), .o(n13122) );
no02f01 g09334 ( .a(n13122), .b(n11515), .o(n13123) );
no02f01 g09335 ( .a(n13123), .b(n13121), .o(n13124) );
in01f01 g09336 ( .a(n12988), .o(n13125) );
na02f01 g09337 ( .a(n12989), .b(n12803), .o(n13126) );
no02f01 g09338 ( .a(n13126), .b(n13125), .o(n13127) );
na02f01 g09339 ( .a(n13126), .b(n13125), .o(n13128) );
in01f01 g09340 ( .a(n13128), .o(n13129) );
no02f01 g09341 ( .a(n13129), .b(n13127), .o(n13130) );
no02f01 g09342 ( .a(n13130), .b(n11515), .o(n13131) );
in01f01 g09343 ( .a(n13131), .o(n13132) );
in01f01 g09344 ( .a(n12999), .o(n13133) );
in01f01 g09345 ( .a(n13003), .o(n13134) );
no02f01 g09346 ( .a(n13134), .b(n13133), .o(n13135) );
in01f01 g09347 ( .a(n13135), .o(n13136) );
na02f01 g09348 ( .a(n13136), .b(n13025), .o(n13137) );
in01f01 g09349 ( .a(n13025), .o(n13138) );
na02f01 g09350 ( .a(n13135), .b(n13138), .o(n13139) );
na02f01 g09351 ( .a(n13139), .b(n13137), .o(n13140) );
na02f01 g09352 ( .a(n13140), .b(n11514), .o(n13141) );
na03f01 g09353 ( .a(n13141), .b(n13132), .c(n13124), .o(n13142) );
ao12f01 g09354 ( .a(n13133), .b(n13003), .c(n13138), .o(n13143) );
in01f01 g09355 ( .a(n13143), .o(n13144) );
in01f01 g09356 ( .a(n13001), .o(n13145) );
no02f01 g09357 ( .a(n13145), .b(n12785), .o(n13146) );
no02f01 g09358 ( .a(n13146), .b(n13144), .o(n13147) );
in01f01 g09359 ( .a(n13146), .o(n13148) );
no02f01 g09360 ( .a(n13148), .b(n13143), .o(n13149) );
no02f01 g09361 ( .a(n13149), .b(n13147), .o(n13150) );
no02f01 g09362 ( .a(n13150), .b(n11515), .o(n13151) );
no02f01 g09363 ( .a(n13026), .b(n12785), .o(n13152) );
no02f01 g09364 ( .a(n13007), .b(n13024), .o(n13153) );
in01f01 g09365 ( .a(n13153), .o(n13154) );
no02f01 g09366 ( .a(n13154), .b(n13152), .o(n13155) );
na02f01 g09367 ( .a(n13154), .b(n13152), .o(n13156) );
in01f01 g09368 ( .a(n13156), .o(n13157) );
no02f01 g09369 ( .a(n13157), .b(n13155), .o(n13158) );
no02f01 g09370 ( .a(n13158), .b(n11515), .o(n13159) );
no03f01 g09371 ( .a(n13159), .b(n13151), .c(n13142), .o(n13160) );
na02f01 g09372 ( .a(n13140), .b(n11515), .o(n13161) );
no02f01 g09373 ( .a(n13130), .b(n11514), .o(n13162) );
in01f01 g09374 ( .a(n13162), .o(n13163) );
na02f01 g09375 ( .a(n13163), .b(n13161), .o(n13164) );
no02f01 g09376 ( .a(n13150), .b(n11514), .o(n13165) );
no02f01 g09377 ( .a(n13165), .b(n13164), .o(n13166) );
oa12f01 g09378 ( .a(n13166), .b(n13158), .c(n11514), .o(n13167) );
no02f01 g09379 ( .a(n13027), .b(n13024), .o(n13168) );
no02f01 g09380 ( .a(n13028), .b(n12761), .o(n13169) );
no02f01 g09381 ( .a(n13169), .b(n13168), .o(n13170) );
na02f01 g09382 ( .a(n13169), .b(n13168), .o(n13171) );
in01f01 g09383 ( .a(n13171), .o(n13172) );
no02f01 g09384 ( .a(n13172), .b(n13170), .o(n13173) );
in01f01 g09385 ( .a(n13173), .o(n13174) );
na02f01 g09386 ( .a(n13174), .b(n11514), .o(n13175) );
oa12f01 g09387 ( .a(n13175), .b(n13167), .c(n13160), .o(n13176) );
no02f01 g09388 ( .a(n13029), .b(n12761), .o(n13177) );
in01f01 g09389 ( .a(n13177), .o(n13178) );
no02f01 g09390 ( .a(n13033), .b(n12747), .o(n13179) );
na02f01 g09391 ( .a(n13179), .b(n13178), .o(n13180) );
in01f01 g09392 ( .a(n13180), .o(n13181) );
no02f01 g09393 ( .a(n13179), .b(n13178), .o(n13182) );
no02f01 g09394 ( .a(n13182), .b(n13181), .o(n13183) );
no02f01 g09395 ( .a(n13183), .b(n11515), .o(n13184) );
no02f01 g09396 ( .a(n13184), .b(n13176), .o(n13185) );
no02f01 g09397 ( .a(n13034), .b(n12747), .o(n13186) );
no02f01 g09398 ( .a(n13016), .b(n12736), .o(n13187) );
na02f01 g09399 ( .a(n13187), .b(n13186), .o(n13188) );
in01f01 g09400 ( .a(n13186), .o(n13189) );
na02f01 g09401 ( .a(n13035), .b(n13023), .o(n13190) );
na02f01 g09402 ( .a(n13190), .b(n13189), .o(n13191) );
na02f01 g09403 ( .a(n13191), .b(n13188), .o(n13192) );
na02f01 g09404 ( .a(n13192), .b(n11514), .o(n13193) );
na02f01 g09405 ( .a(n13193), .b(n13185), .o(n13194) );
no02f01 g09406 ( .a(n13194), .b(n13040), .o(n13195) );
no02f01 g09407 ( .a(n13190), .b(n13189), .o(n13196) );
no02f01 g09408 ( .a(n13187), .b(n13186), .o(n13197) );
no02f01 g09409 ( .a(n13197), .b(n13196), .o(n13198) );
no02f01 g09410 ( .a(n13198), .b(n11514), .o(n13199) );
in01f01 g09411 ( .a(n13182), .o(n13200) );
na02f01 g09412 ( .a(n13200), .b(n13180), .o(n13201) );
na02f01 g09413 ( .a(n13201), .b(n11515), .o(n13202) );
na02f01 g09414 ( .a(n13174), .b(n11515), .o(n13203) );
na02f01 g09415 ( .a(n13203), .b(n13202), .o(n13204) );
no02f01 g09416 ( .a(n13204), .b(n13199), .o(n13205) );
oa12f01 g09417 ( .a(n13205), .b(n13039), .c(n11514), .o(n13206) );
ao12f01 g09418 ( .a(n12722), .b(n13036), .c(n13023), .o(n13207) );
no02f01 g09419 ( .a(n13207), .b(n12725), .o(n13208) );
no02f01 g09420 ( .a(n12419), .b(n11158), .o(n13209) );
in01f01 g09421 ( .a(n13209), .o(n13210) );
no02f01 g09422 ( .a(n12419), .b(n11179), .o(n13211) );
in01f01 g09423 ( .a(n13211), .o(n13212) );
na02f01 g09424 ( .a(n13212), .b(n12397), .o(n13213) );
no02f01 g09425 ( .a(n12404), .b(n12403), .o(n13214) );
no02f01 g09426 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_25_), .b(n11021), .o(n13215) );
in01f01 g09427 ( .a(n13215), .o(n13216) );
na02f01 g09428 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_25_), .b(n11021), .o(n13217) );
na02f01 g09429 ( .a(n13217), .b(n13216), .o(n13218) );
no02f01 g09430 ( .a(n13218), .b(n13214), .o(n13219) );
na02f01 g09431 ( .a(n13218), .b(n13214), .o(n13220) );
in01f01 g09432 ( .a(n13220), .o(n13221) );
no02f01 g09433 ( .a(n13221), .b(n13219), .o(n13222) );
in01f01 g09434 ( .a(n13222), .o(n13223) );
no02f01 g09435 ( .a(n13223), .b(delay_add_ln22_unr2_stage2_stallmux_q_25_), .o(n13224) );
na02f01 g09436 ( .a(n13223), .b(delay_add_ln22_unr2_stage2_stallmux_q_25_), .o(n13225) );
in01f01 g09437 ( .a(n13225), .o(n13226) );
no02f01 g09438 ( .a(n13226), .b(n13224), .o(n13227) );
in01f01 g09439 ( .a(n13227), .o(n13228) );
in01f01 g09440 ( .a(n12412), .o(n13229) );
oa12f01 g09441 ( .a(n12413), .b(n12399), .c(n11938), .o(n13230) );
na02f01 g09442 ( .a(n13230), .b(n13229), .o(n13231) );
na02f01 g09443 ( .a(n13231), .b(n13228), .o(n13232) );
no02f01 g09444 ( .a(n12414), .b(n12400), .o(n13233) );
no02f01 g09445 ( .a(n13233), .b(n12412), .o(n13234) );
na02f01 g09446 ( .a(n13234), .b(n13227), .o(n13235) );
na02f01 g09447 ( .a(n13235), .b(n13232), .o(n13236) );
na02f01 g09448 ( .a(n13236), .b(n11179), .o(n13237) );
na02f01 g09449 ( .a(n13236), .b(n11158), .o(n13238) );
na04f01 g09450 ( .a(n13238), .b(n13237), .c(n13213), .d(n13210), .o(n13239) );
ao12f01 g09451 ( .a(n13211), .b(n12396), .c(n12252), .o(n13240) );
no02f01 g09452 ( .a(n13234), .b(n13227), .o(n13241) );
no02f01 g09453 ( .a(n13231), .b(n13228), .o(n13242) );
no02f01 g09454 ( .a(n13242), .b(n13241), .o(n13243) );
no02f01 g09455 ( .a(n13243), .b(n11158), .o(n13244) );
no02f01 g09456 ( .a(n13243), .b(n11179), .o(n13245) );
oa22f01 g09457 ( .a(n13245), .b(n13244), .c(n13240), .d(n13209), .o(n13246) );
oa12f01 g09458 ( .a(n12713), .b(n12712), .c(n12718), .o(n13247) );
in01f01 g09459 ( .a(n13247), .o(n13248) );
no02f01 g09460 ( .a(n12704), .b(n12702), .o(n13249) );
in01f01 g09461 ( .a(n13249), .o(n13250) );
no02f01 g09462 ( .a(n11021), .b(delay_xor_ln21_unr3_stage2_stallmux_q_21_), .o(n13251) );
in01f01 g09463 ( .a(n13251), .o(n13252) );
na02f01 g09464 ( .a(n11021), .b(delay_xor_ln21_unr3_stage2_stallmux_q_21_), .o(n13253) );
na02f01 g09465 ( .a(n13253), .b(n13252), .o(n13254) );
in01f01 g09466 ( .a(n13254), .o(n13255) );
no02f01 g09467 ( .a(n13255), .b(n13250), .o(n13256) );
no02f01 g09468 ( .a(n13254), .b(n13249), .o(n13257) );
no02f01 g09469 ( .a(n13257), .b(n13256), .o(n13258) );
no02f01 g09470 ( .a(n13258), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_21_), .o(n13259) );
na02f01 g09471 ( .a(n13258), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_21_), .o(n13260) );
in01f01 g09472 ( .a(n13260), .o(n13261) );
no02f01 g09473 ( .a(n13261), .b(n13259), .o(n13262) );
no02f01 g09474 ( .a(n13262), .b(n13248), .o(n13263) );
na02f01 g09475 ( .a(n13262), .b(n13248), .o(n13264) );
in01f01 g09476 ( .a(n13264), .o(n13265) );
no02f01 g09477 ( .a(n13265), .b(n13263), .o(n13266) );
in01f01 g09478 ( .a(n13266), .o(n13267) );
ao12f01 g09479 ( .a(n13267), .b(n13246), .c(n13239), .o(n13268) );
no04f01 g09480 ( .a(n13245), .b(n13244), .c(n13240), .d(n13209), .o(n13269) );
ao22f01 g09481 ( .a(n13238), .b(n13237), .c(n13213), .d(n13210), .o(n13270) );
no03f01 g09482 ( .a(n13266), .b(n13270), .c(n13269), .o(n13271) );
no02f01 g09483 ( .a(n13271), .b(n13268), .o(n13272) );
na02f01 g09484 ( .a(n13272), .b(n13208), .o(n13273) );
in01f01 g09485 ( .a(n13273), .o(n13274) );
no02f01 g09486 ( .a(n13272), .b(n13208), .o(n13275) );
no02f01 g09487 ( .a(n13275), .b(n13274), .o(n13276) );
oa22f01 g09488 ( .a(n13276), .b(n11515), .c(n13206), .d(n13195), .o(n13277) );
in01f01 g09489 ( .a(n13224), .o(n13278) );
in01f01 g09490 ( .a(delay_add_ln22_unr2_stage2_stallmux_q_26_), .o(n13279) );
na02f01 g09491 ( .a(n13216), .b(n13214), .o(n13280) );
no02f01 g09492 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_26_), .b(n11021), .o(n13281) );
in01f01 g09493 ( .a(n13281), .o(n13282) );
na02f01 g09494 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_26_), .b(n11021), .o(n13283) );
na02f01 g09495 ( .a(n13283), .b(n13282), .o(n13284) );
in01f01 g09496 ( .a(n13284), .o(n13285) );
no02f01 g09497 ( .a(n13285), .b(n13280), .o(n13286) );
ao12f01 g09498 ( .a(n13284), .b(n13216), .c(n13214), .o(n13287) );
no02f01 g09499 ( .a(n13287), .b(n13286), .o(n13288) );
no02f01 g09500 ( .a(n13288), .b(n13279), .o(n13289) );
na02f01 g09501 ( .a(n13288), .b(n13279), .o(n13290) );
in01f01 g09502 ( .a(n13290), .o(n13291) );
no02f01 g09503 ( .a(n13291), .b(n13289), .o(n13292) );
in01f01 g09504 ( .a(n13292), .o(n13293) );
na03f01 g09505 ( .a(n13230), .b(n13225), .c(n13229), .o(n13294) );
ao12f01 g09506 ( .a(n13293), .b(n13294), .c(n13278), .o(n13295) );
in01f01 g09507 ( .a(n13295), .o(n13296) );
na03f01 g09508 ( .a(n13294), .b(n13293), .c(n13278), .o(n13297) );
na02f01 g09509 ( .a(n13297), .b(n13296), .o(n13298) );
na02f01 g09510 ( .a(n13298), .b(n11179), .o(n13299) );
na02f01 g09511 ( .a(n13298), .b(n11158), .o(n13300) );
na02f01 g09512 ( .a(n13300), .b(n13299), .o(n13301) );
ao12f01 g09513 ( .a(n11179), .b(n13243), .c(n12419), .o(n13302) );
ao12f01 g09514 ( .a(n13209), .b(n13236), .c(n11179), .o(n13303) );
oa12f01 g09515 ( .a(n13303), .b(n13302), .c(n12431), .o(n13304) );
na02f01 g09516 ( .a(n13304), .b(n13301), .o(n13305) );
in01f01 g09517 ( .a(n13297), .o(n13306) );
no02f01 g09518 ( .a(n13306), .b(n13295), .o(n13307) );
no02f01 g09519 ( .a(n13307), .b(n11158), .o(n13308) );
no02f01 g09520 ( .a(n13307), .b(n11179), .o(n13309) );
no02f01 g09521 ( .a(n13309), .b(n13308), .o(n13310) );
ao12f01 g09522 ( .a(n13211), .b(n13236), .c(n11158), .o(n13311) );
ao12f01 g09523 ( .a(n11158), .b(n13243), .c(n12419), .o(n13312) );
ao12f01 g09524 ( .a(n13312), .b(n13311), .c(n12397), .o(n13313) );
na02f01 g09525 ( .a(n13313), .b(n13310), .o(n13314) );
oa12f01 g09526 ( .a(n13260), .b(n13259), .c(n13248), .o(n13315) );
in01f01 g09527 ( .a(n13315), .o(n13316) );
in01f01 g09528 ( .a(delay_sub_ln21_0_unr2_stage2_stallmux_q_22_), .o(n13317) );
no02f01 g09529 ( .a(n13251), .b(n13250), .o(n13318) );
in01f01 g09530 ( .a(n13318), .o(n13319) );
no02f01 g09531 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_22_), .b(n11021), .o(n13320) );
in01f01 g09532 ( .a(n13320), .o(n13321) );
na02f01 g09533 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_22_), .b(n11021), .o(n13322) );
na02f01 g09534 ( .a(n13322), .b(n13321), .o(n13323) );
in01f01 g09535 ( .a(n13323), .o(n13324) );
no02f01 g09536 ( .a(n13324), .b(n13319), .o(n13325) );
no02f01 g09537 ( .a(n13323), .b(n13318), .o(n13326) );
no02f01 g09538 ( .a(n13326), .b(n13325), .o(n13327) );
in01f01 g09539 ( .a(n13327), .o(n13328) );
no02f01 g09540 ( .a(n13328), .b(n13317), .o(n13329) );
no02f01 g09541 ( .a(n13327), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_22_), .o(n13330) );
no02f01 g09542 ( .a(n13330), .b(n13329), .o(n13331) );
no02f01 g09543 ( .a(n13331), .b(n13316), .o(n13332) );
na02f01 g09544 ( .a(n13331), .b(n13316), .o(n13333) );
in01f01 g09545 ( .a(n13333), .o(n13334) );
no02f01 g09546 ( .a(n13334), .b(n13332), .o(n13335) );
in01f01 g09547 ( .a(n13335), .o(n13336) );
na03f01 g09548 ( .a(n13336), .b(n13314), .c(n13305), .o(n13337) );
no02f01 g09549 ( .a(n13313), .b(n13310), .o(n13338) );
no02f01 g09550 ( .a(n13304), .b(n13301), .o(n13339) );
oa12f01 g09551 ( .a(n13335), .b(n13339), .c(n13338), .o(n13340) );
na02f01 g09552 ( .a(n13340), .b(n13337), .o(n13341) );
no03f01 g09553 ( .a(n13271), .b(n13207), .c(n12725), .o(n13342) );
no02f01 g09554 ( .a(n13342), .b(n13268), .o(n13343) );
no02f01 g09555 ( .a(n13343), .b(n13341), .o(n13344) );
no03f01 g09556 ( .a(n13335), .b(n13339), .c(n13338), .o(n13345) );
ao12f01 g09557 ( .a(n13336), .b(n13314), .c(n13305), .o(n13346) );
no02f01 g09558 ( .a(n13346), .b(n13345), .o(n13347) );
in01f01 g09559 ( .a(n13268), .o(n13348) );
oa12f01 g09560 ( .a(n13020), .b(n13017), .c(n12736), .o(n13349) );
na03f01 g09561 ( .a(n13267), .b(n13246), .c(n13239), .o(n13350) );
na03f01 g09562 ( .a(n13350), .b(n13349), .c(n13021), .o(n13351) );
na02f01 g09563 ( .a(n13351), .b(n13348), .o(n13352) );
no02f01 g09564 ( .a(n13352), .b(n13347), .o(n13353) );
no02f01 g09565 ( .a(n13353), .b(n13344), .o(n13354) );
no02f01 g09566 ( .a(n13354), .b(n11515), .o(n13355) );
no02f01 g09567 ( .a(n13355), .b(n13277), .o(n13356) );
ao12f01 g09568 ( .a(n13309), .b(n13313), .c(n13299), .o(n13357) );
in01f01 g09569 ( .a(delay_add_ln22_unr2_stage2_stallmux_q_27_), .o(n13358) );
no02f01 g09570 ( .a(n13281), .b(n13280), .o(n13359) );
in01f01 g09571 ( .a(n13359), .o(n13360) );
no02f01 g09572 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_27_), .b(n11021), .o(n13361) );
in01f01 g09573 ( .a(n13361), .o(n13362) );
na02f01 g09574 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_27_), .b(n11021), .o(n13363) );
na02f01 g09575 ( .a(n13363), .b(n13362), .o(n13364) );
in01f01 g09576 ( .a(n13364), .o(n13365) );
no02f01 g09577 ( .a(n13365), .b(n13360), .o(n13366) );
no02f01 g09578 ( .a(n13364), .b(n13359), .o(n13367) );
no02f01 g09579 ( .a(n13367), .b(n13366), .o(n13368) );
no02f01 g09580 ( .a(n13368), .b(n13358), .o(n13369) );
na02f01 g09581 ( .a(n13368), .b(n13358), .o(n13370) );
in01f01 g09582 ( .a(n13370), .o(n13371) );
no02f01 g09583 ( .a(n13371), .b(n13369), .o(n13372) );
ao12f01 g09584 ( .a(n13289), .b(n13294), .c(n13278), .o(n13373) );
oa12f01 g09585 ( .a(n13372), .b(n13373), .c(n13291), .o(n13374) );
no03f01 g09586 ( .a(n13373), .b(n13372), .c(n13291), .o(n13375) );
in01f01 g09587 ( .a(n13375), .o(n13376) );
na02f01 g09588 ( .a(n13376), .b(n13374), .o(n13377) );
na02f01 g09589 ( .a(n13377), .b(n11158), .o(n13378) );
na02f01 g09590 ( .a(n13377), .b(n11179), .o(n13379) );
na02f01 g09591 ( .a(n13379), .b(n13378), .o(n13380) );
no02f01 g09592 ( .a(n13380), .b(n13357), .o(n13381) );
oa12f01 g09593 ( .a(n13300), .b(n13304), .c(n13308), .o(n13382) );
ao12f01 g09594 ( .a(n11179), .b(n13376), .c(n13374), .o(n13383) );
in01f01 g09595 ( .a(n13374), .o(n13384) );
no02f01 g09596 ( .a(n13375), .b(n13384), .o(n13385) );
no02f01 g09597 ( .a(n13385), .b(n11158), .o(n13386) );
no02f01 g09598 ( .a(n13386), .b(n13383), .o(n13387) );
no02f01 g09599 ( .a(n13387), .b(n13382), .o(n13388) );
no02f01 g09600 ( .a(n13388), .b(n13381), .o(n13389) );
no02f01 g09601 ( .a(n13329), .b(n13315), .o(n13390) );
no02f01 g09602 ( .a(n13390), .b(n13330), .o(n13391) );
no02f01 g09603 ( .a(n13320), .b(n13319), .o(n13392) );
in01f01 g09604 ( .a(n13392), .o(n13393) );
no02f01 g09605 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_23_), .b(n11021), .o(n13394) );
in01f01 g09606 ( .a(n13394), .o(n13395) );
na02f01 g09607 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_23_), .b(n11021), .o(n13396) );
na02f01 g09608 ( .a(n13396), .b(n13395), .o(n13397) );
in01f01 g09609 ( .a(n13397), .o(n13398) );
no02f01 g09610 ( .a(n13398), .b(n13393), .o(n13399) );
no02f01 g09611 ( .a(n13397), .b(n13392), .o(n13400) );
no02f01 g09612 ( .a(n13400), .b(n13399), .o(n13401) );
no02f01 g09613 ( .a(n13401), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_23_), .o(n13402) );
na02f01 g09614 ( .a(n13401), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_23_), .o(n13403) );
in01f01 g09615 ( .a(n13403), .o(n13404) );
no02f01 g09616 ( .a(n13404), .b(n13402), .o(n13405) );
in01f01 g09617 ( .a(n13405), .o(n13406) );
no02f01 g09618 ( .a(n13406), .b(n13391), .o(n13407) );
na02f01 g09619 ( .a(n13406), .b(n13391), .o(n13408) );
in01f01 g09620 ( .a(n13408), .o(n13409) );
no02f01 g09621 ( .a(n13409), .b(n13407), .o(n13410) );
in01f01 g09622 ( .a(n13410), .o(n13411) );
no02f01 g09623 ( .a(n13411), .b(n13389), .o(n13412) );
na02f01 g09624 ( .a(n13387), .b(n13382), .o(n13413) );
na02f01 g09625 ( .a(n13380), .b(n13357), .o(n13414) );
na03f01 g09626 ( .a(n13411), .b(n13414), .c(n13413), .o(n13415) );
in01f01 g09627 ( .a(n13415), .o(n13416) );
no02f01 g09628 ( .a(n13416), .b(n13412), .o(n13417) );
oa12f01 g09629 ( .a(n13340), .b(n13343), .c(n13345), .o(n13418) );
no02f01 g09630 ( .a(n13418), .b(n13417), .o(n13419) );
oa12f01 g09631 ( .a(n13410), .b(n13388), .c(n13381), .o(n13420) );
na02f01 g09632 ( .a(n13415), .b(n13420), .o(n13421) );
na02f01 g09633 ( .a(n13352), .b(n13337), .o(n13422) );
ao12f01 g09634 ( .a(n13421), .b(n13422), .c(n13340), .o(n13423) );
no02f01 g09635 ( .a(n13423), .b(n13419), .o(n13424) );
oa12f01 g09636 ( .a(n13356), .b(n13424), .c(n11515), .o(n13425) );
na02f01 g09637 ( .a(n13414), .b(n13413), .o(n13426) );
na03f01 g09638 ( .a(n13351), .b(n13340), .c(n13348), .o(n13427) );
na02f01 g09639 ( .a(n13410), .b(n13337), .o(n13428) );
in01f01 g09640 ( .a(n13428), .o(n13429) );
ao12f01 g09641 ( .a(n13426), .b(n13429), .c(n13427), .o(n13430) );
ao12f01 g09642 ( .a(n13410), .b(n13427), .c(n13337), .o(n13431) );
no02f01 g09643 ( .a(n13431), .b(n13430), .o(n13432) );
no02f01 g09644 ( .a(n13302), .b(n13309), .o(n13433) );
na03f01 g09645 ( .a(n13433), .b(n13378), .c(n12428), .o(n13434) );
no02f01 g09646 ( .a(n13312), .b(n13308), .o(n13435) );
in01f01 g09647 ( .a(n13435), .o(n13436) );
no02f01 g09648 ( .a(n13436), .b(n13386), .o(n13437) );
na03f01 g09649 ( .a(n13433), .b(n13378), .c(n12430), .o(n13438) );
na03f01 g09650 ( .a(n13438), .b(n13437), .c(n13434), .o(n13439) );
in01f01 g09651 ( .a(n13289), .o(n13440) );
na03f01 g09652 ( .a(n13294), .b(n13290), .c(n13278), .o(n13441) );
ao12f01 g09653 ( .a(n13371), .b(n13441), .c(n13440), .o(n13442) );
in01f01 g09654 ( .a(delay_add_ln22_unr2_stage2_stallmux_q_28_), .o(n13443) );
no02f01 g09655 ( .a(n13361), .b(n13360), .o(n13444) );
in01f01 g09656 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_28_), .o(n13445) );
no02f01 g09657 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(n13445), .o(n13446) );
no02f01 g09658 ( .a(n11021), .b(delay_xor_ln22_unr3_stage2_stallmux_q_28_), .o(n13447) );
no02f01 g09659 ( .a(n13447), .b(n13446), .o(n13448) );
in01f01 g09660 ( .a(n13448), .o(n13449) );
no02f01 g09661 ( .a(n13449), .b(n13444), .o(n13450) );
in01f01 g09662 ( .a(n13450), .o(n13451) );
na02f01 g09663 ( .a(n13449), .b(n13444), .o(n13452) );
na02f01 g09664 ( .a(n13452), .b(n13451), .o(n13453) );
in01f01 g09665 ( .a(n13453), .o(n13454) );
no02f01 g09666 ( .a(n13454), .b(n13443), .o(n13455) );
no03f01 g09667 ( .a(n13455), .b(n13442), .c(n13369), .o(n13456) );
no02f01 g09668 ( .a(n13453), .b(delay_add_ln22_unr2_stage2_stallmux_q_28_), .o(n13457) );
in01f01 g09669 ( .a(n13457), .o(n13458) );
na02f01 g09670 ( .a(n13458), .b(n13456), .o(n13459) );
oa22f01 g09671 ( .a(n13457), .b(n13455), .c(n13442), .d(n13369), .o(n13460) );
na02f01 g09672 ( .a(n13460), .b(n13459), .o(n13461) );
na02f01 g09673 ( .a(n13461), .b(n11179), .o(n13462) );
in01f01 g09674 ( .a(n13462), .o(n13463) );
na02f01 g09675 ( .a(n13461), .b(n11158), .o(n13464) );
in01f01 g09676 ( .a(n13464), .o(n13465) );
no03f01 g09677 ( .a(n13465), .b(n13463), .c(n13439), .o(n13466) );
na02f01 g09678 ( .a(n13311), .b(n13300), .o(n13467) );
no03f01 g09679 ( .a(n13467), .b(n13383), .c(n12252), .o(n13468) );
na02f01 g09680 ( .a(n13435), .b(n13379), .o(n13469) );
no03f01 g09681 ( .a(n13467), .b(n13383), .c(n12396), .o(n13470) );
no03f01 g09682 ( .a(n13470), .b(n13469), .c(n13468), .o(n13471) );
ao12f01 g09683 ( .a(n13471), .b(n13464), .c(n13462), .o(n13472) );
in01f01 g09684 ( .a(n13402), .o(n13473) );
no02f01 g09685 ( .a(n13404), .b(n13329), .o(n13474) );
oa12f01 g09686 ( .a(n13474), .b(n13330), .c(n13316), .o(n13475) );
no02f01 g09687 ( .a(n13394), .b(n13393), .o(n13476) );
in01f01 g09688 ( .a(n13476), .o(n13477) );
no02f01 g09689 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_24_), .b(n11021), .o(n13478) );
in01f01 g09690 ( .a(n13478), .o(n13479) );
na02f01 g09691 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_24_), .b(n11021), .o(n13480) );
na02f01 g09692 ( .a(n13480), .b(n13479), .o(n13481) );
in01f01 g09693 ( .a(n13481), .o(n13482) );
no02f01 g09694 ( .a(n13482), .b(n13477), .o(n13483) );
no02f01 g09695 ( .a(n13481), .b(n13476), .o(n13484) );
no02f01 g09696 ( .a(n13484), .b(n13483), .o(n13485) );
no02f01 g09697 ( .a(n13485), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_24_), .o(n13486) );
na02f01 g09698 ( .a(n13485), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_24_), .o(n13487) );
in01f01 g09699 ( .a(n13487), .o(n13488) );
no02f01 g09700 ( .a(n13488), .b(n13486), .o(n13489) );
in01f01 g09701 ( .a(n13489), .o(n13490) );
ao12f01 g09702 ( .a(n13490), .b(n13475), .c(n13473), .o(n13491) );
na02f01 g09703 ( .a(n13475), .b(n13473), .o(n13492) );
no02f01 g09704 ( .a(n13489), .b(n13492), .o(n13493) );
no02f01 g09705 ( .a(n13493), .b(n13491), .o(n13494) );
no03f01 g09706 ( .a(n13494), .b(n13472), .c(n13466), .o(n13495) );
na03f01 g09707 ( .a(n13464), .b(n13462), .c(n13471), .o(n13496) );
oa12f01 g09708 ( .a(n13439), .b(n13465), .c(n13463), .o(n13497) );
in01f01 g09709 ( .a(n13494), .o(n13498) );
ao12f01 g09710 ( .a(n13498), .b(n13497), .c(n13496), .o(n13499) );
no02f01 g09711 ( .a(n13499), .b(n13495), .o(n13500) );
na02f01 g09712 ( .a(n13500), .b(n13432), .o(n13501) );
no03f01 g09713 ( .a(n13342), .b(n13346), .c(n13268), .o(n13502) );
oa12f01 g09714 ( .a(n13389), .b(n13428), .c(n13502), .o(n13503) );
oa12f01 g09715 ( .a(n13411), .b(n13502), .c(n13345), .o(n13504) );
na02f01 g09716 ( .a(n13504), .b(n13503), .o(n13505) );
na03f01 g09717 ( .a(n13498), .b(n13497), .c(n13496), .o(n13506) );
oa12f01 g09718 ( .a(n13494), .b(n13472), .c(n13466), .o(n13507) );
na02f01 g09719 ( .a(n13507), .b(n13506), .o(n13508) );
na02f01 g09720 ( .a(n13508), .b(n13505), .o(n13509) );
na02f01 g09721 ( .a(n13509), .b(n13501), .o(n13510) );
ao12f01 g09722 ( .a(n13425), .b(n13510), .c(n11514), .o(n13511) );
no02f01 g09723 ( .a(n13508), .b(n13505), .o(n13512) );
no02f01 g09724 ( .a(n13500), .b(n13432), .o(n13513) );
no02f01 g09725 ( .a(n13513), .b(n13512), .o(n13514) );
na03f01 g09726 ( .a(n13422), .b(n13421), .c(n13340), .o(n13515) );
na02f01 g09727 ( .a(n13418), .b(n13417), .o(n13516) );
na02f01 g09728 ( .a(n13516), .b(n13515), .o(n13517) );
na02f01 g09729 ( .a(n13352), .b(n13347), .o(n13518) );
na02f01 g09730 ( .a(n13343), .b(n13341), .o(n13519) );
na02f01 g09731 ( .a(n13519), .b(n13518), .o(n13520) );
na02f01 g09732 ( .a(n13520), .b(n11515), .o(n13521) );
in01f01 g09733 ( .a(n13275), .o(n13522) );
na02f01 g09734 ( .a(n13522), .b(n13273), .o(n13523) );
na02f01 g09735 ( .a(n13523), .b(n11515), .o(n13524) );
na02f01 g09736 ( .a(n13524), .b(n13521), .o(n13525) );
ao12f01 g09737 ( .a(n13525), .b(n13517), .c(n11515), .o(n13526) );
oa12f01 g09738 ( .a(n13526), .b(n13514), .c(n11514), .o(n13527) );
no02f01 g09739 ( .a(n13527), .b(n13511), .o(n13528) );
na02f01 g09740 ( .a(n13462), .b(n13471), .o(n13529) );
no02f01 g09741 ( .a(n13450), .b(n13446), .o(n13530) );
in01f01 g09742 ( .a(n13530), .o(n13531) );
no02f01 g09743 ( .a(n13531), .b(delay_add_ln22_unr2_stage2_stallmux_q_29_), .o(n13532) );
na02f01 g09744 ( .a(n13531), .b(delay_add_ln22_unr2_stage2_stallmux_q_29_), .o(n13533) );
in01f01 g09745 ( .a(n13533), .o(n13534) );
no02f01 g09746 ( .a(n13534), .b(n13532), .o(n13535) );
oa12f01 g09747 ( .a(n13535), .b(n13457), .c(n13456), .o(n13536) );
no03f01 g09748 ( .a(n13535), .b(n13457), .c(n13456), .o(n13537) );
in01f01 g09749 ( .a(n13537), .o(n13538) );
na02f01 g09750 ( .a(n13538), .b(n13536), .o(n13539) );
na02f01 g09751 ( .a(n13539), .b(n11179), .o(n13540) );
na02f01 g09752 ( .a(n13539), .b(n11158), .o(n13541) );
na02f01 g09753 ( .a(n13541), .b(n13540), .o(n13542) );
na03f01 g09754 ( .a(n13542), .b(n13464), .c(n13529), .o(n13543) );
no02f01 g09755 ( .a(n13463), .b(n13439), .o(n13544) );
in01f01 g09756 ( .a(n13536), .o(n13545) );
no02f01 g09757 ( .a(n13537), .b(n13545), .o(n13546) );
no02f01 g09758 ( .a(n13546), .b(n11158), .o(n13547) );
no02f01 g09759 ( .a(n13546), .b(n11179), .o(n13548) );
no02f01 g09760 ( .a(n13548), .b(n13547), .o(n13549) );
oa12f01 g09761 ( .a(n13549), .b(n13465), .c(n13544), .o(n13550) );
oa12f01 g09762 ( .a(n13487), .b(n13486), .c(n13492), .o(n13551) );
no02f01 g09763 ( .a(n13478), .b(n13477), .o(n13552) );
in01f01 g09764 ( .a(n13552), .o(n13553) );
no02f01 g09765 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_25_), .b(n11021), .o(n13554) );
in01f01 g09766 ( .a(n13554), .o(n13555) );
na02f01 g09767 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_25_), .b(n11021), .o(n13556) );
na02f01 g09768 ( .a(n13556), .b(n13555), .o(n13557) );
in01f01 g09769 ( .a(n13557), .o(n13558) );
no02f01 g09770 ( .a(n13558), .b(n13553), .o(n13559) );
no02f01 g09771 ( .a(n13557), .b(n13552), .o(n13560) );
no02f01 g09772 ( .a(n13560), .b(n13559), .o(n13561) );
no02f01 g09773 ( .a(n13561), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_25_), .o(n13562) );
na02f01 g09774 ( .a(n13561), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_25_), .o(n13563) );
in01f01 g09775 ( .a(n13563), .o(n13564) );
no02f01 g09776 ( .a(n13564), .b(n13562), .o(n13565) );
in01f01 g09777 ( .a(n13565), .o(n13566) );
no02f01 g09778 ( .a(n13566), .b(n13551), .o(n13567) );
in01f01 g09779 ( .a(n13551), .o(n13568) );
no02f01 g09780 ( .a(n13565), .b(n13568), .o(n13569) );
no02f01 g09781 ( .a(n13569), .b(n13567), .o(n13570) );
in01f01 g09782 ( .a(n13570), .o(n13571) );
na03f01 g09783 ( .a(n13571), .b(n13550), .c(n13543), .o(n13572) );
no03f01 g09784 ( .a(n13549), .b(n13465), .c(n13544), .o(n13573) );
ao12f01 g09785 ( .a(n13542), .b(n13464), .c(n13529), .o(n13574) );
oa12f01 g09786 ( .a(n13570), .b(n13574), .c(n13573), .o(n13575) );
na02f01 g09787 ( .a(n13575), .b(n13572), .o(n13576) );
oa12f01 g09788 ( .a(n13507), .b(n13431), .c(n13430), .o(n13577) );
na02f01 g09789 ( .a(n13577), .b(n13506), .o(n13578) );
no02f01 g09790 ( .a(n13578), .b(n13576), .o(n13579) );
no03f01 g09791 ( .a(n13570), .b(n13574), .c(n13573), .o(n13580) );
ao12f01 g09792 ( .a(n13571), .b(n13550), .c(n13543), .o(n13581) );
no02f01 g09793 ( .a(n13581), .b(n13580), .o(n13582) );
ao12f01 g09794 ( .a(n13499), .b(n13504), .c(n13503), .o(n13583) );
no02f01 g09795 ( .a(n13583), .b(n13495), .o(n13584) );
no02f01 g09796 ( .a(n13584), .b(n13582), .o(n13585) );
no02f01 g09797 ( .a(n13585), .b(n13579), .o(n13586) );
no02f01 g09798 ( .a(n13586), .b(n11515), .o(n13587) );
no02f01 g09799 ( .a(n13586), .b(n11514), .o(n13588) );
no02f01 g09800 ( .a(n13588), .b(n13587), .o(n13589) );
no02f01 g09801 ( .a(n13589), .b(n13528), .o(n13590) );
na02f01 g09802 ( .a(n13589), .b(n13528), .o(n13591) );
in01f01 g09803 ( .a(n13591), .o(n13592) );
no02f01 g09804 ( .a(n12735), .b(n11179), .o(n13593) );
no02f01 g09805 ( .a(n12746), .b(n11179), .o(n13594) );
ao12f01 g09806 ( .a(n11179), .b(n12876), .c(n12864), .o(n13595) );
ao12f01 g09807 ( .a(n13595), .b(n12941), .c(n11158), .o(n13596) );
no02f01 g09808 ( .a(n12852), .b(n11179), .o(n13597) );
in01f01 g09809 ( .a(n13597), .o(n13598) );
na02f01 g09810 ( .a(n13598), .b(n13596), .o(n13599) );
no02f01 g09811 ( .a(n12844), .b(n11179), .o(n13600) );
no02f01 g09812 ( .a(n13600), .b(n13599), .o(n13601) );
in01f01 g09813 ( .a(n13601), .o(n13602) );
no02f01 g09814 ( .a(n12831), .b(n11179), .o(n13603) );
no02f01 g09815 ( .a(n13603), .b(n13602), .o(n13604) );
in01f01 g09816 ( .a(n13604), .o(n13605) );
no02f01 g09817 ( .a(n12970), .b(n11179), .o(n13606) );
no02f01 g09818 ( .a(n13606), .b(n13605), .o(n13607) );
no02f01 g09819 ( .a(n12819), .b(n11179), .o(n13608) );
in01f01 g09820 ( .a(n13608), .o(n13609) );
na02f01 g09821 ( .a(n13609), .b(n13607), .o(n13610) );
no02f01 g09822 ( .a(n12814), .b(n11179), .o(n13611) );
no02f01 g09823 ( .a(n13611), .b(n13610), .o(n13612) );
oa12f01 g09824 ( .a(n13612), .b(n12800), .c(n11179), .o(n13613) );
ao12f01 g09825 ( .a(n13613), .b(n13002), .c(n11158), .o(n13614) );
no02f01 g09826 ( .a(n12783), .b(n11179), .o(n13615) );
in01f01 g09827 ( .a(n13615), .o(n13616) );
na02f01 g09828 ( .a(n13616), .b(n13614), .o(n13617) );
oa12f01 g09829 ( .a(n11179), .b(n12985), .c(n12801), .o(n13618) );
in01f01 g09830 ( .a(n13618), .o(n13619) );
ao12f01 g09831 ( .a(n13619), .b(n13002), .c(n11179), .o(n13620) );
in01f01 g09832 ( .a(n13620), .o(n13621) );
ao12f01 g09833 ( .a(n13621), .b(n12784), .c(n11179), .o(n13622) );
na02f01 g09834 ( .a(n13622), .b(n13617), .o(n13623) );
in01f01 g09835 ( .a(n13623), .o(n13624) );
no02f01 g09836 ( .a(n12770), .b(n11179), .o(n13625) );
ao12f01 g09837 ( .a(n13625), .b(n12760), .c(n11158), .o(n13626) );
in01f01 g09838 ( .a(n13626), .o(n13627) );
no04f01 g09839 ( .a(n13627), .b(n13624), .c(n13594), .d(n13593), .o(n13628) );
no02f01 g09840 ( .a(n12770), .b(n11158), .o(n13629) );
ao12f01 g09841 ( .a(n13629), .b(n12760), .c(n11179), .o(n13630) );
in01f01 g09842 ( .a(n13630), .o(n13631) );
ao12f01 g09843 ( .a(n13631), .b(n13032), .c(n11179), .o(n13632) );
oa12f01 g09844 ( .a(n13632), .b(n12735), .c(n11158), .o(n13633) );
no02f01 g09845 ( .a(n13633), .b(n13628), .o(n13634) );
ao12f01 g09846 ( .a(n13634), .b(n12721), .c(n11158), .o(n13635) );
oa12f01 g09847 ( .a(n13635), .b(n13266), .c(n11179), .o(n13636) );
ao12f01 g09848 ( .a(n13636), .b(n13336), .c(n11158), .o(n13637) );
no02f01 g09849 ( .a(n12720), .b(n11158), .o(n13638) );
ao12f01 g09850 ( .a(n13638), .b(n13267), .c(n11179), .o(n13639) );
in01f01 g09851 ( .a(n13639), .o(n13640) );
ao12f01 g09852 ( .a(n13640), .b(n13336), .c(n11179), .o(n13641) );
in01f01 g09853 ( .a(n13641), .o(n13642) );
no02f01 g09854 ( .a(n13642), .b(n13637), .o(n13643) );
no02f01 g09855 ( .a(n13643), .b(n13410), .o(n13644) );
na02f01 g09856 ( .a(n13643), .b(n13410), .o(n13645) );
in01f01 g09857 ( .a(n13645), .o(n13646) );
no02f01 g09858 ( .a(n13646), .b(n13644), .o(n13647) );
no02f01 g09859 ( .a(n13647), .b(n12261), .o(n13648) );
na02f01 g09860 ( .a(n13639), .b(n13636), .o(n13649) );
na02f01 g09861 ( .a(n13649), .b(n13336), .o(n13650) );
in01f01 g09862 ( .a(n13650), .o(n13651) );
no02f01 g09863 ( .a(n13649), .b(n13336), .o(n13652) );
no02f01 g09864 ( .a(n13652), .b(n13651), .o(n13653) );
no02f01 g09865 ( .a(n13653), .b(n12379), .o(n13654) );
in01f01 g09866 ( .a(n13654), .o(n13655) );
no02f01 g09867 ( .a(n13638), .b(n13635), .o(n13656) );
no02f01 g09868 ( .a(n13656), .b(n13266), .o(n13657) );
in01f01 g09869 ( .a(n13657), .o(n13658) );
na02f01 g09870 ( .a(n13656), .b(n13266), .o(n13659) );
na02f01 g09871 ( .a(n13659), .b(n13658), .o(n13660) );
no02f01 g09872 ( .a(n13660), .b(n12787), .o(n13661) );
in01f01 g09873 ( .a(n13661), .o(n13662) );
no02f01 g09874 ( .a(n13634), .b(n12720), .o(n13663) );
na02f01 g09875 ( .a(n13634), .b(n12720), .o(n13664) );
in01f01 g09876 ( .a(n13664), .o(n13665) );
no02f01 g09877 ( .a(n13665), .b(n13663), .o(n13666) );
no02f01 g09878 ( .a(n13666), .b(n12368), .o(n13667) );
in01f01 g09879 ( .a(n13667), .o(n13668) );
in01f01 g09880 ( .a(n13622), .o(n13669) );
no02f01 g09881 ( .a(n13629), .b(n13669), .o(n13670) );
oa12f01 g09882 ( .a(n13670), .b(n13625), .c(n13617), .o(n13671) );
in01f01 g09883 ( .a(n13671), .o(n13672) );
no02f01 g09884 ( .a(n13672), .b(n12759), .o(n13673) );
no02f01 g09885 ( .a(n13671), .b(n12760), .o(n13674) );
no02f01 g09886 ( .a(n13674), .b(n13673), .o(n13675) );
in01f01 g09887 ( .a(n13675), .o(n13676) );
no02f01 g09888 ( .a(n13621), .b(n13614), .o(n13677) );
no02f01 g09889 ( .a(n13677), .b(n12783), .o(n13678) );
na02f01 g09890 ( .a(n13677), .b(n12783), .o(n13679) );
in01f01 g09891 ( .a(n13679), .o(n13680) );
no02f01 g09892 ( .a(n13680), .b(n13678), .o(n13681) );
no02f01 g09893 ( .a(n13681), .b(n12275), .o(n13682) );
na02f01 g09894 ( .a(n13618), .b(n13613), .o(n13683) );
na02f01 g09895 ( .a(n13683), .b(n13002), .o(n13684) );
in01f01 g09896 ( .a(n13684), .o(n13685) );
no02f01 g09897 ( .a(n13683), .b(n13002), .o(n13686) );
no02f01 g09898 ( .a(n13686), .b(n13685), .o(n13687) );
no02f01 g09899 ( .a(n13687), .b(n12327), .o(n13688) );
in01f01 g09900 ( .a(n13688), .o(n13689) );
no03f01 g09901 ( .a(n13611), .b(n13610), .c(n12800), .o(n13690) );
no02f01 g09902 ( .a(n13612), .b(n12801), .o(n13691) );
no02f01 g09903 ( .a(n13691), .b(n13690), .o(n13692) );
na02f01 g09904 ( .a(n13692), .b(n12281), .o(n13693) );
no02f01 g09905 ( .a(n13610), .b(n12814), .o(n13694) );
na02f01 g09906 ( .a(n13610), .b(n12814), .o(n13695) );
in01f01 g09907 ( .a(n13695), .o(n13696) );
no02f01 g09908 ( .a(n13696), .b(n13694), .o(n13697) );
no02f01 g09909 ( .a(n13697), .b(n12319), .o(n13698) );
in01f01 g09910 ( .a(n13698), .o(n13699) );
na02f01 g09911 ( .a(n13607), .b(n12820), .o(n13700) );
in01f01 g09912 ( .a(n13700), .o(n13701) );
no02f01 g09913 ( .a(n13607), .b(n12820), .o(n13702) );
no02f01 g09914 ( .a(n13702), .b(n13701), .o(n13703) );
no02f01 g09915 ( .a(n13703), .b(n12287), .o(n13704) );
no02f01 g09916 ( .a(n13604), .b(n12971), .o(n13705) );
in01f01 g09917 ( .a(n13705), .o(n13706) );
na02f01 g09918 ( .a(n13604), .b(n12971), .o(n13707) );
na02f01 g09919 ( .a(n13707), .b(n13706), .o(n13708) );
na02f01 g09920 ( .a(n13708), .b(n12312), .o(n13709) );
no02f01 g09921 ( .a(n13602), .b(n12831), .o(n13710) );
no02f01 g09922 ( .a(n13601), .b(n12832), .o(n13711) );
no02f01 g09923 ( .a(n13711), .b(n13710), .o(n13712) );
no02f01 g09924 ( .a(n13712), .b(n12303), .o(n13713) );
in01f01 g09925 ( .a(n13596), .o(n13714) );
no02f01 g09926 ( .a(n13714), .b(n12852), .o(n13715) );
no02f01 g09927 ( .a(n13596), .b(n12853), .o(n13716) );
in01f01 g09928 ( .a(n12090), .o(n13717) );
no02f01 g09929 ( .a(n12091), .b(n12071), .o(n13718) );
no02f01 g09930 ( .a(n13718), .b(n13717), .o(n13719) );
na02f01 g09931 ( .a(n13718), .b(n13717), .o(n13720) );
in01f01 g09932 ( .a(n13720), .o(n13721) );
no02f01 g09933 ( .a(n13721), .b(n13719), .o(n13722) );
in01f01 g09934 ( .a(n13722), .o(n13723) );
oa12f01 g09935 ( .a(n13723), .b(n13716), .c(n13715), .o(n13724) );
in01f01 g09936 ( .a(n13724), .o(n13725) );
na03f01 g09937 ( .a(n12877), .b(n12864), .c(n11158), .o(n13726) );
oa12f01 g09938 ( .a(n12865), .b(n12876), .c(n11179), .o(n13727) );
no02f01 g09939 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_0_), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(n13728) );
no02f01 g09940 ( .a(n11873), .b(n11021), .o(n13729) );
no02f01 g09941 ( .a(n13729), .b(n13728), .o(n13730) );
in01f01 g09942 ( .a(n13730), .o(n13731) );
no02f01 g09943 ( .a(n13731), .b(n12876), .o(n13732) );
in01f01 g09944 ( .a(n13732), .o(n13733) );
no03f01 g09945 ( .a(n12077), .b(n12075), .c(delay_add_ln22_unr2_stage2_stallmux_q_1_), .o(n13734) );
no02f01 g09946 ( .a(n13734), .b(n12079), .o(n13735) );
in01f01 g09947 ( .a(n13735), .o(n13736) );
ao22f01 g09948 ( .a(n13736), .b(n13733), .c(n13727), .d(n13726), .o(n13737) );
no02f01 g09949 ( .a(n13736), .b(n13733), .o(n13738) );
in01f01 g09950 ( .a(n12079), .o(n13739) );
no02f01 g09951 ( .a(n12087), .b(delay_add_ln22_unr2_stage2_stallmux_q_2_), .o(n13740) );
in01f01 g09952 ( .a(delay_add_ln22_unr2_stage2_stallmux_q_2_), .o(n13741) );
ao12f01 g09953 ( .a(n13741), .b(n12086), .c(n12085), .o(n13742) );
no02f01 g09954 ( .a(n13742), .b(n13740), .o(n13743) );
no02f01 g09955 ( .a(n13743), .b(n13739), .o(n13744) );
na02f01 g09956 ( .a(n13743), .b(n13739), .o(n13745) );
in01f01 g09957 ( .a(n13745), .o(n13746) );
no02f01 g09958 ( .a(n13746), .b(n13744), .o(n13747) );
in01f01 g09959 ( .a(n13747), .o(n13748) );
no03f01 g09960 ( .a(n13748), .b(n13738), .c(n13737), .o(n13749) );
in01f01 g09961 ( .a(n13595), .o(n13750) );
no02f01 g09962 ( .a(n13750), .b(n12941), .o(n13751) );
no02f01 g09963 ( .a(n13595), .b(n12940), .o(n13752) );
no02f01 g09964 ( .a(n13752), .b(n13751), .o(n13753) );
oa12f01 g09965 ( .a(n13748), .b(n13738), .c(n13737), .o(n13754) );
oa12f01 g09966 ( .a(n13754), .b(n13753), .c(n13749), .o(n13755) );
no03f01 g09967 ( .a(n13723), .b(n13716), .c(n13715), .o(n13756) );
in01f01 g09968 ( .a(n13756), .o(n13757) );
ao12f01 g09969 ( .a(n13725), .b(n13757), .c(n13755), .o(n13758) );
no02f01 g09970 ( .a(n13599), .b(n12844), .o(n13759) );
in01f01 g09971 ( .a(n13759), .o(n13760) );
na02f01 g09972 ( .a(n13599), .b(n12844), .o(n13761) );
na02f01 g09973 ( .a(n13761), .b(n13760), .o(n13762) );
no02f01 g09974 ( .a(n13762), .b(n12296), .o(n13763) );
in01f01 g09975 ( .a(n13761), .o(n13764) );
no02f01 g09976 ( .a(n13764), .b(n13759), .o(n13765) );
no02f01 g09977 ( .a(n13765), .b(n12295), .o(n13766) );
in01f01 g09978 ( .a(n13766), .o(n13767) );
oa12f01 g09979 ( .a(n13767), .b(n13763), .c(n13758), .o(n13768) );
na02f01 g09980 ( .a(n13712), .b(n12303), .o(n13769) );
ao12f01 g09981 ( .a(n13713), .b(n13769), .c(n13768), .o(n13770) );
no02f01 g09982 ( .a(n13708), .b(n12312), .o(n13771) );
oa12f01 g09983 ( .a(n13709), .b(n13771), .c(n13770), .o(n13772) );
no03f01 g09984 ( .a(n13702), .b(n13701), .c(n12879), .o(n13773) );
in01f01 g09985 ( .a(n13773), .o(n13774) );
ao12f01 g09986 ( .a(n13704), .b(n13774), .c(n13772), .o(n13775) );
na02f01 g09987 ( .a(n13697), .b(n12319), .o(n13776) );
in01f01 g09988 ( .a(n13776), .o(n13777) );
oa12f01 g09989 ( .a(n13699), .b(n13777), .c(n13775), .o(n13778) );
no02f01 g09990 ( .a(n13692), .b(n12281), .o(n13779) );
oa12f01 g09991 ( .a(n13693), .b(n13779), .c(n13778), .o(n13780) );
in01f01 g09992 ( .a(n12327), .o(n13781) );
no03f01 g09993 ( .a(n13686), .b(n13685), .c(n13781), .o(n13782) );
oa12f01 g09994 ( .a(n13689), .b(n13782), .c(n13780), .o(n13783) );
na02f01 g09995 ( .a(n13681), .b(n12275), .o(n13784) );
ao12f01 g09996 ( .a(n13682), .b(n13784), .c(n13783), .o(n13785) );
na02f01 g09997 ( .a(n13623), .b(n12771), .o(n13786) );
na02f01 g09998 ( .a(n13624), .b(n12770), .o(n13787) );
na02f01 g09999 ( .a(n13787), .b(n13786), .o(n13788) );
no02f01 g10000 ( .a(n13788), .b(n12337), .o(n13789) );
ao12f01 g10001 ( .a(n12336), .b(n13787), .c(n13786), .o(n13790) );
no02f01 g10002 ( .a(n13790), .b(n12821), .o(n13791) );
oa12f01 g10003 ( .a(n13791), .b(n13789), .c(n13785), .o(n13792) );
in01f01 g10004 ( .a(n13790), .o(n13793) );
oa12f01 g10005 ( .a(n13793), .b(n13789), .c(n13785), .o(n13794) );
ao22f01 g10006 ( .a(n13794), .b(n12821), .c(n13792), .d(n13676), .o(n13795) );
no02f01 g10007 ( .a(n13627), .b(n13617), .o(n13796) );
no02f01 g10008 ( .a(n13631), .b(n13669), .o(n13797) );
in01f01 g10009 ( .a(n13797), .o(n13798) );
no02f01 g10010 ( .a(n13798), .b(n13796), .o(n13799) );
no02f01 g10011 ( .a(n13799), .b(n12746), .o(n13800) );
in01f01 g10012 ( .a(n13800), .o(n13801) );
na02f01 g10013 ( .a(n13799), .b(n12746), .o(n13802) );
na02f01 g10014 ( .a(n13802), .b(n13801), .o(n13803) );
no02f01 g10015 ( .a(n13803), .b(n12350), .o(n13804) );
in01f01 g10016 ( .a(n13594), .o(n13805) );
oa12f01 g10017 ( .a(n13797), .b(n12746), .c(n11158), .o(n13806) );
ao12f01 g10018 ( .a(n13806), .b(n13796), .c(n13805), .o(n13807) );
no02f01 g10019 ( .a(n13807), .b(n12735), .o(n13808) );
na02f01 g10020 ( .a(n13807), .b(n12735), .o(n13809) );
in01f01 g10021 ( .a(n13809), .o(n13810) );
no02f01 g10022 ( .a(n13810), .b(n13808), .o(n13811) );
no02f01 g10023 ( .a(n13811), .b(n12356), .o(n13812) );
ao12f01 g10024 ( .a(n12349), .b(n13802), .c(n13801), .o(n13813) );
no02f01 g10025 ( .a(n13813), .b(n13812), .o(n13814) );
oa12f01 g10026 ( .a(n13814), .b(n13804), .c(n13795), .o(n13815) );
in01f01 g10027 ( .a(n13811), .o(n13816) );
no02f01 g10028 ( .a(n13816), .b(n12358), .o(n13817) );
in01f01 g10029 ( .a(n13817), .o(n13818) );
na02f01 g10030 ( .a(n13666), .b(n12368), .o(n13819) );
na03f01 g10031 ( .a(n13819), .b(n13818), .c(n13815), .o(n13820) );
ao12f01 g10032 ( .a(n12268), .b(n13659), .c(n13658), .o(n13821) );
in01f01 g10033 ( .a(n13821), .o(n13822) );
na03f01 g10034 ( .a(n13822), .b(n13820), .c(n13668), .o(n13823) );
no03f01 g10035 ( .a(n13652), .b(n13651), .c(n12385), .o(n13824) );
in01f01 g10036 ( .a(n13824), .o(n13825) );
na03f01 g10037 ( .a(n13825), .b(n13823), .c(n13662), .o(n13826) );
no03f01 g10038 ( .a(n13646), .b(n13644), .c(n12773), .o(n13827) );
ao12f01 g10039 ( .a(n13827), .b(n13826), .c(n13655), .o(n13828) );
no02f01 g10040 ( .a(n13828), .b(n13648), .o(n13829) );
oa12f01 g10041 ( .a(n13637), .b(n13410), .c(n11179), .o(n13830) );
in01f01 g10042 ( .a(n13830), .o(n13831) );
oa12f01 g10043 ( .a(n13641), .b(n13410), .c(n11158), .o(n13832) );
no02f01 g10044 ( .a(n13832), .b(n13831), .o(n13833) );
no02f01 g10045 ( .a(n13833), .b(n13494), .o(n13834) );
na02f01 g10046 ( .a(n13833), .b(n13494), .o(n13835) );
in01f01 g10047 ( .a(n13835), .o(n13836) );
no02f01 g10048 ( .a(n13836), .b(n13834), .o(n13837) );
no02f01 g10049 ( .a(n13837), .b(n12235), .o(n13838) );
na02f01 g10050 ( .a(n13837), .b(n12235), .o(n13839) );
in01f01 g10051 ( .a(n13839), .o(n13840) );
no02f01 g10052 ( .a(n13840), .b(n13838), .o(n13841) );
na02f01 g10053 ( .a(n13841), .b(n13829), .o(n13842) );
in01f01 g10054 ( .a(n13648), .o(n13843) );
in01f01 g10055 ( .a(n13682), .o(n13844) );
in01f01 g10056 ( .a(n13693), .o(n13845) );
in01f01 g10057 ( .a(n13704), .o(n13846) );
in01f01 g10058 ( .a(n13709), .o(n13847) );
in01f01 g10059 ( .a(n13713), .o(n13848) );
no03f01 g10060 ( .a(n12876), .b(n12865), .c(n11179), .o(n13849) );
ao12f01 g10061 ( .a(n12864), .b(n12877), .c(n11158), .o(n13850) );
oa22f01 g10062 ( .a(n13735), .b(n13732), .c(n13850), .d(n13849), .o(n13851) );
in01f01 g10063 ( .a(n13738), .o(n13852) );
na03f01 g10064 ( .a(n13747), .b(n13852), .c(n13851), .o(n13853) );
in01f01 g10065 ( .a(n13753), .o(n13854) );
ao12f01 g10066 ( .a(n13747), .b(n13852), .c(n13851), .o(n13855) );
ao12f01 g10067 ( .a(n13855), .b(n13854), .c(n13853), .o(n13856) );
oa12f01 g10068 ( .a(n13724), .b(n13756), .c(n13856), .o(n13857) );
na02f01 g10069 ( .a(n13765), .b(n12295), .o(n13858) );
ao12f01 g10070 ( .a(n13766), .b(n13858), .c(n13857), .o(n13859) );
in01f01 g10071 ( .a(n13769), .o(n13860) );
oa12f01 g10072 ( .a(n13848), .b(n13860), .c(n13859), .o(n13861) );
in01f01 g10073 ( .a(n13771), .o(n13862) );
ao12f01 g10074 ( .a(n13847), .b(n13862), .c(n13861), .o(n13863) );
oa12f01 g10075 ( .a(n13846), .b(n13773), .c(n13863), .o(n13864) );
ao12f01 g10076 ( .a(n13698), .b(n13776), .c(n13864), .o(n13865) );
in01f01 g10077 ( .a(n13779), .o(n13866) );
ao12f01 g10078 ( .a(n13845), .b(n13866), .c(n13865), .o(n13867) );
in01f01 g10079 ( .a(n13782), .o(n13868) );
ao12f01 g10080 ( .a(n13688), .b(n13868), .c(n13867), .o(n13869) );
in01f01 g10081 ( .a(n13784), .o(n13870) );
oa12f01 g10082 ( .a(n13844), .b(n13870), .c(n13869), .o(n13871) );
in01f01 g10083 ( .a(n13789), .o(n13872) );
in01f01 g10084 ( .a(n13791), .o(n13873) );
ao12f01 g10085 ( .a(n13873), .b(n13872), .c(n13871), .o(n13874) );
ao12f01 g10086 ( .a(n13790), .b(n13872), .c(n13871), .o(n13875) );
oa22f01 g10087 ( .a(n13875), .b(n12343), .c(n13874), .d(n13675), .o(n13876) );
in01f01 g10088 ( .a(n13804), .o(n13877) );
in01f01 g10089 ( .a(n13814), .o(n13878) );
ao12f01 g10090 ( .a(n13878), .b(n13877), .c(n13876), .o(n13879) );
in01f01 g10091 ( .a(n13819), .o(n13880) );
no03f01 g10092 ( .a(n13880), .b(n13817), .c(n13879), .o(n13881) );
no03f01 g10093 ( .a(n13821), .b(n13881), .c(n13667), .o(n13882) );
no03f01 g10094 ( .a(n13824), .b(n13882), .c(n13661), .o(n13883) );
in01f01 g10095 ( .a(n13827), .o(n13884) );
oa12f01 g10096 ( .a(n13884), .b(n13883), .c(n13654), .o(n13885) );
na02f01 g10097 ( .a(n13885), .b(n13843), .o(n13886) );
in01f01 g10098 ( .a(n13841), .o(n13887) );
na02f01 g10099 ( .a(n13887), .b(n13886), .o(n13888) );
na02f01 g10100 ( .a(n13888), .b(n13842), .o(n13889) );
oa12f01 g10101 ( .a(n13889), .b(n13592), .c(n13590), .o(n13890) );
in01f01 g10102 ( .a(n13890), .o(n13891) );
na02f01 g10103 ( .a(n13526), .b(n13425), .o(n13892) );
in01f01 g10104 ( .a(n13892), .o(n13893) );
no02f01 g10105 ( .a(n13514), .b(n11515), .o(n13894) );
no02f01 g10106 ( .a(n13514), .b(n11514), .o(n13895) );
no02f01 g10107 ( .a(n13895), .b(n13894), .o(n13896) );
na02f01 g10108 ( .a(n13896), .b(n13893), .o(n13897) );
no02f01 g10109 ( .a(n13896), .b(n13893), .o(n13898) );
in01f01 g10110 ( .a(n13898), .o(n13899) );
na02f01 g10111 ( .a(n13899), .b(n13897), .o(n13900) );
no02f01 g10112 ( .a(n13883), .b(n13654), .o(n13901) );
no02f01 g10113 ( .a(n13827), .b(n13648), .o(n13902) );
no02f01 g10114 ( .a(n13902), .b(n13901), .o(n13903) );
na02f01 g10115 ( .a(n13902), .b(n13901), .o(n13904) );
in01f01 g10116 ( .a(n13904), .o(n13905) );
no02f01 g10117 ( .a(n13905), .b(n13903), .o(n13906) );
in01f01 g10118 ( .a(n13906), .o(n13907) );
no02f01 g10119 ( .a(n13907), .b(n13900), .o(n13908) );
in01f01 g10120 ( .a(n13908), .o(n13909) );
na02f01 g10121 ( .a(n13907), .b(n13900), .o(n13910) );
no02f01 g10122 ( .a(n13525), .b(n13356), .o(n13911) );
no02f01 g10123 ( .a(n13424), .b(n11515), .o(n13912) );
no02f01 g10124 ( .a(n13424), .b(n11514), .o(n13913) );
no02f01 g10125 ( .a(n13913), .b(n13912), .o(n13914) );
no02f01 g10126 ( .a(n13914), .b(n13911), .o(n13915) );
na02f01 g10127 ( .a(n13914), .b(n13911), .o(n13916) );
in01f01 g10128 ( .a(n13916), .o(n13917) );
no02f01 g10129 ( .a(n13917), .b(n13915), .o(n13918) );
no02f01 g10130 ( .a(n13882), .b(n13661), .o(n13919) );
no02f01 g10131 ( .a(n13824), .b(n13654), .o(n13920) );
in01f01 g10132 ( .a(n13920), .o(n13921) );
no02f01 g10133 ( .a(n13921), .b(n13919), .o(n13922) );
na02f01 g10134 ( .a(n13921), .b(n13919), .o(n13923) );
in01f01 g10135 ( .a(n13923), .o(n13924) );
no02f01 g10136 ( .a(n13924), .b(n13922), .o(n13925) );
no02f01 g10137 ( .a(n13925), .b(n13918), .o(n13926) );
in01f01 g10138 ( .a(n13521), .o(n13927) );
no02f01 g10139 ( .a(n13927), .b(n13355), .o(n13928) );
na02f01 g10140 ( .a(n13524), .b(n13277), .o(n13929) );
in01f01 g10141 ( .a(n13929), .o(n13930) );
no02f01 g10142 ( .a(n13930), .b(n13928), .o(n13931) );
in01f01 g10143 ( .a(n13931), .o(n13932) );
na02f01 g10144 ( .a(n13930), .b(n13928), .o(n13933) );
na02f01 g10145 ( .a(n13933), .b(n13932), .o(n13934) );
na02f01 g10146 ( .a(n13820), .b(n13668), .o(n13935) );
no02f01 g10147 ( .a(n13821), .b(n13661), .o(n13936) );
in01f01 g10148 ( .a(n13936), .o(n13937) );
no02f01 g10149 ( .a(n13937), .b(n13935), .o(n13938) );
na02f01 g10150 ( .a(n13937), .b(n13935), .o(n13939) );
in01f01 g10151 ( .a(n13939), .o(n13940) );
no02f01 g10152 ( .a(n13940), .b(n13938), .o(n13941) );
in01f01 g10153 ( .a(n13941), .o(n13942) );
no02f01 g10154 ( .a(n13942), .b(n13934), .o(n13943) );
na02f01 g10155 ( .a(n13942), .b(n13934), .o(n13944) );
no02f01 g10156 ( .a(n13206), .b(n13195), .o(n13945) );
no02f01 g10157 ( .a(n13276), .b(n11515), .o(n13946) );
in01f01 g10158 ( .a(n13524), .o(n13947) );
no02f01 g10159 ( .a(n13947), .b(n13946), .o(n13948) );
no02f01 g10160 ( .a(n13948), .b(n13945), .o(n13949) );
na02f01 g10161 ( .a(n13948), .b(n13945), .o(n13950) );
in01f01 g10162 ( .a(n13950), .o(n13951) );
no02f01 g10163 ( .a(n13951), .b(n13949), .o(n13952) );
no02f01 g10164 ( .a(n13817), .b(n13879), .o(n13953) );
in01f01 g10165 ( .a(n13953), .o(n13954) );
no02f01 g10166 ( .a(n13880), .b(n13667), .o(n13955) );
no02f01 g10167 ( .a(n13955), .b(n13954), .o(n13956) );
na02f01 g10168 ( .a(n13955), .b(n13954), .o(n13957) );
in01f01 g10169 ( .a(n13957), .o(n13958) );
no02f01 g10170 ( .a(n13958), .b(n13956), .o(n13959) );
no02f01 g10171 ( .a(n13959), .b(n13952), .o(n13960) );
in01f01 g10172 ( .a(n13960), .o(n13961) );
ao12f01 g10173 ( .a(n13943), .b(n13961), .c(n13944), .o(n13962) );
na02f01 g10174 ( .a(n13925), .b(n13918), .o(n13963) );
ao12f01 g10175 ( .a(n13926), .b(n13963), .c(n13962), .o(n13964) );
na02f01 g10176 ( .a(n13964), .b(n13910), .o(n13965) );
in01f01 g10177 ( .a(n13943), .o(n13966) );
no02f01 g10178 ( .a(n13039), .b(n11514), .o(n13967) );
no02f01 g10179 ( .a(n13967), .b(n13040), .o(n13968) );
in01f01 g10180 ( .a(n13968), .o(n13969) );
in01f01 g10181 ( .a(n13193), .o(n13970) );
in01f01 g10182 ( .a(n13199), .o(n13971) );
no02f01 g10183 ( .a(n13204), .b(n13185), .o(n13972) );
ao12f01 g10184 ( .a(n13970), .b(n13972), .c(n13971), .o(n13973) );
no02f01 g10185 ( .a(n13973), .b(n13969), .o(n13974) );
na02f01 g10186 ( .a(n13973), .b(n13969), .o(n13975) );
in01f01 g10187 ( .a(n13975), .o(n13976) );
no02f01 g10188 ( .a(n13976), .b(n13974), .o(n13977) );
in01f01 g10189 ( .a(n13977), .o(n13978) );
oa12f01 g10190 ( .a(n13877), .b(n13813), .c(n13876), .o(n13979) );
no02f01 g10191 ( .a(n13817), .b(n13812), .o(n13980) );
no02f01 g10192 ( .a(n13980), .b(n13979), .o(n13981) );
na02f01 g10193 ( .a(n13980), .b(n13979), .o(n13982) );
in01f01 g10194 ( .a(n13982), .o(n13983) );
no02f01 g10195 ( .a(n13983), .b(n13981), .o(n13984) );
in01f01 g10196 ( .a(n13984), .o(n13985) );
no02f01 g10197 ( .a(n13985), .b(n13978), .o(n13986) );
na02f01 g10198 ( .a(n13203), .b(n13176), .o(n13987) );
in01f01 g10199 ( .a(n13202), .o(n13988) );
no02f01 g10200 ( .a(n13988), .b(n13184), .o(n13989) );
in01f01 g10201 ( .a(n13989), .o(n13990) );
no02f01 g10202 ( .a(n13990), .b(n13987), .o(n13991) );
na02f01 g10203 ( .a(n13990), .b(n13987), .o(n13992) );
in01f01 g10204 ( .a(n13992), .o(n13993) );
no02f01 g10205 ( .a(n13993), .b(n13991), .o(n13994) );
in01f01 g10206 ( .a(n13994), .o(n13995) );
ao12f01 g10207 ( .a(n13789), .b(n13793), .c(n13785), .o(n13996) );
no02f01 g10208 ( .a(n13676), .b(n12821), .o(n13997) );
no02f01 g10209 ( .a(n13675), .b(n12343), .o(n13998) );
no02f01 g10210 ( .a(n13998), .b(n13997), .o(n13999) );
in01f01 g10211 ( .a(n13999), .o(n14000) );
no02f01 g10212 ( .a(n14000), .b(n13996), .o(n14001) );
na02f01 g10213 ( .a(n14000), .b(n13996), .o(n14002) );
in01f01 g10214 ( .a(n14002), .o(n14003) );
no02f01 g10215 ( .a(n14003), .b(n14001), .o(n14004) );
in01f01 g10216 ( .a(n14004), .o(n14005) );
no02f01 g10217 ( .a(n14005), .b(n13995), .o(n14006) );
in01f01 g10218 ( .a(n14006), .o(n14007) );
no02f01 g10219 ( .a(n13167), .b(n13160), .o(n14008) );
in01f01 g10220 ( .a(n14008), .o(n14009) );
na02f01 g10221 ( .a(n13203), .b(n13175), .o(n14010) );
no02f01 g10222 ( .a(n14010), .b(n14009), .o(n14011) );
na02f01 g10223 ( .a(n14010), .b(n14009), .o(n14012) );
in01f01 g10224 ( .a(n14012), .o(n14013) );
no02f01 g10225 ( .a(n14013), .b(n14011), .o(n14014) );
no02f01 g10226 ( .a(n13790), .b(n13789), .o(n14015) );
no02f01 g10227 ( .a(n14015), .b(n13785), .o(n14016) );
na02f01 g10228 ( .a(n14015), .b(n13785), .o(n14017) );
in01f01 g10229 ( .a(n14017), .o(n14018) );
no02f01 g10230 ( .a(n14018), .b(n14016), .o(n14019) );
no02f01 g10231 ( .a(n14019), .b(n14014), .o(n14020) );
in01f01 g10232 ( .a(n14020), .o(n14021) );
oa12f01 g10233 ( .a(n13166), .b(n13151), .c(n13142), .o(n14022) );
in01f01 g10234 ( .a(n14022), .o(n14023) );
no02f01 g10235 ( .a(n13158), .b(n11514), .o(n14024) );
no02f01 g10236 ( .a(n14024), .b(n13159), .o(n14025) );
no02f01 g10237 ( .a(n14025), .b(n14023), .o(n14026) );
na02f01 g10238 ( .a(n14025), .b(n14023), .o(n14027) );
in01f01 g10239 ( .a(n14027), .o(n14028) );
no02f01 g10240 ( .a(n14028), .b(n14026), .o(n14029) );
in01f01 g10241 ( .a(n14029), .o(n14030) );
no03f01 g10242 ( .a(n13870), .b(n13783), .c(n13682), .o(n14031) );
ao12f01 g10243 ( .a(n13869), .b(n13784), .c(n13844), .o(n14032) );
no02f01 g10244 ( .a(n14032), .b(n14031), .o(n14033) );
in01f01 g10245 ( .a(n14033), .o(n14034) );
no02f01 g10246 ( .a(n14034), .b(n14030), .o(n14035) );
in01f01 g10247 ( .a(n14035), .o(n14036) );
na02f01 g10248 ( .a(n13132), .b(n13124), .o(n14037) );
in01f01 g10249 ( .a(n14037), .o(n14038) );
ao12f01 g10250 ( .a(n13164), .b(n13141), .c(n14038), .o(n14039) );
no02f01 g10251 ( .a(n13165), .b(n13151), .o(n14040) );
no02f01 g10252 ( .a(n14040), .b(n14039), .o(n14041) );
na02f01 g10253 ( .a(n14040), .b(n14039), .o(n14042) );
in01f01 g10254 ( .a(n14042), .o(n14043) );
no02f01 g10255 ( .a(n14043), .b(n14041), .o(n14044) );
no03f01 g10256 ( .a(n13782), .b(n13867), .c(n13688), .o(n14045) );
ao12f01 g10257 ( .a(n13780), .b(n13868), .c(n13689), .o(n14046) );
no02f01 g10258 ( .a(n14046), .b(n14045), .o(n14047) );
no02f01 g10259 ( .a(n14047), .b(n14044), .o(n14048) );
in01f01 g10260 ( .a(n14048), .o(n14049) );
na02f01 g10261 ( .a(n13163), .b(n14037), .o(n14050) );
na02f01 g10262 ( .a(n13161), .b(n13141), .o(n14051) );
na02f01 g10263 ( .a(n14051), .b(n14050), .o(n14052) );
no02f01 g10264 ( .a(n14051), .b(n14050), .o(n14053) );
in01f01 g10265 ( .a(n14053), .o(n14054) );
na02f01 g10266 ( .a(n14054), .b(n14052), .o(n14055) );
no03f01 g10267 ( .a(n13779), .b(n13778), .c(n13845), .o(n14056) );
ao12f01 g10268 ( .a(n13865), .b(n13866), .c(n13693), .o(n14057) );
no02f01 g10269 ( .a(n14057), .b(n14056), .o(n14058) );
in01f01 g10270 ( .a(n14058), .o(n14059) );
no02f01 g10271 ( .a(n14059), .b(n14055), .o(n14060) );
in01f01 g10272 ( .a(n14060), .o(n14061) );
in01f01 g10273 ( .a(n13124), .o(n14062) );
no02f01 g10274 ( .a(n13162), .b(n13131), .o(n14063) );
no02f01 g10275 ( .a(n14063), .b(n14062), .o(n14064) );
na02f01 g10276 ( .a(n14063), .b(n14062), .o(n14065) );
in01f01 g10277 ( .a(n14065), .o(n14066) );
no02f01 g10278 ( .a(n14066), .b(n14064), .o(n14067) );
no03f01 g10279 ( .a(n13777), .b(n13864), .c(n13698), .o(n14068) );
ao12f01 g10280 ( .a(n13775), .b(n13776), .c(n13699), .o(n14069) );
no02f01 g10281 ( .a(n14069), .b(n14068), .o(n14070) );
no02f01 g10282 ( .a(n14070), .b(n14067), .o(n14071) );
in01f01 g10283 ( .a(n14071), .o(n14072) );
in01f01 g10284 ( .a(n13086), .o(n14073) );
ao12f01 g10285 ( .a(n13108), .b(n14073), .c(n13080), .o(n14074) );
in01f01 g10286 ( .a(n14074), .o(n14075) );
no02f01 g10287 ( .a(n13109), .b(n13093), .o(n14076) );
in01f01 g10288 ( .a(n14076), .o(n14077) );
no02f01 g10289 ( .a(n14077), .b(n14075), .o(n14078) );
no02f01 g10290 ( .a(n14076), .b(n14074), .o(n14079) );
no02f01 g10291 ( .a(n14079), .b(n14078), .o(n14080) );
in01f01 g10292 ( .a(n14080), .o(n14081) );
no02f01 g10293 ( .a(n13860), .b(n13713), .o(n14082) );
no02f01 g10294 ( .a(n14082), .b(n13859), .o(n14083) );
na02f01 g10295 ( .a(n14082), .b(n13859), .o(n14084) );
in01f01 g10296 ( .a(n14084), .o(n14085) );
no02f01 g10297 ( .a(n14085), .b(n14083), .o(n14086) );
in01f01 g10298 ( .a(n14086), .o(n14087) );
no02f01 g10299 ( .a(n14087), .b(n14081), .o(n14088) );
in01f01 g10300 ( .a(n13080), .o(n14089) );
no02f01 g10301 ( .a(n13108), .b(n13086), .o(n14090) );
no02f01 g10302 ( .a(n14090), .b(n14089), .o(n14091) );
na02f01 g10303 ( .a(n14090), .b(n14089), .o(n14092) );
in01f01 g10304 ( .a(n14092), .o(n14093) );
no02f01 g10305 ( .a(n14093), .b(n14091), .o(n14094) );
no02f01 g10306 ( .a(n13766), .b(n13763), .o(n14095) );
no02f01 g10307 ( .a(n14095), .b(n13758), .o(n14096) );
na02f01 g10308 ( .a(n14095), .b(n13758), .o(n14097) );
in01f01 g10309 ( .a(n14097), .o(n14098) );
no02f01 g10310 ( .a(n14098), .b(n14096), .o(n14099) );
no02f01 g10311 ( .a(n14099), .b(n14094), .o(n14100) );
no02f01 g10312 ( .a(n13077), .b(n13076), .o(n14101) );
in01f01 g10313 ( .a(n13078), .o(n14102) );
na02f01 g10314 ( .a(n14102), .b(n13067), .o(n14103) );
in01f01 g10315 ( .a(n14103), .o(n14104) );
no02f01 g10316 ( .a(n14104), .b(n14101), .o(n14105) );
in01f01 g10317 ( .a(n14105), .o(n14106) );
na02f01 g10318 ( .a(n14104), .b(n14101), .o(n14107) );
na02f01 g10319 ( .a(n14107), .b(n14106), .o(n14108) );
no02f01 g10320 ( .a(n13756), .b(n13725), .o(n14109) );
no02f01 g10321 ( .a(n14109), .b(n13856), .o(n14110) );
na02f01 g10322 ( .a(n14109), .b(n13856), .o(n14111) );
in01f01 g10323 ( .a(n14111), .o(n14112) );
no02f01 g10324 ( .a(n14112), .b(n14110), .o(n14113) );
in01f01 g10325 ( .a(n14113), .o(n14114) );
no02f01 g10326 ( .a(n14114), .b(n14108), .o(n14115) );
na02f01 g10327 ( .a(n14102), .b(n13066), .o(n14116) );
no02f01 g10328 ( .a(n14116), .b(n13055), .o(n14117) );
na02f01 g10329 ( .a(n14116), .b(n13055), .o(n14118) );
in01f01 g10330 ( .a(n14118), .o(n14119) );
no02f01 g10331 ( .a(n14119), .b(n14117), .o(n14120) );
no02f01 g10332 ( .a(n13738), .b(n13737), .o(n14121) );
no02f01 g10333 ( .a(n13854), .b(n13748), .o(n14122) );
no02f01 g10334 ( .a(n13753), .b(n13747), .o(n14123) );
no02f01 g10335 ( .a(n14123), .b(n14122), .o(n14124) );
no02f01 g10336 ( .a(n14124), .b(n14121), .o(n14125) );
na02f01 g10337 ( .a(n14124), .b(n14121), .o(n14126) );
in01f01 g10338 ( .a(n14126), .o(n14127) );
no02f01 g10339 ( .a(n14127), .b(n14125), .o(n14128) );
no02f01 g10340 ( .a(n14128), .b(n14120), .o(n14129) );
na02f01 g10341 ( .a(n14128), .b(n14120), .o(n14130) );
na03f01 g10342 ( .a(n13053), .b(n13047), .c(n11514), .o(n14131) );
oa12f01 g10343 ( .a(n13054), .b(n13046), .c(n11515), .o(n14132) );
na02f01 g10344 ( .a(n14132), .b(n14131), .o(n14133) );
no03f01 g10345 ( .a(n13735), .b(n13850), .c(n13849), .o(n14134) );
ao12f01 g10346 ( .a(n13736), .b(n13727), .c(n13726), .o(n14135) );
no02f01 g10347 ( .a(n14135), .b(n14134), .o(n14136) );
no02f01 g10348 ( .a(n14136), .b(n13733), .o(n14137) );
na02f01 g10349 ( .a(n14136), .b(n13733), .o(n14138) );
in01f01 g10350 ( .a(n14138), .o(n14139) );
no02f01 g10351 ( .a(n14139), .b(n14137), .o(n14140) );
in01f01 g10352 ( .a(n14140), .o(n14141) );
no02f01 g10353 ( .a(n14141), .b(n14133), .o(n14142) );
no02f01 g10354 ( .a(n13047), .b(n11515), .o(n14143) );
no02f01 g10355 ( .a(n13047), .b(n11514), .o(n14144) );
no02f01 g10356 ( .a(n14144), .b(n14143), .o(n14145) );
no02f01 g10357 ( .a(n13731), .b(n12877), .o(n14146) );
no02f01 g10358 ( .a(n13730), .b(n12876), .o(n14147) );
no02f01 g10359 ( .a(n14147), .b(n14146), .o(n14148) );
in01f01 g10360 ( .a(n14148), .o(n14149) );
na02f01 g10361 ( .a(n14149), .b(n14145), .o(n14150) );
na02f01 g10362 ( .a(n14141), .b(n14133), .o(n14151) );
oa12f01 g10363 ( .a(n14151), .b(n14150), .c(n14142), .o(n14152) );
ao12f01 g10364 ( .a(n14129), .b(n14152), .c(n14130), .o(n14153) );
na02f01 g10365 ( .a(n14114), .b(n14108), .o(n14154) );
ao12f01 g10366 ( .a(n14115), .b(n14154), .c(n14153), .o(n14155) );
na02f01 g10367 ( .a(n14099), .b(n14094), .o(n14156) );
ao12f01 g10368 ( .a(n14100), .b(n14156), .c(n14155), .o(n14157) );
no02f01 g10369 ( .a(n14086), .b(n14080), .o(n14158) );
in01f01 g10370 ( .a(n14158), .o(n14159) );
ao12f01 g10371 ( .a(n14088), .b(n14159), .c(n14157), .o(n14160) );
in01f01 g10372 ( .a(n13110), .o(n14161) );
no02f01 g10373 ( .a(n14161), .b(n13096), .o(n14162) );
no02f01 g10374 ( .a(n13111), .b(n13106), .o(n14163) );
na02f01 g10375 ( .a(n14163), .b(n14162), .o(n14164) );
no02f01 g10376 ( .a(n14163), .b(n14162), .o(n14165) );
in01f01 g10377 ( .a(n14165), .o(n14166) );
na02f01 g10378 ( .a(n14166), .b(n14164), .o(n14167) );
no02f01 g10379 ( .a(n13771), .b(n13847), .o(n14168) );
no02f01 g10380 ( .a(n14168), .b(n13770), .o(n14169) );
na02f01 g10381 ( .a(n14168), .b(n13770), .o(n14170) );
in01f01 g10382 ( .a(n14170), .o(n14171) );
no02f01 g10383 ( .a(n14171), .b(n14169), .o(n14172) );
in01f01 g10384 ( .a(n14172), .o(n14173) );
no02f01 g10385 ( .a(n14173), .b(n14167), .o(n14174) );
in01f01 g10386 ( .a(n14174), .o(n14175) );
in01f01 g10387 ( .a(n13123), .o(n14176) );
na02f01 g10388 ( .a(n14176), .b(n13119), .o(n14177) );
ao12f01 g10389 ( .a(n13111), .b(n14161), .c(n13107), .o(n14178) );
oa12f01 g10390 ( .a(n14178), .b(n13106), .c(n13095), .o(n14179) );
na02f01 g10391 ( .a(n14179), .b(n14177), .o(n14180) );
in01f01 g10392 ( .a(n14177), .o(n14181) );
in01f01 g10393 ( .a(n14179), .o(n14182) );
na02f01 g10394 ( .a(n14182), .b(n14181), .o(n14183) );
na02f01 g10395 ( .a(n14183), .b(n14180), .o(n14184) );
no03f01 g10396 ( .a(n13773), .b(n13772), .c(n13704), .o(n14185) );
ao12f01 g10397 ( .a(n13863), .b(n13774), .c(n13846), .o(n14186) );
no02f01 g10398 ( .a(n14186), .b(n14185), .o(n14187) );
in01f01 g10399 ( .a(n14187), .o(n14188) );
na02f01 g10400 ( .a(n14188), .b(n14184), .o(n14189) );
ao12f01 g10401 ( .a(n14172), .b(n14166), .c(n14164), .o(n14190) );
in01f01 g10402 ( .a(n14190), .o(n14191) );
na02f01 g10403 ( .a(n14191), .b(n14189), .o(n14192) );
ao12f01 g10404 ( .a(n14192), .b(n14175), .c(n14160), .o(n14193) );
no02f01 g10405 ( .a(n14188), .b(n14184), .o(n14194) );
no02f01 g10406 ( .a(n14194), .b(n14193), .o(n14195) );
in01f01 g10407 ( .a(n14070), .o(n14196) );
no03f01 g10408 ( .a(n14196), .b(n14066), .c(n14064), .o(n14197) );
in01f01 g10409 ( .a(n14197), .o(n14198) );
na02f01 g10410 ( .a(n14198), .b(n14195), .o(n14199) );
na02f01 g10411 ( .a(n14059), .b(n14055), .o(n14200) );
na03f01 g10412 ( .a(n14200), .b(n14199), .c(n14072), .o(n14201) );
in01f01 g10413 ( .a(n14047), .o(n14202) );
no03f01 g10414 ( .a(n14202), .b(n14043), .c(n14041), .o(n14203) );
in01f01 g10415 ( .a(n14203), .o(n14204) );
na03f01 g10416 ( .a(n14204), .b(n14201), .c(n14061), .o(n14205) );
no02f01 g10417 ( .a(n14033), .b(n14029), .o(n14206) );
in01f01 g10418 ( .a(n14206), .o(n14207) );
na03f01 g10419 ( .a(n14207), .b(n14205), .c(n14049), .o(n14208) );
na02f01 g10420 ( .a(n14019), .b(n14014), .o(n14209) );
na03f01 g10421 ( .a(n14209), .b(n14208), .c(n14036), .o(n14210) );
no02f01 g10422 ( .a(n14004), .b(n13994), .o(n14211) );
in01f01 g10423 ( .a(n14211), .o(n14212) );
na03f01 g10424 ( .a(n14212), .b(n14210), .c(n14021), .o(n14213) );
no02f01 g10425 ( .a(n13199), .b(n13970), .o(n14214) );
no02f01 g10426 ( .a(n14214), .b(n13972), .o(n14215) );
na02f01 g10427 ( .a(n14214), .b(n13972), .o(n14216) );
in01f01 g10428 ( .a(n14216), .o(n14217) );
no02f01 g10429 ( .a(n14217), .b(n14215), .o(n14218) );
in01f01 g10430 ( .a(n14218), .o(n14219) );
no02f01 g10431 ( .a(n13813), .b(n13804), .o(n14220) );
na02f01 g10432 ( .a(n14220), .b(n13795), .o(n14221) );
in01f01 g10433 ( .a(n14221), .o(n14222) );
no02f01 g10434 ( .a(n14220), .b(n13795), .o(n14223) );
no02f01 g10435 ( .a(n14223), .b(n14222), .o(n14224) );
in01f01 g10436 ( .a(n14224), .o(n14225) );
no02f01 g10437 ( .a(n14225), .b(n14219), .o(n14226) );
in01f01 g10438 ( .a(n14226), .o(n14227) );
na03f01 g10439 ( .a(n14227), .b(n14213), .c(n14007), .o(n14228) );
no02f01 g10440 ( .a(n13984), .b(n13977), .o(n14229) );
no02f01 g10441 ( .a(n14224), .b(n14218), .o(n14230) );
no02f01 g10442 ( .a(n14230), .b(n14229), .o(n14231) );
ao12f01 g10443 ( .a(n13986), .b(n14231), .c(n14228), .o(n14232) );
in01f01 g10444 ( .a(n13952), .o(n14233) );
in01f01 g10445 ( .a(n13959), .o(n14234) );
no02f01 g10446 ( .a(n14234), .b(n14233), .o(n14235) );
in01f01 g10447 ( .a(n14235), .o(n14236) );
in01f01 g10448 ( .a(n13963), .o(n14237) );
no02f01 g10449 ( .a(n14237), .b(n13908), .o(n14238) );
na04f01 g10450 ( .a(n14238), .b(n14236), .c(n14232), .d(n13966), .o(n14239) );
in01f01 g10451 ( .a(n14239), .o(n14240) );
ao12f01 g10452 ( .a(n14240), .b(n13965), .c(n13909), .o(n14241) );
in01f01 g10453 ( .a(n14241), .o(n14242) );
in01f01 g10454 ( .a(n13590), .o(n14243) );
no02f01 g10455 ( .a(n13887), .b(n13886), .o(n14244) );
no02f01 g10456 ( .a(n13841), .b(n13829), .o(n14245) );
no02f01 g10457 ( .a(n14245), .b(n14244), .o(n14246) );
na03f01 g10458 ( .a(n14246), .b(n13591), .c(n14243), .o(n14247) );
ao12f01 g10459 ( .a(n13891), .b(n14247), .c(n14242), .o(n14248) );
na02f01 g10460 ( .a(n13584), .b(n13582), .o(n14249) );
in01f01 g10461 ( .a(n13585), .o(n14250) );
na02f01 g10462 ( .a(n14250), .b(n14249), .o(n14251) );
na02f01 g10463 ( .a(n14251), .b(n11515), .o(n14252) );
oa22f01 g10464 ( .a(n13586), .b(n11515), .c(n13527), .d(n13511), .o(n14253) );
na02f01 g10465 ( .a(n14253), .b(n14252), .o(n14254) );
oa12f01 g10466 ( .a(n13575), .b(n13583), .c(n13495), .o(n14255) );
na02f01 g10467 ( .a(n14255), .b(n13572), .o(n14256) );
no02f01 g10468 ( .a(n13548), .b(n13465), .o(n14257) );
na02f01 g10469 ( .a(n13540), .b(n13544), .o(n14258) );
no02f01 g10470 ( .a(n13531), .b(delay_add_ln22_unr2_stage2_stallmux_q_30_), .o(n14259) );
na02f01 g10471 ( .a(n13531), .b(delay_add_ln22_unr2_stage2_stallmux_q_30_), .o(n14260) );
in01f01 g10472 ( .a(n14260), .o(n14261) );
no02f01 g10473 ( .a(n14261), .b(n14259), .o(n14262) );
no04f01 g10474 ( .a(n13534), .b(n13455), .c(n13442), .d(n13369), .o(n14263) );
no02f01 g10475 ( .a(n13532), .b(n13457), .o(n14264) );
in01f01 g10476 ( .a(n14264), .o(n14265) );
oa12f01 g10477 ( .a(n14262), .b(n14265), .c(n14263), .o(n14266) );
in01f01 g10478 ( .a(n14266), .o(n14267) );
no03f01 g10479 ( .a(n14265), .b(n14263), .c(n14262), .o(n14268) );
no02f01 g10480 ( .a(n14268), .b(n14267), .o(n14269) );
no02f01 g10481 ( .a(n14269), .b(n11179), .o(n14270) );
no02f01 g10482 ( .a(n14269), .b(n11158), .o(n14271) );
no02f01 g10483 ( .a(n14271), .b(n14270), .o(n14272) );
in01f01 g10484 ( .a(n14272), .o(n14273) );
na03f01 g10485 ( .a(n14273), .b(n14258), .c(n14257), .o(n14274) );
na02f01 g10486 ( .a(n13541), .b(n13464), .o(n14275) );
no02f01 g10487 ( .a(n13547), .b(n13529), .o(n14276) );
oa12f01 g10488 ( .a(n14272), .b(n14276), .c(n14275), .o(n14277) );
ao12f01 g10489 ( .a(n13562), .b(n13563), .c(n13568), .o(n14278) );
no02f01 g10490 ( .a(n13554), .b(n13553), .o(n14279) );
no02f01 g10491 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_26_), .b(n11021), .o(n14280) );
in01f01 g10492 ( .a(n14280), .o(n14281) );
na02f01 g10493 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_26_), .b(n11021), .o(n14282) );
na02f01 g10494 ( .a(n14282), .b(n14281), .o(n14283) );
no02f01 g10495 ( .a(n14283), .b(n14279), .o(n14284) );
na02f01 g10496 ( .a(n14283), .b(n14279), .o(n14285) );
in01f01 g10497 ( .a(n14285), .o(n14286) );
no02f01 g10498 ( .a(n14286), .b(n14284), .o(n14287) );
no02f01 g10499 ( .a(n14287), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_26_), .o(n14288) );
na02f01 g10500 ( .a(n14287), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_26_), .o(n14289) );
in01f01 g10501 ( .a(n14289), .o(n14290) );
no02f01 g10502 ( .a(n14290), .b(n14288), .o(n14291) );
in01f01 g10503 ( .a(n14291), .o(n14292) );
no02f01 g10504 ( .a(n14292), .b(n14278), .o(n14293) );
in01f01 g10505 ( .a(n14278), .o(n14294) );
no02f01 g10506 ( .a(n14291), .b(n14294), .o(n14295) );
no02f01 g10507 ( .a(n14295), .b(n14293), .o(n14296) );
in01f01 g10508 ( .a(n14296), .o(n14297) );
na03f01 g10509 ( .a(n14297), .b(n14277), .c(n14274), .o(n14298) );
no03f01 g10510 ( .a(n14272), .b(n14276), .c(n14275), .o(n14299) );
ao12f01 g10511 ( .a(n14273), .b(n14258), .c(n14257), .o(n14300) );
oa12f01 g10512 ( .a(n14296), .b(n14300), .c(n14299), .o(n14301) );
na02f01 g10513 ( .a(n14301), .b(n14298), .o(n14302) );
no02f01 g10514 ( .a(n14302), .b(n14256), .o(n14303) );
no03f01 g10515 ( .a(n14296), .b(n14300), .c(n14299), .o(n14304) );
ao12f01 g10516 ( .a(n14297), .b(n14277), .c(n14274), .o(n14305) );
no02f01 g10517 ( .a(n14305), .b(n14304), .o(n14306) );
ao12f01 g10518 ( .a(n14306), .b(n14255), .c(n13572), .o(n14307) );
no02f01 g10519 ( .a(n14307), .b(n14303), .o(n14308) );
no02f01 g10520 ( .a(n14308), .b(n11515), .o(n14309) );
no02f01 g10521 ( .a(n14308), .b(n11514), .o(n14310) );
oa12f01 g10522 ( .a(n14254), .b(n14310), .c(n14309), .o(n14311) );
no03f01 g10523 ( .a(n14310), .b(n14309), .c(n14254), .o(n14312) );
in01f01 g10524 ( .a(n14312), .o(n14313) );
ao12f01 g10525 ( .a(n13840), .b(n13885), .c(n13843), .o(n14314) );
no02f01 g10526 ( .a(n14314), .b(n13838), .o(n14315) );
no02f01 g10527 ( .a(n13494), .b(n11179), .o(n14316) );
no02f01 g10528 ( .a(n13494), .b(n11158), .o(n14317) );
no02f01 g10529 ( .a(n14317), .b(n13832), .o(n14318) );
oa12f01 g10530 ( .a(n14318), .b(n14316), .c(n13830), .o(n14319) );
no02f01 g10531 ( .a(n14319), .b(n13571), .o(n14320) );
na02f01 g10532 ( .a(n14319), .b(n13571), .o(n14321) );
in01f01 g10533 ( .a(n14321), .o(n14322) );
no02f01 g10534 ( .a(n14322), .b(n14320), .o(n14323) );
na02f01 g10535 ( .a(n14323), .b(n12254), .o(n14324) );
in01f01 g10536 ( .a(n14324), .o(n14325) );
no02f01 g10537 ( .a(n14323), .b(n12254), .o(n14326) );
no02f01 g10538 ( .a(n14326), .b(n14325), .o(n14327) );
no02f01 g10539 ( .a(n14327), .b(n14315), .o(n14328) );
na02f01 g10540 ( .a(n14327), .b(n14315), .o(n14329) );
in01f01 g10541 ( .a(n14329), .o(n14330) );
no02f01 g10542 ( .a(n14330), .b(n14328), .o(n14331) );
ao12f01 g10543 ( .a(n14331), .b(n14313), .c(n14311), .o(n14332) );
in01f01 g10544 ( .a(n14311), .o(n14333) );
in01f01 g10545 ( .a(n14328), .o(n14334) );
na02f01 g10546 ( .a(n14329), .b(n14334), .o(n14335) );
no03f01 g10547 ( .a(n14335), .b(n14312), .c(n14333), .o(n14336) );
no02f01 g10548 ( .a(n14336), .b(n14332), .o(n14337) );
no02f01 g10549 ( .a(n14337), .b(n14248), .o(n14338) );
na02f01 g10550 ( .a(n14337), .b(n14248), .o(n14339) );
in01f01 g10551 ( .a(n14339), .o(n14340) );
no02f01 g10552 ( .a(n14340), .b(n14338), .o(n14341) );
in01f01 g10553 ( .a(n14341), .o(n3747) );
na02f01 g10554 ( .a(n3747), .b(n4116), .o(n14343) );
in01f01 g10555 ( .a(n11526), .o(n14344) );
na02f01 g10556 ( .a(n11868), .b(n11861), .o(n14345) );
na02f01 g10557 ( .a(n14345), .b(n14344), .o(n2589) );
na02f01 g10558 ( .a(n14341), .b(n2589), .o(n14347) );
na02f01 g10559 ( .a(n14347), .b(n14343), .o(n253) );
no02f01 g10560 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_7_), .b(delay_sub_ln22_unr24_stage9_stallmux_q_7_), .o(n14349) );
in01f01 g10561 ( .a(n14349), .o(n14350) );
no02f01 g10562 ( .a(delay_sub_ln22_unr24_stage9_stallmux_q_5_), .b(delay_add_ln22_unr23_stage9_stallmux_q_5_), .o(n14351) );
na02f01 g10563 ( .a(delay_sub_ln22_unr24_stage9_stallmux_q_4_), .b(delay_add_ln22_unr23_stage9_stallmux_q_4_), .o(n14352) );
in01f01 g10564 ( .a(n14352), .o(n14353) );
na02f01 g10565 ( .a(delay_sub_ln22_unr24_stage9_stallmux_q_5_), .b(delay_add_ln22_unr23_stage9_stallmux_q_5_), .o(n14354) );
in01f01 g10566 ( .a(n14354), .o(n14355) );
no02f01 g10567 ( .a(n14355), .b(n14353), .o(n14356) );
no02f01 g10568 ( .a(n14356), .b(n14351), .o(n14357) );
na02f01 g10569 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_3_), .b(delay_sub_ln22_unr24_stage9_stallmux_q_3_), .o(n14358) );
in01f01 g10570 ( .a(delay_sub_ln22_unr24_stage9_stallmux_q_2_), .o(n14359) );
in01f01 g10571 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_2_), .o(n14360) );
no02f01 g10572 ( .a(n14360), .b(n14359), .o(n14361) );
no02f01 g10573 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_2_), .b(delay_sub_ln22_unr24_stage9_stallmux_q_2_), .o(n14362) );
in01f01 g10574 ( .a(n14362), .o(n14363) );
na02f01 g10575 ( .a(delay_sub_ln22_unr24_stage9_stallmux_q_1_), .b(delay_add_ln22_unr23_stage9_stallmux_q_1_), .o(n14364) );
no02f01 g10576 ( .a(delay_sub_ln22_unr24_stage9_stallmux_q_1_), .b(delay_add_ln22_unr23_stage9_stallmux_q_1_), .o(n14365) );
na02f01 g10577 ( .a(delay_sub_ln22_unr24_stage9_stallmux_q_0_), .b(delay_add_ln22_unr23_stage9_stallmux_q_0_), .o(n14366) );
oa12f01 g10578 ( .a(n14364), .b(n14366), .c(n14365), .o(n14367) );
ao12f01 g10579 ( .a(n14361), .b(n14367), .c(n14363), .o(n14368) );
no02f01 g10580 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_3_), .b(delay_sub_ln22_unr24_stage9_stallmux_q_3_), .o(n14369) );
oa12f01 g10581 ( .a(n14358), .b(n14369), .c(n14368), .o(n14370) );
no02f01 g10582 ( .a(delay_sub_ln22_unr24_stage9_stallmux_q_4_), .b(delay_add_ln22_unr23_stage9_stallmux_q_4_), .o(n14371) );
no02f01 g10583 ( .a(n14371), .b(n14351), .o(n14372) );
ao12f01 g10584 ( .a(n14357), .b(n14372), .c(n14370), .o(n14373) );
no02f01 g10585 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_6_), .b(delay_sub_ln22_unr24_stage9_stallmux_q_6_), .o(n14374) );
no02f01 g10586 ( .a(n14374), .b(n14373), .o(n14375) );
na02f01 g10587 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_6_), .b(delay_sub_ln22_unr24_stage9_stallmux_q_6_), .o(n14376) );
in01f01 g10588 ( .a(n14376), .o(n14377) );
na02f01 g10589 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_7_), .b(delay_sub_ln22_unr24_stage9_stallmux_q_7_), .o(n14378) );
in01f01 g10590 ( .a(n14378), .o(n14379) );
no02f01 g10591 ( .a(n14379), .b(n14377), .o(n14380) );
in01f01 g10592 ( .a(n14380), .o(n14381) );
oa12f01 g10593 ( .a(n14350), .b(n14381), .c(n14375), .o(n14382) );
ao12f01 g10594 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_9_), .c(delay_add_ln22_unr23_stage9_stallmux_q_8_), .o(n14383) );
no02f01 g10595 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_10_), .b(n_46254), .o(n14384) );
no02f01 g10596 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_11_), .o(n14385) );
no03f01 g10597 ( .a(n14385), .b(n14384), .c(n14383), .o(n14386) );
in01f01 g10598 ( .a(n14386), .o(n14387) );
no02f01 g10599 ( .a(n14387), .b(n14382), .o(n14388) );
no02f01 g10600 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_13_), .o(n14389) );
no02f01 g10601 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_12_), .o(n14390) );
no02f01 g10602 ( .a(n14390), .b(n14389), .o(n14391) );
in01f01 g10603 ( .a(n14391), .o(n14392) );
no02f01 g10604 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_14_), .b(n_46254), .o(n14393) );
no02f01 g10605 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_15_), .b(n_46254), .o(n14394) );
no03f01 g10606 ( .a(n14394), .b(n14393), .c(n14392), .o(n14395) );
in01f01 g10607 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_11_), .o(n14396) );
in01f01 g10608 ( .a(n_46254), .o(n14397) );
in01f01 g10609 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_10_), .o(n14398) );
ao12f01 g10610 ( .a(n14397), .b(n14398), .c(n14396), .o(n14399) );
in01f01 g10611 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_8_), .o(n14400) );
in01f01 g10612 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_9_), .o(n14401) );
ao12f01 g10613 ( .a(n14397), .b(n14401), .c(n14400), .o(n14402) );
no02f01 g10614 ( .a(n14402), .b(n14399), .o(n14403) );
in01f01 g10615 ( .a(n14403), .o(n14404) );
in01f01 g10616 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_12_), .o(n14405) );
in01f01 g10617 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_13_), .o(n14406) );
ao12f01 g10618 ( .a(n14397), .b(n14406), .c(n14405), .o(n14407) );
no02f01 g10619 ( .a(n14407), .b(n14404), .o(n14408) );
in01f01 g10620 ( .a(n14408), .o(n14409) );
in01f01 g10621 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_15_), .o(n14410) );
in01f01 g10622 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_14_), .o(n14411) );
ao12f01 g10623 ( .a(n14397), .b(n14411), .c(n14410), .o(n14412) );
no02f01 g10624 ( .a(n14412), .b(n14409), .o(n14413) );
in01f01 g10625 ( .a(n14413), .o(n14414) );
ao12f01 g10626 ( .a(n14414), .b(n14395), .c(n14388), .o(n14415) );
ao12f01 g10627 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_17_), .c(delay_add_ln22_unr23_stage9_stallmux_q_16_), .o(n14416) );
no02f01 g10628 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_18_), .o(n14417) );
no02f01 g10629 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_19_), .o(n14418) );
no03f01 g10630 ( .a(n14418), .b(n14417), .c(n14416), .o(n14419) );
in01f01 g10631 ( .a(n14419), .o(n14420) );
no02f01 g10632 ( .a(n14420), .b(n14415), .o(n14421) );
no02f01 g10633 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_21_), .o(n14422) );
no02f01 g10634 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_20_), .o(n14423) );
no02f01 g10635 ( .a(n14423), .b(n14422), .o(n14424) );
in01f01 g10636 ( .a(n14424), .o(n14425) );
no02f01 g10637 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_23_), .o(n14426) );
no02f01 g10638 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_22_), .o(n14427) );
no03f01 g10639 ( .a(n14427), .b(n14426), .c(n14425), .o(n14428) );
na02f01 g10640 ( .a(n14428), .b(n14421), .o(n14429) );
in01f01 g10641 ( .a(n14429), .o(n14430) );
no02f01 g10642 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_25_), .b(n_46254), .o(n14431) );
no02f01 g10643 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_24_), .o(n14432) );
no02f01 g10644 ( .a(n14432), .b(n14431), .o(n14433) );
in01f01 g10645 ( .a(n14433), .o(n14434) );
no02f01 g10646 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_27_), .o(n14435) );
no02f01 g10647 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_26_), .o(n14436) );
no03f01 g10648 ( .a(n14436), .b(n14435), .c(n14434), .o(n14437) );
na02f01 g10649 ( .a(n14437), .b(n14430), .o(n14438) );
no02f01 g10650 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_28_), .o(n14439) );
no02f01 g10651 ( .a(n14439), .b(n14438), .o(n14440) );
in01f01 g10652 ( .a(n14440), .o(n14441) );
no02f01 g10653 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_29_), .o(n14442) );
no02f01 g10654 ( .a(n14442), .b(n14441), .o(n14443) );
in01f01 g10655 ( .a(n14443), .o(n14444) );
no02f01 g10656 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_30_), .o(n14445) );
in01f01 g10657 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_16_), .o(n14446) );
in01f01 g10658 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_17_), .o(n14447) );
ao12f01 g10659 ( .a(n14397), .b(n14447), .c(n14446), .o(n14448) );
in01f01 g10660 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_19_), .o(n14449) );
in01f01 g10661 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_18_), .o(n14450) );
ao12f01 g10662 ( .a(n14397), .b(n14450), .c(n14449), .o(n14451) );
no02f01 g10663 ( .a(n14451), .b(n14448), .o(n14452) );
in01f01 g10664 ( .a(n14452), .o(n14453) );
in01f01 g10665 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_21_), .o(n14454) );
in01f01 g10666 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_20_), .o(n14455) );
ao12f01 g10667 ( .a(n14397), .b(n14455), .c(n14454), .o(n14456) );
no02f01 g10668 ( .a(n14456), .b(n14453), .o(n14457) );
in01f01 g10669 ( .a(n14457), .o(n14458) );
in01f01 g10670 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_23_), .o(n14459) );
in01f01 g10671 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_22_), .o(n14460) );
ao12f01 g10672 ( .a(n14397), .b(n14460), .c(n14459), .o(n14461) );
no02f01 g10673 ( .a(n14461), .b(n14458), .o(n14462) );
in01f01 g10674 ( .a(n14462), .o(n14463) );
in01f01 g10675 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_24_), .o(n14464) );
in01f01 g10676 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_25_), .o(n14465) );
ao12f01 g10677 ( .a(n14397), .b(n14465), .c(n14464), .o(n14466) );
no02f01 g10678 ( .a(n14466), .b(n14463), .o(n14467) );
in01f01 g10679 ( .a(n14467), .o(n14468) );
in01f01 g10680 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_26_), .o(n14469) );
in01f01 g10681 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_27_), .o(n14470) );
ao12f01 g10682 ( .a(n14397), .b(n14470), .c(n14469), .o(n14471) );
no02f01 g10683 ( .a(n14471), .b(n14468), .o(n14472) );
in01f01 g10684 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_28_), .o(n14473) );
no02f01 g10685 ( .a(n14397), .b(n14473), .o(n14474) );
in01f01 g10686 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_29_), .o(n14475) );
no02f01 g10687 ( .a(n14397), .b(n14475), .o(n14476) );
no02f01 g10688 ( .a(n14476), .b(n14474), .o(n14477) );
na02f01 g10689 ( .a(n14477), .b(n14472), .o(n14478) );
na02f01 g10690 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_30_), .o(n14479) );
in01f01 g10691 ( .a(n14479), .o(n14480) );
no02f01 g10692 ( .a(n14480), .b(n14478), .o(n14481) );
oa12f01 g10693 ( .a(n14481), .b(n14445), .c(n14444), .o(n14482) );
in01f01 g10694 ( .a(n14482), .o(n14483) );
no02f01 g10695 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_31_), .o(n14484) );
na02f01 g10696 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_31_), .o(n14485) );
in01f01 g10697 ( .a(n14485), .o(n14486) );
no02f01 g10698 ( .a(n14486), .b(n14484), .o(n14487) );
no02f01 g10699 ( .a(n14487), .b(n14483), .o(n14488) );
na02f01 g10700 ( .a(n14487), .b(n14483), .o(n14489) );
in01f01 g10701 ( .a(n14489), .o(n14490) );
no02f01 g10702 ( .a(n14490), .b(n14488), .o(n14491) );
in01f01 g10703 ( .a(delay_sub_ln23_0_unr24_stage9_stallmux_q), .o(n14492) );
no02f01 g10704 ( .a(n14491), .b(n14492), .o(n14493) );
in01f01 g10705 ( .a(n14472), .o(n14494) );
no03f01 g10706 ( .a(n14474), .b(n14494), .c(n14440), .o(n14495) );
no02f01 g10707 ( .a(n14476), .b(n14442), .o(n14496) );
no02f01 g10708 ( .a(n14496), .b(n14495), .o(n14497) );
na02f01 g10709 ( .a(n14496), .b(n14495), .o(n14498) );
in01f01 g10710 ( .a(n14498), .o(n14499) );
no02f01 g10711 ( .a(n14499), .b(n14497), .o(n14500) );
no02f01 g10712 ( .a(n14500), .b(n14492), .o(n14501) );
na02f01 g10713 ( .a(n14472), .b(n14438), .o(n14502) );
in01f01 g10714 ( .a(n14502), .o(n14503) );
no02f01 g10715 ( .a(n14474), .b(n14439), .o(n14504) );
no02f01 g10716 ( .a(n14504), .b(n14503), .o(n14505) );
na02f01 g10717 ( .a(n14504), .b(n14503), .o(n14506) );
in01f01 g10718 ( .a(n14506), .o(n14507) );
no02f01 g10719 ( .a(n14507), .b(n14505), .o(n14508) );
no02f01 g10720 ( .a(n14508), .b(n14492), .o(n14509) );
no02f01 g10721 ( .a(n14465), .b(n14397), .o(n14510) );
no02f01 g10722 ( .a(n14510), .b(n14431), .o(n14511) );
in01f01 g10723 ( .a(n14511), .o(n14512) );
no02f01 g10724 ( .a(n14397), .b(n14464), .o(n14513) );
no02f01 g10725 ( .a(n14513), .b(n14463), .o(n14514) );
oa12f01 g10726 ( .a(n14514), .b(n14432), .c(n14429), .o(n14515) );
no02f01 g10727 ( .a(n14515), .b(n14512), .o(n14516) );
na02f01 g10728 ( .a(n14515), .b(n14512), .o(n14517) );
in01f01 g10729 ( .a(n14517), .o(n14518) );
no02f01 g10730 ( .a(n14518), .b(n14516), .o(n14519) );
no02f01 g10731 ( .a(n14397), .b(n14469), .o(n14520) );
no02f01 g10732 ( .a(n14520), .b(n14436), .o(n14521) );
in01f01 g10733 ( .a(n14521), .o(n14522) );
no02f01 g10734 ( .a(n14434), .b(n14429), .o(n14523) );
in01f01 g10735 ( .a(n14523), .o(n14524) );
na02f01 g10736 ( .a(n14524), .b(n14467), .o(n14525) );
no02f01 g10737 ( .a(n14522), .b(n14468), .o(n14526) );
ao22f01 g10738 ( .a(n14526), .b(n14524), .c(n14525), .d(n14522), .o(n14527) );
ao12f01 g10739 ( .a(n14492), .b(n14527), .c(n14519), .o(n14528) );
in01f01 g10740 ( .a(n14528), .o(n14529) );
no02f01 g10741 ( .a(n14397), .b(n14470), .o(n14530) );
no02f01 g10742 ( .a(n14530), .b(n14435), .o(n14531) );
in01f01 g10743 ( .a(n14531), .o(n14532) );
no02f01 g10744 ( .a(n14520), .b(n14468), .o(n14533) );
oa12f01 g10745 ( .a(n14533), .b(n14524), .c(n14436), .o(n14534) );
no02f01 g10746 ( .a(n14534), .b(n14532), .o(n14535) );
na02f01 g10747 ( .a(n14534), .b(n14532), .o(n14536) );
in01f01 g10748 ( .a(n14536), .o(n14537) );
no02f01 g10749 ( .a(n14537), .b(n14535), .o(n14538) );
oa12f01 g10750 ( .a(n14529), .b(n14538), .c(n14492), .o(n14539) );
no02f01 g10751 ( .a(n14539), .b(n14509), .o(n14540) );
in01f01 g10752 ( .a(n14540), .o(n14541) );
no02f01 g10753 ( .a(n14541), .b(n14501), .o(n14542) );
in01f01 g10754 ( .a(n14542), .o(n14543) );
no02f01 g10755 ( .a(n14478), .b(n14443), .o(n14544) );
no02f01 g10756 ( .a(n14480), .b(n14445), .o(n14545) );
no02f01 g10757 ( .a(n14545), .b(n14544), .o(n14546) );
na02f01 g10758 ( .a(n14545), .b(n14544), .o(n14547) );
in01f01 g10759 ( .a(n14547), .o(n14548) );
no02f01 g10760 ( .a(n14548), .b(n14546), .o(n14549) );
no02f01 g10761 ( .a(n14549), .b(n14492), .o(n14550) );
no02f01 g10762 ( .a(n14550), .b(n14543), .o(n14551) );
ao12f01 g10763 ( .a(n14493), .b(n14551), .c(n14491), .o(n14552) );
in01f01 g10764 ( .a(n14552), .o(n14553) );
in01f01 g10765 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_31_), .o(n14554) );
no02f01 g10766 ( .a(n14554), .b(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .o(n14555) );
in01f01 g10767 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .o(n14556) );
no02f01 g10768 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_31_), .b(n14556), .o(n14557) );
no02f01 g10769 ( .a(n14557), .b(n14555), .o(n14558) );
in01f01 g10770 ( .a(n14558), .o(n14559) );
in01f01 g10771 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_7_), .o(n14560) );
no02f01 g10772 ( .a(n14560), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_7_), .o(n14561) );
in01f01 g10773 ( .a(n14561), .o(n14562) );
in01f01 g10774 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_1_), .o(n14563) );
no02f01 g10775 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_1_), .b(n14563), .o(n14564) );
in01f01 g10776 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_0_), .o(n14565) );
na02f01 g10777 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_24_), .b(n14565), .o(n14566) );
na02f01 g10778 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_1_), .b(n14563), .o(n14567) );
ao12f01 g10779 ( .a(n14564), .b(n14567), .c(n14566), .o(n14568) );
in01f01 g10780 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_2_), .o(n14569) );
no02f01 g10781 ( .a(n14569), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_2_), .o(n14570) );
no02f01 g10782 ( .a(n14570), .b(n14568), .o(n14571) );
in01f01 g10783 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_2_), .o(n14572) );
no02f01 g10784 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_2_), .b(n14572), .o(n14573) );
in01f01 g10785 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_3_), .o(n14574) );
no02f01 g10786 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_3_), .b(n14574), .o(n14575) );
no03f01 g10787 ( .a(n14575), .b(n14573), .c(n14571), .o(n14576) );
in01f01 g10788 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_5_), .o(n14577) );
no02f01 g10789 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_5_), .b(n14577), .o(n14578) );
in01f01 g10790 ( .a(n14578), .o(n14579) );
in01f01 g10791 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_6_), .o(n14580) );
na02f01 g10792 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_6_), .b(n14580), .o(n14581) );
na02f01 g10793 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_3_), .b(n14574), .o(n14582) );
in01f01 g10794 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_4_), .o(n14583) );
no02f01 g10795 ( .a(n14583), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_4_), .o(n14584) );
in01f01 g10796 ( .a(n14584), .o(n14585) );
na04f01 g10797 ( .a(n14585), .b(n14582), .c(n14581), .d(n14579), .o(n14586) );
no02f01 g10798 ( .a(n14586), .b(n14576), .o(n14587) );
na02f01 g10799 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_5_), .b(n14577), .o(n14588) );
na02f01 g10800 ( .a(n14583), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_4_), .o(n14589) );
ao12f01 g10801 ( .a(n14578), .b(n14589), .c(n14588), .o(n14590) );
na02f01 g10802 ( .a(n14590), .b(n14581), .o(n14591) );
na02f01 g10803 ( .a(n14560), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_7_), .o(n14592) );
no02f01 g10804 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_6_), .b(n14580), .o(n14593) );
in01f01 g10805 ( .a(n14593), .o(n14594) );
na03f01 g10806 ( .a(n14594), .b(n14592), .c(n14591), .o(n14595) );
oa12f01 g10807 ( .a(n14562), .b(n14595), .c(n14587), .o(n14596) );
ao12f01 g10808 ( .a(n14556), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_9_), .c(delay_sub_ln21_0_unr23_stage9_stallmux_q_8_), .o(n14597) );
no02f01 g10809 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_15_), .b(n14556), .o(n14598) );
no02f01 g10810 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_14_), .b(n14556), .o(n14599) );
no03f01 g10811 ( .a(n14599), .b(n14598), .c(n14597), .o(n14600) );
no02f01 g10812 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_12_), .b(n14556), .o(n14601) );
no02f01 g10813 ( .a(n14556), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_13_), .o(n14602) );
no02f01 g10814 ( .a(n14602), .b(n14601), .o(n14603) );
no02f01 g10815 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_11_), .b(n14556), .o(n14604) );
no02f01 g10816 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_10_), .b(n14556), .o(n14605) );
no02f01 g10817 ( .a(n14605), .b(n14604), .o(n14606) );
na03f01 g10818 ( .a(n14606), .b(n14603), .c(n14600), .o(n14607) );
in01f01 g10819 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_14_), .o(n14608) );
in01f01 g10820 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_15_), .o(n14609) );
ao12f01 g10821 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(n14609), .c(n14608), .o(n14610) );
in01f01 g10822 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_8_), .o(n14611) );
in01f01 g10823 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_9_), .o(n14612) );
ao12f01 g10824 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(n14612), .c(n14611), .o(n14613) );
in01f01 g10825 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_10_), .o(n14614) );
in01f01 g10826 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_11_), .o(n14615) );
ao12f01 g10827 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(n14615), .c(n14614), .o(n14616) );
no02f01 g10828 ( .a(n14616), .b(n14613), .o(n14617) );
in01f01 g10829 ( .a(n14617), .o(n14618) );
in01f01 g10830 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_13_), .o(n14619) );
in01f01 g10831 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_12_), .o(n14620) );
ao12f01 g10832 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(n14620), .c(n14619), .o(n14621) );
no02f01 g10833 ( .a(n14621), .b(n14618), .o(n14622) );
in01f01 g10834 ( .a(n14622), .o(n14623) );
no02f01 g10835 ( .a(n14623), .b(n14610), .o(n14624) );
oa12f01 g10836 ( .a(n14624), .b(n14607), .c(n14596), .o(n14625) );
ao12f01 g10837 ( .a(n14556), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_16_), .c(delay_sub_ln21_0_unr23_stage9_stallmux_q_17_), .o(n14626) );
in01f01 g10838 ( .a(n14626), .o(n14627) );
no02f01 g10839 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_19_), .b(n14556), .o(n14628) );
no02f01 g10840 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_18_), .b(n14556), .o(n14629) );
no02f01 g10841 ( .a(n14629), .b(n14628), .o(n14630) );
na02f01 g10842 ( .a(n14630), .b(n14627), .o(n14631) );
in01f01 g10843 ( .a(n14631), .o(n14632) );
ao12f01 g10844 ( .a(n14556), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_20_), .c(delay_sub_ln21_0_unr23_stage9_stallmux_q_21_), .o(n14633) );
in01f01 g10845 ( .a(n14633), .o(n14634) );
in01f01 g10846 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_23_), .o(n14635) );
in01f01 g10847 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_22_), .o(n14636) );
oa12f01 g10848 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(n14636), .c(n14635), .o(n14637) );
na03f01 g10849 ( .a(n14637), .b(n14634), .c(n14632), .o(n14638) );
in01f01 g10850 ( .a(n14638), .o(n14639) );
na02f01 g10851 ( .a(n14639), .b(n14625), .o(n14640) );
in01f01 g10852 ( .a(n14640), .o(n14641) );
no02f01 g10853 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_25_), .b(n14556), .o(n14642) );
no02f01 g10854 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_24_), .b(n14556), .o(n14643) );
no02f01 g10855 ( .a(n14643), .b(n14642), .o(n14644) );
no02f01 g10856 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_26_), .b(n14556), .o(n14645) );
no02f01 g10857 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_27_), .b(n14556), .o(n14646) );
no02f01 g10858 ( .a(n14646), .b(n14645), .o(n14647) );
na02f01 g10859 ( .a(n14647), .b(n14644), .o(n14648) );
no02f01 g10860 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_29_), .b(n14556), .o(n14649) );
no02f01 g10861 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_28_), .b(n14556), .o(n14650) );
no03f01 g10862 ( .a(n14650), .b(n14649), .c(n14648), .o(n14651) );
na02f01 g10863 ( .a(n14651), .b(n14641), .o(n14652) );
no02f01 g10864 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_30_), .b(n14556), .o(n14653) );
in01f01 g10865 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_18_), .o(n14654) );
in01f01 g10866 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_19_), .o(n14655) );
ao12f01 g10867 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(n14655), .c(n14654), .o(n14656) );
in01f01 g10868 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_17_), .o(n14657) );
in01f01 g10869 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_16_), .o(n14658) );
ao12f01 g10870 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(n14658), .c(n14657), .o(n14659) );
no02f01 g10871 ( .a(n14659), .b(n14656), .o(n14660) );
in01f01 g10872 ( .a(n14660), .o(n14661) );
in01f01 g10873 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_21_), .o(n14662) );
in01f01 g10874 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_20_), .o(n14663) );
ao12f01 g10875 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(n14663), .c(n14662), .o(n14664) );
no02f01 g10876 ( .a(n14664), .b(n14661), .o(n14665) );
in01f01 g10877 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_24_), .o(n14666) );
in01f01 g10878 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_25_), .o(n14667) );
ao12f01 g10879 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(n14667), .c(n14666), .o(n14668) );
ao12f01 g10880 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(n14636), .c(n14635), .o(n14669) );
in01f01 g10881 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_27_), .o(n14670) );
in01f01 g10882 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_26_), .o(n14671) );
ao12f01 g10883 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(n14671), .c(n14670), .o(n14672) );
no03f01 g10884 ( .a(n14672), .b(n14669), .c(n14668), .o(n14673) );
na02f01 g10885 ( .a(n14673), .b(n14665), .o(n14674) );
na02f01 g10886 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_28_), .b(n14556), .o(n14675) );
in01f01 g10887 ( .a(n14675), .o(n14676) );
no02f01 g10888 ( .a(n14676), .b(n14674), .o(n14677) );
in01f01 g10889 ( .a(n14677), .o(n14678) );
na02f01 g10890 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_29_), .b(n14556), .o(n14679) );
in01f01 g10891 ( .a(n14679), .o(n14680) );
no02f01 g10892 ( .a(n14680), .b(n14678), .o(n14681) );
in01f01 g10893 ( .a(n14681), .o(n14682) );
na02f01 g10894 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_30_), .b(n14556), .o(n14683) );
in01f01 g10895 ( .a(n14683), .o(n14684) );
no02f01 g10896 ( .a(n14684), .b(n14682), .o(n14685) );
oa12f01 g10897 ( .a(n14685), .b(n14653), .c(n14652), .o(n14686) );
no02f01 g10898 ( .a(n14686), .b(n14559), .o(n14687) );
na02f01 g10899 ( .a(n14686), .b(n14559), .o(n14688) );
in01f01 g10900 ( .a(n14688), .o(n14689) );
no02f01 g10901 ( .a(n14689), .b(n14687), .o(n14690) );
in01f01 g10902 ( .a(n14690), .o(n14691) );
no02f01 g10903 ( .a(n14691), .b(n14553), .o(n14692) );
no02f01 g10904 ( .a(n14690), .b(n14552), .o(n14693) );
no02f01 g10905 ( .a(n14693), .b(n14692), .o(n14694) );
in01f01 g10906 ( .a(n14694), .o(n14695) );
no02f01 g10907 ( .a(n14658), .b(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .o(n14696) );
no02f01 g10908 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_16_), .b(n14556), .o(n14697) );
in01f01 g10909 ( .a(n14697), .o(n14698) );
ao12f01 g10910 ( .a(n14696), .b(n14698), .c(n14625), .o(n14699) );
in01f01 g10911 ( .a(n14699), .o(n14700) );
no02f01 g10912 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(n14657), .o(n14701) );
no02f01 g10913 ( .a(n14556), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_17_), .o(n14702) );
no02f01 g10914 ( .a(n14702), .b(n14701), .o(n14703) );
in01f01 g10915 ( .a(n14703), .o(n14704) );
no02f01 g10916 ( .a(n14704), .b(n14700), .o(n14705) );
no02f01 g10917 ( .a(n14703), .b(n14699), .o(n14706) );
no02f01 g10918 ( .a(n14706), .b(n14705), .o(n14707) );
no02f01 g10919 ( .a(n14697), .b(n14696), .o(n14708) );
in01f01 g10920 ( .a(n14708), .o(n14709) );
no02f01 g10921 ( .a(n14709), .b(n14625), .o(n14710) );
in01f01 g10922 ( .a(n14625), .o(n14711) );
no02f01 g10923 ( .a(n14708), .b(n14711), .o(n14712) );
no02f01 g10924 ( .a(n14712), .b(n14710), .o(n14713) );
ao12f01 g10925 ( .a(n14552), .b(n14713), .c(n14707), .o(n14714) );
no02f01 g10926 ( .a(n14626), .b(n14711), .o(n14715) );
no02f01 g10927 ( .a(n14654), .b(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .o(n14716) );
no02f01 g10928 ( .a(n14716), .b(n14629), .o(n14717) );
in01f01 g10929 ( .a(n14717), .o(n14718) );
no03f01 g10930 ( .a(n14718), .b(n14715), .c(n14659), .o(n14719) );
no02f01 g10931 ( .a(n14715), .b(n14659), .o(n14720) );
no02f01 g10932 ( .a(n14717), .b(n14720), .o(n14721) );
no02f01 g10933 ( .a(n14721), .b(n14719), .o(n14722) );
no03f01 g10934 ( .a(n14629), .b(n14626), .c(n14711), .o(n14723) );
no03f01 g10935 ( .a(n14723), .b(n14659), .c(n14716), .o(n14724) );
in01f01 g10936 ( .a(n14724), .o(n14725) );
no02f01 g10937 ( .a(n14655), .b(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .o(n14726) );
no02f01 g10938 ( .a(n14726), .b(n14628), .o(n14727) );
in01f01 g10939 ( .a(n14727), .o(n14728) );
no02f01 g10940 ( .a(n14728), .b(n14725), .o(n14729) );
no02f01 g10941 ( .a(n14727), .b(n14724), .o(n14730) );
no02f01 g10942 ( .a(n14730), .b(n14729), .o(n14731) );
ao12f01 g10943 ( .a(n14552), .b(n14731), .c(n14722), .o(n14732) );
in01f01 g10944 ( .a(n14665), .o(n14733) );
no02f01 g10945 ( .a(n14631), .b(n14711), .o(n14734) );
ao12f01 g10946 ( .a(n14733), .b(n14734), .c(n14634), .o(n14735) );
no02f01 g10947 ( .a(n14636), .b(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .o(n14736) );
no02f01 g10948 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_22_), .b(n14556), .o(n14737) );
no02f01 g10949 ( .a(n14737), .b(n14736), .o(n14738) );
no02f01 g10950 ( .a(n14738), .b(n14735), .o(n14739) );
na02f01 g10951 ( .a(n14738), .b(n14735), .o(n14740) );
in01f01 g10952 ( .a(n14740), .o(n14741) );
no02f01 g10953 ( .a(n14741), .b(n14739), .o(n14742) );
no04f01 g10954 ( .a(n14737), .b(n14633), .c(n14631), .d(n14711), .o(n14743) );
no03f01 g10955 ( .a(n14743), .b(n14736), .c(n14733), .o(n14744) );
in01f01 g10956 ( .a(n14744), .o(n14745) );
no02f01 g10957 ( .a(n14635), .b(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .o(n14746) );
no02f01 g10958 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_23_), .b(n14556), .o(n14747) );
no02f01 g10959 ( .a(n14747), .b(n14746), .o(n14748) );
in01f01 g10960 ( .a(n14748), .o(n14749) );
no02f01 g10961 ( .a(n14749), .b(n14745), .o(n14750) );
no02f01 g10962 ( .a(n14748), .b(n14744), .o(n14751) );
no02f01 g10963 ( .a(n14751), .b(n14750), .o(n14752) );
in01f01 g10964 ( .a(n14752), .o(n14753) );
no02f01 g10965 ( .a(n14663), .b(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .o(n14754) );
no02f01 g10966 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_20_), .b(n14556), .o(n14755) );
no03f01 g10967 ( .a(n14755), .b(n14631), .c(n14711), .o(n14756) );
no03f01 g10968 ( .a(n14756), .b(n14754), .c(n14661), .o(n14757) );
no02f01 g10969 ( .a(n14662), .b(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .o(n14758) );
no02f01 g10970 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_21_), .b(n14556), .o(n14759) );
no02f01 g10971 ( .a(n14759), .b(n14758), .o(n14760) );
no02f01 g10972 ( .a(n14760), .b(n14757), .o(n14761) );
na02f01 g10973 ( .a(n14760), .b(n14757), .o(n14762) );
in01f01 g10974 ( .a(n14762), .o(n14763) );
no02f01 g10975 ( .a(n14763), .b(n14761), .o(n14764) );
in01f01 g10976 ( .a(n14764), .o(n14765) );
no02f01 g10977 ( .a(n14734), .b(n14661), .o(n14766) );
no02f01 g10978 ( .a(n14755), .b(n14754), .o(n14767) );
no02f01 g10979 ( .a(n14767), .b(n14766), .o(n14768) );
na02f01 g10980 ( .a(n14767), .b(n14766), .o(n14769) );
in01f01 g10981 ( .a(n14769), .o(n14770) );
no02f01 g10982 ( .a(n14770), .b(n14768), .o(n14771) );
in01f01 g10983 ( .a(n14771), .o(n14772) );
no03f01 g10984 ( .a(n14772), .b(n14765), .c(n14753), .o(n14773) );
ao12f01 g10985 ( .a(n14552), .b(n14773), .c(n14742), .o(n14774) );
no03f01 g10986 ( .a(n14774), .b(n14732), .c(n14714), .o(n14775) );
in01f01 g10987 ( .a(n14775), .o(n14776) );
no02f01 g10988 ( .a(n14549), .b(n14543), .o(n14777) );
in01f01 g10989 ( .a(n14549), .o(n14778) );
no02f01 g10990 ( .a(n14778), .b(n14542), .o(n14779) );
no02f01 g10991 ( .a(n14779), .b(n14777), .o(n14780) );
in01f01 g10992 ( .a(n14589), .o(n14781) );
in01f01 g10993 ( .a(n14582), .o(n14782) );
no02f01 g10994 ( .a(n14782), .b(n14576), .o(n14783) );
in01f01 g10995 ( .a(n14783), .o(n14784) );
no02f01 g10996 ( .a(n14784), .b(n14584), .o(n14785) );
no02f01 g10997 ( .a(n14785), .b(n14781), .o(n14786) );
in01f01 g10998 ( .a(n14588), .o(n14787) );
no02f01 g10999 ( .a(n14787), .b(n14578), .o(n14788) );
no02f01 g11000 ( .a(n14788), .b(n14786), .o(n14789) );
na02f01 g11001 ( .a(n14788), .b(n14786), .o(n14790) );
in01f01 g11002 ( .a(n14790), .o(n14791) );
no02f01 g11003 ( .a(n14791), .b(n14789), .o(n14792) );
in01f01 g11004 ( .a(n14792), .o(n14793) );
no02f01 g11005 ( .a(n14793), .b(n14780), .o(n14794) );
in01f01 g11006 ( .a(n14500), .o(n14795) );
no02f01 g11007 ( .a(n14540), .b(n14795), .o(n14796) );
no02f01 g11008 ( .a(n14541), .b(n14500), .o(n14797) );
no02f01 g11009 ( .a(n14797), .b(n14796), .o(n14798) );
in01f01 g11010 ( .a(n14798), .o(n14799) );
no02f01 g11011 ( .a(n14781), .b(n14584), .o(n14800) );
no02f01 g11012 ( .a(n14800), .b(n14784), .o(n14801) );
na02f01 g11013 ( .a(n14800), .b(n14784), .o(n14802) );
in01f01 g11014 ( .a(n14802), .o(n14803) );
no02f01 g11015 ( .a(n14803), .b(n14801), .o(n14804) );
no02f01 g11016 ( .a(n14804), .b(n14799), .o(n14805) );
in01f01 g11017 ( .a(n14805), .o(n14806) );
na02f01 g11018 ( .a(n14539), .b(n14508), .o(n14807) );
no02f01 g11019 ( .a(n14539), .b(n14508), .o(n14808) );
in01f01 g11020 ( .a(n14808), .o(n14809) );
na02f01 g11021 ( .a(n14809), .b(n14807), .o(n14810) );
no02f01 g11022 ( .a(n14573), .b(n14571), .o(n14811) );
no02f01 g11023 ( .a(n14782), .b(n14575), .o(n14812) );
no02f01 g11024 ( .a(n14812), .b(n14811), .o(n14813) );
na02f01 g11025 ( .a(n14812), .b(n14811), .o(n14814) );
in01f01 g11026 ( .a(n14814), .o(n14815) );
no02f01 g11027 ( .a(n14815), .b(n14813), .o(n14816) );
no02f01 g11028 ( .a(n14816), .b(n14810), .o(n14817) );
in01f01 g11029 ( .a(n14817), .o(n14818) );
na02f01 g11030 ( .a(n14538), .b(n14528), .o(n14819) );
no02f01 g11031 ( .a(n14538), .b(n14528), .o(n14820) );
in01f01 g11032 ( .a(n14820), .o(n14821) );
na02f01 g11033 ( .a(n14821), .b(n14819), .o(n14822) );
in01f01 g11034 ( .a(n14568), .o(n14823) );
no02f01 g11035 ( .a(n14573), .b(n14570), .o(n14824) );
in01f01 g11036 ( .a(n14824), .o(n14825) );
no02f01 g11037 ( .a(n14825), .b(n14823), .o(n14826) );
no02f01 g11038 ( .a(n14824), .b(n14568), .o(n14827) );
no02f01 g11039 ( .a(n14827), .b(n14826), .o(n14828) );
no02f01 g11040 ( .a(n14828), .b(n14822), .o(n14829) );
in01f01 g11041 ( .a(n14829), .o(n14830) );
na02f01 g11042 ( .a(n14828), .b(n14822), .o(n14831) );
in01f01 g11043 ( .a(n14567), .o(n14832) );
no03f01 g11044 ( .a(n14832), .b(n14566), .c(n14564), .o(n14833) );
in01f01 g11045 ( .a(n14564), .o(n14834) );
in01f01 g11046 ( .a(n14566), .o(n14835) );
ao12f01 g11047 ( .a(n14835), .b(n14567), .c(n14834), .o(n14836) );
no02f01 g11048 ( .a(n14836), .b(n14833), .o(n14837) );
no02f01 g11049 ( .a(n14464), .b(n14565), .o(n14838) );
no02f01 g11050 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_24_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_0_), .o(n14839) );
no02f01 g11051 ( .a(n14839), .b(n14838), .o(n14840) );
no02f01 g11052 ( .a(n14840), .b(n14519), .o(n14841) );
no02f01 g11053 ( .a(n14841), .b(n14837), .o(n14842) );
in01f01 g11054 ( .a(n14842), .o(n14843) );
na02f01 g11055 ( .a(n14841), .b(n14837), .o(n14844) );
in01f01 g11056 ( .a(n14519), .o(n14845) );
ao12f01 g11057 ( .a(n14527), .b(n14845), .c(delay_sub_ln23_0_unr24_stage9_stallmux_q), .o(n14846) );
in01f01 g11058 ( .a(n14527), .o(n14847) );
no03f01 g11059 ( .a(n14847), .b(n14519), .c(n14492), .o(n14848) );
no02f01 g11060 ( .a(n14848), .b(n14846), .o(n14849) );
na02f01 g11061 ( .a(n14849), .b(n14844), .o(n14850) );
na02f01 g11062 ( .a(n14850), .b(n14843), .o(n14851) );
na02f01 g11063 ( .a(n14851), .b(n14831), .o(n14852) );
na02f01 g11064 ( .a(n14852), .b(n14830), .o(n14853) );
na02f01 g11065 ( .a(n14816), .b(n14810), .o(n14854) );
na02f01 g11066 ( .a(n14854), .b(n14853), .o(n14855) );
na02f01 g11067 ( .a(n14855), .b(n14818), .o(n14856) );
na02f01 g11068 ( .a(n14804), .b(n14799), .o(n14857) );
na02f01 g11069 ( .a(n14857), .b(n14856), .o(n14858) );
na02f01 g11070 ( .a(n14858), .b(n14806), .o(n14859) );
in01f01 g11071 ( .a(n14859), .o(n14860) );
na02f01 g11072 ( .a(n14793), .b(n14780), .o(n14861) );
ao12f01 g11073 ( .a(n14794), .b(n14861), .c(n14860), .o(n14862) );
no03f01 g11074 ( .a(n14550), .b(n14543), .c(n14491), .o(n14863) );
in01f01 g11075 ( .a(n14491), .o(n14864) );
no02f01 g11076 ( .a(n14551), .b(n14864), .o(n14865) );
no02f01 g11077 ( .a(n14865), .b(n14863), .o(n14866) );
ao12f01 g11078 ( .a(n14590), .b(n14785), .c(n14579), .o(n14867) );
in01f01 g11079 ( .a(n14581), .o(n14868) );
no02f01 g11080 ( .a(n14593), .b(n14868), .o(n14869) );
no02f01 g11081 ( .a(n14869), .b(n14867), .o(n14870) );
na02f01 g11082 ( .a(n14869), .b(n14867), .o(n14871) );
in01f01 g11083 ( .a(n14871), .o(n14872) );
no02f01 g11084 ( .a(n14872), .b(n14870), .o(n14873) );
in01f01 g11085 ( .a(n14873), .o(n14874) );
no02f01 g11086 ( .a(n14874), .b(n14866), .o(n14875) );
in01f01 g11087 ( .a(n14875), .o(n14876) );
na02f01 g11088 ( .a(n14594), .b(n14591), .o(n14877) );
no02f01 g11089 ( .a(n14877), .b(n14587), .o(n14878) );
in01f01 g11090 ( .a(n14878), .o(n14879) );
na02f01 g11091 ( .a(n14592), .b(n14562), .o(n14880) );
no02f01 g11092 ( .a(n14880), .b(n14879), .o(n14881) );
na02f01 g11093 ( .a(n14880), .b(n14879), .o(n14882) );
in01f01 g11094 ( .a(n14882), .o(n14883) );
no02f01 g11095 ( .a(n14883), .b(n14881), .o(n14884) );
no02f01 g11096 ( .a(n14884), .b(n14552), .o(n14885) );
na02f01 g11097 ( .a(n14874), .b(n14866), .o(n14886) );
in01f01 g11098 ( .a(n14886), .o(n14887) );
no02f01 g11099 ( .a(n14887), .b(n14885), .o(n14888) );
in01f01 g11100 ( .a(n14888), .o(n14889) );
ao12f01 g11101 ( .a(n14889), .b(n14876), .c(n14862), .o(n14890) );
na02f01 g11102 ( .a(n14884), .b(n14552), .o(n14891) );
in01f01 g11103 ( .a(n14891), .o(n14892) );
no02f01 g11104 ( .a(n14892), .b(n14890), .o(n14893) );
no02f01 g11105 ( .a(n14597), .b(n14596), .o(n14894) );
no02f01 g11106 ( .a(n14894), .b(n14613), .o(n14895) );
no02f01 g11107 ( .a(n14614), .b(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .o(n14896) );
no02f01 g11108 ( .a(n14896), .b(n14605), .o(n14897) );
no02f01 g11109 ( .a(n14897), .b(n14895), .o(n14898) );
na02f01 g11110 ( .a(n14897), .b(n14895), .o(n14899) );
in01f01 g11111 ( .a(n14899), .o(n14900) );
no02f01 g11112 ( .a(n14900), .b(n14898), .o(n14901) );
in01f01 g11113 ( .a(n14901), .o(n14902) );
no02f01 g11114 ( .a(n14902), .b(n14553), .o(n14903) );
no02f01 g11115 ( .a(n14611), .b(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .o(n14904) );
no02f01 g11116 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_8_), .b(n14556), .o(n14905) );
no02f01 g11117 ( .a(n14905), .b(n14596), .o(n14906) );
no02f01 g11118 ( .a(n14906), .b(n14904), .o(n14907) );
no02f01 g11119 ( .a(n14612), .b(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .o(n14908) );
no02f01 g11120 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_9_), .b(n14556), .o(n14909) );
no02f01 g11121 ( .a(n14909), .b(n14908), .o(n14910) );
no02f01 g11122 ( .a(n14910), .b(n14907), .o(n14911) );
na02f01 g11123 ( .a(n14910), .b(n14907), .o(n14912) );
in01f01 g11124 ( .a(n14912), .o(n14913) );
no02f01 g11125 ( .a(n14913), .b(n14911), .o(n14914) );
in01f01 g11126 ( .a(n14914), .o(n14915) );
no02f01 g11127 ( .a(n14905), .b(n14904), .o(n14916) );
no02f01 g11128 ( .a(n14916), .b(n14596), .o(n14917) );
na02f01 g11129 ( .a(n14916), .b(n14596), .o(n14918) );
in01f01 g11130 ( .a(n14918), .o(n14919) );
no02f01 g11131 ( .a(n14919), .b(n14917), .o(n14920) );
in01f01 g11132 ( .a(n14920), .o(n14921) );
ao12f01 g11133 ( .a(n14553), .b(n14921), .c(n14915), .o(n14922) );
no03f01 g11134 ( .a(n14605), .b(n14597), .c(n14596), .o(n14923) );
no03f01 g11135 ( .a(n14923), .b(n14896), .c(n14613), .o(n14924) );
no02f01 g11136 ( .a(n14615), .b(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .o(n14925) );
no02f01 g11137 ( .a(n14925), .b(n14604), .o(n14926) );
no02f01 g11138 ( .a(n14926), .b(n14924), .o(n14927) );
na02f01 g11139 ( .a(n14926), .b(n14924), .o(n14928) );
in01f01 g11140 ( .a(n14928), .o(n14929) );
no02f01 g11141 ( .a(n14929), .b(n14927), .o(n14930) );
in01f01 g11142 ( .a(n14930), .o(n14931) );
no02f01 g11143 ( .a(n14931), .b(n14553), .o(n14932) );
no03f01 g11144 ( .a(n14932), .b(n14922), .c(n14903), .o(n14933) );
na02f01 g11145 ( .a(n14933), .b(n14893), .o(n14934) );
in01f01 g11146 ( .a(n14934), .o(n14935) );
no02f01 g11147 ( .a(n14620), .b(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .o(n14936) );
na02f01 g11148 ( .a(n14894), .b(n14606), .o(n14937) );
no02f01 g11149 ( .a(n14937), .b(n14601), .o(n14938) );
no03f01 g11150 ( .a(n14938), .b(n14936), .c(n14618), .o(n14939) );
no02f01 g11151 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(n14619), .o(n14940) );
no02f01 g11152 ( .a(n14940), .b(n14602), .o(n14941) );
no02f01 g11153 ( .a(n14941), .b(n14939), .o(n14942) );
na02f01 g11154 ( .a(n14941), .b(n14939), .o(n14943) );
in01f01 g11155 ( .a(n14943), .o(n14944) );
no02f01 g11156 ( .a(n14944), .b(n14942), .o(n14945) );
in01f01 g11157 ( .a(n14937), .o(n14946) );
no02f01 g11158 ( .a(n14946), .b(n14618), .o(n14947) );
no02f01 g11159 ( .a(n14936), .b(n14601), .o(n14948) );
no02f01 g11160 ( .a(n14948), .b(n14947), .o(n14949) );
na02f01 g11161 ( .a(n14948), .b(n14947), .o(n14950) );
in01f01 g11162 ( .a(n14950), .o(n14951) );
no02f01 g11163 ( .a(n14951), .b(n14949), .o(n14952) );
no02f01 g11164 ( .a(n14952), .b(n14945), .o(n14953) );
no02f01 g11165 ( .a(n14953), .b(n14553), .o(n14954) );
ao12f01 g11166 ( .a(n14623), .b(n14946), .c(n14603), .o(n14955) );
no02f01 g11167 ( .a(n14608), .b(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .o(n14956) );
no02f01 g11168 ( .a(n14956), .b(n14599), .o(n14957) );
no02f01 g11169 ( .a(n14957), .b(n14955), .o(n14958) );
na02f01 g11170 ( .a(n14957), .b(n14955), .o(n14959) );
in01f01 g11171 ( .a(n14959), .o(n14960) );
no02f01 g11172 ( .a(n14960), .b(n14958), .o(n14961) );
in01f01 g11173 ( .a(n14961), .o(n14962) );
no02f01 g11174 ( .a(n14962), .b(n14553), .o(n14963) );
in01f01 g11175 ( .a(n14603), .o(n14964) );
no03f01 g11176 ( .a(n14937), .b(n14964), .c(n14599), .o(n14965) );
no03f01 g11177 ( .a(n14965), .b(n14623), .c(n14956), .o(n14966) );
in01f01 g11178 ( .a(n14966), .o(n14967) );
no02f01 g11179 ( .a(n14609), .b(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .o(n14968) );
no02f01 g11180 ( .a(n14968), .b(n14598), .o(n14969) );
in01f01 g11181 ( .a(n14969), .o(n14970) );
no02f01 g11182 ( .a(n14970), .b(n14967), .o(n14971) );
no02f01 g11183 ( .a(n14969), .b(n14966), .o(n14972) );
no02f01 g11184 ( .a(n14972), .b(n14971), .o(n14973) );
in01f01 g11185 ( .a(n14973), .o(n14974) );
no02f01 g11186 ( .a(n14974), .b(n14553), .o(n14975) );
no03f01 g11187 ( .a(n14975), .b(n14963), .c(n14954), .o(n14976) );
na02f01 g11188 ( .a(n14976), .b(n14935), .o(n14977) );
ao12f01 g11189 ( .a(n14552), .b(n14930), .c(n14901), .o(n14978) );
ao12f01 g11190 ( .a(n14552), .b(n14920), .c(n14914), .o(n14979) );
no02f01 g11191 ( .a(n14979), .b(n14978), .o(n14980) );
in01f01 g11192 ( .a(n14980), .o(n14981) );
ao12f01 g11193 ( .a(n14552), .b(n14952), .c(n14945), .o(n14982) );
ao12f01 g11194 ( .a(n14552), .b(n14973), .c(n14961), .o(n14983) );
no03f01 g11195 ( .a(n14983), .b(n14982), .c(n14981), .o(n14984) );
na02f01 g11196 ( .a(n14722), .b(n14552), .o(n14985) );
in01f01 g11197 ( .a(n14985), .o(n14986) );
in01f01 g11198 ( .a(n14731), .o(n14987) );
no02f01 g11199 ( .a(n14987), .b(n14553), .o(n14988) );
in01f01 g11200 ( .a(n14707), .o(n14989) );
in01f01 g11201 ( .a(n14713), .o(n14990) );
ao12f01 g11202 ( .a(n14553), .b(n14990), .c(n14989), .o(n14991) );
no03f01 g11203 ( .a(n14991), .b(n14988), .c(n14986), .o(n14992) );
na02f01 g11204 ( .a(n14742), .b(n14552), .o(n14993) );
in01f01 g11205 ( .a(n14993), .o(n14994) );
no02f01 g11206 ( .a(n14771), .b(n14764), .o(n14995) );
no02f01 g11207 ( .a(n14995), .b(n14553), .o(n14996) );
no02f01 g11208 ( .a(n14753), .b(n14553), .o(n14997) );
no03f01 g11209 ( .a(n14997), .b(n14996), .c(n14994), .o(n14998) );
na02f01 g11210 ( .a(n14998), .b(n14992), .o(n14999) );
ao12f01 g11211 ( .a(n14999), .b(n14984), .c(n14977), .o(n15000) );
no02f01 g11212 ( .a(n14669), .b(n14733), .o(n15001) );
in01f01 g11213 ( .a(n15001), .o(n15002) );
no02f01 g11214 ( .a(n15002), .b(n14641), .o(n15003) );
no02f01 g11215 ( .a(n14666), .b(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .o(n15004) );
no02f01 g11216 ( .a(n15004), .b(n14643), .o(n15005) );
no02f01 g11217 ( .a(n15005), .b(n15003), .o(n15006) );
na02f01 g11218 ( .a(n15005), .b(n15003), .o(n15007) );
in01f01 g11219 ( .a(n15007), .o(n15008) );
no02f01 g11220 ( .a(n15008), .b(n15006), .o(n15009) );
in01f01 g11221 ( .a(n15009), .o(n15010) );
no02f01 g11222 ( .a(n14643), .b(n14638), .o(n15011) );
na02f01 g11223 ( .a(n15011), .b(n14625), .o(n15012) );
no02f01 g11224 ( .a(n14667), .b(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .o(n15013) );
no02f01 g11225 ( .a(n15013), .b(n14642), .o(n15014) );
in01f01 g11226 ( .a(n15014), .o(n15015) );
no02f01 g11227 ( .a(n15002), .b(n15004), .o(n15016) );
in01f01 g11228 ( .a(n15016), .o(n15017) );
no02f01 g11229 ( .a(n15015), .b(n15017), .o(n15018) );
na02f01 g11230 ( .a(n15016), .b(n15012), .o(n15019) );
ao22f01 g11231 ( .a(n15019), .b(n15015), .c(n15018), .d(n15012), .o(n15020) );
in01f01 g11232 ( .a(n15020), .o(n15021) );
ao12f01 g11233 ( .a(n14553), .b(n15021), .c(n15010), .o(n15022) );
no02f01 g11234 ( .a(n14670), .b(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .o(n15023) );
no02f01 g11235 ( .a(n15023), .b(n14646), .o(n15024) );
in01f01 g11236 ( .a(n15024), .o(n15025) );
in01f01 g11237 ( .a(n14644), .o(n15026) );
no03f01 g11238 ( .a(n14645), .b(n15026), .c(n14638), .o(n15027) );
na02f01 g11239 ( .a(n15027), .b(n14625), .o(n15028) );
no02f01 g11240 ( .a(n14671), .b(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .o(n15029) );
no02f01 g11241 ( .a(n15002), .b(n14668), .o(n15030) );
in01f01 g11242 ( .a(n15030), .o(n15031) );
no02f01 g11243 ( .a(n15031), .b(n15029), .o(n15032) );
na02f01 g11244 ( .a(n15032), .b(n15028), .o(n15033) );
no02f01 g11245 ( .a(n15033), .b(n15025), .o(n15034) );
na02f01 g11246 ( .a(n15033), .b(n15025), .o(n15035) );
in01f01 g11247 ( .a(n15035), .o(n15036) );
no02f01 g11248 ( .a(n15036), .b(n15034), .o(n15037) );
in01f01 g11249 ( .a(n15037), .o(n15038) );
no02f01 g11250 ( .a(n15038), .b(n14553), .o(n15039) );
no02f01 g11251 ( .a(n15029), .b(n14645), .o(n15040) );
no02f01 g11252 ( .a(n15026), .b(n14640), .o(n15041) );
no02f01 g11253 ( .a(n15041), .b(n15031), .o(n15042) );
in01f01 g11254 ( .a(n15040), .o(n15043) );
no02f01 g11255 ( .a(n15043), .b(n15031), .o(n15044) );
in01f01 g11256 ( .a(n15044), .o(n15045) );
oa22f01 g11257 ( .a(n15045), .b(n15041), .c(n15042), .d(n15040), .o(n15046) );
no02f01 g11258 ( .a(n15046), .b(n14553), .o(n15047) );
no03f01 g11259 ( .a(n15047), .b(n15039), .c(n15022), .o(n15048) );
oa12f01 g11260 ( .a(n15048), .b(n15000), .c(n14776), .o(n15049) );
in01f01 g11261 ( .a(n15046), .o(n15050) );
ao12f01 g11262 ( .a(n14552), .b(n15050), .c(n15037), .o(n15051) );
ao12f01 g11263 ( .a(n14552), .b(n15020), .c(n15009), .o(n15052) );
no02f01 g11264 ( .a(n15052), .b(n15051), .o(n15053) );
na02f01 g11265 ( .a(n15053), .b(n15049), .o(n15054) );
in01f01 g11266 ( .a(n14650), .o(n15055) );
no02f01 g11267 ( .a(n14648), .b(n14640), .o(n15056) );
ao12f01 g11268 ( .a(n14678), .b(n15056), .c(n15055), .o(n15057) );
in01f01 g11269 ( .a(n15057), .o(n15058) );
no02f01 g11270 ( .a(n14680), .b(n14649), .o(n15059) );
in01f01 g11271 ( .a(n15059), .o(n15060) );
no02f01 g11272 ( .a(n15060), .b(n15058), .o(n15061) );
no02f01 g11273 ( .a(n15059), .b(n15057), .o(n15062) );
no02f01 g11274 ( .a(n15062), .b(n15061), .o(n15063) );
no02f01 g11275 ( .a(n15056), .b(n14674), .o(n15064) );
no02f01 g11276 ( .a(n14676), .b(n14650), .o(n15065) );
no02f01 g11277 ( .a(n15065), .b(n15064), .o(n15066) );
na02f01 g11278 ( .a(n15065), .b(n15064), .o(n15067) );
in01f01 g11279 ( .a(n15067), .o(n15068) );
no02f01 g11280 ( .a(n15068), .b(n15066), .o(n15069) );
no02f01 g11281 ( .a(n15069), .b(n15063), .o(n15070) );
oa12f01 g11282 ( .a(n15054), .b(n15070), .c(n14553), .o(n15071) );
no02f01 g11283 ( .a(n14684), .b(n14653), .o(n15072) );
in01f01 g11284 ( .a(n15072), .o(n15073) );
ao12f01 g11285 ( .a(n14682), .b(n14651), .c(n14641), .o(n15074) );
in01f01 g11286 ( .a(n15074), .o(n15075) );
no02f01 g11287 ( .a(n15073), .b(n14682), .o(n15076) );
ao22f01 g11288 ( .a(n15076), .b(n14652), .c(n15075), .d(n15073), .o(n15077) );
in01f01 g11289 ( .a(n15077), .o(n15078) );
no02f01 g11290 ( .a(n15078), .b(n14553), .o(n15079) );
no02f01 g11291 ( .a(n15077), .b(n14552), .o(n15080) );
ao12f01 g11292 ( .a(n14552), .b(n15069), .c(n15063), .o(n15081) );
no02f01 g11293 ( .a(n15081), .b(n15080), .o(n15082) );
oa12f01 g11294 ( .a(n15082), .b(n15079), .c(n15071), .o(n15083) );
no02f01 g11295 ( .a(n15083), .b(n14695), .o(n15084) );
na02f01 g11296 ( .a(n15083), .b(n14695), .o(n15085) );
in01f01 g11297 ( .a(n15085), .o(n15086) );
no02f01 g11298 ( .a(n15086), .b(n15084), .o(n15087) );
no02f01 g11299 ( .a(n15087), .b(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n15088) );
in01f01 g11300 ( .a(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n15089) );
in01f01 g11301 ( .a(n15087), .o(n15090) );
no02f01 g11302 ( .a(n15090), .b(n15089), .o(n15091) );
no02f01 g11303 ( .a(n15091), .b(n15088), .o(n15092) );
in01f01 g11304 ( .a(n15047), .o(n15093) );
no02f01 g11305 ( .a(n15037), .b(n14552), .o(n15094) );
no02f01 g11306 ( .a(n15094), .b(n15039), .o(n15095) );
in01f01 g11307 ( .a(n15095), .o(n15096) );
no02f01 g11308 ( .a(n15050), .b(n14552), .o(n15097) );
in01f01 g11309 ( .a(n15097), .o(n15098) );
na02f01 g11310 ( .a(n14984), .b(n14977), .o(n15099) );
in01f01 g11311 ( .a(n15022), .o(n15100) );
na04f01 g11312 ( .a(n15100), .b(n14998), .c(n14992), .d(n15099), .o(n15101) );
no02f01 g11313 ( .a(n15052), .b(n14776), .o(n15102) );
na03f01 g11314 ( .a(n15102), .b(n15101), .c(n15098), .o(n15103) );
ao12f01 g11315 ( .a(n15096), .b(n15103), .c(n15093), .o(n15104) );
na03f01 g11316 ( .a(n15103), .b(n15096), .c(n15093), .o(n15105) );
in01f01 g11317 ( .a(n15105), .o(n15106) );
no02f01 g11318 ( .a(n15106), .b(n15104), .o(n15107) );
na02f01 g11319 ( .a(n15102), .b(n15101), .o(n15108) );
no02f01 g11320 ( .a(n15097), .b(n15047), .o(n15109) );
in01f01 g11321 ( .a(n15109), .o(n15110) );
no02f01 g11322 ( .a(n15110), .b(n15108), .o(n15111) );
na02f01 g11323 ( .a(n15110), .b(n15108), .o(n15112) );
in01f01 g11324 ( .a(n15112), .o(n15113) );
no02f01 g11325 ( .a(n15113), .b(n15111), .o(n15114) );
ao12f01 g11326 ( .a(n15089), .b(n15114), .c(n15107), .o(n15115) );
no02f01 g11327 ( .a(n15069), .b(n14552), .o(n15116) );
in01f01 g11328 ( .a(n15069), .o(n15117) );
no02f01 g11329 ( .a(n15117), .b(n14553), .o(n15118) );
no02f01 g11330 ( .a(n15118), .b(n15116), .o(n15119) );
na03f01 g11331 ( .a(n15119), .b(n15053), .c(n15049), .o(n15120) );
in01f01 g11332 ( .a(n15119), .o(n15121) );
na02f01 g11333 ( .a(n15121), .b(n15054), .o(n15122) );
na02f01 g11334 ( .a(n15122), .b(n15120), .o(n15123) );
na02f01 g11335 ( .a(n15123), .b(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n15124) );
in01f01 g11336 ( .a(n15124), .o(n15125) );
no02f01 g11337 ( .a(n15125), .b(n15115), .o(n15126) );
no02f01 g11338 ( .a(n15063), .b(n14552), .o(n15127) );
in01f01 g11339 ( .a(n15063), .o(n15128) );
no02f01 g11340 ( .a(n15128), .b(n14553), .o(n15129) );
no02f01 g11341 ( .a(n15129), .b(n15127), .o(n15130) );
in01f01 g11342 ( .a(n15130), .o(n15131) );
ao12f01 g11343 ( .a(n15118), .b(n15053), .c(n15049), .o(n15132) );
no03f01 g11344 ( .a(n15132), .b(n15131), .c(n15116), .o(n15133) );
no02f01 g11345 ( .a(n15132), .b(n15116), .o(n15134) );
no02f01 g11346 ( .a(n15134), .b(n15130), .o(n15135) );
no02f01 g11347 ( .a(n15135), .b(n15133), .o(n15136) );
no02f01 g11348 ( .a(n15136), .b(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n15137) );
in01f01 g11349 ( .a(n15133), .o(n15138) );
oa12f01 g11350 ( .a(n15131), .b(n15132), .c(n15116), .o(n15139) );
na02f01 g11351 ( .a(n15139), .b(n15138), .o(n15140) );
no02f01 g11352 ( .a(n15140), .b(n15089), .o(n15141) );
oa12f01 g11353 ( .a(n15126), .b(n15141), .c(n15137), .o(n15142) );
na02f01 g11354 ( .a(n15140), .b(n15089), .o(n15143) );
na02f01 g11355 ( .a(n15136), .b(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n15144) );
na02f01 g11356 ( .a(n15123), .b(n15089), .o(n15145) );
na03f01 g11357 ( .a(n15145), .b(n15144), .c(n15143), .o(n15146) );
oa12f01 g11358 ( .a(n15089), .b(n15146), .c(n15126), .o(n15147) );
in01f01 g11359 ( .a(n15081), .o(n15148) );
na02f01 g11360 ( .a(n15148), .b(n15071), .o(n15149) );
in01f01 g11361 ( .a(n15149), .o(n15150) );
no02f01 g11362 ( .a(n15080), .b(n15079), .o(n15151) );
no02f01 g11363 ( .a(n15151), .b(n15150), .o(n15152) );
in01f01 g11364 ( .a(n15151), .o(n15153) );
no02f01 g11365 ( .a(n15153), .b(n15149), .o(n15154) );
no02f01 g11366 ( .a(n15154), .b(n15152), .o(n15155) );
no02f01 g11367 ( .a(n15155), .b(n15089), .o(n15156) );
ao12f01 g11368 ( .a(n15156), .b(n15147), .c(n15142), .o(n15157) );
in01f01 g11369 ( .a(n15142), .o(n15158) );
in01f01 g11370 ( .a(n15104), .o(n15159) );
na02f01 g11371 ( .a(n15105), .b(n15159), .o(n15160) );
in01f01 g11372 ( .a(n15111), .o(n15161) );
na02f01 g11373 ( .a(n15112), .b(n15161), .o(n15162) );
oa12f01 g11374 ( .a(delay_sub_ln23_0_unr25_stage9_stallmux_q), .b(n15162), .c(n15160), .o(n15163) );
na02f01 g11375 ( .a(n15124), .b(n15163), .o(n15164) );
in01f01 g11376 ( .a(n15145), .o(n15165) );
no03f01 g11377 ( .a(n15165), .b(n15141), .c(n15137), .o(n15166) );
ao12f01 g11378 ( .a(delay_sub_ln23_0_unr25_stage9_stallmux_q), .b(n15166), .c(n15164), .o(n15167) );
in01f01 g11379 ( .a(n15156), .o(n15168) );
oa12f01 g11380 ( .a(n15168), .b(n15167), .c(n15158), .o(n15169) );
no02f01 g11381 ( .a(n15155), .b(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n15170) );
in01f01 g11382 ( .a(n15170), .o(n15171) );
na03f01 g11383 ( .a(n15171), .b(n15169), .c(n15089), .o(n15172) );
ao22f01 g11384 ( .a(n15172), .b(n15092), .c(n15157), .d(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n15173) );
no02f01 g11385 ( .a(n14690), .b(n14492), .o(n15174) );
no02f01 g11386 ( .a(n15063), .b(n14492), .o(n15175) );
no02f01 g11387 ( .a(n15077), .b(n14492), .o(n15176) );
oa12f01 g11388 ( .a(delay_sub_ln23_0_unr24_stage9_stallmux_q), .b(n15046), .c(n15021), .o(n15177) );
na02f01 g11389 ( .a(n15038), .b(delay_sub_ln23_0_unr24_stage9_stallmux_q), .o(n15178) );
no02f01 g11390 ( .a(n15069), .b(n14492), .o(n15179) );
in01f01 g11391 ( .a(n15179), .o(n15180) );
na03f01 g11392 ( .a(n15180), .b(n15178), .c(n15177), .o(n15181) );
no03f01 g11393 ( .a(n15181), .b(n15176), .c(n15175), .o(n15182) );
ao12f01 g11394 ( .a(delay_sub_ln23_0_unr24_stage9_stallmux_q), .b(n15077), .c(n15063), .o(n15183) );
oa12f01 g11395 ( .a(n14690), .b(n15183), .c(n15182), .o(n15184) );
in01f01 g11396 ( .a(n15184), .o(n15185) );
no02f01 g11397 ( .a(n15185), .b(n15174), .o(n15186) );
in01f01 g11398 ( .a(n15186), .o(n15187) );
no02f01 g11399 ( .a(n14513), .b(n14432), .o(n15188) );
in01f01 g11400 ( .a(n15188), .o(n15189) );
no03f01 g11401 ( .a(n15189), .b(n14463), .c(n14430), .o(n15190) );
ao12f01 g11402 ( .a(n15188), .b(n14462), .c(n14429), .o(n15191) );
no02f01 g11403 ( .a(n15191), .b(n15190), .o(n15192) );
ao12f01 g11404 ( .a(n15187), .b(n15192), .c(n14519), .o(n15193) );
no02f01 g11405 ( .a(n15187), .b(n14527), .o(n15194) );
no02f01 g11406 ( .a(n15194), .b(n15193), .o(n15195) );
ao12f01 g11407 ( .a(n15187), .b(n15195), .c(n14538), .o(n15196) );
no02f01 g11408 ( .a(n14377), .b(n14375), .o(n15197) );
no02f01 g11409 ( .a(n14379), .b(n14349), .o(n15198) );
no02f01 g11410 ( .a(n15198), .b(n15197), .o(n15199) );
na02f01 g11411 ( .a(n15198), .b(n15197), .o(n15200) );
in01f01 g11412 ( .a(n15200), .o(n15201) );
no02f01 g11413 ( .a(n15201), .b(n15199), .o(n15202) );
in01f01 g11414 ( .a(n15202), .o(n15203) );
no02f01 g11415 ( .a(n15203), .b(n15186), .o(n15204) );
no04f01 g11416 ( .a(n15181), .b(n15176), .c(n15175), .d(n14690), .o(n15205) );
no02f01 g11417 ( .a(n15182), .b(n14691), .o(n15206) );
no02f01 g11418 ( .a(n15206), .b(n15205), .o(n15207) );
in01f01 g11419 ( .a(n14373), .o(n15208) );
no02f01 g11420 ( .a(n14377), .b(n14374), .o(n15209) );
in01f01 g11421 ( .a(n15209), .o(n15210) );
no02f01 g11422 ( .a(n15210), .b(n15208), .o(n15211) );
no02f01 g11423 ( .a(n15209), .b(n14373), .o(n15212) );
no02f01 g11424 ( .a(n15212), .b(n15211), .o(n15213) );
no02f01 g11425 ( .a(n15213), .b(n15207), .o(n15214) );
na02f01 g11426 ( .a(n15178), .b(n15177), .o(n15215) );
no03f01 g11427 ( .a(n15215), .b(n15179), .c(n15175), .o(n15216) );
no02f01 g11428 ( .a(n15216), .b(n15078), .o(n15217) );
na02f01 g11429 ( .a(n15216), .b(n15078), .o(n15218) );
in01f01 g11430 ( .a(n15218), .o(n15219) );
in01f01 g11431 ( .a(n14371), .o(n15220) );
ao12f01 g11432 ( .a(n14353), .b(n15220), .c(n14370), .o(n15221) );
no02f01 g11433 ( .a(n14355), .b(n14351), .o(n15222) );
no02f01 g11434 ( .a(n15222), .b(n15221), .o(n15223) );
na02f01 g11435 ( .a(n15222), .b(n15221), .o(n15224) );
in01f01 g11436 ( .a(n15224), .o(n15225) );
no02f01 g11437 ( .a(n15225), .b(n15223), .o(n15226) );
in01f01 g11438 ( .a(n15226), .o(n15227) );
no03f01 g11439 ( .a(n15227), .b(n15219), .c(n15217), .o(n15228) );
na02f01 g11440 ( .a(n15215), .b(n15069), .o(n15229) );
in01f01 g11441 ( .a(n15229), .o(n15230) );
no02f01 g11442 ( .a(n15215), .b(n15069), .o(n15231) );
in01f01 g11443 ( .a(n14368), .o(n15232) );
in01f01 g11444 ( .a(n14358), .o(n15233) );
no02f01 g11445 ( .a(n14369), .b(n15233), .o(n15234) );
in01f01 g11446 ( .a(n15234), .o(n15235) );
no02f01 g11447 ( .a(n15235), .b(n15232), .o(n15236) );
no02f01 g11448 ( .a(n15234), .b(n14368), .o(n15237) );
no02f01 g11449 ( .a(n15237), .b(n15236), .o(n15238) );
in01f01 g11450 ( .a(n15238), .o(n15239) );
no03f01 g11451 ( .a(n15239), .b(n15231), .c(n15230), .o(n15240) );
no02f01 g11452 ( .a(n15177), .b(n15038), .o(n15241) );
na02f01 g11453 ( .a(n15177), .b(n15038), .o(n15242) );
in01f01 g11454 ( .a(n15242), .o(n15243) );
no02f01 g11455 ( .a(n15243), .b(n15241), .o(n15244) );
in01f01 g11456 ( .a(n14367), .o(n15245) );
no02f01 g11457 ( .a(n14362), .b(n14361), .o(n15246) );
na02f01 g11458 ( .a(n15246), .b(n15245), .o(n15247) );
in01f01 g11459 ( .a(n15247), .o(n15248) );
no02f01 g11460 ( .a(n15246), .b(n15245), .o(n15249) );
no02f01 g11461 ( .a(n15249), .b(n15248), .o(n15250) );
na02f01 g11462 ( .a(n15250), .b(n15244), .o(n15251) );
no02f01 g11463 ( .a(n15020), .b(n14492), .o(n15252) );
in01f01 g11464 ( .a(n15252), .o(n15253) );
na02f01 g11465 ( .a(n15253), .b(n15046), .o(n15254) );
na02f01 g11466 ( .a(n15252), .b(n15050), .o(n15255) );
na02f01 g11467 ( .a(n15255), .b(n15254), .o(n15256) );
in01f01 g11468 ( .a(n14364), .o(n15257) );
in01f01 g11469 ( .a(n14366), .o(n15258) );
no03f01 g11470 ( .a(n15258), .b(n14365), .c(n15257), .o(n15259) );
in01f01 g11471 ( .a(n14365), .o(n15260) );
ao12f01 g11472 ( .a(n14366), .b(n15260), .c(n14364), .o(n15261) );
no02f01 g11473 ( .a(n15261), .b(n15259), .o(n15262) );
in01f01 g11474 ( .a(n15262), .o(n15263) );
na02f01 g11475 ( .a(n15263), .b(n15256), .o(n15264) );
no02f01 g11476 ( .a(n15263), .b(n15256), .o(n15265) );
in01f01 g11477 ( .a(delay_sub_ln22_unr24_stage9_stallmux_q_0_), .o(n15266) );
no02f01 g11478 ( .a(n15266), .b(delay_add_ln22_unr23_stage9_stallmux_q_0_), .o(n15267) );
na02f01 g11479 ( .a(n15266), .b(delay_add_ln22_unr23_stage9_stallmux_q_0_), .o(n15268) );
in01f01 g11480 ( .a(n15268), .o(n15269) );
no02f01 g11481 ( .a(n15269), .b(n15267), .o(n15270) );
no02f01 g11482 ( .a(n15270), .b(n15020), .o(n15271) );
in01f01 g11483 ( .a(n15271), .o(n15272) );
oa12f01 g11484 ( .a(n15264), .b(n15272), .c(n15265), .o(n15273) );
no02f01 g11485 ( .a(n15250), .b(n15244), .o(n15274) );
ao12f01 g11486 ( .a(n15274), .b(n15273), .c(n15251), .o(n15275) );
in01f01 g11487 ( .a(n15231), .o(n15276) );
ao12f01 g11488 ( .a(n15238), .b(n15276), .c(n15229), .o(n15277) );
in01f01 g11489 ( .a(n15277), .o(n15278) );
ao12f01 g11490 ( .a(n15240), .b(n15278), .c(n15275), .o(n15279) );
no02f01 g11491 ( .a(n15181), .b(n15063), .o(n15280) );
na02f01 g11492 ( .a(n15181), .b(n15063), .o(n15281) );
in01f01 g11493 ( .a(n15281), .o(n15282) );
no02f01 g11494 ( .a(n15282), .b(n15280), .o(n15283) );
no02f01 g11495 ( .a(n14371), .b(n14353), .o(n15284) );
in01f01 g11496 ( .a(n15284), .o(n15285) );
no02f01 g11497 ( .a(n15285), .b(n14370), .o(n15286) );
in01f01 g11498 ( .a(n14370), .o(n15287) );
no02f01 g11499 ( .a(n15284), .b(n15287), .o(n15288) );
no02f01 g11500 ( .a(n15288), .b(n15286), .o(n15289) );
na02f01 g11501 ( .a(n15289), .b(n15283), .o(n15290) );
na02f01 g11502 ( .a(n15290), .b(n15279), .o(n15291) );
in01f01 g11503 ( .a(n15217), .o(n15292) );
ao12f01 g11504 ( .a(n15226), .b(n15218), .c(n15292), .o(n15293) );
no02f01 g11505 ( .a(n15289), .b(n15283), .o(n15294) );
no02f01 g11506 ( .a(n15294), .b(n15293), .o(n15295) );
ao12f01 g11507 ( .a(n15228), .b(n15295), .c(n15291), .o(n15296) );
na02f01 g11508 ( .a(n15213), .b(n15207), .o(n15297) );
ao12f01 g11509 ( .a(n15214), .b(n15297), .c(n15296), .o(n15298) );
no02f01 g11510 ( .a(n15202), .b(n15187), .o(n15299) );
in01f01 g11511 ( .a(n15299), .o(n15300) );
ao12f01 g11512 ( .a(n15204), .b(n15300), .c(n15298), .o(n15301) );
no02f01 g11513 ( .a(n14383), .b(n14382), .o(n15302) );
no02f01 g11514 ( .a(n15302), .b(n14402), .o(n15303) );
no02f01 g11515 ( .a(n14398), .b(n14397), .o(n15304) );
no02f01 g11516 ( .a(n15304), .b(n14384), .o(n15305) );
no02f01 g11517 ( .a(n15305), .b(n15303), .o(n15306) );
na02f01 g11518 ( .a(n15305), .b(n15303), .o(n15307) );
in01f01 g11519 ( .a(n15307), .o(n15308) );
no02f01 g11520 ( .a(n15308), .b(n15306), .o(n15309) );
in01f01 g11521 ( .a(n15309), .o(n15310) );
no02f01 g11522 ( .a(n15310), .b(n15186), .o(n15311) );
in01f01 g11523 ( .a(n15311), .o(n15312) );
in01f01 g11524 ( .a(n14382), .o(n15313) );
no02f01 g11525 ( .a(n14397), .b(n14400), .o(n15314) );
no02f01 g11526 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_8_), .o(n15315) );
in01f01 g11527 ( .a(n15315), .o(n15316) );
ao12f01 g11528 ( .a(n15314), .b(n15316), .c(n15313), .o(n15317) );
in01f01 g11529 ( .a(n15317), .o(n15318) );
no02f01 g11530 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_9_), .b(n_46254), .o(n15319) );
no02f01 g11531 ( .a(n14401), .b(n14397), .o(n15320) );
no02f01 g11532 ( .a(n15320), .b(n15319), .o(n15321) );
in01f01 g11533 ( .a(n15321), .o(n15322) );
no02f01 g11534 ( .a(n15322), .b(n15318), .o(n15323) );
no02f01 g11535 ( .a(n15321), .b(n15317), .o(n15324) );
no02f01 g11536 ( .a(n15324), .b(n15323), .o(n15325) );
in01f01 g11537 ( .a(n15325), .o(n15326) );
no02f01 g11538 ( .a(n15315), .b(n15314), .o(n15327) );
in01f01 g11539 ( .a(n15327), .o(n15328) );
no02f01 g11540 ( .a(n15328), .b(n15313), .o(n15329) );
no02f01 g11541 ( .a(n15327), .b(n14382), .o(n15330) );
no02f01 g11542 ( .a(n15330), .b(n15329), .o(n15331) );
in01f01 g11543 ( .a(n15331), .o(n15332) );
ao12f01 g11544 ( .a(n15186), .b(n15332), .c(n15326), .o(n15333) );
no03f01 g11545 ( .a(n14384), .b(n14383), .c(n14382), .o(n15334) );
no03f01 g11546 ( .a(n15334), .b(n14402), .c(n15304), .o(n15335) );
in01f01 g11547 ( .a(n15335), .o(n15336) );
no02f01 g11548 ( .a(n14397), .b(n14396), .o(n15337) );
no02f01 g11549 ( .a(n15337), .b(n14385), .o(n15338) );
in01f01 g11550 ( .a(n15338), .o(n15339) );
no02f01 g11551 ( .a(n15339), .b(n15336), .o(n15340) );
no02f01 g11552 ( .a(n15338), .b(n15335), .o(n15341) );
no02f01 g11553 ( .a(n15341), .b(n15340), .o(n15342) );
in01f01 g11554 ( .a(n15342), .o(n15343) );
no02f01 g11555 ( .a(n15343), .b(n15186), .o(n15344) );
no02f01 g11556 ( .a(n15344), .b(n15333), .o(n15345) );
na02f01 g11557 ( .a(n15345), .b(n15312), .o(n15346) );
no02f01 g11558 ( .a(n14397), .b(n14405), .o(n15347) );
in01f01 g11559 ( .a(n14388), .o(n15348) );
no02f01 g11560 ( .a(n14390), .b(n15348), .o(n15349) );
no03f01 g11561 ( .a(n15349), .b(n15347), .c(n14404), .o(n15350) );
in01f01 g11562 ( .a(n15350), .o(n15351) );
no02f01 g11563 ( .a(n14397), .b(n14406), .o(n15352) );
no02f01 g11564 ( .a(n15352), .b(n14389), .o(n15353) );
in01f01 g11565 ( .a(n15353), .o(n15354) );
no02f01 g11566 ( .a(n15354), .b(n15351), .o(n15355) );
no02f01 g11567 ( .a(n15353), .b(n15350), .o(n15356) );
no02f01 g11568 ( .a(n15356), .b(n15355), .o(n15357) );
in01f01 g11569 ( .a(n15357), .o(n15358) );
no02f01 g11570 ( .a(n15358), .b(n15186), .o(n15359) );
no02f01 g11571 ( .a(n15347), .b(n14390), .o(n15360) );
in01f01 g11572 ( .a(n15360), .o(n15361) );
no03f01 g11573 ( .a(n15361), .b(n14404), .c(n14388), .o(n15362) );
ao12f01 g11574 ( .a(n15360), .b(n14403), .c(n15348), .o(n15363) );
no02f01 g11575 ( .a(n15363), .b(n15362), .o(n15364) );
in01f01 g11576 ( .a(n15364), .o(n15365) );
no02f01 g11577 ( .a(n15365), .b(n15186), .o(n15366) );
no02f01 g11578 ( .a(n15366), .b(n15359), .o(n15367) );
in01f01 g11579 ( .a(n15367), .o(n15368) );
no02f01 g11580 ( .a(n14392), .b(n15348), .o(n15369) );
no02f01 g11581 ( .a(n15369), .b(n14409), .o(n15370) );
no02f01 g11582 ( .a(n14411), .b(n14397), .o(n15371) );
no02f01 g11583 ( .a(n15371), .b(n14393), .o(n15372) );
no02f01 g11584 ( .a(n15372), .b(n15370), .o(n15373) );
na02f01 g11585 ( .a(n15372), .b(n15370), .o(n15374) );
in01f01 g11586 ( .a(n15374), .o(n15375) );
no02f01 g11587 ( .a(n15375), .b(n15373), .o(n15376) );
in01f01 g11588 ( .a(n15376), .o(n15377) );
no02f01 g11589 ( .a(n15377), .b(n15186), .o(n15378) );
in01f01 g11590 ( .a(n15369), .o(n15379) );
no02f01 g11591 ( .a(n15371), .b(n14409), .o(n15380) );
oa12f01 g11592 ( .a(n15380), .b(n15379), .c(n14393), .o(n15381) );
no02f01 g11593 ( .a(n14410), .b(n14397), .o(n15382) );
no02f01 g11594 ( .a(n15382), .b(n14394), .o(n15383) );
in01f01 g11595 ( .a(n15383), .o(n15384) );
no02f01 g11596 ( .a(n15384), .b(n15381), .o(n15385) );
na02f01 g11597 ( .a(n15384), .b(n15381), .o(n15386) );
in01f01 g11598 ( .a(n15386), .o(n15387) );
no02f01 g11599 ( .a(n15387), .b(n15385), .o(n15388) );
in01f01 g11600 ( .a(n15388), .o(n15389) );
no02f01 g11601 ( .a(n15389), .b(n15186), .o(n15390) );
no04f01 g11602 ( .a(n15390), .b(n15378), .c(n15368), .d(n15346), .o(n15391) );
na02f01 g11603 ( .a(n15391), .b(n15301), .o(n15392) );
ao12f01 g11604 ( .a(n15187), .b(n15331), .c(n15325), .o(n15393) );
ao12f01 g11605 ( .a(n15187), .b(n15342), .c(n15309), .o(n15394) );
ao12f01 g11606 ( .a(n15187), .b(n15388), .c(n15376), .o(n15395) );
ao12f01 g11607 ( .a(n15187), .b(n15364), .c(n15357), .o(n15396) );
no04f01 g11608 ( .a(n15396), .b(n15395), .c(n15394), .d(n15393), .o(n15397) );
na02f01 g11609 ( .a(n15397), .b(n15392), .o(n15398) );
no03f01 g11610 ( .a(n14417), .b(n14416), .c(n14415), .o(n15399) );
no02f01 g11611 ( .a(n14397), .b(n14450), .o(n15400) );
no03f01 g11612 ( .a(n15400), .b(n15399), .c(n14448), .o(n15401) );
in01f01 g11613 ( .a(n15401), .o(n15402) );
no02f01 g11614 ( .a(n14397), .b(n14449), .o(n15403) );
no02f01 g11615 ( .a(n15403), .b(n14418), .o(n15404) );
in01f01 g11616 ( .a(n15404), .o(n15405) );
no02f01 g11617 ( .a(n15405), .b(n15402), .o(n15406) );
no02f01 g11618 ( .a(n15404), .b(n15401), .o(n15407) );
no02f01 g11619 ( .a(n15407), .b(n15406), .o(n15408) );
in01f01 g11620 ( .a(n15408), .o(n15409) );
no02f01 g11621 ( .a(n15409), .b(n15186), .o(n15410) );
in01f01 g11622 ( .a(n14415), .o(n15411) );
no02f01 g11623 ( .a(n14397), .b(n14446), .o(n15412) );
no02f01 g11624 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_16_), .o(n15413) );
in01f01 g11625 ( .a(n15413), .o(n15414) );
ao12f01 g11626 ( .a(n15412), .b(n15414), .c(n15411), .o(n15415) );
in01f01 g11627 ( .a(n15415), .o(n15416) );
no02f01 g11628 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_17_), .o(n15417) );
no02f01 g11629 ( .a(n14397), .b(n14447), .o(n15418) );
no02f01 g11630 ( .a(n15418), .b(n15417), .o(n15419) );
in01f01 g11631 ( .a(n15419), .o(n15420) );
no02f01 g11632 ( .a(n15420), .b(n15416), .o(n15421) );
no02f01 g11633 ( .a(n15419), .b(n15415), .o(n15422) );
no02f01 g11634 ( .a(n15422), .b(n15421), .o(n15423) );
in01f01 g11635 ( .a(n15423), .o(n15424) );
no02f01 g11636 ( .a(n15413), .b(n15412), .o(n15425) );
in01f01 g11637 ( .a(n15425), .o(n15426) );
no02f01 g11638 ( .a(n15426), .b(n15411), .o(n15427) );
no02f01 g11639 ( .a(n15425), .b(n14415), .o(n15428) );
no02f01 g11640 ( .a(n15428), .b(n15427), .o(n15429) );
in01f01 g11641 ( .a(n15429), .o(n15430) );
ao12f01 g11642 ( .a(n15186), .b(n15430), .c(n15424), .o(n15431) );
no02f01 g11643 ( .a(n14416), .b(n14415), .o(n15432) );
no02f01 g11644 ( .a(n15432), .b(n14448), .o(n15433) );
no02f01 g11645 ( .a(n15400), .b(n14417), .o(n15434) );
no02f01 g11646 ( .a(n15434), .b(n15433), .o(n15435) );
na02f01 g11647 ( .a(n15434), .b(n15433), .o(n15436) );
in01f01 g11648 ( .a(n15436), .o(n15437) );
no02f01 g11649 ( .a(n15437), .b(n15435), .o(n15438) );
in01f01 g11650 ( .a(n15438), .o(n15439) );
no02f01 g11651 ( .a(n15439), .b(n15186), .o(n15440) );
no03f01 g11652 ( .a(n15440), .b(n15431), .c(n15410), .o(n15441) );
in01f01 g11653 ( .a(n14421), .o(n15442) );
no02f01 g11654 ( .a(n14423), .b(n15442), .o(n15443) );
no02f01 g11655 ( .a(n14397), .b(n14455), .o(n15444) );
no03f01 g11656 ( .a(n15444), .b(n15443), .c(n14453), .o(n15445) );
no02f01 g11657 ( .a(n14397), .b(n14454), .o(n15446) );
no02f01 g11658 ( .a(n15446), .b(n14422), .o(n15447) );
no02f01 g11659 ( .a(n15447), .b(n15445), .o(n15448) );
na02f01 g11660 ( .a(n15447), .b(n15445), .o(n15449) );
in01f01 g11661 ( .a(n15449), .o(n15450) );
no02f01 g11662 ( .a(n15450), .b(n15448), .o(n15451) );
in01f01 g11663 ( .a(n15451), .o(n15452) );
no02f01 g11664 ( .a(n15452), .b(n15186), .o(n15453) );
no02f01 g11665 ( .a(n15444), .b(n14423), .o(n15454) );
in01f01 g11666 ( .a(n15454), .o(n15455) );
no03f01 g11667 ( .a(n15455), .b(n14453), .c(n14421), .o(n15456) );
ao12f01 g11668 ( .a(n15454), .b(n14452), .c(n15442), .o(n15457) );
no02f01 g11669 ( .a(n15457), .b(n15456), .o(n15458) );
in01f01 g11670 ( .a(n15458), .o(n15459) );
no02f01 g11671 ( .a(n15459), .b(n15186), .o(n15460) );
no02f01 g11672 ( .a(n15460), .b(n15453), .o(n15461) );
no02f01 g11673 ( .a(n14397), .b(n14460), .o(n15462) );
no03f01 g11674 ( .a(n14427), .b(n14425), .c(n15442), .o(n15463) );
no03f01 g11675 ( .a(n15463), .b(n15462), .c(n14458), .o(n15464) );
in01f01 g11676 ( .a(n15464), .o(n15465) );
no02f01 g11677 ( .a(n14397), .b(n14459), .o(n15466) );
no02f01 g11678 ( .a(n15466), .b(n14426), .o(n15467) );
in01f01 g11679 ( .a(n15467), .o(n15468) );
no02f01 g11680 ( .a(n15468), .b(n15465), .o(n15469) );
no02f01 g11681 ( .a(n15467), .b(n15464), .o(n15470) );
no02f01 g11682 ( .a(n15470), .b(n15469), .o(n15471) );
in01f01 g11683 ( .a(n15471), .o(n15472) );
no02f01 g11684 ( .a(n14425), .b(n15442), .o(n15473) );
no02f01 g11685 ( .a(n15462), .b(n14427), .o(n15474) );
in01f01 g11686 ( .a(n15474), .o(n15475) );
no03f01 g11687 ( .a(n15475), .b(n15473), .c(n14458), .o(n15476) );
no02f01 g11688 ( .a(n15473), .b(n14458), .o(n15477) );
no02f01 g11689 ( .a(n15474), .b(n15477), .o(n15478) );
no02f01 g11690 ( .a(n15478), .b(n15476), .o(n15479) );
in01f01 g11691 ( .a(n15479), .o(n15480) );
ao12f01 g11692 ( .a(n15186), .b(n15480), .c(n15472), .o(n15481) );
in01f01 g11693 ( .a(n15481), .o(n15482) );
na04f01 g11694 ( .a(n15482), .b(n15461), .c(n15441), .d(n15398), .o(n15483) );
in01f01 g11695 ( .a(n15483), .o(n15484) );
ao12f01 g11696 ( .a(n15187), .b(n15458), .c(n15451), .o(n15485) );
ao12f01 g11697 ( .a(n15187), .b(n15479), .c(n15471), .o(n15486) );
no02f01 g11698 ( .a(n15439), .b(n15409), .o(n15487) );
no02f01 g11699 ( .a(n15430), .b(n15424), .o(n15488) );
ao12f01 g11700 ( .a(n15187), .b(n15488), .c(n15487), .o(n15489) );
no03f01 g11701 ( .a(n15489), .b(n15486), .c(n15485), .o(n15490) );
in01f01 g11702 ( .a(n15490), .o(n15491) );
no02f01 g11703 ( .a(n15491), .b(n15484), .o(n15492) );
in01f01 g11704 ( .a(n15492), .o(n15493) );
in01f01 g11705 ( .a(n15192), .o(n15494) );
ao12f01 g11706 ( .a(n15186), .b(n15494), .c(n14845), .o(n15495) );
no02f01 g11707 ( .a(n15186), .b(n14847), .o(n15496) );
in01f01 g11708 ( .a(n14538), .o(n15497) );
no02f01 g11709 ( .a(n15186), .b(n15497), .o(n15498) );
no03f01 g11710 ( .a(n15498), .b(n15496), .c(n15495), .o(n15499) );
ao12f01 g11711 ( .a(n15196), .b(n15499), .c(n15493), .o(n15500) );
no02f01 g11712 ( .a(n15187), .b(n14508), .o(n15501) );
in01f01 g11713 ( .a(n14508), .o(n15502) );
no02f01 g11714 ( .a(n15186), .b(n15502), .o(n15503) );
no02f01 g11715 ( .a(n15503), .b(n15501), .o(n15504) );
na02f01 g11716 ( .a(n15504), .b(n15500), .o(n15505) );
in01f01 g11717 ( .a(n15505), .o(n15506) );
no02f01 g11718 ( .a(n15504), .b(n15500), .o(n15507) );
no02f01 g11719 ( .a(n15507), .b(n15506), .o(n15508) );
in01f01 g11720 ( .a(n15508), .o(n15509) );
no02f01 g11721 ( .a(n15509), .b(n15173), .o(n15510) );
no02f01 g11722 ( .a(n15087), .b(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n15511) );
no02f01 g11723 ( .a(n15087), .b(n15089), .o(n15512) );
no02f01 g11724 ( .a(n15512), .b(n15511), .o(n15513) );
na03f01 g11725 ( .a(n15513), .b(n15171), .c(n15169), .o(n15514) );
in01f01 g11726 ( .a(n15513), .o(n15515) );
oa12f01 g11727 ( .a(n15515), .b(n15170), .c(n15157), .o(n15516) );
in01f01 g11728 ( .a(n15294), .o(n15517) );
na02f01 g11729 ( .a(n15517), .b(n15291), .o(n15518) );
in01f01 g11730 ( .a(n15518), .o(n15519) );
no02f01 g11731 ( .a(n15293), .b(n15228), .o(n15520) );
no02f01 g11732 ( .a(n15520), .b(n15519), .o(n15521) );
na02f01 g11733 ( .a(n15520), .b(n15519), .o(n15522) );
in01f01 g11734 ( .a(n15522), .o(n15523) );
no02f01 g11735 ( .a(n15523), .b(n15521), .o(n15524) );
ao12f01 g11736 ( .a(n15524), .b(n15516), .c(n15514), .o(n15525) );
no02f01 g11737 ( .a(n15170), .b(n15156), .o(n15526) );
na03f01 g11738 ( .a(n15526), .b(n15147), .c(n15142), .o(n15527) );
in01f01 g11739 ( .a(n15526), .o(n15528) );
oa12f01 g11740 ( .a(n15528), .b(n15167), .c(n15158), .o(n15529) );
na02f01 g11741 ( .a(n15517), .b(n15290), .o(n15530) );
no02f01 g11742 ( .a(n15530), .b(n15279), .o(n15531) );
na02f01 g11743 ( .a(n15530), .b(n15279), .o(n15532) );
in01f01 g11744 ( .a(n15532), .o(n15533) );
no02f01 g11745 ( .a(n15533), .b(n15531), .o(n15534) );
ao12f01 g11746 ( .a(n15534), .b(n15529), .c(n15527), .o(n15535) );
no02f01 g11747 ( .a(n15136), .b(n15089), .o(n15536) );
no02f01 g11748 ( .a(n15136), .b(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n15537) );
no02f01 g11749 ( .a(n15537), .b(n15536), .o(n15538) );
na02f01 g11750 ( .a(n15538), .b(n15164), .o(n15539) );
in01f01 g11751 ( .a(n15539), .o(n15540) );
no02f01 g11752 ( .a(n15538), .b(n15164), .o(n15541) );
in01f01 g11753 ( .a(n15275), .o(n15542) );
no03f01 g11754 ( .a(n15277), .b(n15542), .c(n15240), .o(n15543) );
no02f01 g11755 ( .a(n15277), .b(n15240), .o(n15544) );
no02f01 g11756 ( .a(n15544), .b(n15275), .o(n15545) );
no02f01 g11757 ( .a(n15545), .b(n15543), .o(n15546) );
in01f01 g11758 ( .a(n15546), .o(n15547) );
oa12f01 g11759 ( .a(n15547), .b(n15541), .c(n15540), .o(n15548) );
na02f01 g11760 ( .a(n15145), .b(n15124), .o(n15549) );
in01f01 g11761 ( .a(n15549), .o(n15550) );
na02f01 g11762 ( .a(n15550), .b(n15115), .o(n15551) );
na02f01 g11763 ( .a(n15549), .b(n15163), .o(n15552) );
in01f01 g11764 ( .a(n15273), .o(n15553) );
in01f01 g11765 ( .a(n15251), .o(n15554) );
no02f01 g11766 ( .a(n15274), .b(n15554), .o(n15555) );
no02f01 g11767 ( .a(n15555), .b(n15553), .o(n15556) );
na02f01 g11768 ( .a(n15555), .b(n15553), .o(n15557) );
in01f01 g11769 ( .a(n15557), .o(n15558) );
no02f01 g11770 ( .a(n15558), .b(n15556), .o(n15559) );
ao12f01 g11771 ( .a(n15559), .b(n15552), .c(n15551), .o(n15560) );
in01f01 g11772 ( .a(n15264), .o(n15561) );
no02f01 g11773 ( .a(n15265), .b(n15561), .o(n15562) );
no02f01 g11774 ( .a(n15562), .b(n15272), .o(n15563) );
na02f01 g11775 ( .a(n15562), .b(n15272), .o(n15564) );
in01f01 g11776 ( .a(n15564), .o(n15565) );
no02f01 g11777 ( .a(n15565), .b(n15563), .o(n15566) );
in01f01 g11778 ( .a(n15566), .o(n15567) );
no02f01 g11779 ( .a(n15162), .b(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n15568) );
no02f01 g11780 ( .a(n15162), .b(n15089), .o(n15569) );
in01f01 g11781 ( .a(n15270), .o(n15570) );
no02f01 g11782 ( .a(n15570), .b(n15020), .o(n15571) );
no02f01 g11783 ( .a(n15270), .b(n15021), .o(n15572) );
no02f01 g11784 ( .a(n15572), .b(n15571), .o(n15573) );
no03f01 g11785 ( .a(n15573), .b(n15569), .c(n15568), .o(n15574) );
na02f01 g11786 ( .a(n15574), .b(n15567), .o(n15575) );
no02f01 g11787 ( .a(n15574), .b(n15567), .o(n15576) );
no03f01 g11788 ( .a(n15114), .b(n15160), .c(n15089), .o(n15577) );
ao12f01 g11789 ( .a(n15107), .b(n15162), .c(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n15578) );
no02f01 g11790 ( .a(n15578), .b(n15577), .o(n15579) );
oa12f01 g11791 ( .a(n15575), .b(n15579), .c(n15576), .o(n15580) );
na03f01 g11792 ( .a(n15559), .b(n15552), .c(n15551), .o(n15581) );
ao12f01 g11793 ( .a(n15560), .b(n15581), .c(n15580), .o(n15582) );
no03f01 g11794 ( .a(n15547), .b(n15541), .c(n15540), .o(n15583) );
oa12f01 g11795 ( .a(n15548), .b(n15583), .c(n15582), .o(n15584) );
na03f01 g11796 ( .a(n15534), .b(n15529), .c(n15527), .o(n15585) );
ao12f01 g11797 ( .a(n15535), .b(n15585), .c(n15584), .o(n15586) );
no03f01 g11798 ( .a(n15515), .b(n15170), .c(n15157), .o(n15587) );
ao12f01 g11799 ( .a(n15513), .b(n15171), .c(n15169), .o(n15588) );
in01f01 g11800 ( .a(n15524), .o(n15589) );
no03f01 g11801 ( .a(n15589), .b(n15588), .c(n15587), .o(n15590) );
no02f01 g11802 ( .a(n15590), .b(n15586), .o(n15591) );
in01f01 g11803 ( .a(n15092), .o(n15592) );
no03f01 g11804 ( .a(n15170), .b(n15157), .c(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n15593) );
oa22f01 g11805 ( .a(n15593), .b(n15592), .c(n15169), .d(n15089), .o(n15594) );
in01f01 g11806 ( .a(n15298), .o(n15595) );
no02f01 g11807 ( .a(n15299), .b(n15204), .o(n15596) );
in01f01 g11808 ( .a(n15596), .o(n15597) );
no02f01 g11809 ( .a(n15597), .b(n15595), .o(n15598) );
no02f01 g11810 ( .a(n15596), .b(n15298), .o(n15599) );
no02f01 g11811 ( .a(n15599), .b(n15598), .o(n15600) );
in01f01 g11812 ( .a(n15297), .o(n15601) );
no02f01 g11813 ( .a(n15601), .b(n15214), .o(n15602) );
in01f01 g11814 ( .a(n15602), .o(n15603) );
no02f01 g11815 ( .a(n15603), .b(n15296), .o(n15604) );
na02f01 g11816 ( .a(n15603), .b(n15296), .o(n15605) );
in01f01 g11817 ( .a(n15605), .o(n15606) );
no02f01 g11818 ( .a(n15606), .b(n15604), .o(n15607) );
ao12f01 g11819 ( .a(n15594), .b(n15607), .c(n15600), .o(n15608) );
no03f01 g11820 ( .a(n15608), .b(n15591), .c(n15525), .o(n15609) );
in01f01 g11821 ( .a(n15600), .o(n15610) );
in01f01 g11822 ( .a(n15607), .o(n15611) );
ao12f01 g11823 ( .a(n15173), .b(n15611), .c(n15610), .o(n15612) );
in01f01 g11824 ( .a(n15301), .o(n15613) );
no02f01 g11825 ( .a(n15333), .b(n15613), .o(n15614) );
no02f01 g11826 ( .a(n15309), .b(n15187), .o(n15615) );
no02f01 g11827 ( .a(n15615), .b(n15311), .o(n15616) );
in01f01 g11828 ( .a(n15616), .o(n15617) );
no03f01 g11829 ( .a(n15617), .b(n15614), .c(n15393), .o(n15618) );
no02f01 g11830 ( .a(n15614), .b(n15393), .o(n15619) );
no02f01 g11831 ( .a(n15616), .b(n15619), .o(n15620) );
no02f01 g11832 ( .a(n15620), .b(n15618), .o(n15621) );
na02f01 g11833 ( .a(n15621), .b(n15594), .o(n15622) );
no02f01 g11834 ( .a(n15331), .b(n15187), .o(n15623) );
no02f01 g11835 ( .a(n15332), .b(n15186), .o(n15624) );
in01f01 g11836 ( .a(n15624), .o(n15625) );
ao12f01 g11837 ( .a(n15623), .b(n15625), .c(n15301), .o(n15626) );
no02f01 g11838 ( .a(n15325), .b(n15187), .o(n15627) );
no02f01 g11839 ( .a(n15326), .b(n15186), .o(n15628) );
no02f01 g11840 ( .a(n15628), .b(n15627), .o(n15629) );
no02f01 g11841 ( .a(n15629), .b(n15626), .o(n15630) );
na02f01 g11842 ( .a(n15629), .b(n15626), .o(n15631) );
in01f01 g11843 ( .a(n15631), .o(n15632) );
no02f01 g11844 ( .a(n15632), .b(n15630), .o(n15633) );
no02f01 g11845 ( .a(n15624), .b(n15623), .o(n15634) );
in01f01 g11846 ( .a(n15634), .o(n15635) );
no02f01 g11847 ( .a(n15635), .b(n15301), .o(n15636) );
no02f01 g11848 ( .a(n15634), .b(n15613), .o(n15637) );
no02f01 g11849 ( .a(n15637), .b(n15636), .o(n15638) );
oa12f01 g11850 ( .a(n15594), .b(n15638), .c(n15633), .o(n15639) );
na02f01 g11851 ( .a(n15614), .b(n15312), .o(n15640) );
no02f01 g11852 ( .a(n15615), .b(n15393), .o(n15641) );
na02f01 g11853 ( .a(n15641), .b(n15640), .o(n15642) );
in01f01 g11854 ( .a(n15642), .o(n15643) );
no02f01 g11855 ( .a(n15342), .b(n15187), .o(n15644) );
no02f01 g11856 ( .a(n15644), .b(n15344), .o(n15645) );
no02f01 g11857 ( .a(n15645), .b(n15643), .o(n15646) );
na02f01 g11858 ( .a(n15645), .b(n15643), .o(n15647) );
in01f01 g11859 ( .a(n15647), .o(n15648) );
no02f01 g11860 ( .a(n15648), .b(n15646), .o(n15649) );
na02f01 g11861 ( .a(n15649), .b(n15594), .o(n15650) );
na03f01 g11862 ( .a(n15650), .b(n15639), .c(n15622), .o(n15651) );
in01f01 g11863 ( .a(n15378), .o(n15652) );
no02f01 g11864 ( .a(n15394), .b(n15393), .o(n15653) );
oa12f01 g11865 ( .a(n15653), .b(n15346), .c(n15613), .o(n15654) );
in01f01 g11866 ( .a(n15654), .o(n15655) );
no02f01 g11867 ( .a(n15376), .b(n15187), .o(n15656) );
no02f01 g11868 ( .a(n15396), .b(n15656), .o(n15657) );
oa12f01 g11869 ( .a(n15657), .b(n15655), .c(n15368), .o(n15658) );
na02f01 g11870 ( .a(n15658), .b(n15652), .o(n15659) );
no02f01 g11871 ( .a(n15388), .b(n15187), .o(n15660) );
no02f01 g11872 ( .a(n15660), .b(n15390), .o(n15661) );
no02f01 g11873 ( .a(n15661), .b(n15659), .o(n15662) );
na02f01 g11874 ( .a(n15661), .b(n15659), .o(n15663) );
in01f01 g11875 ( .a(n15663), .o(n15664) );
no02f01 g11876 ( .a(n15664), .b(n15662), .o(n15665) );
na02f01 g11877 ( .a(n15665), .b(n15594), .o(n15666) );
no02f01 g11878 ( .a(n15364), .b(n15187), .o(n15667) );
no02f01 g11879 ( .a(n15667), .b(n15654), .o(n15668) );
no02f01 g11880 ( .a(n15668), .b(n15366), .o(n15669) );
in01f01 g11881 ( .a(n15669), .o(n15670) );
no02f01 g11882 ( .a(n15357), .b(n15187), .o(n15671) );
no02f01 g11883 ( .a(n15671), .b(n15359), .o(n15672) );
no02f01 g11884 ( .a(n15672), .b(n15670), .o(n15673) );
na02f01 g11885 ( .a(n15672), .b(n15670), .o(n15674) );
in01f01 g11886 ( .a(n15674), .o(n15675) );
no02f01 g11887 ( .a(n15675), .b(n15673), .o(n15676) );
no02f01 g11888 ( .a(n15667), .b(n15366), .o(n15677) );
no02f01 g11889 ( .a(n15677), .b(n15655), .o(n15678) );
na02f01 g11890 ( .a(n15677), .b(n15655), .o(n15679) );
in01f01 g11891 ( .a(n15679), .o(n15680) );
no02f01 g11892 ( .a(n15680), .b(n15678), .o(n15681) );
oa12f01 g11893 ( .a(n15594), .b(n15681), .c(n15676), .o(n15682) );
oa12f01 g11894 ( .a(n15367), .b(n15654), .c(n15396), .o(n15683) );
in01f01 g11895 ( .a(n15683), .o(n15684) );
no02f01 g11896 ( .a(n15656), .b(n15378), .o(n15685) );
in01f01 g11897 ( .a(n15685), .o(n15686) );
no02f01 g11898 ( .a(n15686), .b(n15684), .o(n15687) );
no02f01 g11899 ( .a(n15685), .b(n15683), .o(n15688) );
no02f01 g11900 ( .a(n15688), .b(n15687), .o(n15689) );
na02f01 g11901 ( .a(n15689), .b(n15594), .o(n15690) );
na03f01 g11902 ( .a(n15690), .b(n15682), .c(n15666), .o(n15691) );
no04f01 g11903 ( .a(n15691), .b(n15651), .c(n15612), .d(n15609), .o(n15692) );
ao12f01 g11904 ( .a(n15594), .b(n15649), .c(n15621), .o(n15693) );
ao12f01 g11905 ( .a(n15594), .b(n15638), .c(n15633), .o(n15694) );
no02f01 g11906 ( .a(n15694), .b(n15693), .o(n15695) );
ao12f01 g11907 ( .a(n15594), .b(n15681), .c(n15676), .o(n15696) );
in01f01 g11908 ( .a(n15696), .o(n15697) );
ao12f01 g11909 ( .a(n15594), .b(n15689), .c(n15665), .o(n15698) );
in01f01 g11910 ( .a(n15698), .o(n15699) );
na03f01 g11911 ( .a(n15699), .b(n15697), .c(n15695), .o(n15700) );
no02f01 g11912 ( .a(n15700), .b(n15692), .o(n15701) );
no02f01 g11913 ( .a(n15488), .b(n15187), .o(n15702) );
in01f01 g11914 ( .a(n15398), .o(n15703) );
no02f01 g11915 ( .a(n15431), .b(n15703), .o(n15704) );
no02f01 g11916 ( .a(n15438), .b(n15187), .o(n15705) );
no02f01 g11917 ( .a(n15705), .b(n15440), .o(n15706) );
in01f01 g11918 ( .a(n15706), .o(n15707) );
no03f01 g11919 ( .a(n15707), .b(n15704), .c(n15702), .o(n15708) );
no02f01 g11920 ( .a(n15704), .b(n15702), .o(n15709) );
no02f01 g11921 ( .a(n15706), .b(n15709), .o(n15710) );
no02f01 g11922 ( .a(n15710), .b(n15708), .o(n15711) );
in01f01 g11923 ( .a(n15711), .o(n15712) );
no02f01 g11924 ( .a(n15712), .b(n15173), .o(n15713) );
no03f01 g11925 ( .a(n15440), .b(n15431), .c(n15703), .o(n15714) );
no03f01 g11926 ( .a(n15714), .b(n15705), .c(n15702), .o(n15715) );
no02f01 g11927 ( .a(n15408), .b(n15187), .o(n15716) );
no02f01 g11928 ( .a(n15716), .b(n15410), .o(n15717) );
no02f01 g11929 ( .a(n15717), .b(n15715), .o(n15718) );
na02f01 g11930 ( .a(n15717), .b(n15715), .o(n15719) );
in01f01 g11931 ( .a(n15719), .o(n15720) );
no02f01 g11932 ( .a(n15720), .b(n15718), .o(n15721) );
in01f01 g11933 ( .a(n15721), .o(n15722) );
no02f01 g11934 ( .a(n15722), .b(n15173), .o(n15723) );
no02f01 g11935 ( .a(n15429), .b(n15187), .o(n15724) );
no02f01 g11936 ( .a(n15430), .b(n15186), .o(n15725) );
in01f01 g11937 ( .a(n15725), .o(n15726) );
ao12f01 g11938 ( .a(n15724), .b(n15726), .c(n15398), .o(n15727) );
no02f01 g11939 ( .a(n15424), .b(n15186), .o(n15728) );
no02f01 g11940 ( .a(n15423), .b(n15187), .o(n15729) );
no02f01 g11941 ( .a(n15729), .b(n15728), .o(n15730) );
no02f01 g11942 ( .a(n15730), .b(n15727), .o(n15731) );
na02f01 g11943 ( .a(n15730), .b(n15727), .o(n15732) );
in01f01 g11944 ( .a(n15732), .o(n15733) );
no02f01 g11945 ( .a(n15733), .b(n15731), .o(n15734) );
in01f01 g11946 ( .a(n15734), .o(n15735) );
no02f01 g11947 ( .a(n15725), .b(n15724), .o(n15736) );
no02f01 g11948 ( .a(n15736), .b(n15703), .o(n15737) );
na02f01 g11949 ( .a(n15736), .b(n15703), .o(n15738) );
in01f01 g11950 ( .a(n15738), .o(n15739) );
no02f01 g11951 ( .a(n15739), .b(n15737), .o(n15740) );
in01f01 g11952 ( .a(n15740), .o(n15741) );
ao12f01 g11953 ( .a(n15173), .b(n15741), .c(n15735), .o(n15742) );
no03f01 g11954 ( .a(n15742), .b(n15723), .c(n15713), .o(n15743) );
in01f01 g11955 ( .a(n15743), .o(n15744) );
na02f01 g11956 ( .a(n15441), .b(n15398), .o(n15745) );
in01f01 g11957 ( .a(n15745), .o(n15746) );
no02f01 g11958 ( .a(n15489), .b(n15746), .o(n15747) );
in01f01 g11959 ( .a(n15747), .o(n15748) );
ao12f01 g11960 ( .a(n15485), .b(n15748), .c(n15461), .o(n15749) );
no02f01 g11961 ( .a(n15479), .b(n15187), .o(n15750) );
no02f01 g11962 ( .a(n15480), .b(n15186), .o(n15751) );
no02f01 g11963 ( .a(n15751), .b(n15750), .o(n15752) );
no02f01 g11964 ( .a(n15752), .b(n15749), .o(n15753) );
na02f01 g11965 ( .a(n15752), .b(n15749), .o(n15754) );
in01f01 g11966 ( .a(n15754), .o(n15755) );
no02f01 g11967 ( .a(n15755), .b(n15753), .o(n15756) );
in01f01 g11968 ( .a(n15756), .o(n15757) );
no02f01 g11969 ( .a(n15757), .b(n15173), .o(n15758) );
no02f01 g11970 ( .a(n15458), .b(n15187), .o(n15759) );
no02f01 g11971 ( .a(n15489), .b(n15759), .o(n15760) );
oa12f01 g11972 ( .a(n15760), .b(n15460), .c(n15745), .o(n15761) );
in01f01 g11973 ( .a(n15761), .o(n15762) );
no02f01 g11974 ( .a(n15451), .b(n15187), .o(n15763) );
no02f01 g11975 ( .a(n15763), .b(n15453), .o(n15764) );
no02f01 g11976 ( .a(n15764), .b(n15762), .o(n15765) );
na02f01 g11977 ( .a(n15764), .b(n15762), .o(n15766) );
in01f01 g11978 ( .a(n15766), .o(n15767) );
no02f01 g11979 ( .a(n15767), .b(n15765), .o(n15768) );
in01f01 g11980 ( .a(n15768), .o(n15769) );
no02f01 g11981 ( .a(n15759), .b(n15460), .o(n15770) );
no02f01 g11982 ( .a(n15770), .b(n15747), .o(n15771) );
na02f01 g11983 ( .a(n15770), .b(n15747), .o(n15772) );
in01f01 g11984 ( .a(n15772), .o(n15773) );
no02f01 g11985 ( .a(n15773), .b(n15771), .o(n15774) );
in01f01 g11986 ( .a(n15774), .o(n15775) );
ao12f01 g11987 ( .a(n15173), .b(n15775), .c(n15769), .o(n15776) );
in01f01 g11988 ( .a(n15750), .o(n15777) );
ao12f01 g11989 ( .a(n15751), .b(n15749), .c(n15777), .o(n15778) );
in01f01 g11990 ( .a(n15778), .o(n15779) );
no02f01 g11991 ( .a(n15472), .b(n15186), .o(n15780) );
no02f01 g11992 ( .a(n15471), .b(n15187), .o(n15781) );
no02f01 g11993 ( .a(n15781), .b(n15780), .o(n15782) );
no02f01 g11994 ( .a(n15782), .b(n15779), .o(n15783) );
na02f01 g11995 ( .a(n15782), .b(n15779), .o(n15784) );
in01f01 g11996 ( .a(n15784), .o(n15785) );
no02f01 g11997 ( .a(n15785), .b(n15783), .o(n15786) );
in01f01 g11998 ( .a(n15786), .o(n15787) );
no02f01 g11999 ( .a(n15787), .b(n15173), .o(n15788) );
no03f01 g12000 ( .a(n15788), .b(n15776), .c(n15758), .o(n15789) );
in01f01 g12001 ( .a(n15193), .o(n15790) );
ao12f01 g12002 ( .a(n15495), .b(n15492), .c(n15790), .o(n15791) );
in01f01 g12003 ( .a(n15791), .o(n15792) );
no02f01 g12004 ( .a(n15496), .b(n15194), .o(n15793) );
no02f01 g12005 ( .a(n15793), .b(n15792), .o(n15794) );
na02f01 g12006 ( .a(n15793), .b(n15792), .o(n15795) );
in01f01 g12007 ( .a(n15795), .o(n15796) );
no02f01 g12008 ( .a(n15796), .b(n15794), .o(n15797) );
in01f01 g12009 ( .a(n15797), .o(n15798) );
no02f01 g12010 ( .a(n15798), .b(n15173), .o(n15799) );
no02f01 g12011 ( .a(n15192), .b(n15187), .o(n15800) );
in01f01 g12012 ( .a(n15800), .o(n15801) );
no02f01 g12013 ( .a(n15494), .b(n15186), .o(n15802) );
ao12f01 g12014 ( .a(n15802), .b(n15492), .c(n15801), .o(n15803) );
in01f01 g12015 ( .a(n15803), .o(n15804) );
no02f01 g12016 ( .a(n15186), .b(n14845), .o(n15805) );
no02f01 g12017 ( .a(n15187), .b(n14519), .o(n15806) );
no02f01 g12018 ( .a(n15806), .b(n15805), .o(n15807) );
no02f01 g12019 ( .a(n15807), .b(n15804), .o(n15808) );
na02f01 g12020 ( .a(n15807), .b(n15804), .o(n15809) );
in01f01 g12021 ( .a(n15809), .o(n15810) );
no02f01 g12022 ( .a(n15810), .b(n15808), .o(n15811) );
in01f01 g12023 ( .a(n15811), .o(n15812) );
no02f01 g12024 ( .a(n15802), .b(n15800), .o(n15813) );
no02f01 g12025 ( .a(n15813), .b(n15492), .o(n15814) );
na02f01 g12026 ( .a(n15813), .b(n15492), .o(n15815) );
in01f01 g12027 ( .a(n15815), .o(n15816) );
no02f01 g12028 ( .a(n15816), .b(n15814), .o(n15817) );
in01f01 g12029 ( .a(n15817), .o(n15818) );
ao12f01 g12030 ( .a(n15173), .b(n15818), .c(n15812), .o(n15819) );
no02f01 g12031 ( .a(n15187), .b(n14538), .o(n15820) );
no02f01 g12032 ( .a(n15820), .b(n15498), .o(n15821) );
in01f01 g12033 ( .a(n15821), .o(n15822) );
no02f01 g12034 ( .a(n15496), .b(n15495), .o(n15823) );
na02f01 g12035 ( .a(n15490), .b(n15195), .o(n15824) );
ao12f01 g12036 ( .a(n15824), .b(n15823), .c(n15484), .o(n15825) );
in01f01 g12037 ( .a(n15825), .o(n15826) );
no02f01 g12038 ( .a(n15826), .b(n15822), .o(n15827) );
no02f01 g12039 ( .a(n15825), .b(n15821), .o(n15828) );
no02f01 g12040 ( .a(n15828), .b(n15827), .o(n15829) );
in01f01 g12041 ( .a(n15829), .o(n15830) );
no02f01 g12042 ( .a(n15830), .b(n15173), .o(n15831) );
no03f01 g12043 ( .a(n15831), .b(n15819), .c(n15799), .o(n15832) );
na02f01 g12044 ( .a(n15832), .b(n15789), .o(n15833) );
no03f01 g12045 ( .a(n15833), .b(n15744), .c(n15701), .o(n15834) );
ao12f01 g12046 ( .a(n15594), .b(n15721), .c(n15711), .o(n15835) );
no02f01 g12047 ( .a(n15741), .b(n15735), .o(n15836) );
no02f01 g12048 ( .a(n15836), .b(n15594), .o(n15837) );
no02f01 g12049 ( .a(n15837), .b(n15835), .o(n15838) );
no02f01 g12050 ( .a(n15775), .b(n15769), .o(n15839) );
no02f01 g12051 ( .a(n15839), .b(n15594), .o(n15840) );
in01f01 g12052 ( .a(n15840), .o(n15841) );
oa12f01 g12053 ( .a(n15173), .b(n15787), .c(n15757), .o(n15842) );
na03f01 g12054 ( .a(n15842), .b(n15841), .c(n15838), .o(n15843) );
ao12f01 g12055 ( .a(n15594), .b(n15817), .c(n15811), .o(n15844) );
ao12f01 g12056 ( .a(n15594), .b(n15829), .c(n15797), .o(n15845) );
no02f01 g12057 ( .a(n15845), .b(n15844), .o(n15846) );
in01f01 g12058 ( .a(n15846), .o(n15847) );
no02f01 g12059 ( .a(n15847), .b(n15843), .o(n15848) );
in01f01 g12060 ( .a(n15848), .o(n15849) );
no02f01 g12061 ( .a(n15508), .b(n15594), .o(n15850) );
no03f01 g12062 ( .a(n15850), .b(n15849), .c(n15834), .o(n15851) );
no02f01 g12063 ( .a(n15186), .b(n14795), .o(n15852) );
no02f01 g12064 ( .a(n15187), .b(n14500), .o(n15853) );
no02f01 g12065 ( .a(n15853), .b(n15852), .o(n15854) );
in01f01 g12066 ( .a(n15500), .o(n15855) );
in01f01 g12067 ( .a(n15503), .o(n15856) );
oa12f01 g12068 ( .a(n15856), .b(n15501), .c(n15855), .o(n15857) );
na02f01 g12069 ( .a(n15857), .b(n15854), .o(n15858) );
in01f01 g12070 ( .a(n15858), .o(n15859) );
no02f01 g12071 ( .a(n15857), .b(n15854), .o(n15860) );
no02f01 g12072 ( .a(n15860), .b(n15859), .o(n15861) );
no02f01 g12073 ( .a(n15861), .b(n15594), .o(n15862) );
in01f01 g12074 ( .a(n15861), .o(n15863) );
no02f01 g12075 ( .a(n15863), .b(n15173), .o(n15864) );
no02f01 g12076 ( .a(n15864), .b(n15862), .o(n15865) );
no03f01 g12077 ( .a(n15865), .b(n15851), .c(n15510), .o(n15866) );
in01f01 g12078 ( .a(n15510), .o(n15867) );
in01f01 g12079 ( .a(n15525), .o(n15868) );
in01f01 g12080 ( .a(n15541), .o(n15869) );
ao12f01 g12081 ( .a(n15546), .b(n15869), .c(n15539), .o(n15870) );
no02f01 g12082 ( .a(n15549), .b(n15163), .o(n15871) );
no02f01 g12083 ( .a(n15550), .b(n15115), .o(n15872) );
in01f01 g12084 ( .a(n15559), .o(n15873) );
oa12f01 g12085 ( .a(n15873), .b(n15872), .c(n15871), .o(n15874) );
na02f01 g12086 ( .a(n15114), .b(n15089), .o(n15875) );
na02f01 g12087 ( .a(n15114), .b(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n15876) );
in01f01 g12088 ( .a(n15573), .o(n15877) );
na03f01 g12089 ( .a(n15877), .b(n15876), .c(n15875), .o(n15878) );
no02f01 g12090 ( .a(n15878), .b(n15566), .o(n15879) );
na02f01 g12091 ( .a(n15878), .b(n15566), .o(n15880) );
na03f01 g12092 ( .a(n15162), .b(n15107), .c(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n15881) );
in01f01 g12093 ( .a(n15578), .o(n15882) );
na02f01 g12094 ( .a(n15882), .b(n15881), .o(n15883) );
ao12f01 g12095 ( .a(n15879), .b(n15883), .c(n15880), .o(n15884) );
no03f01 g12096 ( .a(n15873), .b(n15872), .c(n15871), .o(n15885) );
oa12f01 g12097 ( .a(n15874), .b(n15885), .c(n15884), .o(n15886) );
na03f01 g12098 ( .a(n15546), .b(n15869), .c(n15539), .o(n15887) );
ao12f01 g12099 ( .a(n15870), .b(n15887), .c(n15886), .o(n15888) );
no03f01 g12100 ( .a(n15528), .b(n15167), .c(n15158), .o(n15889) );
ao12f01 g12101 ( .a(n15526), .b(n15147), .c(n15142), .o(n15890) );
in01f01 g12102 ( .a(n15534), .o(n15891) );
no03f01 g12103 ( .a(n15891), .b(n15890), .c(n15889), .o(n15892) );
no02f01 g12104 ( .a(n15892), .b(n15888), .o(n15893) );
na03f01 g12105 ( .a(n15524), .b(n15516), .c(n15514), .o(n15894) );
oa12f01 g12106 ( .a(n15894), .b(n15893), .c(n15535), .o(n15895) );
oa12f01 g12107 ( .a(n15173), .b(n15611), .c(n15610), .o(n15896) );
na03f01 g12108 ( .a(n15896), .b(n15895), .c(n15868), .o(n15897) );
in01f01 g12109 ( .a(n15612), .o(n15898) );
in01f01 g12110 ( .a(n15621), .o(n15899) );
no02f01 g12111 ( .a(n15899), .b(n15173), .o(n15900) );
in01f01 g12112 ( .a(n15633), .o(n15901) );
in01f01 g12113 ( .a(n15638), .o(n15902) );
ao12f01 g12114 ( .a(n15173), .b(n15902), .c(n15901), .o(n15903) );
in01f01 g12115 ( .a(n15649), .o(n15904) );
no02f01 g12116 ( .a(n15904), .b(n15173), .o(n15905) );
no03f01 g12117 ( .a(n15905), .b(n15903), .c(n15900), .o(n15906) );
in01f01 g12118 ( .a(n15665), .o(n15907) );
no02f01 g12119 ( .a(n15907), .b(n15173), .o(n15908) );
in01f01 g12120 ( .a(n15676), .o(n15909) );
in01f01 g12121 ( .a(n15681), .o(n15910) );
ao12f01 g12122 ( .a(n15173), .b(n15910), .c(n15909), .o(n15911) );
in01f01 g12123 ( .a(n15689), .o(n15912) );
no02f01 g12124 ( .a(n15912), .b(n15173), .o(n15913) );
no03f01 g12125 ( .a(n15913), .b(n15911), .c(n15908), .o(n15914) );
na04f01 g12126 ( .a(n15914), .b(n15906), .c(n15898), .d(n15897), .o(n15915) );
in01f01 g12127 ( .a(n15700), .o(n15916) );
na02f01 g12128 ( .a(n15916), .b(n15915), .o(n15917) );
in01f01 g12129 ( .a(n15833), .o(n15918) );
na03f01 g12130 ( .a(n15918), .b(n15743), .c(n15917), .o(n15919) );
in01f01 g12131 ( .a(n15850), .o(n15920) );
na03f01 g12132 ( .a(n15920), .b(n15848), .c(n15919), .o(n15921) );
in01f01 g12133 ( .a(n15865), .o(n15922) );
ao12f01 g12134 ( .a(n15922), .b(n15921), .c(n15867), .o(n15923) );
oa12f01 g12135 ( .a(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .b(n15923), .c(n15866), .o(n15924) );
in01f01 g12136 ( .a(n15799), .o(n15925) );
in01f01 g12137 ( .a(n15789), .o(n15926) );
no02f01 g12138 ( .a(n15819), .b(n15926), .o(n15927) );
na04f01 g12139 ( .a(n15927), .b(n15925), .c(n15743), .d(n15917), .o(n15928) );
no02f01 g12140 ( .a(n15797), .b(n15594), .o(n15929) );
in01f01 g12141 ( .a(n15929), .o(n15930) );
no02f01 g12142 ( .a(n15844), .b(n15843), .o(n15931) );
na02f01 g12143 ( .a(n15931), .b(n15930), .o(n15932) );
in01f01 g12144 ( .a(n15932), .o(n15933) );
no02f01 g12145 ( .a(n15829), .b(n15594), .o(n15934) );
no02f01 g12146 ( .a(n15934), .b(n15831), .o(n15935) );
na03f01 g12147 ( .a(n15935), .b(n15933), .c(n15928), .o(n15936) );
in01f01 g12148 ( .a(n15927), .o(n15937) );
no04f01 g12149 ( .a(n15937), .b(n15799), .c(n15744), .d(n15701), .o(n15938) );
in01f01 g12150 ( .a(n15935), .o(n15939) );
oa12f01 g12151 ( .a(n15939), .b(n15932), .c(n15938), .o(n15940) );
na02f01 g12152 ( .a(n15940), .b(n15936), .o(n15941) );
no02f01 g12153 ( .a(n15850), .b(n15510), .o(n15942) );
in01f01 g12154 ( .a(n15942), .o(n15943) );
oa12f01 g12155 ( .a(n15943), .b(n15849), .c(n15834), .o(n15944) );
na03f01 g12156 ( .a(n15942), .b(n15848), .c(n15919), .o(n15945) );
na02f01 g12157 ( .a(n15945), .b(n15944), .o(n15946) );
oa12f01 g12158 ( .a(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .b(n15946), .c(n15941), .o(n15947) );
na02f01 g12159 ( .a(n15947), .b(n15924), .o(n15948) );
in01f01 g12160 ( .a(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .o(n15949) );
no02f01 g12161 ( .a(n15187), .b(n14549), .o(n15950) );
no02f01 g12162 ( .a(n15186), .b(n14778), .o(n15951) );
no02f01 g12163 ( .a(n15951), .b(n15950), .o(n15952) );
in01f01 g12164 ( .a(n15952), .o(n15953) );
no02f01 g12165 ( .a(n15852), .b(n15503), .o(n15954) );
in01f01 g12166 ( .a(n15954), .o(n15955) );
no02f01 g12167 ( .a(n15955), .b(n15500), .o(n15956) );
ao12f01 g12168 ( .a(n15187), .b(n14508), .c(n14500), .o(n15957) );
no03f01 g12169 ( .a(n15957), .b(n15956), .c(n15953), .o(n15958) );
no02f01 g12170 ( .a(n15957), .b(n15956), .o(n15959) );
no02f01 g12171 ( .a(n15959), .b(n15952), .o(n15960) );
no02f01 g12172 ( .a(n15960), .b(n15958), .o(n15961) );
in01f01 g12173 ( .a(n15961), .o(n15962) );
no02f01 g12174 ( .a(n15962), .b(n15173), .o(n15963) );
no02f01 g12175 ( .a(n15961), .b(n15594), .o(n15964) );
no02f01 g12176 ( .a(n15964), .b(n15963), .o(n15965) );
ao12f01 g12177 ( .a(n15594), .b(n15861), .c(n15508), .o(n15966) );
in01f01 g12178 ( .a(n15966), .o(n15967) );
no02f01 g12179 ( .a(n15861), .b(n15508), .o(n15968) );
no02f01 g12180 ( .a(n15968), .b(n15173), .o(n15969) );
in01f01 g12181 ( .a(n15969), .o(n15970) );
oa12f01 g12182 ( .a(n15970), .b(n15849), .c(n15834), .o(n15971) );
ao12f01 g12183 ( .a(n15965), .b(n15971), .c(n15967), .o(n15972) );
in01f01 g12184 ( .a(n15972), .o(n15973) );
na03f01 g12185 ( .a(n15971), .b(n15967), .c(n15965), .o(n15974) );
ao12f01 g12186 ( .a(n15949), .b(n15974), .c(n15973), .o(n15975) );
ao12f01 g12187 ( .a(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .b(n15974), .c(n15973), .o(n15976) );
no02f01 g12188 ( .a(n15976), .b(n15975), .o(n15977) );
no02f01 g12189 ( .a(n15977), .b(n15948), .o(n15978) );
na03f01 g12190 ( .a(n15922), .b(n15921), .c(n15867), .o(n15979) );
oa12f01 g12191 ( .a(n15865), .b(n15851), .c(n15510), .o(n15980) );
ao12f01 g12192 ( .a(n15949), .b(n15980), .c(n15979), .o(n15981) );
no03f01 g12193 ( .a(n15939), .b(n15932), .c(n15938), .o(n15982) );
ao12f01 g12194 ( .a(n15935), .b(n15933), .c(n15928), .o(n15983) );
no02f01 g12195 ( .a(n15983), .b(n15982), .o(n15984) );
ao12f01 g12196 ( .a(n15942), .b(n15848), .c(n15919), .o(n15985) );
no03f01 g12197 ( .a(n15943), .b(n15849), .c(n15834), .o(n15986) );
no02f01 g12198 ( .a(n15986), .b(n15985), .o(n15987) );
ao12f01 g12199 ( .a(n15949), .b(n15987), .c(n15984), .o(n15988) );
no02f01 g12200 ( .a(n15988), .b(n15981), .o(n15989) );
in01f01 g12201 ( .a(n15974), .o(n15990) );
oa12f01 g12202 ( .a(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .b(n15990), .c(n15972), .o(n15991) );
oa12f01 g12203 ( .a(n15949), .b(n15990), .c(n15972), .o(n15992) );
na02f01 g12204 ( .a(n15992), .b(n15991), .o(n15993) );
no02f01 g12205 ( .a(n15993), .b(n15989), .o(n15994) );
oa12f01 g12206 ( .a(delay_sub_ln23_0_unr25_stage9_stallmux_q), .b(n15830), .c(n15798), .o(n15995) );
in01f01 g12207 ( .a(n15995), .o(n15996) );
no02f01 g12208 ( .a(n15508), .b(n15089), .o(n15997) );
no02f01 g12209 ( .a(n15508), .b(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n15998) );
no02f01 g12210 ( .a(n15998), .b(n15997), .o(n15999) );
no02f01 g12211 ( .a(n15999), .b(n15996), .o(n16000) );
no03f01 g12212 ( .a(n15998), .b(n15997), .c(n15995), .o(n16001) );
in01f01 g12213 ( .a(n14851), .o(n16002) );
ao12f01 g12214 ( .a(n16002), .b(n14831), .c(n14830), .o(n16003) );
in01f01 g12215 ( .a(n14831), .o(n16004) );
no03f01 g12216 ( .a(n14851), .b(n16004), .c(n14829), .o(n16005) );
no02f01 g12217 ( .a(n16005), .b(n16003), .o(n16006) );
no03f01 g12218 ( .a(n16006), .b(n16001), .c(n16000), .o(n16007) );
ao12f01 g12219 ( .a(n15829), .b(n15798), .c(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n16008) );
no03f01 g12220 ( .a(n15830), .b(n15797), .c(n15089), .o(n16009) );
no03f01 g12221 ( .a(n14848), .b(n14846), .c(n14837), .o(n16010) );
in01f01 g12222 ( .a(n14837), .o(n16011) );
no02f01 g12223 ( .a(n14849), .b(n16011), .o(n16012) );
no02f01 g12224 ( .a(n16012), .b(n16010), .o(n16013) );
no02f01 g12225 ( .a(n16013), .b(n14841), .o(n16014) );
na02f01 g12226 ( .a(n16013), .b(n14841), .o(n16015) );
in01f01 g12227 ( .a(n16015), .o(n16016) );
no02f01 g12228 ( .a(n16016), .b(n16014), .o(n16017) );
no03f01 g12229 ( .a(n16017), .b(n16009), .c(n16008), .o(n16018) );
in01f01 g12230 ( .a(n16018), .o(n16019) );
oa12f01 g12231 ( .a(n16017), .b(n16009), .c(n16008), .o(n16020) );
in01f01 g12232 ( .a(n16020), .o(n16021) );
no02f01 g12233 ( .a(n15798), .b(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n16022) );
no02f01 g12234 ( .a(n15798), .b(n15089), .o(n16023) );
no02f01 g12235 ( .a(n16023), .b(n16022), .o(n16024) );
in01f01 g12236 ( .a(n16024), .o(n16025) );
no02f01 g12237 ( .a(n14840), .b(n14845), .o(n16026) );
na02f01 g12238 ( .a(n14840), .b(n14845), .o(n16027) );
in01f01 g12239 ( .a(n16027), .o(n16028) );
no02f01 g12240 ( .a(n16028), .b(n16026), .o(n16029) );
no02f01 g12241 ( .a(n16029), .b(n16025), .o(n16030) );
oa12f01 g12242 ( .a(n16019), .b(n16030), .c(n16021), .o(n16031) );
oa12f01 g12243 ( .a(n16006), .b(n16001), .c(n16000), .o(n16032) );
ao12f01 g12244 ( .a(n16007), .b(n16032), .c(n16031), .o(n16033) );
in01f01 g12245 ( .a(n15998), .o(n16034) );
in01f01 g12246 ( .a(n15997), .o(n16035) );
na02f01 g12247 ( .a(n16035), .b(n15995), .o(n16036) );
na02f01 g12248 ( .a(n16036), .b(n16034), .o(n16037) );
no02f01 g12249 ( .a(n15861), .b(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n16038) );
no02f01 g12250 ( .a(n15861), .b(n15089), .o(n16039) );
oa12f01 g12251 ( .a(n16037), .b(n16039), .c(n16038), .o(n16040) );
in01f01 g12252 ( .a(n16040), .o(n16041) );
no03f01 g12253 ( .a(n16039), .b(n16038), .c(n16037), .o(n16042) );
ao22f01 g12254 ( .a(n14854), .b(n14818), .c(n14852), .d(n14830), .o(n16043) );
in01f01 g12255 ( .a(n14854), .o(n16044) );
no03f01 g12256 ( .a(n16044), .b(n14853), .c(n14817), .o(n16045) );
no02f01 g12257 ( .a(n16045), .b(n16043), .o(n16046) );
no03f01 g12258 ( .a(n16046), .b(n16042), .c(n16041), .o(n16047) );
in01f01 g12259 ( .a(n16042), .o(n16048) );
in01f01 g12260 ( .a(n16046), .o(n16049) );
ao12f01 g12261 ( .a(n16049), .b(n16048), .c(n16040), .o(n16050) );
no02f01 g12262 ( .a(n16050), .b(n16047), .o(n16051) );
no02f01 g12263 ( .a(n16051), .b(n16033), .o(n16052) );
na02f01 g12264 ( .a(n16051), .b(n16033), .o(n16053) );
in01f01 g12265 ( .a(n16053), .o(n16054) );
no02f01 g12266 ( .a(n16054), .b(n16052), .o(n16055) );
no03f01 g12267 ( .a(n16055), .b(n15994), .c(n15978), .o(n16056) );
ao12f01 g12268 ( .a(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .b(n15980), .c(n15979), .o(n16057) );
oa12f01 g12269 ( .a(n15947), .b(n16057), .c(n15981), .o(n16058) );
oa12f01 g12270 ( .a(n15949), .b(n15923), .c(n15866), .o(n16059) );
na03f01 g12271 ( .a(n16059), .b(n15988), .c(n15924), .o(n16060) );
in01f01 g12272 ( .a(n16031), .o(n16061) );
in01f01 g12273 ( .a(n16032), .o(n16062) );
no02f01 g12274 ( .a(n16062), .b(n16007), .o(n16063) );
no02f01 g12275 ( .a(n16063), .b(n16061), .o(n16064) );
na02f01 g12276 ( .a(n16063), .b(n16061), .o(n16065) );
in01f01 g12277 ( .a(n16065), .o(n16066) );
no02f01 g12278 ( .a(n16066), .b(n16064), .o(n16067) );
in01f01 g12279 ( .a(n16067), .o(n16068) );
na03f01 g12280 ( .a(n16068), .b(n16060), .c(n16058), .o(n16069) );
ao12f01 g12281 ( .a(n16068), .b(n16060), .c(n16058), .o(n16070) );
ao12f01 g12282 ( .a(n15987), .b(n15941), .c(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .o(n16071) );
no03f01 g12283 ( .a(n15946), .b(n15984), .c(n15949), .o(n16072) );
no04f01 g12284 ( .a(n16029), .b(n16025), .c(n16021), .d(n16018), .o(n16073) );
ao12f01 g12285 ( .a(n16030), .b(n16020), .c(n16019), .o(n16074) );
no02f01 g12286 ( .a(n16074), .b(n16073), .o(n16075) );
oa12f01 g12287 ( .a(n16075), .b(n16072), .c(n16071), .o(n16076) );
na02f01 g12288 ( .a(n15984), .b(n15949), .o(n16077) );
na02f01 g12289 ( .a(n15984), .b(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .o(n16078) );
no02f01 g12290 ( .a(n16029), .b(n16024), .o(n16079) );
in01f01 g12291 ( .a(n16029), .o(n16080) );
no02f01 g12292 ( .a(n16080), .b(n16025), .o(n16081) );
no02f01 g12293 ( .a(n16081), .b(n16079), .o(n16082) );
in01f01 g12294 ( .a(n16082), .o(n16083) );
na03f01 g12295 ( .a(n16083), .b(n16078), .c(n16077), .o(n16084) );
no03f01 g12296 ( .a(n16075), .b(n16072), .c(n16071), .o(n16085) );
ao12f01 g12297 ( .a(n16085), .b(n16084), .c(n16076), .o(n16086) );
oa12f01 g12298 ( .a(n16069), .b(n16086), .c(n16070), .o(n16087) );
oa12f01 g12299 ( .a(n16055), .b(n15994), .c(n15978), .o(n16088) );
ao12f01 g12300 ( .a(n16056), .b(n16088), .c(n16087), .o(n16089) );
na02f01 g12301 ( .a(n15991), .b(n15989), .o(n16090) );
no02f01 g12302 ( .a(n15186), .b(n14864), .o(n16091) );
no02f01 g12303 ( .a(n15187), .b(n14491), .o(n16092) );
no02f01 g12304 ( .a(n16092), .b(n16091), .o(n16093) );
in01f01 g12305 ( .a(n16093), .o(n16094) );
no03f01 g12306 ( .a(n15955), .b(n15951), .c(n15500), .o(n16095) );
no02f01 g12307 ( .a(n15957), .b(n15950), .o(n16096) );
in01f01 g12308 ( .a(n16096), .o(n16097) );
no03f01 g12309 ( .a(n16097), .b(n16095), .c(n16094), .o(n16098) );
no02f01 g12310 ( .a(n16097), .b(n16095), .o(n16099) );
no02f01 g12311 ( .a(n16099), .b(n16093), .o(n16100) );
no02f01 g12312 ( .a(n16100), .b(n16098), .o(n16101) );
no02f01 g12313 ( .a(n16101), .b(n15594), .o(n16102) );
in01f01 g12314 ( .a(n16101), .o(n16103) );
no02f01 g12315 ( .a(n16103), .b(n15173), .o(n16104) );
no02f01 g12316 ( .a(n16104), .b(n16102), .o(n16105) );
in01f01 g12317 ( .a(n16105), .o(n16106) );
no02f01 g12318 ( .a(n15744), .b(n15701), .o(n16107) );
ao12f01 g12319 ( .a(n15843), .b(n15789), .c(n16107), .o(n16108) );
no02f01 g12320 ( .a(n15969), .b(n15963), .o(n16109) );
na02f01 g12321 ( .a(n16109), .b(n15832), .o(n16110) );
no02f01 g12322 ( .a(n16110), .b(n16108), .o(n16111) );
na02f01 g12323 ( .a(n15967), .b(n15961), .o(n16112) );
ao12f01 g12324 ( .a(n15847), .b(n16112), .c(n15173), .o(n16113) );
in01f01 g12325 ( .a(n16113), .o(n16114) );
no03f01 g12326 ( .a(n16114), .b(n16111), .c(n16106), .o(n16115) );
in01f01 g12327 ( .a(n16115), .o(n16116) );
oa12f01 g12328 ( .a(n16106), .b(n16114), .c(n16111), .o(n16117) );
ao12f01 g12329 ( .a(n15949), .b(n16117), .c(n16116), .o(n16118) );
ao12f01 g12330 ( .a(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .b(n16117), .c(n16116), .o(n16119) );
no02f01 g12331 ( .a(n16119), .b(n16118), .o(n16120) );
no02f01 g12332 ( .a(n16120), .b(n16090), .o(n16121) );
no02f01 g12333 ( .a(n15975), .b(n15948), .o(n16122) );
no03f01 g12334 ( .a(n16119), .b(n16118), .c(n16122), .o(n16123) );
no02f01 g12335 ( .a(n16050), .b(n16033), .o(n16124) );
no02f01 g12336 ( .a(n16124), .b(n16047), .o(n16125) );
na02f01 g12337 ( .a(n15863), .b(n15089), .o(n16126) );
na02f01 g12338 ( .a(n15861), .b(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n16127) );
ao22f01 g12339 ( .a(n16127), .b(n16126), .c(n16036), .d(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n16128) );
ao12f01 g12340 ( .a(n16128), .b(n16037), .c(n15089), .o(n16129) );
no02f01 g12341 ( .a(n15961), .b(n15089), .o(n16130) );
no02f01 g12342 ( .a(n15961), .b(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n16131) );
no02f01 g12343 ( .a(n16131), .b(n16130), .o(n16132) );
na02f01 g12344 ( .a(n16132), .b(n16129), .o(n16133) );
in01f01 g12345 ( .a(n16133), .o(n16134) );
no02f01 g12346 ( .a(n16132), .b(n16129), .o(n16135) );
ao22f01 g12347 ( .a(n14857), .b(n14806), .c(n14855), .d(n14818), .o(n16136) );
in01f01 g12348 ( .a(n14857), .o(n16137) );
no03f01 g12349 ( .a(n16137), .b(n14856), .c(n14805), .o(n16138) );
no02f01 g12350 ( .a(n16138), .b(n16136), .o(n16139) );
no03f01 g12351 ( .a(n16139), .b(n16135), .c(n16134), .o(n16140) );
in01f01 g12352 ( .a(n16135), .o(n16141) );
in01f01 g12353 ( .a(n16139), .o(n16142) );
ao12f01 g12354 ( .a(n16142), .b(n16141), .c(n16133), .o(n16143) );
no02f01 g12355 ( .a(n16143), .b(n16140), .o(n16144) );
no02f01 g12356 ( .a(n16144), .b(n16125), .o(n16145) );
na02f01 g12357 ( .a(n16144), .b(n16125), .o(n16146) );
in01f01 g12358 ( .a(n16146), .o(n16147) );
no02f01 g12359 ( .a(n16147), .b(n16145), .o(n16148) );
oa12f01 g12360 ( .a(n16148), .b(n16123), .c(n16121), .o(n16149) );
in01f01 g12361 ( .a(n16149), .o(n16150) );
no03f01 g12362 ( .a(n16119), .b(n16118), .c(n16122), .o(n16151) );
na02f01 g12363 ( .a(n16117), .b(n16116), .o(n16152) );
in01f01 g12364 ( .a(n16152), .o(n16153) );
no03f01 g12365 ( .a(n16153), .b(n16090), .c(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .o(n16154) );
no02f01 g12366 ( .a(n16154), .b(n16151), .o(n16155) );
no02f01 g12367 ( .a(n16143), .b(n16125), .o(n16156) );
no02f01 g12368 ( .a(n16156), .b(n16140), .o(n16157) );
in01f01 g12369 ( .a(n16131), .o(n16158) );
no02f01 g12370 ( .a(n16130), .b(n16129), .o(n16159) );
in01f01 g12371 ( .a(n16159), .o(n16160) );
no02f01 g12372 ( .a(n16101), .b(n15089), .o(n16161) );
no02f01 g12373 ( .a(n16101), .b(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n16162) );
no02f01 g12374 ( .a(n16162), .b(n16161), .o(n16163) );
ao12f01 g12375 ( .a(n16163), .b(n16160), .c(n16158), .o(n16164) );
in01f01 g12376 ( .a(n16163), .o(n16165) );
no03f01 g12377 ( .a(n16165), .b(n16159), .c(n16131), .o(n16166) );
no02f01 g12378 ( .a(n16166), .b(n16164), .o(n16167) );
in01f01 g12379 ( .a(n14861), .o(n16168) );
no02f01 g12380 ( .a(n16168), .b(n14794), .o(n16169) );
no02f01 g12381 ( .a(n16169), .b(n14860), .o(n16170) );
na02f01 g12382 ( .a(n16169), .b(n14860), .o(n16171) );
in01f01 g12383 ( .a(n16171), .o(n16172) );
no02f01 g12384 ( .a(n16172), .b(n16170), .o(n16173) );
in01f01 g12385 ( .a(n16173), .o(n16174) );
no02f01 g12386 ( .a(n16174), .b(n16167), .o(n16175) );
na02f01 g12387 ( .a(n16174), .b(n16167), .o(n16176) );
in01f01 g12388 ( .a(n16176), .o(n16177) );
no02f01 g12389 ( .a(n16177), .b(n16175), .o(n16178) );
no02f01 g12390 ( .a(n16178), .b(n16157), .o(n16179) );
na02f01 g12391 ( .a(n16178), .b(n16157), .o(n16180) );
in01f01 g12392 ( .a(n16180), .o(n16181) );
no02f01 g12393 ( .a(n16181), .b(n16179), .o(n16182) );
in01f01 g12394 ( .a(n16182), .o(n16183) );
no02f01 g12395 ( .a(n16183), .b(n16155), .o(n16184) );
oa22f01 g12396 ( .a(n16174), .b(n16167), .c(n16156), .d(n16140), .o(n16185) );
in01f01 g12397 ( .a(n16185), .o(n16186) );
no02f01 g12398 ( .a(n16186), .b(n16177), .o(n16187) );
in01f01 g12399 ( .a(n16187), .o(n16188) );
no02f01 g12400 ( .a(n16101), .b(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n16189) );
no02f01 g12401 ( .a(n16103), .b(n15089), .o(n16190) );
no02f01 g12402 ( .a(n16190), .b(n16189), .o(n16191) );
na03f01 g12403 ( .a(n16129), .b(n15961), .c(n15089), .o(n16192) );
ao22f01 g12404 ( .a(n16192), .b(n16191), .c(n16159), .d(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n16193) );
in01f01 g12405 ( .a(n16193), .o(n16194) );
no02f01 g12406 ( .a(n14887), .b(n14875), .o(n16195) );
in01f01 g12407 ( .a(n16195), .o(n16196) );
no02f01 g12408 ( .a(n16196), .b(n14862), .o(n16197) );
in01f01 g12409 ( .a(n14862), .o(n16198) );
no02f01 g12410 ( .a(n16195), .b(n16198), .o(n16199) );
no02f01 g12411 ( .a(n16199), .b(n16197), .o(n16200) );
in01f01 g12412 ( .a(n16200), .o(n16201) );
no02f01 g12413 ( .a(n16201), .b(n16194), .o(n16202) );
no02f01 g12414 ( .a(n16200), .b(n16193), .o(n16203) );
no02f01 g12415 ( .a(n16203), .b(n16202), .o(n16204) );
in01f01 g12416 ( .a(n16204), .o(n16205) );
no02f01 g12417 ( .a(n16205), .b(n16188), .o(n16206) );
no02f01 g12418 ( .a(n16204), .b(n16187), .o(n16207) );
no02f01 g12419 ( .a(n16207), .b(n16206), .o(n16208) );
in01f01 g12420 ( .a(n16208), .o(n16209) );
in01f01 g12421 ( .a(n16202), .o(n16210) );
ao12f01 g12422 ( .a(n16203), .b(n16210), .c(n16188), .o(n16211) );
in01f01 g12423 ( .a(n16211), .o(n16212) );
ao12f01 g12424 ( .a(n14875), .b(n14886), .c(n16198), .o(n16213) );
no02f01 g12425 ( .a(n14892), .b(n14885), .o(n16214) );
in01f01 g12426 ( .a(n16214), .o(n16215) );
no02f01 g12427 ( .a(n16215), .b(n16213), .o(n16216) );
na02f01 g12428 ( .a(n16215), .b(n16213), .o(n16217) );
in01f01 g12429 ( .a(n16217), .o(n16218) );
no02f01 g12430 ( .a(n16218), .b(n16216), .o(n16219) );
in01f01 g12431 ( .a(n16219), .o(n16220) );
no02f01 g12432 ( .a(n16220), .b(n16194), .o(n16221) );
no02f01 g12433 ( .a(n16219), .b(n16193), .o(n16222) );
no02f01 g12434 ( .a(n16222), .b(n16221), .o(n16223) );
in01f01 g12435 ( .a(n16223), .o(n16224) );
no02f01 g12436 ( .a(n16224), .b(n16212), .o(n16225) );
no02f01 g12437 ( .a(n16223), .b(n16211), .o(n16226) );
no02f01 g12438 ( .a(n16226), .b(n16225), .o(n16227) );
in01f01 g12439 ( .a(n16227), .o(n16228) );
ao12f01 g12440 ( .a(n16155), .b(n16228), .c(n16209), .o(n16229) );
no04f01 g12441 ( .a(n16229), .b(n16184), .c(n16150), .d(n16089), .o(n16230) );
no03f01 g12442 ( .a(n16182), .b(n16154), .c(n16151), .o(n16231) );
no03f01 g12443 ( .a(n16148), .b(n16123), .c(n16121), .o(n16232) );
no02f01 g12444 ( .a(n16232), .b(n16231), .o(n16233) );
oa12f01 g12445 ( .a(n16155), .b(n16228), .c(n16209), .o(n16234) );
na02f01 g12446 ( .a(n16234), .b(n16233), .o(n16235) );
no02f01 g12447 ( .a(n16235), .b(n16230), .o(n16236) );
no02f01 g12448 ( .a(n14920), .b(n14552), .o(n16237) );
no02f01 g12449 ( .a(n14921), .b(n14553), .o(n16238) );
in01f01 g12450 ( .a(n16238), .o(n16239) );
ao12f01 g12451 ( .a(n16237), .b(n16239), .c(n14893), .o(n16240) );
no02f01 g12452 ( .a(n14915), .b(n14553), .o(n16241) );
no02f01 g12453 ( .a(n14914), .b(n14552), .o(n16242) );
no02f01 g12454 ( .a(n16242), .b(n16241), .o(n16243) );
no02f01 g12455 ( .a(n16243), .b(n16240), .o(n16244) );
na02f01 g12456 ( .a(n16243), .b(n16240), .o(n16245) );
in01f01 g12457 ( .a(n16245), .o(n16246) );
no02f01 g12458 ( .a(n16246), .b(n16244), .o(n16247) );
no02f01 g12459 ( .a(n16238), .b(n16237), .o(n16248) );
in01f01 g12460 ( .a(n16248), .o(n16249) );
no02f01 g12461 ( .a(n16249), .b(n14893), .o(n16250) );
in01f01 g12462 ( .a(n14893), .o(n16251) );
no02f01 g12463 ( .a(n16248), .b(n16251), .o(n16252) );
no02f01 g12464 ( .a(n16252), .b(n16250), .o(n16253) );
ao12f01 g12465 ( .a(n16193), .b(n16253), .c(n16247), .o(n16254) );
in01f01 g12466 ( .a(n16247), .o(n16255) );
in01f01 g12467 ( .a(n16253), .o(n16256) );
ao12f01 g12468 ( .a(n16194), .b(n16256), .c(n16255), .o(n16257) );
ao12f01 g12469 ( .a(n16193), .b(n16219), .c(n16200), .o(n16258) );
in01f01 g12470 ( .a(n16258), .o(n16259) );
na03f01 g12471 ( .a(n16259), .b(n16185), .c(n16176), .o(n16260) );
in01f01 g12472 ( .a(n16260), .o(n16261) );
ao12f01 g12473 ( .a(n16194), .b(n16220), .c(n16201), .o(n16262) );
no02f01 g12474 ( .a(n16262), .b(n16261), .o(n16263) );
in01f01 g12475 ( .a(n16263), .o(n16264) );
no02f01 g12476 ( .a(n16264), .b(n16257), .o(n16265) );
in01f01 g12477 ( .a(n14922), .o(n16266) );
ao12f01 g12478 ( .a(n14979), .b(n16266), .c(n14893), .o(n16267) );
no02f01 g12479 ( .a(n14901), .b(n14552), .o(n16268) );
no02f01 g12480 ( .a(n16268), .b(n14903), .o(n16269) );
no02f01 g12481 ( .a(n16269), .b(n16267), .o(n16270) );
na02f01 g12482 ( .a(n16269), .b(n16267), .o(n16271) );
in01f01 g12483 ( .a(n16271), .o(n16272) );
no02f01 g12484 ( .a(n16272), .b(n16270), .o(n16273) );
na02f01 g12485 ( .a(n16273), .b(n16193), .o(n16274) );
in01f01 g12486 ( .a(n16274), .o(n16275) );
no02f01 g12487 ( .a(n16273), .b(n16193), .o(n16276) );
no02f01 g12488 ( .a(n16276), .b(n16275), .o(n16277) );
in01f01 g12489 ( .a(n16277), .o(n16278) );
no03f01 g12490 ( .a(n16278), .b(n16265), .c(n16254), .o(n16279) );
no02f01 g12491 ( .a(n16265), .b(n16254), .o(n16280) );
no02f01 g12492 ( .a(n16277), .b(n16280), .o(n16281) );
no02f01 g12493 ( .a(n16281), .b(n16279), .o(n16282) );
in01f01 g12494 ( .a(n16282), .o(n16283) );
no02f01 g12495 ( .a(n16283), .b(n16155), .o(n16284) );
no02f01 g12496 ( .a(n16253), .b(n16193), .o(n16285) );
no02f01 g12497 ( .a(n16256), .b(n16194), .o(n16286) );
in01f01 g12498 ( .a(n16286), .o(n16287) );
ao12f01 g12499 ( .a(n16285), .b(n16287), .c(n16263), .o(n16288) );
no02f01 g12500 ( .a(n16255), .b(n16194), .o(n16289) );
no02f01 g12501 ( .a(n16247), .b(n16193), .o(n16290) );
no02f01 g12502 ( .a(n16290), .b(n16289), .o(n16291) );
no02f01 g12503 ( .a(n16291), .b(n16288), .o(n16292) );
na02f01 g12504 ( .a(n16291), .b(n16288), .o(n16293) );
in01f01 g12505 ( .a(n16293), .o(n16294) );
no02f01 g12506 ( .a(n16294), .b(n16292), .o(n16295) );
no02f01 g12507 ( .a(n16286), .b(n16285), .o(n16296) );
in01f01 g12508 ( .a(n16296), .o(n16297) );
no02f01 g12509 ( .a(n16297), .b(n16263), .o(n16298) );
no02f01 g12510 ( .a(n16296), .b(n16264), .o(n16299) );
no02f01 g12511 ( .a(n16299), .b(n16298), .o(n16300) );
no02f01 g12512 ( .a(n16300), .b(n16295), .o(n16301) );
no02f01 g12513 ( .a(n16301), .b(n16155), .o(n16302) );
na02f01 g12514 ( .a(n16274), .b(n16265), .o(n16303) );
no02f01 g12515 ( .a(n16276), .b(n16254), .o(n16304) );
na02f01 g12516 ( .a(n16304), .b(n16303), .o(n16305) );
in01f01 g12517 ( .a(n16305), .o(n16306) );
no03f01 g12518 ( .a(n14922), .b(n14903), .c(n16251), .o(n16307) );
no03f01 g12519 ( .a(n16307), .b(n14979), .c(n16268), .o(n16308) );
no02f01 g12520 ( .a(n14930), .b(n14552), .o(n16309) );
no02f01 g12521 ( .a(n16309), .b(n14932), .o(n16310) );
no02f01 g12522 ( .a(n16310), .b(n16308), .o(n16311) );
na02f01 g12523 ( .a(n16310), .b(n16308), .o(n16312) );
in01f01 g12524 ( .a(n16312), .o(n16313) );
no02f01 g12525 ( .a(n16313), .b(n16311), .o(n16314) );
in01f01 g12526 ( .a(n16314), .o(n16315) );
no02f01 g12527 ( .a(n16315), .b(n16194), .o(n16316) );
no02f01 g12528 ( .a(n16314), .b(n16193), .o(n16317) );
no02f01 g12529 ( .a(n16317), .b(n16316), .o(n16318) );
no02f01 g12530 ( .a(n16318), .b(n16306), .o(n16319) );
na02f01 g12531 ( .a(n16318), .b(n16306), .o(n16320) );
in01f01 g12532 ( .a(n16320), .o(n16321) );
no02f01 g12533 ( .a(n16321), .b(n16319), .o(n16322) );
in01f01 g12534 ( .a(n16322), .o(n16323) );
no02f01 g12535 ( .a(n16323), .b(n16155), .o(n16324) );
no03f01 g12536 ( .a(n16324), .b(n16302), .c(n16284), .o(n16325) );
in01f01 g12537 ( .a(n16325), .o(n16326) );
oa12f01 g12538 ( .a(n16120), .b(n16118), .c(n16090), .o(n16327) );
na03f01 g12539 ( .a(n16152), .b(n16122), .c(n15949), .o(n16328) );
na02f01 g12540 ( .a(n16328), .b(n16327), .o(n16329) );
no03f01 g12541 ( .a(n16316), .b(n16275), .c(n16257), .o(n16330) );
in01f01 g12542 ( .a(n16330), .o(n16331) );
no02f01 g12543 ( .a(n16331), .b(n16264), .o(n16332) );
ao12f01 g12544 ( .a(n16193), .b(n16314), .c(n16273), .o(n16333) );
no02f01 g12545 ( .a(n16333), .b(n16254), .o(n16334) );
in01f01 g12546 ( .a(n16334), .o(n16335) );
no02f01 g12547 ( .a(n16335), .b(n16332), .o(n16336) );
no02f01 g12548 ( .a(n14981), .b(n14935), .o(n16337) );
in01f01 g12549 ( .a(n16337), .o(n16338) );
no02f01 g12550 ( .a(n14952), .b(n14552), .o(n16339) );
na02f01 g12551 ( .a(n14952), .b(n14552), .o(n16340) );
in01f01 g12552 ( .a(n16340), .o(n16341) );
no02f01 g12553 ( .a(n16341), .b(n16339), .o(n16342) );
in01f01 g12554 ( .a(n16342), .o(n16343) );
no02f01 g12555 ( .a(n16343), .b(n16338), .o(n16344) );
no02f01 g12556 ( .a(n16342), .b(n16337), .o(n16345) );
no02f01 g12557 ( .a(n16345), .b(n16344), .o(n16346) );
na02f01 g12558 ( .a(n16346), .b(n16193), .o(n16347) );
in01f01 g12559 ( .a(n16347), .o(n16348) );
no02f01 g12560 ( .a(n16346), .b(n16193), .o(n16349) );
no02f01 g12561 ( .a(n16349), .b(n16348), .o(n16350) );
no02f01 g12562 ( .a(n16350), .b(n16336), .o(n16351) );
na02f01 g12563 ( .a(n16350), .b(n16336), .o(n16352) );
in01f01 g12564 ( .a(n16352), .o(n16353) );
no02f01 g12565 ( .a(n16353), .b(n16351), .o(n16354) );
na02f01 g12566 ( .a(n16354), .b(n16329), .o(n16355) );
in01f01 g12567 ( .a(n16355), .o(n16356) );
na02f01 g12568 ( .a(n16347), .b(n16332), .o(n16357) );
no02f01 g12569 ( .a(n16349), .b(n16335), .o(n16358) );
na02f01 g12570 ( .a(n16358), .b(n16357), .o(n16359) );
in01f01 g12571 ( .a(n16359), .o(n16360) );
ao12f01 g12572 ( .a(n16339), .b(n16340), .c(n16338), .o(n16361) );
in01f01 g12573 ( .a(n14945), .o(n16362) );
no02f01 g12574 ( .a(n16362), .b(n14553), .o(n16363) );
no02f01 g12575 ( .a(n14945), .b(n14552), .o(n16364) );
no02f01 g12576 ( .a(n16364), .b(n16363), .o(n16365) );
no02f01 g12577 ( .a(n16365), .b(n16361), .o(n16366) );
na02f01 g12578 ( .a(n16365), .b(n16361), .o(n16367) );
in01f01 g12579 ( .a(n16367), .o(n16368) );
no02f01 g12580 ( .a(n16368), .b(n16366), .o(n16369) );
in01f01 g12581 ( .a(n16369), .o(n16370) );
no02f01 g12582 ( .a(n16370), .b(n16194), .o(n16371) );
no02f01 g12583 ( .a(n16369), .b(n16193), .o(n16372) );
no02f01 g12584 ( .a(n16372), .b(n16371), .o(n16373) );
no02f01 g12585 ( .a(n16373), .b(n16360), .o(n16374) );
na02f01 g12586 ( .a(n16373), .b(n16360), .o(n16375) );
in01f01 g12587 ( .a(n16375), .o(n16376) );
no02f01 g12588 ( .a(n16376), .b(n16374), .o(n16377) );
na02f01 g12589 ( .a(n16377), .b(n16329), .o(n16378) );
in01f01 g12590 ( .a(n16378), .o(n16379) );
no02f01 g12591 ( .a(n16379), .b(n16356), .o(n16380) );
in01f01 g12592 ( .a(n16380), .o(n16381) );
ao12f01 g12593 ( .a(n16193), .b(n16369), .c(n16346), .o(n16382) );
no02f01 g12594 ( .a(n16382), .b(n16335), .o(n16383) );
oa12f01 g12595 ( .a(n16383), .b(n16371), .c(n16357), .o(n16384) );
no02f01 g12596 ( .a(n16337), .b(n14954), .o(n16385) );
no02f01 g12597 ( .a(n16385), .b(n14982), .o(n16386) );
no02f01 g12598 ( .a(n14961), .b(n14552), .o(n16387) );
no02f01 g12599 ( .a(n16387), .b(n14963), .o(n16388) );
no02f01 g12600 ( .a(n16388), .b(n16386), .o(n16389) );
na02f01 g12601 ( .a(n16388), .b(n16386), .o(n16390) );
in01f01 g12602 ( .a(n16390), .o(n16391) );
no02f01 g12603 ( .a(n16391), .b(n16389), .o(n16392) );
in01f01 g12604 ( .a(n16392), .o(n16393) );
no02f01 g12605 ( .a(n16393), .b(n16194), .o(n16394) );
no02f01 g12606 ( .a(n16392), .b(n16193), .o(n16395) );
no02f01 g12607 ( .a(n16395), .b(n16394), .o(n16396) );
in01f01 g12608 ( .a(n16396), .o(n16397) );
no02f01 g12609 ( .a(n16397), .b(n16384), .o(n16398) );
in01f01 g12610 ( .a(n16384), .o(n16399) );
no02f01 g12611 ( .a(n16396), .b(n16399), .o(n16400) );
no02f01 g12612 ( .a(n16400), .b(n16398), .o(n16401) );
in01f01 g12613 ( .a(n16401), .o(n16402) );
no02f01 g12614 ( .a(n16402), .b(n16155), .o(n16403) );
no02f01 g12615 ( .a(n16395), .b(n16384), .o(n16404) );
no02f01 g12616 ( .a(n16404), .b(n16394), .o(n16405) );
in01f01 g12617 ( .a(n16387), .o(n16406) );
ao12f01 g12618 ( .a(n14963), .b(n16386), .c(n16406), .o(n16407) );
no02f01 g12619 ( .a(n14973), .b(n14552), .o(n16408) );
no02f01 g12620 ( .a(n16408), .b(n14975), .o(n16409) );
in01f01 g12621 ( .a(n16409), .o(n16410) );
no02f01 g12622 ( .a(n16410), .b(n16407), .o(n16411) );
na02f01 g12623 ( .a(n16410), .b(n16407), .o(n16412) );
in01f01 g12624 ( .a(n16412), .o(n16413) );
no02f01 g12625 ( .a(n16413), .b(n16411), .o(n16414) );
in01f01 g12626 ( .a(n16414), .o(n16415) );
no02f01 g12627 ( .a(n16415), .b(n16194), .o(n16416) );
no02f01 g12628 ( .a(n16414), .b(n16193), .o(n16417) );
no02f01 g12629 ( .a(n16417), .b(n16416), .o(n16418) );
in01f01 g12630 ( .a(n16418), .o(n16419) );
no02f01 g12631 ( .a(n16419), .b(n16405), .o(n16420) );
na02f01 g12632 ( .a(n16419), .b(n16405), .o(n16421) );
in01f01 g12633 ( .a(n16421), .o(n16422) );
no02f01 g12634 ( .a(n16422), .b(n16420), .o(n16423) );
na02f01 g12635 ( .a(n16423), .b(n16329), .o(n16424) );
in01f01 g12636 ( .a(n16424), .o(n16425) );
no02f01 g12637 ( .a(n16425), .b(n16403), .o(n16426) );
in01f01 g12638 ( .a(n16426), .o(n16427) );
no04f01 g12639 ( .a(n16427), .b(n16381), .c(n16326), .d(n16236), .o(n16428) );
in01f01 g12640 ( .a(n16295), .o(n16429) );
in01f01 g12641 ( .a(n16300), .o(n16430) );
no02f01 g12642 ( .a(n16430), .b(n16429), .o(n16431) );
in01f01 g12643 ( .a(n16431), .o(n16432) );
na02f01 g12644 ( .a(n16432), .b(n16155), .o(n16433) );
oa12f01 g12645 ( .a(n16155), .b(n16323), .c(n16283), .o(n16434) );
na02f01 g12646 ( .a(n16434), .b(n16433), .o(n16435) );
ao12f01 g12647 ( .a(n16329), .b(n16377), .c(n16354), .o(n16436) );
no02f01 g12648 ( .a(n16436), .b(n16435), .o(n16437) );
ao12f01 g12649 ( .a(n16329), .b(n16423), .c(n16401), .o(n16438) );
in01f01 g12650 ( .a(n16438), .o(n16439) );
na02f01 g12651 ( .a(n16439), .b(n16437), .o(n16440) );
no02f01 g12652 ( .a(n16440), .b(n16428), .o(n16441) );
no02f01 g12653 ( .a(n14990), .b(n14553), .o(n16442) );
no02f01 g12654 ( .a(n14713), .b(n14552), .o(n16443) );
no02f01 g12655 ( .a(n16443), .b(n16442), .o(n16444) );
in01f01 g12656 ( .a(n16444), .o(n16445) );
no02f01 g12657 ( .a(n16445), .b(n15099), .o(n16446) );
in01f01 g12658 ( .a(n15099), .o(n16447) );
no02f01 g12659 ( .a(n16444), .b(n16447), .o(n16448) );
no02f01 g12660 ( .a(n16448), .b(n16446), .o(n16449) );
no02f01 g12661 ( .a(n16449), .b(n16193), .o(n16450) );
in01f01 g12662 ( .a(n16262), .o(n16451) );
no04f01 g12663 ( .a(n16416), .b(n16394), .c(n16371), .d(n16348), .o(n16452) );
na04f01 g12664 ( .a(n16452), .b(n16330), .c(n16451), .d(n16260), .o(n16453) );
ao12f01 g12665 ( .a(n16193), .b(n16414), .c(n16392), .o(n16454) );
no03f01 g12666 ( .a(n16454), .b(n16382), .c(n16335), .o(n16455) );
na02f01 g12667 ( .a(n16455), .b(n16453), .o(n16456) );
in01f01 g12668 ( .a(n16449), .o(n16457) );
no02f01 g12669 ( .a(n16457), .b(n16194), .o(n16458) );
in01f01 g12670 ( .a(n16458), .o(n16459) );
ao12f01 g12671 ( .a(n16450), .b(n16459), .c(n16456), .o(n16460) );
in01f01 g12672 ( .a(n16460), .o(n16461) );
in01f01 g12673 ( .a(n16442), .o(n16462) );
ao12f01 g12674 ( .a(n16443), .b(n16462), .c(n15099), .o(n16463) );
in01f01 g12675 ( .a(n16463), .o(n16464) );
no02f01 g12676 ( .a(n14989), .b(n14553), .o(n16465) );
no02f01 g12677 ( .a(n14707), .b(n14552), .o(n16466) );
no02f01 g12678 ( .a(n16466), .b(n16465), .o(n16467) );
in01f01 g12679 ( .a(n16467), .o(n16468) );
no02f01 g12680 ( .a(n16468), .b(n16464), .o(n16469) );
no02f01 g12681 ( .a(n16467), .b(n16463), .o(n16470) );
no02f01 g12682 ( .a(n16470), .b(n16469), .o(n16471) );
in01f01 g12683 ( .a(n16471), .o(n16472) );
no02f01 g12684 ( .a(n16472), .b(n16194), .o(n16473) );
no02f01 g12685 ( .a(n16471), .b(n16193), .o(n16474) );
no02f01 g12686 ( .a(n16474), .b(n16473), .o(n16475) );
in01f01 g12687 ( .a(n16475), .o(n16476) );
no02f01 g12688 ( .a(n16476), .b(n16461), .o(n16477) );
no02f01 g12689 ( .a(n16475), .b(n16460), .o(n16478) );
no02f01 g12690 ( .a(n16478), .b(n16477), .o(n16479) );
in01f01 g12691 ( .a(n16479), .o(n16480) );
in01f01 g12692 ( .a(n16456), .o(n16481) );
no02f01 g12693 ( .a(n16458), .b(n16450), .o(n16482) );
no02f01 g12694 ( .a(n16482), .b(n16481), .o(n16483) );
na02f01 g12695 ( .a(n16482), .b(n16481), .o(n16484) );
in01f01 g12696 ( .a(n16484), .o(n16485) );
no02f01 g12697 ( .a(n16485), .b(n16483), .o(n16486) );
in01f01 g12698 ( .a(n16486), .o(n16487) );
ao12f01 g12699 ( .a(n16155), .b(n16487), .c(n16480), .o(n16488) );
no02f01 g12700 ( .a(n16488), .b(n16441), .o(n16489) );
no02f01 g12701 ( .a(n16473), .b(n16458), .o(n16490) );
in01f01 g12702 ( .a(n16490), .o(n16491) );
no02f01 g12703 ( .a(n16491), .b(n16481), .o(n16492) );
ao12f01 g12704 ( .a(n16193), .b(n16471), .c(n16449), .o(n16493) );
no02f01 g12705 ( .a(n16493), .b(n16492), .o(n16494) );
no02f01 g12706 ( .a(n14991), .b(n16447), .o(n16495) );
no02f01 g12707 ( .a(n16495), .b(n14714), .o(n16496) );
no02f01 g12708 ( .a(n14722), .b(n14552), .o(n16497) );
no02f01 g12709 ( .a(n14986), .b(n16497), .o(n16498) );
no02f01 g12710 ( .a(n16498), .b(n16496), .o(n16499) );
na02f01 g12711 ( .a(n16498), .b(n16496), .o(n16500) );
in01f01 g12712 ( .a(n16500), .o(n16501) );
no02f01 g12713 ( .a(n16501), .b(n16499), .o(n16502) );
na02f01 g12714 ( .a(n16502), .b(n16193), .o(n16503) );
in01f01 g12715 ( .a(n16503), .o(n16504) );
no02f01 g12716 ( .a(n16502), .b(n16193), .o(n16505) );
no02f01 g12717 ( .a(n16505), .b(n16504), .o(n16506) );
no02f01 g12718 ( .a(n16506), .b(n16494), .o(n16507) );
na02f01 g12719 ( .a(n16506), .b(n16494), .o(n16508) );
in01f01 g12720 ( .a(n16508), .o(n16509) );
no02f01 g12721 ( .a(n16509), .b(n16507), .o(n16510) );
in01f01 g12722 ( .a(n16510), .o(n16511) );
no02f01 g12723 ( .a(n16511), .b(n16155), .o(n16512) );
in01f01 g12724 ( .a(n16512), .o(n16513) );
na02f01 g12725 ( .a(n16513), .b(n16489), .o(n16514) );
ao12f01 g12726 ( .a(n16329), .b(n16486), .c(n16479), .o(n16515) );
no02f01 g12727 ( .a(n16510), .b(n16329), .o(n16516) );
no02f01 g12728 ( .a(n16516), .b(n16515), .o(n16517) );
na02f01 g12729 ( .a(n16503), .b(n16492), .o(n16518) );
no02f01 g12730 ( .a(n16505), .b(n16493), .o(n16519) );
na02f01 g12731 ( .a(n16519), .b(n16518), .o(n16520) );
na02f01 g12732 ( .a(n16495), .b(n14985), .o(n16521) );
no02f01 g12733 ( .a(n16497), .b(n14714), .o(n16522) );
na02f01 g12734 ( .a(n16522), .b(n16521), .o(n16523) );
in01f01 g12735 ( .a(n16523), .o(n16524) );
no02f01 g12736 ( .a(n14731), .b(n14552), .o(n16525) );
no02f01 g12737 ( .a(n16525), .b(n14988), .o(n16526) );
no02f01 g12738 ( .a(n16526), .b(n16524), .o(n16527) );
na02f01 g12739 ( .a(n16526), .b(n16524), .o(n16528) );
in01f01 g12740 ( .a(n16528), .o(n16529) );
no02f01 g12741 ( .a(n16529), .b(n16527), .o(n16530) );
in01f01 g12742 ( .a(n16530), .o(n16531) );
no02f01 g12743 ( .a(n16531), .b(n16194), .o(n16532) );
no02f01 g12744 ( .a(n16530), .b(n16193), .o(n16533) );
no02f01 g12745 ( .a(n16533), .b(n16532), .o(n16534) );
in01f01 g12746 ( .a(n16534), .o(n16535) );
no02f01 g12747 ( .a(n16535), .b(n16520), .o(n16536) );
na02f01 g12748 ( .a(n16535), .b(n16520), .o(n16537) );
in01f01 g12749 ( .a(n16537), .o(n16538) );
no02f01 g12750 ( .a(n16538), .b(n16536), .o(n16539) );
no02f01 g12751 ( .a(n16539), .b(n16329), .o(n16540) );
in01f01 g12752 ( .a(n16539), .o(n16541) );
no02f01 g12753 ( .a(n16541), .b(n16155), .o(n16542) );
no02f01 g12754 ( .a(n16542), .b(n16540), .o(n16543) );
na03f01 g12755 ( .a(n16543), .b(n16517), .c(n16514), .o(n16544) );
na02f01 g12756 ( .a(n16517), .b(n16514), .o(n16545) );
in01f01 g12757 ( .a(n16543), .o(n16546) );
na02f01 g12758 ( .a(n16546), .b(n16545), .o(n16547) );
na02f01 g12759 ( .a(n16547), .b(n16544), .o(n258) );
in01f01 g12760 ( .a(n_44365), .o(n16549) );
no02f01 g12761 ( .a(n16549), .b(delay_xor_ln21_unr12_stage5_stallmux_q_14_), .o(n16550) );
no02f01 g12762 ( .a(n16549), .b(delay_xor_ln21_unr12_stage5_stallmux_q_6_), .o(n16551) );
no02f01 g12763 ( .a(n16549), .b(delay_xor_ln21_unr12_stage5_stallmux_q_5_), .o(n16552) );
in01f01 g12764 ( .a(n16552), .o(n16553) );
in01f01 g12765 ( .a(n_44847), .o(n16554) );
na02f01 g12766 ( .a(n_44365), .b(n16554), .o(n16555) );
in01f01 g12767 ( .a(n_44721), .o(n16556) );
na02f01 g12768 ( .a(n_44365), .b(n16556), .o(n16557) );
no02f01 g12769 ( .a(n16549), .b(delay_xor_ln21_unr12_stage5_stallmux_q_2_), .o(n16558) );
in01f01 g12770 ( .a(n16558), .o(n16559) );
na03f01 g12771 ( .a(n16559), .b(n16557), .c(n16555), .o(n16560) );
no02f01 g12772 ( .a(n16549), .b(delay_xor_ln21_unr12_stage5_stallmux_q_4_), .o(n16561) );
no02f01 g12773 ( .a(n16549), .b(delay_xor_ln21_unr12_stage5_stallmux_q_3_), .o(n16562) );
no03f01 g12774 ( .a(n16562), .b(n16561), .c(n16560), .o(n16563) );
na02f01 g12775 ( .a(n16563), .b(n16553), .o(n16564) );
no02f01 g12776 ( .a(n16564), .b(n16551), .o(n16565) );
in01f01 g12777 ( .a(n16565), .o(n16566) );
no02f01 g12778 ( .a(n16549), .b(delay_xor_ln21_unr12_stage5_stallmux_q_7_), .o(n16567) );
no02f01 g12779 ( .a(n16567), .b(n16566), .o(n16568) );
in01f01 g12780 ( .a(n16568), .o(n16569) );
no02f01 g12781 ( .a(n16549), .b(delay_xor_ln21_unr12_stage5_stallmux_q_8_), .o(n16570) );
no02f01 g12782 ( .a(n16570), .b(n16569), .o(n16571) );
no02f01 g12783 ( .a(n16549), .b(delay_xor_ln21_unr12_stage5_stallmux_q_11_), .o(n16572) );
no02f01 g12784 ( .a(delay_xor_ln21_unr12_stage5_stallmux_q_9_), .b(n16549), .o(n16573) );
no02f01 g12785 ( .a(n16549), .b(delay_xor_ln21_unr12_stage5_stallmux_q_10_), .o(n16574) );
no02f01 g12786 ( .a(n16574), .b(n16573), .o(n16575) );
in01f01 g12787 ( .a(n16575), .o(n16576) );
no02f01 g12788 ( .a(n16576), .b(n16572), .o(n16577) );
na02f01 g12789 ( .a(n16577), .b(n16571), .o(n16578) );
no02f01 g12790 ( .a(n16549), .b(delay_xor_ln21_unr12_stage5_stallmux_q_13_), .o(n16579) );
no02f01 g12791 ( .a(n16549), .b(delay_xor_ln21_unr12_stage5_stallmux_q_12_), .o(n16580) );
no02f01 g12792 ( .a(n16580), .b(n16579), .o(n16581) );
in01f01 g12793 ( .a(n16581), .o(n16582) );
no02f01 g12794 ( .a(n16582), .b(n16578), .o(n16583) );
in01f01 g12795 ( .a(n16583), .o(n16584) );
no02f01 g12796 ( .a(n16584), .b(n16550), .o(n16585) );
in01f01 g12797 ( .a(n16585), .o(n16586) );
no02f01 g12798 ( .a(n16549), .b(delay_xor_ln21_unr12_stage5_stallmux_q_15_), .o(n16587) );
in01f01 g12799 ( .a(n16587), .o(n16588) );
na02f01 g12800 ( .a(n16549), .b(delay_xor_ln21_unr12_stage5_stallmux_q_15_), .o(n16589) );
na02f01 g12801 ( .a(n16589), .b(n16588), .o(n16590) );
in01f01 g12802 ( .a(n16590), .o(n16591) );
no02f01 g12803 ( .a(n16591), .b(n16586), .o(n16592) );
no02f01 g12804 ( .a(n16590), .b(n16585), .o(n16593) );
no02f01 g12805 ( .a(n16593), .b(n16592), .o(n16594) );
no02f01 g12806 ( .a(n16594), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_15_), .o(n16595) );
in01f01 g12807 ( .a(n16595), .o(n16596) );
na02f01 g12808 ( .a(n16549), .b(delay_xor_ln21_unr12_stage5_stallmux_q_13_), .o(n16597) );
in01f01 g12809 ( .a(n16597), .o(n16598) );
no02f01 g12810 ( .a(n16598), .b(n16579), .o(n16599) );
no02f01 g12811 ( .a(n16580), .b(n16578), .o(n16600) );
in01f01 g12812 ( .a(n16600), .o(n16601) );
in01f01 g12813 ( .a(n16571), .o(n16602) );
no02f01 g12814 ( .a(n16576), .b(n16602), .o(n16603) );
no03f01 g12815 ( .a(n16599), .b(n16580), .c(n16572), .o(n16604) );
ao22f01 g12816 ( .a(n16604), .b(n16603), .c(n16601), .d(n16599), .o(n16605) );
no02f01 g12817 ( .a(n16605), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_13_), .o(n16606) );
in01f01 g12818 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_12_), .o(n16607) );
na02f01 g12819 ( .a(n16549), .b(delay_xor_ln21_unr12_stage5_stallmux_q_12_), .o(n16608) );
in01f01 g12820 ( .a(n16608), .o(n16609) );
no02f01 g12821 ( .a(n16609), .b(n16580), .o(n16610) );
no02f01 g12822 ( .a(n16610), .b(n16578), .o(n16611) );
na02f01 g12823 ( .a(n16610), .b(n16578), .o(n16612) );
in01f01 g12824 ( .a(n16612), .o(n16613) );
no02f01 g12825 ( .a(n16613), .b(n16611), .o(n16614) );
in01f01 g12826 ( .a(n16614), .o(n16615) );
no02f01 g12827 ( .a(n16615), .b(n16607), .o(n16616) );
in01f01 g12828 ( .a(n16603), .o(n16617) );
na02f01 g12829 ( .a(n16549), .b(delay_xor_ln21_unr12_stage5_stallmux_q_11_), .o(n16618) );
in01f01 g12830 ( .a(n16618), .o(n16619) );
no02f01 g12831 ( .a(n16619), .b(n16572), .o(n16620) );
no02f01 g12832 ( .a(n16620), .b(n16617), .o(n16621) );
na02f01 g12833 ( .a(n16620), .b(n16617), .o(n16622) );
in01f01 g12834 ( .a(n16622), .o(n16623) );
no02f01 g12835 ( .a(n16623), .b(n16621), .o(n16624) );
no02f01 g12836 ( .a(n16624), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_11_), .o(n16625) );
in01f01 g12837 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_10_), .o(n16626) );
in01f01 g12838 ( .a(n16573), .o(n16627) );
na02f01 g12839 ( .a(n16549), .b(delay_xor_ln21_unr12_stage5_stallmux_q_10_), .o(n16628) );
in01f01 g12840 ( .a(n16628), .o(n16629) );
no02f01 g12841 ( .a(n16629), .b(n16574), .o(n16630) );
in01f01 g12842 ( .a(n16630), .o(n16631) );
no03f01 g12843 ( .a(n16570), .b(n16567), .c(n16566), .o(n16632) );
ao12f01 g12844 ( .a(n16631), .b(n16632), .c(n16627), .o(n16633) );
no03f01 g12845 ( .a(n16630), .b(n16573), .c(n16602), .o(n16634) );
no02f01 g12846 ( .a(n16634), .b(n16633), .o(n16635) );
in01f01 g12847 ( .a(n16635), .o(n16636) );
no02f01 g12848 ( .a(n16636), .b(n16626), .o(n16637) );
na02f01 g12849 ( .a(delay_xor_ln21_unr12_stage5_stallmux_q_9_), .b(n16549), .o(n16638) );
na02f01 g12850 ( .a(n16638), .b(n16627), .o(n16639) );
no02f01 g12851 ( .a(n16639), .b(n16632), .o(n16640) );
ao12f01 g12852 ( .a(n16640), .b(n16639), .c(n16571), .o(n16641) );
no02f01 g12853 ( .a(n16641), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_9_), .o(n16642) );
in01f01 g12854 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_8_), .o(n16643) );
na02f01 g12855 ( .a(n16549), .b(delay_xor_ln21_unr12_stage5_stallmux_q_8_), .o(n16644) );
in01f01 g12856 ( .a(n16644), .o(n16645) );
no02f01 g12857 ( .a(n16645), .b(n16570), .o(n16646) );
no02f01 g12858 ( .a(n16646), .b(n16567), .o(n16647) );
ao22f01 g12859 ( .a(n16647), .b(n16565), .c(n16646), .d(n16569), .o(n16648) );
in01f01 g12860 ( .a(n16648), .o(n16649) );
no02f01 g12861 ( .a(n16649), .b(n16643), .o(n16650) );
na02f01 g12862 ( .a(n16549), .b(delay_xor_ln21_unr12_stage5_stallmux_q_7_), .o(n16651) );
in01f01 g12863 ( .a(n16651), .o(n16652) );
no02f01 g12864 ( .a(n16652), .b(n16567), .o(n16653) );
no03f01 g12865 ( .a(n16653), .b(n16552), .c(n16551), .o(n16654) );
ao22f01 g12866 ( .a(n16654), .b(n16563), .c(n16653), .d(n16566), .o(n16655) );
no02f01 g12867 ( .a(n16655), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_7_), .o(n16656) );
in01f01 g12868 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_6_), .o(n16657) );
na02f01 g12869 ( .a(n16549), .b(delay_xor_ln21_unr12_stage5_stallmux_q_6_), .o(n16658) );
in01f01 g12870 ( .a(n16658), .o(n16659) );
no02f01 g12871 ( .a(n16659), .b(n16551), .o(n16660) );
na02f01 g12872 ( .a(n16660), .b(n16564), .o(n16661) );
no02f01 g12873 ( .a(n16660), .b(n16564), .o(n16662) );
in01f01 g12874 ( .a(n16662), .o(n16663) );
na02f01 g12875 ( .a(n16663), .b(n16661), .o(n16664) );
no02f01 g12876 ( .a(n16664), .b(n16657), .o(n16665) );
na02f01 g12877 ( .a(n16549), .b(delay_xor_ln21_unr12_stage5_stallmux_q_5_), .o(n16666) );
na02f01 g12878 ( .a(n16666), .b(n16553), .o(n16667) );
no02f01 g12879 ( .a(n16667), .b(n16563), .o(n16668) );
na02f01 g12880 ( .a(n16667), .b(n16563), .o(n16669) );
in01f01 g12881 ( .a(n16669), .o(n16670) );
no02f01 g12882 ( .a(n16670), .b(n16668), .o(n16671) );
no02f01 g12883 ( .a(n16671), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_5_), .o(n16672) );
na02f01 g12884 ( .a(n16549), .b(delay_xor_ln21_unr12_stage5_stallmux_q_4_), .o(n16673) );
in01f01 g12885 ( .a(n16673), .o(n16674) );
no02f01 g12886 ( .a(n16674), .b(n16561), .o(n16675) );
no02f01 g12887 ( .a(n16549), .b(n_44847), .o(n16676) );
no02f01 g12888 ( .a(n16549), .b(n_44721), .o(n16677) );
no02f01 g12889 ( .a(n16677), .b(n16676), .o(n16678) );
in01f01 g12890 ( .a(n16678), .o(n16679) );
no02f01 g12891 ( .a(n16679), .b(n16558), .o(n16680) );
in01f01 g12892 ( .a(n16562), .o(n16681) );
na02f01 g12893 ( .a(n16680), .b(n16681), .o(n16682) );
no02f01 g12894 ( .a(n16675), .b(n16562), .o(n16683) );
ao22f01 g12895 ( .a(n16683), .b(n16680), .c(n16682), .d(n16675), .o(n16684) );
na02f01 g12896 ( .a(n16684), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_4_), .o(n16685) );
in01f01 g12897 ( .a(n16685), .o(n16686) );
in01f01 g12898 ( .a(n16680), .o(n16687) );
in01f01 g12899 ( .a(delay_xor_ln21_unr12_stage5_stallmux_q_3_), .o(n16688) );
no02f01 g12900 ( .a(n_44365), .b(n16688), .o(n16689) );
no02f01 g12901 ( .a(n16689), .b(n16562), .o(n16690) );
no02f01 g12902 ( .a(n16690), .b(n16560), .o(n16691) );
ao12f01 g12903 ( .a(n16691), .b(n16690), .c(n16687), .o(n16692) );
no02f01 g12904 ( .a(n16692), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_3_), .o(n16693) );
in01f01 g12905 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_2_), .o(n16694) );
na02f01 g12906 ( .a(n16549), .b(delay_xor_ln21_unr12_stage5_stallmux_q_2_), .o(n16695) );
in01f01 g12907 ( .a(n16695), .o(n16696) );
no02f01 g12908 ( .a(n16696), .b(n16558), .o(n16697) );
na02f01 g12909 ( .a(n16697), .b(n16679), .o(n16698) );
na02f01 g12910 ( .a(n16695), .b(n16559), .o(n16699) );
na02f01 g12911 ( .a(n16699), .b(n16678), .o(n16700) );
na02f01 g12912 ( .a(n16700), .b(n16698), .o(n16701) );
no02f01 g12913 ( .a(n16701), .b(n16694), .o(n16702) );
in01f01 g12914 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_1_), .o(n16703) );
no02f01 g12915 ( .a(n_44365), .b(n16556), .o(n16704) );
oa12f01 g12916 ( .a(n16555), .b(n16704), .c(n16677), .o(n16705) );
oa12f01 g12917 ( .a(n16705), .b(n16677), .c(n16555), .o(n16706) );
no02f01 g12918 ( .a(n16706), .b(n16703), .o(n16707) );
na02f01 g12919 ( .a(n16706), .b(n16703), .o(n16708) );
no02f01 g12920 ( .a(n_44365), .b(n_44847), .o(n16709) );
no02f01 g12921 ( .a(n16549), .b(n16554), .o(n16710) );
no02f01 g12922 ( .a(n16710), .b(n16709), .o(n16711) );
in01f01 g12923 ( .a(n16711), .o(n16712) );
no02f01 g12924 ( .a(n16712), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_0_), .o(n16713) );
in01f01 g12925 ( .a(n16713), .o(n16714) );
ao12f01 g12926 ( .a(n16707), .b(n16714), .c(n16708), .o(n16715) );
ao12f01 g12927 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_2_), .b(n16700), .c(n16698), .o(n16716) );
no02f01 g12928 ( .a(n16716), .b(n16715), .o(n16717) );
in01f01 g12929 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_3_), .o(n16718) );
no03f01 g12930 ( .a(n16689), .b(n16680), .c(n16562), .o(n16719) );
no03f01 g12931 ( .a(n16691), .b(n16719), .c(n16718), .o(n16720) );
no03f01 g12932 ( .a(n16720), .b(n16717), .c(n16702), .o(n16721) );
no02f01 g12933 ( .a(n16684), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_4_), .o(n16722) );
no03f01 g12934 ( .a(n16722), .b(n16721), .c(n16693), .o(n16723) );
in01f01 g12935 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_5_), .o(n16724) );
no03f01 g12936 ( .a(n16670), .b(n16668), .c(n16724), .o(n16725) );
no03f01 g12937 ( .a(n16725), .b(n16723), .c(n16686), .o(n16726) );
ao12f01 g12938 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_6_), .b(n16663), .c(n16661), .o(n16727) );
no03f01 g12939 ( .a(n16727), .b(n16726), .c(n16672), .o(n16728) );
na02f01 g12940 ( .a(n16655), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_7_), .o(n16729) );
in01f01 g12941 ( .a(n16729), .o(n16730) );
no03f01 g12942 ( .a(n16730), .b(n16728), .c(n16665), .o(n16731) );
no02f01 g12943 ( .a(n16648), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_8_), .o(n16732) );
no03f01 g12944 ( .a(n16732), .b(n16731), .c(n16656), .o(n16733) );
na02f01 g12945 ( .a(n16641), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_9_), .o(n16734) );
in01f01 g12946 ( .a(n16734), .o(n16735) );
no03f01 g12947 ( .a(n16735), .b(n16733), .c(n16650), .o(n16736) );
no02f01 g12948 ( .a(n16635), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_10_), .o(n16737) );
no03f01 g12949 ( .a(n16737), .b(n16736), .c(n16642), .o(n16738) );
in01f01 g12950 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_11_), .o(n16739) );
no03f01 g12951 ( .a(n16623), .b(n16621), .c(n16739), .o(n16740) );
no03f01 g12952 ( .a(n16740), .b(n16738), .c(n16637), .o(n16741) );
no02f01 g12953 ( .a(n16614), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_12_), .o(n16742) );
no03f01 g12954 ( .a(n16742), .b(n16741), .c(n16625), .o(n16743) );
na02f01 g12955 ( .a(n16605), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_13_), .o(n16744) );
in01f01 g12956 ( .a(n16744), .o(n16745) );
no03f01 g12957 ( .a(n16745), .b(n16743), .c(n16616), .o(n16746) );
na02f01 g12958 ( .a(n16549), .b(delay_xor_ln21_unr12_stage5_stallmux_q_14_), .o(n16747) );
in01f01 g12959 ( .a(n16747), .o(n16748) );
no02f01 g12960 ( .a(n16748), .b(n16550), .o(n16749) );
no03f01 g12961 ( .a(n16749), .b(n16582), .c(n16578), .o(n16750) );
ao12f01 g12962 ( .a(n16750), .b(n16749), .c(n16584), .o(n16751) );
no02f01 g12963 ( .a(n16751), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_14_), .o(n16752) );
no03f01 g12964 ( .a(n16752), .b(n16746), .c(n16606), .o(n16753) );
na02f01 g12965 ( .a(n16594), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_15_), .o(n16754) );
in01f01 g12966 ( .a(n16754), .o(n16755) );
na02f01 g12967 ( .a(n16751), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_14_), .o(n16756) );
in01f01 g12968 ( .a(n16756), .o(n16757) );
no02f01 g12969 ( .a(n16757), .b(n16755), .o(n16758) );
in01f01 g12970 ( .a(n16758), .o(n16759) );
oa12f01 g12971 ( .a(n16596), .b(n16759), .c(n16753), .o(n16760) );
no02f01 g12972 ( .a(n16587), .b(n16586), .o(n16761) );
no02f01 g12973 ( .a(n16549), .b(delay_xor_ln21_unr12_stage5_stallmux_q_16_), .o(n16762) );
in01f01 g12974 ( .a(n16762), .o(n16763) );
na02f01 g12975 ( .a(n16549), .b(delay_xor_ln21_unr12_stage5_stallmux_q_16_), .o(n16764) );
na02f01 g12976 ( .a(n16764), .b(n16763), .o(n16765) );
no02f01 g12977 ( .a(n16765), .b(n16761), .o(n16766) );
na02f01 g12978 ( .a(n16765), .b(n16761), .o(n16767) );
in01f01 g12979 ( .a(n16767), .o(n16768) );
no02f01 g12980 ( .a(n16768), .b(n16766), .o(n16769) );
no02f01 g12981 ( .a(n16769), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_16_), .o(n16770) );
no02f01 g12982 ( .a(n16770), .b(n16760), .o(n16771) );
na02f01 g12983 ( .a(n16769), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_16_), .o(n16772) );
in01f01 g12984 ( .a(n16772), .o(n16773) );
no02f01 g12985 ( .a(n16773), .b(n16771), .o(n16774) );
na02f01 g12986 ( .a(n16763), .b(n16761), .o(n16775) );
no02f01 g12987 ( .a(n16549), .b(delay_xor_ln21_unr12_stage5_stallmux_q_17_), .o(n16776) );
in01f01 g12988 ( .a(n16776), .o(n16777) );
na02f01 g12989 ( .a(n16549), .b(delay_xor_ln21_unr12_stage5_stallmux_q_17_), .o(n16778) );
na02f01 g12990 ( .a(n16778), .b(n16777), .o(n16779) );
in01f01 g12991 ( .a(n16779), .o(n16780) );
no02f01 g12992 ( .a(n16780), .b(n16775), .o(n16781) );
na02f01 g12993 ( .a(n16780), .b(n16775), .o(n16782) );
in01f01 g12994 ( .a(n16782), .o(n16783) );
no02f01 g12995 ( .a(n16783), .b(n16781), .o(n16784) );
no02f01 g12996 ( .a(n16784), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_17_), .o(n16785) );
na02f01 g12997 ( .a(n16784), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_17_), .o(n16786) );
in01f01 g12998 ( .a(n16786), .o(n16787) );
no02f01 g12999 ( .a(n16787), .b(n16785), .o(n16788) );
in01f01 g13000 ( .a(n16606), .o(n16789) );
in01f01 g13001 ( .a(n16616), .o(n16790) );
in01f01 g13002 ( .a(n16625), .o(n16791) );
in01f01 g13003 ( .a(n16637), .o(n16792) );
in01f01 g13004 ( .a(n16642), .o(n16793) );
in01f01 g13005 ( .a(n16650), .o(n16794) );
in01f01 g13006 ( .a(n16656), .o(n16795) );
in01f01 g13007 ( .a(n16665), .o(n16796) );
in01f01 g13008 ( .a(n16672), .o(n16797) );
in01f01 g13009 ( .a(n16693), .o(n16798) );
in01f01 g13010 ( .a(n16702), .o(n16799) );
na02f01 g13011 ( .a(n16549), .b(n_44721), .o(n16800) );
ao12f01 g13012 ( .a(n16676), .b(n16800), .c(n16557), .o(n16801) );
ao12f01 g13013 ( .a(n16801), .b(n16557), .c(n16676), .o(n16802) );
na02f01 g13014 ( .a(n16802), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_1_), .o(n16803) );
no02f01 g13015 ( .a(n16802), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_1_), .o(n16804) );
oa12f01 g13016 ( .a(n16803), .b(n16713), .c(n16804), .o(n16805) );
in01f01 g13017 ( .a(n16716), .o(n16806) );
na02f01 g13018 ( .a(n16806), .b(n16805), .o(n16807) );
in01f01 g13019 ( .a(n16720), .o(n16808) );
na03f01 g13020 ( .a(n16808), .b(n16807), .c(n16799), .o(n16809) );
in01f01 g13021 ( .a(n16722), .o(n16810) );
na03f01 g13022 ( .a(n16810), .b(n16809), .c(n16798), .o(n16811) );
in01f01 g13023 ( .a(n16725), .o(n16812) );
na03f01 g13024 ( .a(n16812), .b(n16811), .c(n16685), .o(n16813) );
in01f01 g13025 ( .a(n16727), .o(n16814) );
na03f01 g13026 ( .a(n16814), .b(n16813), .c(n16797), .o(n16815) );
na03f01 g13027 ( .a(n16729), .b(n16815), .c(n16796), .o(n16816) );
in01f01 g13028 ( .a(n16732), .o(n16817) );
na03f01 g13029 ( .a(n16817), .b(n16816), .c(n16795), .o(n16818) );
na03f01 g13030 ( .a(n16734), .b(n16818), .c(n16794), .o(n16819) );
in01f01 g13031 ( .a(n16737), .o(n16820) );
na03f01 g13032 ( .a(n16820), .b(n16819), .c(n16793), .o(n16821) );
in01f01 g13033 ( .a(n16740), .o(n16822) );
na03f01 g13034 ( .a(n16822), .b(n16821), .c(n16792), .o(n16823) );
in01f01 g13035 ( .a(n16742), .o(n16824) );
na03f01 g13036 ( .a(n16824), .b(n16823), .c(n16791), .o(n16825) );
na03f01 g13037 ( .a(n16744), .b(n16825), .c(n16790), .o(n16826) );
in01f01 g13038 ( .a(n16752), .o(n16827) );
na03f01 g13039 ( .a(n16827), .b(n16826), .c(n16789), .o(n16828) );
ao12f01 g13040 ( .a(n16595), .b(n16758), .c(n16828), .o(n16829) );
in01f01 g13041 ( .a(n16770), .o(n16830) );
na02f01 g13042 ( .a(n16830), .b(n16829), .o(n16831) );
in01f01 g13043 ( .a(n16788), .o(n16832) );
no02f01 g13044 ( .a(n16832), .b(n16773), .o(n16833) );
na02f01 g13045 ( .a(n16833), .b(n16831), .o(n16834) );
oa12f01 g13046 ( .a(n16834), .b(n16788), .c(n16774), .o(n16835) );
no02f01 g13047 ( .a(n16549), .b(delay_xor_ln22_unr12_stage5_stallmux_q_4_), .o(n16836) );
no02f01 g13048 ( .a(n16549), .b(delay_xor_ln22_unr12_stage5_stallmux_q_2_), .o(n16837) );
no02f01 g13049 ( .a(n16549), .b(delay_xor_ln22_unr12_stage5_stallmux_q_0_), .o(n16838) );
no02f01 g13050 ( .a(n16549), .b(delay_xor_ln22_unr12_stage5_stallmux_q_1_), .o(n16839) );
no02f01 g13051 ( .a(n16839), .b(n16838), .o(n16840) );
in01f01 g13052 ( .a(n16840), .o(n16841) );
no02f01 g13053 ( .a(n16841), .b(n16837), .o(n16842) );
no02f01 g13054 ( .a(n16549), .b(delay_xor_ln22_unr12_stage5_stallmux_q_3_), .o(n16843) );
in01f01 g13055 ( .a(n16843), .o(n16844) );
na02f01 g13056 ( .a(n16844), .b(n16842), .o(n16845) );
no02f01 g13057 ( .a(n16845), .b(n16836), .o(n16846) );
no02f01 g13058 ( .a(n16549), .b(delay_xor_ln22_unr12_stage5_stallmux_q_5_), .o(n16847) );
no02f01 g13059 ( .a(n16549), .b(delay_xor_ln22_unr12_stage5_stallmux_q_6_), .o(n16848) );
no02f01 g13060 ( .a(n16848), .b(n16847), .o(n16849) );
na02f01 g13061 ( .a(n16849), .b(n16846), .o(n16850) );
in01f01 g13062 ( .a(n16850), .o(n16851) );
no02f01 g13063 ( .a(n16549), .b(delay_xor_ln22_unr12_stage5_stallmux_q_7_), .o(n16852) );
no02f01 g13064 ( .a(n16549), .b(delay_xor_ln22_unr12_stage5_stallmux_q_8_), .o(n16853) );
no02f01 g13065 ( .a(n16853), .b(n16852), .o(n16854) );
na02f01 g13066 ( .a(n16854), .b(n16851), .o(n16855) );
no02f01 g13067 ( .a(n16549), .b(delay_xor_ln22_unr12_stage5_stallmux_q_9_), .o(n16856) );
no02f01 g13068 ( .a(n16856), .b(n16855), .o(n16857) );
no02f01 g13069 ( .a(n16549), .b(delay_xor_ln22_unr12_stage5_stallmux_q_12_), .o(n16858) );
no02f01 g13070 ( .a(n16549), .b(delay_xor_ln22_unr12_stage5_stallmux_q_11_), .o(n16859) );
no02f01 g13071 ( .a(n16549), .b(delay_xor_ln22_unr12_stage5_stallmux_q_10_), .o(n16860) );
no03f01 g13072 ( .a(n16860), .b(n16859), .c(n16858), .o(n16861) );
no02f01 g13073 ( .a(delay_xor_ln22_unr12_stage5_stallmux_q_15_), .b(n16549), .o(n16862) );
no02f01 g13074 ( .a(n16549), .b(delay_xor_ln22_unr12_stage5_stallmux_q_13_), .o(n16863) );
no02f01 g13075 ( .a(n16549), .b(delay_xor_ln22_unr12_stage5_stallmux_q_14_), .o(n16864) );
no03f01 g13076 ( .a(n16864), .b(n16863), .c(n16862), .o(n16865) );
na03f01 g13077 ( .a(n16865), .b(n16861), .c(n16857), .o(n16866) );
no02f01 g13078 ( .a(n16549), .b(delay_xor_ln22_unr12_stage5_stallmux_q_16_), .o(n16867) );
no02f01 g13079 ( .a(n16867), .b(n16866), .o(n16868) );
in01f01 g13080 ( .a(n16868), .o(n16869) );
no02f01 g13081 ( .a(n16549), .b(delay_xor_ln22_unr12_stage5_stallmux_q_17_), .o(n16870) );
no02f01 g13082 ( .a(n16870), .b(n16869), .o(n16871) );
in01f01 g13083 ( .a(n16871), .o(n16872) );
no02f01 g13084 ( .a(n16549), .b(delay_xor_ln22_unr12_stage5_stallmux_q_18_), .o(n16873) );
no02f01 g13085 ( .a(n16873), .b(n16872), .o(n16874) );
in01f01 g13086 ( .a(delay_xor_ln22_unr12_stage5_stallmux_q_19_), .o(n16875) );
no02f01 g13087 ( .a(n_44365), .b(n16875), .o(n16876) );
in01f01 g13088 ( .a(n16876), .o(n16877) );
no02f01 g13089 ( .a(n16549), .b(delay_xor_ln22_unr12_stage5_stallmux_q_19_), .o(n16878) );
ao12f01 g13090 ( .a(n16878), .b(n16877), .c(n16874), .o(n16879) );
no02f01 g13091 ( .a(n16879), .b(delay_add_ln22_unr11_stage5_stallmux_q_21_), .o(n16880) );
in01f01 g13092 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_21_), .o(n16881) );
in01f01 g13093 ( .a(n16879), .o(n16882) );
no02f01 g13094 ( .a(n16882), .b(n16881), .o(n16883) );
no02f01 g13095 ( .a(n16883), .b(n16880), .o(n16884) );
in01f01 g13096 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_20_), .o(n16885) );
no02f01 g13097 ( .a(n16882), .b(n16885), .o(n16886) );
in01f01 g13098 ( .a(n16874), .o(n16887) );
no02f01 g13099 ( .a(n16878), .b(n16876), .o(n16888) );
no02f01 g13100 ( .a(n16888), .b(n16887), .o(n16889) );
na02f01 g13101 ( .a(n16888), .b(n16887), .o(n16890) );
in01f01 g13102 ( .a(n16890), .o(n16891) );
no02f01 g13103 ( .a(n16891), .b(n16889), .o(n16892) );
in01f01 g13104 ( .a(n16892), .o(n16893) );
no02f01 g13105 ( .a(n16893), .b(delay_add_ln22_unr11_stage5_stallmux_q_19_), .o(n16894) );
na02f01 g13106 ( .a(n16549), .b(delay_xor_ln22_unr12_stage5_stallmux_q_17_), .o(n16895) );
in01f01 g13107 ( .a(n16895), .o(n16896) );
no02f01 g13108 ( .a(n16896), .b(n16870), .o(n16897) );
in01f01 g13109 ( .a(n16897), .o(n16898) );
no02f01 g13110 ( .a(n16898), .b(n16868), .o(n16899) );
no02f01 g13111 ( .a(n16897), .b(n16869), .o(n16900) );
no02f01 g13112 ( .a(n16900), .b(n16899), .o(n16901) );
in01f01 g13113 ( .a(n16901), .o(n16902) );
no02f01 g13114 ( .a(n16902), .b(delay_add_ln22_unr11_stage5_stallmux_q_17_), .o(n16903) );
in01f01 g13115 ( .a(n16903), .o(n16904) );
in01f01 g13116 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_15_), .o(n16905) );
na02f01 g13117 ( .a(n16861), .b(n16857), .o(n16906) );
no02f01 g13118 ( .a(n16863), .b(n16906), .o(n16907) );
in01f01 g13119 ( .a(n16907), .o(n16908) );
no02f01 g13120 ( .a(n16908), .b(n16864), .o(n16909) );
in01f01 g13121 ( .a(n16909), .o(n16910) );
na02f01 g13122 ( .a(delay_xor_ln22_unr12_stage5_stallmux_q_15_), .b(n16549), .o(n16911) );
in01f01 g13123 ( .a(n16911), .o(n16912) );
no02f01 g13124 ( .a(n16912), .b(n16862), .o(n16913) );
no02f01 g13125 ( .a(n16913), .b(n16910), .o(n16914) );
na02f01 g13126 ( .a(n16913), .b(n16910), .o(n16915) );
in01f01 g13127 ( .a(n16915), .o(n16916) );
no02f01 g13128 ( .a(n16916), .b(n16914), .o(n16917) );
no02f01 g13129 ( .a(n16917), .b(n16905), .o(n16918) );
in01f01 g13130 ( .a(n16918), .o(n16919) );
in01f01 g13131 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_14_), .o(n16920) );
na02f01 g13132 ( .a(n16549), .b(delay_xor_ln22_unr12_stage5_stallmux_q_14_), .o(n16921) );
in01f01 g13133 ( .a(n16921), .o(n16922) );
no02f01 g13134 ( .a(n16922), .b(n16864), .o(n16923) );
no02f01 g13135 ( .a(n16923), .b(n16908), .o(n16924) );
na02f01 g13136 ( .a(n16923), .b(n16908), .o(n16925) );
in01f01 g13137 ( .a(n16925), .o(n16926) );
no02f01 g13138 ( .a(n16926), .b(n16924), .o(n16927) );
no02f01 g13139 ( .a(n16927), .b(n16920), .o(n16928) );
na02f01 g13140 ( .a(n16549), .b(delay_xor_ln22_unr12_stage5_stallmux_q_13_), .o(n16929) );
in01f01 g13141 ( .a(n16929), .o(n16930) );
no02f01 g13142 ( .a(n16930), .b(n16863), .o(n16931) );
no02f01 g13143 ( .a(n16931), .b(n16906), .o(n16932) );
na02f01 g13144 ( .a(n16931), .b(n16906), .o(n16933) );
in01f01 g13145 ( .a(n16933), .o(n16934) );
no02f01 g13146 ( .a(n16934), .b(n16932), .o(n16935) );
in01f01 g13147 ( .a(n16935), .o(n16936) );
no02f01 g13148 ( .a(n16936), .b(delay_add_ln22_unr11_stage5_stallmux_q_13_), .o(n16937) );
in01f01 g13149 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_12_), .o(n16938) );
na02f01 g13150 ( .a(n16549), .b(delay_xor_ln22_unr12_stage5_stallmux_q_12_), .o(n16939) );
in01f01 g13151 ( .a(n16939), .o(n16940) );
no02f01 g13152 ( .a(n16940), .b(n16858), .o(n16941) );
in01f01 g13153 ( .a(n16941), .o(n16942) );
in01f01 g13154 ( .a(n16857), .o(n16943) );
no02f01 g13155 ( .a(n16860), .b(n16943), .o(n16944) );
in01f01 g13156 ( .a(n16944), .o(n16945) );
no02f01 g13157 ( .a(n16945), .b(n16859), .o(n16946) );
no02f01 g13158 ( .a(n16946), .b(n16942), .o(n16947) );
na02f01 g13159 ( .a(n16946), .b(n16942), .o(n16948) );
in01f01 g13160 ( .a(n16948), .o(n16949) );
no02f01 g13161 ( .a(n16949), .b(n16947), .o(n16950) );
no02f01 g13162 ( .a(n16950), .b(n16938), .o(n16951) );
na02f01 g13163 ( .a(n16549), .b(delay_xor_ln22_unr12_stage5_stallmux_q_11_), .o(n16952) );
in01f01 g13164 ( .a(n16952), .o(n16953) );
no02f01 g13165 ( .a(n16953), .b(n16859), .o(n16954) );
in01f01 g13166 ( .a(n16954), .o(n16955) );
no02f01 g13167 ( .a(n16955), .b(n16944), .o(n16956) );
no02f01 g13168 ( .a(n16954), .b(n16945), .o(n16957) );
no02f01 g13169 ( .a(n16957), .b(n16956), .o(n16958) );
in01f01 g13170 ( .a(n16958), .o(n16959) );
no02f01 g13171 ( .a(n16959), .b(delay_add_ln22_unr11_stage5_stallmux_q_11_), .o(n16960) );
in01f01 g13172 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_10_), .o(n16961) );
na02f01 g13173 ( .a(n16549), .b(delay_xor_ln22_unr12_stage5_stallmux_q_10_), .o(n16962) );
in01f01 g13174 ( .a(n16962), .o(n16963) );
no02f01 g13175 ( .a(n16963), .b(n16860), .o(n16964) );
no02f01 g13176 ( .a(n16964), .b(n16943), .o(n16965) );
na02f01 g13177 ( .a(n16964), .b(n16943), .o(n16966) );
in01f01 g13178 ( .a(n16966), .o(n16967) );
no02f01 g13179 ( .a(n16967), .b(n16965), .o(n16968) );
no02f01 g13180 ( .a(n16968), .b(n16961), .o(n16969) );
na02f01 g13181 ( .a(n16549), .b(delay_xor_ln22_unr12_stage5_stallmux_q_9_), .o(n16970) );
in01f01 g13182 ( .a(n16970), .o(n16971) );
no02f01 g13183 ( .a(n16971), .b(n16856), .o(n16972) );
in01f01 g13184 ( .a(n16972), .o(n16973) );
ao12f01 g13185 ( .a(n16973), .b(n16854), .c(n16851), .o(n16974) );
no02f01 g13186 ( .a(n16972), .b(n16855), .o(n16975) );
no02f01 g13187 ( .a(n16975), .b(n16974), .o(n16976) );
in01f01 g13188 ( .a(n16976), .o(n16977) );
no02f01 g13189 ( .a(n16977), .b(delay_add_ln22_unr11_stage5_stallmux_q_9_), .o(n16978) );
in01f01 g13190 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_8_), .o(n16979) );
na02f01 g13191 ( .a(n16549), .b(delay_xor_ln22_unr12_stage5_stallmux_q_8_), .o(n16980) );
in01f01 g13192 ( .a(n16980), .o(n16981) );
no02f01 g13193 ( .a(n16981), .b(n16853), .o(n16982) );
no02f01 g13194 ( .a(n16852), .b(n16850), .o(n16983) );
in01f01 g13195 ( .a(n16983), .o(n16984) );
no02f01 g13196 ( .a(n16984), .b(n16982), .o(n16985) );
na02f01 g13197 ( .a(n16984), .b(n16982), .o(n16986) );
in01f01 g13198 ( .a(n16986), .o(n16987) );
no02f01 g13199 ( .a(n16987), .b(n16985), .o(n16988) );
no02f01 g13200 ( .a(n16988), .b(n16979), .o(n16989) );
na02f01 g13201 ( .a(n16549), .b(delay_xor_ln22_unr12_stage5_stallmux_q_7_), .o(n16990) );
in01f01 g13202 ( .a(n16990), .o(n16991) );
no02f01 g13203 ( .a(n16991), .b(n16852), .o(n16992) );
in01f01 g13204 ( .a(n16992), .o(n16993) );
no02f01 g13205 ( .a(n16993), .b(n16851), .o(n16994) );
no02f01 g13206 ( .a(n16992), .b(n16850), .o(n16995) );
no02f01 g13207 ( .a(n16995), .b(n16994), .o(n16996) );
in01f01 g13208 ( .a(n16996), .o(n16997) );
no02f01 g13209 ( .a(n16997), .b(delay_add_ln22_unr11_stage5_stallmux_q_7_), .o(n16998) );
in01f01 g13210 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_7_), .o(n16999) );
no02f01 g13211 ( .a(n16996), .b(n16999), .o(n17000) );
in01f01 g13212 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_6_), .o(n17001) );
in01f01 g13213 ( .a(n16847), .o(n17002) );
na02f01 g13214 ( .a(n16549), .b(delay_xor_ln22_unr12_stage5_stallmux_q_6_), .o(n17003) );
in01f01 g13215 ( .a(n17003), .o(n17004) );
no02f01 g13216 ( .a(n17004), .b(n16848), .o(n17005) );
in01f01 g13217 ( .a(n17005), .o(n17006) );
ao12f01 g13218 ( .a(n17006), .b(n17002), .c(n16846), .o(n17007) );
in01f01 g13219 ( .a(n16846), .o(n17008) );
no03f01 g13220 ( .a(n17005), .b(n16847), .c(n17008), .o(n17009) );
no02f01 g13221 ( .a(n17009), .b(n17007), .o(n17010) );
no02f01 g13222 ( .a(n17010), .b(n17001), .o(n17011) );
na02f01 g13223 ( .a(n16549), .b(delay_xor_ln22_unr12_stage5_stallmux_q_5_), .o(n17012) );
na02f01 g13224 ( .a(n17012), .b(n17002), .o(n17013) );
na02f01 g13225 ( .a(n17013), .b(n16846), .o(n17014) );
in01f01 g13226 ( .a(n17013), .o(n17015) );
na02f01 g13227 ( .a(n17015), .b(n17008), .o(n17016) );
na02f01 g13228 ( .a(n17016), .b(n17014), .o(n17017) );
no02f01 g13229 ( .a(n17017), .b(delay_add_ln22_unr11_stage5_stallmux_q_5_), .o(n17018) );
in01f01 g13230 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_4_), .o(n17019) );
in01f01 g13231 ( .a(n16836), .o(n17020) );
na02f01 g13232 ( .a(n16549), .b(delay_xor_ln22_unr12_stage5_stallmux_q_4_), .o(n17021) );
na02f01 g13233 ( .a(n17021), .b(n17020), .o(n17022) );
ao12f01 g13234 ( .a(n17022), .b(n16844), .c(n16842), .o(n17023) );
in01f01 g13235 ( .a(n17022), .o(n17024) );
no02f01 g13236 ( .a(n17024), .b(n16845), .o(n17025) );
no02f01 g13237 ( .a(n17025), .b(n17023), .o(n17026) );
no02f01 g13238 ( .a(n17026), .b(n17019), .o(n17027) );
na02f01 g13239 ( .a(n16549), .b(delay_xor_ln22_unr12_stage5_stallmux_q_3_), .o(n17028) );
na02f01 g13240 ( .a(n17028), .b(n16844), .o(n17029) );
na02f01 g13241 ( .a(n17029), .b(n16842), .o(n17030) );
no02f01 g13242 ( .a(n17029), .b(n16842), .o(n17031) );
in01f01 g13243 ( .a(n17031), .o(n17032) );
na02f01 g13244 ( .a(n17032), .b(n17030), .o(n17033) );
no02f01 g13245 ( .a(n17033), .b(delay_add_ln22_unr11_stage5_stallmux_q_3_), .o(n17034) );
in01f01 g13246 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_2_), .o(n17035) );
na02f01 g13247 ( .a(n16549), .b(delay_xor_ln22_unr12_stage5_stallmux_q_2_), .o(n17036) );
in01f01 g13248 ( .a(n17036), .o(n17037) );
no02f01 g13249 ( .a(n17037), .b(n16837), .o(n17038) );
no02f01 g13250 ( .a(n17038), .b(n16841), .o(n17039) );
na02f01 g13251 ( .a(n17038), .b(n16841), .o(n17040) );
in01f01 g13252 ( .a(n17040), .o(n17041) );
no02f01 g13253 ( .a(n17041), .b(n17039), .o(n17042) );
no02f01 g13254 ( .a(n17042), .b(n17035), .o(n17043) );
in01f01 g13255 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_1_), .o(n17044) );
in01f01 g13256 ( .a(n16838), .o(n17045) );
in01f01 g13257 ( .a(delay_xor_ln22_unr12_stage5_stallmux_q_1_), .o(n17046) );
na02f01 g13258 ( .a(n_44365), .b(n17046), .o(n17047) );
na02f01 g13259 ( .a(n16549), .b(delay_xor_ln22_unr12_stage5_stallmux_q_1_), .o(n17048) );
na02f01 g13260 ( .a(n17048), .b(n17047), .o(n17049) );
no02f01 g13261 ( .a(n17049), .b(n17045), .o(n17050) );
no02f01 g13262 ( .a(n_44365), .b(n17046), .o(n17051) );
no02f01 g13263 ( .a(n17051), .b(n16839), .o(n17052) );
no02f01 g13264 ( .a(n17052), .b(n16838), .o(n17053) );
no02f01 g13265 ( .a(n17053), .b(n17050), .o(n17054) );
no02f01 g13266 ( .a(n17054), .b(n17044), .o(n17055) );
na02f01 g13267 ( .a(n17054), .b(n17044), .o(n17056) );
in01f01 g13268 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_0_), .o(n17057) );
no02f01 g13269 ( .a(n_44365), .b(delay_xor_ln22_unr12_stage5_stallmux_q_0_), .o(n17058) );
na02f01 g13270 ( .a(n_44365), .b(delay_xor_ln22_unr12_stage5_stallmux_q_0_), .o(n17059) );
in01f01 g13271 ( .a(n17059), .o(n17060) );
no02f01 g13272 ( .a(n17060), .b(n17058), .o(n17061) );
in01f01 g13273 ( .a(n17061), .o(n17062) );
no02f01 g13274 ( .a(n17062), .b(n17057), .o(n17063) );
ao12f01 g13275 ( .a(n17055), .b(n17063), .c(n17056), .o(n17064) );
no03f01 g13276 ( .a(n17041), .b(n17039), .c(delay_add_ln22_unr11_stage5_stallmux_q_2_), .o(n17065) );
no02f01 g13277 ( .a(n17065), .b(n17064), .o(n17066) );
in01f01 g13278 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_3_), .o(n17067) );
ao12f01 g13279 ( .a(n17067), .b(n17032), .c(n17030), .o(n17068) );
no03f01 g13280 ( .a(n17068), .b(n17066), .c(n17043), .o(n17069) );
na02f01 g13281 ( .a(n17026), .b(n17019), .o(n17070) );
in01f01 g13282 ( .a(n17070), .o(n17071) );
no03f01 g13283 ( .a(n17071), .b(n17069), .c(n17034), .o(n17072) );
in01f01 g13284 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_5_), .o(n17073) );
ao12f01 g13285 ( .a(n17073), .b(n17016), .c(n17014), .o(n17074) );
no03f01 g13286 ( .a(n17074), .b(n17072), .c(n17027), .o(n17075) );
na02f01 g13287 ( .a(n17010), .b(n17001), .o(n17076) );
in01f01 g13288 ( .a(n17076), .o(n17077) );
no03f01 g13289 ( .a(n17077), .b(n17075), .c(n17018), .o(n17078) );
no03f01 g13290 ( .a(n17078), .b(n17011), .c(n17000), .o(n17079) );
no03f01 g13291 ( .a(n16987), .b(n16985), .c(delay_add_ln22_unr11_stage5_stallmux_q_8_), .o(n17080) );
no03f01 g13292 ( .a(n17080), .b(n17079), .c(n16998), .o(n17081) );
na02f01 g13293 ( .a(n16977), .b(delay_add_ln22_unr11_stage5_stallmux_q_9_), .o(n17082) );
in01f01 g13294 ( .a(n17082), .o(n17083) );
no03f01 g13295 ( .a(n17083), .b(n17081), .c(n16989), .o(n17084) );
na02f01 g13296 ( .a(n16968), .b(n16961), .o(n17085) );
in01f01 g13297 ( .a(n17085), .o(n17086) );
no03f01 g13298 ( .a(n17086), .b(n17084), .c(n16978), .o(n17087) );
na02f01 g13299 ( .a(n16959), .b(delay_add_ln22_unr11_stage5_stallmux_q_11_), .o(n17088) );
in01f01 g13300 ( .a(n17088), .o(n17089) );
no03f01 g13301 ( .a(n17089), .b(n17087), .c(n16969), .o(n17090) );
na02f01 g13302 ( .a(n16950), .b(n16938), .o(n17091) );
in01f01 g13303 ( .a(n17091), .o(n17092) );
no03f01 g13304 ( .a(n17092), .b(n17090), .c(n16960), .o(n17093) );
na02f01 g13305 ( .a(n16936), .b(delay_add_ln22_unr11_stage5_stallmux_q_13_), .o(n17094) );
in01f01 g13306 ( .a(n17094), .o(n17095) );
no03f01 g13307 ( .a(n17095), .b(n17093), .c(n16951), .o(n17096) );
na02f01 g13308 ( .a(n16927), .b(n16920), .o(n17097) );
in01f01 g13309 ( .a(n17097), .o(n17098) );
no03f01 g13310 ( .a(n17098), .b(n17096), .c(n16937), .o(n17099) );
na02f01 g13311 ( .a(n16917), .b(n16905), .o(n17100) );
oa12f01 g13312 ( .a(n17100), .b(n17099), .c(n16928), .o(n17101) );
na02f01 g13313 ( .a(n16549), .b(delay_xor_ln22_unr12_stage5_stallmux_q_16_), .o(n17102) );
in01f01 g13314 ( .a(n17102), .o(n17103) );
no02f01 g13315 ( .a(n17103), .b(n16867), .o(n17104) );
no02f01 g13316 ( .a(n17104), .b(n16866), .o(n17105) );
na02f01 g13317 ( .a(n17104), .b(n16866), .o(n17106) );
in01f01 g13318 ( .a(n17106), .o(n17107) );
no02f01 g13319 ( .a(n17107), .b(n17105), .o(n17108) );
in01f01 g13320 ( .a(n17108), .o(n17109) );
no02f01 g13321 ( .a(n17109), .b(delay_add_ln22_unr11_stage5_stallmux_q_16_), .o(n17110) );
ao12f01 g13322 ( .a(n17110), .b(n17101), .c(n16919), .o(n17111) );
na02f01 g13323 ( .a(n16902), .b(delay_add_ln22_unr11_stage5_stallmux_q_17_), .o(n17112) );
in01f01 g13324 ( .a(n17112), .o(n17113) );
na02f01 g13325 ( .a(n17109), .b(delay_add_ln22_unr11_stage5_stallmux_q_16_), .o(n17114) );
in01f01 g13326 ( .a(n17114), .o(n17115) );
no02f01 g13327 ( .a(n17115), .b(n17113), .o(n17116) );
in01f01 g13328 ( .a(n17116), .o(n17117) );
oa12f01 g13329 ( .a(n16904), .b(n17117), .c(n17111), .o(n17118) );
na02f01 g13330 ( .a(n16549), .b(delay_xor_ln22_unr12_stage5_stallmux_q_18_), .o(n17119) );
in01f01 g13331 ( .a(n17119), .o(n17120) );
no02f01 g13332 ( .a(n17120), .b(n16873), .o(n17121) );
no02f01 g13333 ( .a(n17121), .b(n16872), .o(n17122) );
na02f01 g13334 ( .a(n17121), .b(n16872), .o(n17123) );
in01f01 g13335 ( .a(n17123), .o(n17124) );
no02f01 g13336 ( .a(n17124), .b(n17122), .o(n17125) );
in01f01 g13337 ( .a(n17125), .o(n17126) );
no02f01 g13338 ( .a(n17126), .b(delay_add_ln22_unr11_stage5_stallmux_q_18_), .o(n17127) );
na02f01 g13339 ( .a(n17126), .b(delay_add_ln22_unr11_stage5_stallmux_q_18_), .o(n17128) );
oa12f01 g13340 ( .a(n17128), .b(n17127), .c(n17118), .o(n17129) );
na02f01 g13341 ( .a(n16893), .b(delay_add_ln22_unr11_stage5_stallmux_q_19_), .o(n17130) );
in01f01 g13342 ( .a(n17130), .o(n17131) );
no02f01 g13343 ( .a(n17131), .b(n17129), .o(n17132) );
no02f01 g13344 ( .a(n17132), .b(n16894), .o(n17133) );
no02f01 g13345 ( .a(n16879), .b(delay_add_ln22_unr11_stage5_stallmux_q_20_), .o(n17134) );
in01f01 g13346 ( .a(n17134), .o(n17135) );
ao12f01 g13347 ( .a(n16886), .b(n17135), .c(n17133), .o(n17136) );
na02f01 g13348 ( .a(n17136), .b(n16884), .o(n17137) );
in01f01 g13349 ( .a(n16884), .o(n17138) );
in01f01 g13350 ( .a(n16894), .o(n17139) );
in01f01 g13351 ( .a(n16928), .o(n17140) );
in01f01 g13352 ( .a(n16937), .o(n17141) );
in01f01 g13353 ( .a(n16951), .o(n17142) );
in01f01 g13354 ( .a(n16960), .o(n17143) );
in01f01 g13355 ( .a(n16969), .o(n17144) );
in01f01 g13356 ( .a(n16978), .o(n17145) );
in01f01 g13357 ( .a(n16989), .o(n17146) );
in01f01 g13358 ( .a(n16998), .o(n17147) );
in01f01 g13359 ( .a(n17000), .o(n17148) );
in01f01 g13360 ( .a(n17011), .o(n17149) );
in01f01 g13361 ( .a(n17018), .o(n17150) );
in01f01 g13362 ( .a(n17027), .o(n17151) );
in01f01 g13363 ( .a(n17034), .o(n17152) );
in01f01 g13364 ( .a(n17043), .o(n17153) );
na02f01 g13365 ( .a(n17052), .b(n16838), .o(n17154) );
na02f01 g13366 ( .a(n17049), .b(n17045), .o(n17155) );
na02f01 g13367 ( .a(n17155), .b(n17154), .o(n17156) );
na02f01 g13368 ( .a(n17156), .b(delay_add_ln22_unr11_stage5_stallmux_q_1_), .o(n17157) );
no02f01 g13369 ( .a(n17156), .b(delay_add_ln22_unr11_stage5_stallmux_q_1_), .o(n17158) );
in01f01 g13370 ( .a(n17063), .o(n17159) );
oa12f01 g13371 ( .a(n17157), .b(n17159), .c(n17158), .o(n17160) );
in01f01 g13372 ( .a(n17065), .o(n17161) );
na02f01 g13373 ( .a(n17161), .b(n17160), .o(n17162) );
na02f01 g13374 ( .a(n17033), .b(delay_add_ln22_unr11_stage5_stallmux_q_3_), .o(n17163) );
na03f01 g13375 ( .a(n17163), .b(n17162), .c(n17153), .o(n17164) );
na03f01 g13376 ( .a(n17070), .b(n17164), .c(n17152), .o(n17165) );
in01f01 g13377 ( .a(n17074), .o(n17166) );
na03f01 g13378 ( .a(n17166), .b(n17165), .c(n17151), .o(n17167) );
na03f01 g13379 ( .a(n17076), .b(n17167), .c(n17150), .o(n17168) );
na03f01 g13380 ( .a(n17168), .b(n17149), .c(n17148), .o(n17169) );
in01f01 g13381 ( .a(n17080), .o(n17170) );
na03f01 g13382 ( .a(n17170), .b(n17169), .c(n17147), .o(n17171) );
na03f01 g13383 ( .a(n17082), .b(n17171), .c(n17146), .o(n17172) );
na03f01 g13384 ( .a(n17085), .b(n17172), .c(n17145), .o(n17173) );
na03f01 g13385 ( .a(n17088), .b(n17173), .c(n17144), .o(n17174) );
na03f01 g13386 ( .a(n17091), .b(n17174), .c(n17143), .o(n17175) );
na03f01 g13387 ( .a(n17094), .b(n17175), .c(n17142), .o(n17176) );
na03f01 g13388 ( .a(n17097), .b(n17176), .c(n17141), .o(n17177) );
in01f01 g13389 ( .a(n17100), .o(n17178) );
ao12f01 g13390 ( .a(n17178), .b(n17177), .c(n17140), .o(n17179) );
in01f01 g13391 ( .a(n17110), .o(n17180) );
oa12f01 g13392 ( .a(n17180), .b(n17179), .c(n16918), .o(n17181) );
na02f01 g13393 ( .a(n17116), .b(n17181), .o(n17182) );
in01f01 g13394 ( .a(n17127), .o(n17183) );
na03f01 g13395 ( .a(n17183), .b(n17182), .c(n16904), .o(n17184) );
na03f01 g13396 ( .a(n17130), .b(n17128), .c(n17184), .o(n17185) );
na02f01 g13397 ( .a(n17185), .b(n17139), .o(n17186) );
no02f01 g13398 ( .a(n17134), .b(n17186), .o(n17187) );
oa12f01 g13399 ( .a(n17138), .b(n17187), .c(n16886), .o(n17188) );
na02f01 g13400 ( .a(n17188), .b(n17137), .o(n17189) );
na02f01 g13401 ( .a(n17189), .b(n_17093), .o(n17190) );
no02f01 g13402 ( .a(n17134), .b(n16886), .o(n17191) );
in01f01 g13403 ( .a(n17191), .o(n17192) );
na03f01 g13404 ( .a(n17192), .b(n17185), .c(n17139), .o(n17193) );
oa12f01 g13405 ( .a(n17191), .b(n17132), .c(n16894), .o(n17194) );
na02f01 g13406 ( .a(n17194), .b(n17193), .o(n17195) );
no02f01 g13407 ( .a(n17113), .b(n16903), .o(n17196) );
na03f01 g13408 ( .a(n17196), .b(n17114), .c(n17181), .o(n17197) );
in01f01 g13409 ( .a(n17196), .o(n17198) );
oa12f01 g13410 ( .a(n17198), .b(n17115), .c(n17111), .o(n17199) );
na02f01 g13411 ( .a(n17199), .b(n17197), .o(n17200) );
na02f01 g13412 ( .a(n17101), .b(n16919), .o(n17201) );
no02f01 g13413 ( .a(n17115), .b(n17110), .o(n17202) );
in01f01 g13414 ( .a(n17202), .o(n17203) );
no02f01 g13415 ( .a(n17203), .b(n17201), .o(n17204) );
no02f01 g13416 ( .a(n17179), .b(n16918), .o(n17205) );
no02f01 g13417 ( .a(n17202), .b(n17205), .o(n17206) );
no02f01 g13418 ( .a(n17206), .b(n17204), .o(n17207) );
no02f01 g13419 ( .a(n17178), .b(n16918), .o(n17208) );
ao12f01 g13420 ( .a(n16928), .b(n17176), .c(n17141), .o(n17209) );
oa12f01 g13421 ( .a(n17208), .b(n17209), .c(n17098), .o(n17210) );
in01f01 g13422 ( .a(n17208), .o(n17211) );
oa12f01 g13423 ( .a(n17140), .b(n17096), .c(n16937), .o(n17212) );
na03f01 g13424 ( .a(n17212), .b(n17211), .c(n17097), .o(n17213) );
na02f01 g13425 ( .a(n17213), .b(n17210), .o(n17214) );
no02f01 g13426 ( .a(n17098), .b(n16928), .o(n17215) );
no03f01 g13427 ( .a(n17215), .b(n17096), .c(n16937), .o(n17216) );
in01f01 g13428 ( .a(n17215), .o(n17217) );
ao12f01 g13429 ( .a(n17217), .b(n17176), .c(n17141), .o(n17218) );
no02f01 g13430 ( .a(n17218), .b(n17216), .o(n17219) );
no02f01 g13431 ( .a(n17093), .b(n16951), .o(n17220) );
no02f01 g13432 ( .a(n17095), .b(n16937), .o(n17221) );
na02f01 g13433 ( .a(n17221), .b(n17220), .o(n17222) );
in01f01 g13434 ( .a(n17222), .o(n17223) );
no02f01 g13435 ( .a(n17221), .b(n17220), .o(n17224) );
no02f01 g13436 ( .a(n17224), .b(n17223), .o(n17225) );
ao12f01 g13437 ( .a(n7550), .b(n17225), .c(n17219), .o(n17226) );
ao12f01 g13438 ( .a(n17226), .b(n17214), .c(n_17093), .o(n17227) );
oa12f01 g13439 ( .a(n17227), .b(n17207), .c(n7550), .o(n17228) );
ao12f01 g13440 ( .a(n17228), .b(n17200), .c(n_17093), .o(n17229) );
in01f01 g13441 ( .a(n17128), .o(n17230) );
no02f01 g13442 ( .a(n17230), .b(n17127), .o(n17231) );
no02f01 g13443 ( .a(n17231), .b(n17118), .o(n17232) );
ao12f01 g13444 ( .a(n16903), .b(n17116), .c(n17181), .o(n17233) );
in01f01 g13445 ( .a(n17231), .o(n17234) );
no02f01 g13446 ( .a(n17234), .b(n17233), .o(n17235) );
no02f01 g13447 ( .a(n17235), .b(n17232), .o(n17236) );
oa12f01 g13448 ( .a(n17229), .b(n17236), .c(n7550), .o(n17237) );
no02f01 g13449 ( .a(n17131), .b(n16894), .o(n17238) );
in01f01 g13450 ( .a(n17238), .o(n17239) );
na02f01 g13451 ( .a(n17239), .b(n17129), .o(n17240) );
na03f01 g13452 ( .a(n17238), .b(n17128), .c(n17184), .o(n17241) );
ao12f01 g13453 ( .a(n7550), .b(n17241), .c(n17240), .o(n17242) );
ao12f01 g13454 ( .a(n17238), .b(n17128), .c(n17184), .o(n17243) );
no02f01 g13455 ( .a(n17127), .b(n17118), .o(n17244) );
no03f01 g13456 ( .a(n17239), .b(n17230), .c(n17244), .o(n17245) );
oa12f01 g13457 ( .a(n7550), .b(n17245), .c(n17243), .o(n17246) );
oa12f01 g13458 ( .a(n17246), .b(n17242), .c(n17237), .o(n17247) );
oa12f01 g13459 ( .a(n7550), .b(n17247), .c(n17195), .o(n17248) );
no03f01 g13460 ( .a(n17198), .b(n17115), .c(n17111), .o(n17249) );
ao12f01 g13461 ( .a(n17196), .b(n17114), .c(n17181), .o(n17250) );
no02f01 g13462 ( .a(n17250), .b(n17249), .o(n17251) );
ao12f01 g13463 ( .a(n_17093), .b(n17236), .c(n17251), .o(n17252) );
in01f01 g13464 ( .a(n17252), .o(n17253) );
no03f01 g13465 ( .a(n17191), .b(n17132), .c(n16894), .o(n17254) );
ao12f01 g13466 ( .a(n17192), .b(n17185), .c(n17139), .o(n17255) );
no03f01 g13467 ( .a(n17255), .b(n17254), .c(n7550), .o(n17256) );
ao12f01 g13468 ( .a(n_17093), .b(n17194), .c(n17193), .o(n17257) );
na02f01 g13469 ( .a(n17202), .b(n17205), .o(n17258) );
na02f01 g13470 ( .a(n17203), .b(n17201), .o(n17259) );
na02f01 g13471 ( .a(n17259), .b(n17258), .o(n17260) );
ao12f01 g13472 ( .a(n17211), .b(n17212), .c(n17097), .o(n17261) );
no03f01 g13473 ( .a(n17209), .b(n17208), .c(n17098), .o(n17262) );
no02f01 g13474 ( .a(n17262), .b(n17261), .o(n17263) );
na03f01 g13475 ( .a(n17217), .b(n17176), .c(n17141), .o(n17264) );
oa12f01 g13476 ( .a(n17215), .b(n17096), .c(n16937), .o(n17265) );
na02f01 g13477 ( .a(n17265), .b(n17264), .o(n17266) );
in01f01 g13478 ( .a(n17224), .o(n17267) );
na02f01 g13479 ( .a(n17267), .b(n17222), .o(n17268) );
oa12f01 g13480 ( .a(n_17093), .b(n17268), .c(n17266), .o(n17269) );
oa12f01 g13481 ( .a(n17269), .b(n17263), .c(n7550), .o(n17270) );
ao12f01 g13482 ( .a(n17270), .b(n17260), .c(n_17093), .o(n17271) );
oa12f01 g13483 ( .a(n17271), .b(n17251), .c(n7550), .o(n17272) );
na02f01 g13484 ( .a(n17234), .b(n17233), .o(n17273) );
na02f01 g13485 ( .a(n17231), .b(n17118), .o(n17274) );
ao12f01 g13486 ( .a(n7550), .b(n17274), .c(n17273), .o(n17275) );
no02f01 g13487 ( .a(n17275), .b(n17272), .o(n17276) );
oa12f01 g13488 ( .a(n_17093), .b(n17245), .c(n17243), .o(n17277) );
na02f01 g13489 ( .a(n17277), .b(n17276), .o(n17278) );
in01f01 g13490 ( .a(n17278), .o(n17279) );
oa12f01 g13491 ( .a(n17279), .b(n17257), .c(n17256), .o(n17280) );
na03f01 g13492 ( .a(n17280), .b(n17253), .c(n17248), .o(n17281) );
ao12f01 g13493 ( .a(n16882), .b(n16885), .c(n16881), .o(n17282) );
no02f01 g13494 ( .a(n17134), .b(n16880), .o(n17283) );
ao12f01 g13495 ( .a(n17282), .b(n17283), .c(n17133), .o(n17284) );
in01f01 g13496 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_22_), .o(n17285) );
no02f01 g13497 ( .a(n16882), .b(n17285), .o(n17286) );
no02f01 g13498 ( .a(n16879), .b(delay_add_ln22_unr11_stage5_stallmux_q_22_), .o(n17287) );
no02f01 g13499 ( .a(n17287), .b(n17286), .o(n17288) );
na02f01 g13500 ( .a(n17288), .b(n17284), .o(n17289) );
in01f01 g13501 ( .a(n17282), .o(n17290) );
in01f01 g13502 ( .a(n17283), .o(n17291) );
oa12f01 g13503 ( .a(n17290), .b(n17291), .c(n17186), .o(n17292) );
in01f01 g13504 ( .a(n17288), .o(n17293) );
na02f01 g13505 ( .a(n17293), .b(n17292), .o(n17294) );
na02f01 g13506 ( .a(n17294), .b(n17289), .o(n17295) );
na02f01 g13507 ( .a(n17295), .b(n_17093), .o(n17296) );
no02f01 g13508 ( .a(n17286), .b(n17282), .o(n17297) );
in01f01 g13509 ( .a(n17287), .o(n17298) );
na02f01 g13510 ( .a(n17298), .b(n17283), .o(n17299) );
oa12f01 g13511 ( .a(n17297), .b(n17299), .c(n17186), .o(n17300) );
in01f01 g13512 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_23_), .o(n17301) );
no02f01 g13513 ( .a(n16882), .b(n17301), .o(n17302) );
no02f01 g13514 ( .a(n16879), .b(delay_add_ln22_unr11_stage5_stallmux_q_23_), .o(n17303) );
no02f01 g13515 ( .a(n17303), .b(n17302), .o(n17304) );
in01f01 g13516 ( .a(n17304), .o(n17305) );
na02f01 g13517 ( .a(n17305), .b(n17300), .o(n17306) );
in01f01 g13518 ( .a(n17306), .o(n17307) );
no02f01 g13519 ( .a(n17305), .b(n17300), .o(n17308) );
oa12f01 g13520 ( .a(n_17093), .b(n17308), .c(n17307), .o(n17309) );
na04f01 g13521 ( .a(n17309), .b(n17296), .c(n17281), .d(n17190), .o(n17310) );
no03f01 g13522 ( .a(n17303), .b(n17299), .c(n17186), .o(n17311) );
no03f01 g13523 ( .a(n17302), .b(n17286), .c(n17282), .o(n17312) );
in01f01 g13524 ( .a(n17312), .o(n17313) );
no02f01 g13525 ( .a(n16879), .b(delay_add_ln22_unr11_stage5_stallmux_q_24_), .o(n17314) );
in01f01 g13526 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_24_), .o(n17315) );
no02f01 g13527 ( .a(n16882), .b(n17315), .o(n17316) );
no02f01 g13528 ( .a(n17316), .b(n17314), .o(n17317) );
in01f01 g13529 ( .a(n17317), .o(n17318) );
no03f01 g13530 ( .a(n17318), .b(n17313), .c(n17311), .o(n17319) );
oa12f01 g13531 ( .a(n17318), .b(n17313), .c(n17311), .o(n17320) );
in01f01 g13532 ( .a(n17320), .o(n17321) );
no03f01 g13533 ( .a(n17321), .b(n17319), .c(n7550), .o(n17322) );
in01f01 g13534 ( .a(n17319), .o(n17323) );
ao12f01 g13535 ( .a(n_17093), .b(n17320), .c(n17323), .o(n17324) );
no02f01 g13536 ( .a(n17308), .b(n17307), .o(n17325) );
no02f01 g13537 ( .a(n17325), .b(n_17093), .o(n17326) );
no03f01 g13538 ( .a(n17326), .b(n17324), .c(n17322), .o(n17327) );
ao12f01 g13539 ( .a(n_17093), .b(n17327), .c(n17310), .o(n17328) );
no02f01 g13540 ( .a(n17324), .b(n17322), .o(n17329) );
no03f01 g13541 ( .a(n17187), .b(n16886), .c(n17138), .o(n17330) );
no02f01 g13542 ( .a(n17136), .b(n16884), .o(n17331) );
no02f01 g13543 ( .a(n17331), .b(n17330), .o(n17332) );
no02f01 g13544 ( .a(n17293), .b(n17292), .o(n17333) );
no02f01 g13545 ( .a(n17288), .b(n17284), .o(n17334) );
no02f01 g13546 ( .a(n17334), .b(n17333), .o(n17335) );
ao12f01 g13547 ( .a(n_17093), .b(n17335), .c(n17332), .o(n17336) );
in01f01 g13548 ( .a(n17336), .o(n17337) );
oa12f01 g13549 ( .a(n17337), .b(n17329), .c(n17310), .o(n17338) );
no02f01 g13550 ( .a(n16879), .b(delay_add_ln22_unr11_stage5_stallmux_q_25_), .o(n17339) );
in01f01 g13551 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_25_), .o(n17340) );
no02f01 g13552 ( .a(n16882), .b(n17340), .o(n17341) );
no02f01 g13553 ( .a(n17341), .b(n17339), .o(n17342) );
no02f01 g13554 ( .a(n17313), .b(n17311), .o(n17343) );
no02f01 g13555 ( .a(n17314), .b(n17343), .o(n17344) );
no02f01 g13556 ( .a(n17344), .b(n17316), .o(n17345) );
na02f01 g13557 ( .a(n17345), .b(n17342), .o(n17346) );
no02f01 g13558 ( .a(n17345), .b(n17342), .o(n17347) );
in01f01 g13559 ( .a(n17347), .o(n17348) );
na02f01 g13560 ( .a(n17348), .b(n17346), .o(n17349) );
na02f01 g13561 ( .a(n17349), .b(n_17093), .o(n17350) );
oa12f01 g13562 ( .a(n17350), .b(n17338), .c(n17328), .o(n17351) );
no02f01 g13563 ( .a(n17339), .b(n17314), .o(n17352) );
in01f01 g13564 ( .a(n17352), .o(n17353) );
no02f01 g13565 ( .a(n17353), .b(n17343), .o(n17354) );
ao12f01 g13566 ( .a(n16882), .b(n17315), .c(n17340), .o(n17355) );
no02f01 g13567 ( .a(n17355), .b(n17354), .o(n17356) );
no02f01 g13568 ( .a(n16879), .b(delay_add_ln22_unr11_stage5_stallmux_q_26_), .o(n17357) );
in01f01 g13569 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_26_), .o(n17358) );
no02f01 g13570 ( .a(n16882), .b(n17358), .o(n17359) );
no02f01 g13571 ( .a(n17359), .b(n17357), .o(n17360) );
no02f01 g13572 ( .a(n17360), .b(n17356), .o(n17361) );
na02f01 g13573 ( .a(n17360), .b(n17356), .o(n17362) );
in01f01 g13574 ( .a(n17362), .o(n17363) );
no02f01 g13575 ( .a(n17363), .b(n17361), .o(n17364) );
no02f01 g13576 ( .a(n17364), .b(n7550), .o(n17365) );
no02f01 g13577 ( .a(n17365), .b(n17351), .o(n17366) );
no03f01 g13578 ( .a(n17357), .b(n17353), .c(n17343), .o(n17367) );
in01f01 g13579 ( .a(n17367), .o(n17368) );
no02f01 g13580 ( .a(n16879), .b(delay_add_ln22_unr11_stage5_stallmux_q_27_), .o(n17369) );
no02f01 g13581 ( .a(n17369), .b(n17368), .o(n17370) );
in01f01 g13582 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_27_), .o(n17371) );
ao12f01 g13583 ( .a(n16882), .b(n17371), .c(n17358), .o(n17372) );
no02f01 g13584 ( .a(n17372), .b(n17355), .o(n17373) );
in01f01 g13585 ( .a(n17373), .o(n17374) );
no02f01 g13586 ( .a(n17374), .b(n17370), .o(n17375) );
in01f01 g13587 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_28_), .o(n17376) );
no02f01 g13588 ( .a(n16882), .b(n17376), .o(n17377) );
no02f01 g13589 ( .a(n16879), .b(delay_add_ln22_unr11_stage5_stallmux_q_28_), .o(n17378) );
no02f01 g13590 ( .a(n17378), .b(n17377), .o(n17379) );
na02f01 g13591 ( .a(n17379), .b(n17375), .o(n17380) );
no02f01 g13592 ( .a(n17379), .b(n17375), .o(n17381) );
in01f01 g13593 ( .a(n17381), .o(n17382) );
na02f01 g13594 ( .a(n17382), .b(n17380), .o(n17383) );
na02f01 g13595 ( .a(n17383), .b(n_17093), .o(n17384) );
no02f01 g13596 ( .a(n17359), .b(n17355), .o(n17385) );
na02f01 g13597 ( .a(n17385), .b(n17368), .o(n17386) );
no02f01 g13598 ( .a(n16882), .b(n17371), .o(n17387) );
no02f01 g13599 ( .a(n17387), .b(n17369), .o(n17388) );
in01f01 g13600 ( .a(n17388), .o(n17389) );
na02f01 g13601 ( .a(n17389), .b(n17386), .o(n17390) );
in01f01 g13602 ( .a(n17390), .o(n17391) );
no02f01 g13603 ( .a(n17389), .b(n17386), .o(n17392) );
no02f01 g13604 ( .a(n17392), .b(n17391), .o(n17393) );
no02f01 g13605 ( .a(n17393), .b(n7550), .o(n17394) );
in01f01 g13606 ( .a(n17394), .o(n17395) );
na03f01 g13607 ( .a(n17395), .b(n17384), .c(n17366), .o(n17396) );
in01f01 g13608 ( .a(n17346), .o(n17397) );
no02f01 g13609 ( .a(n17347), .b(n17397), .o(n17398) );
ao12f01 g13610 ( .a(n_17093), .b(n17364), .c(n17398), .o(n17399) );
in01f01 g13611 ( .a(n17380), .o(n17400) );
no02f01 g13612 ( .a(n17381), .b(n17400), .o(n17401) );
no02f01 g13613 ( .a(n17401), .b(n_17093), .o(n17402) );
no02f01 g13614 ( .a(n17393), .b(n_17093), .o(n17403) );
no03f01 g13615 ( .a(n17403), .b(n17402), .c(n17399), .o(n17404) );
no02f01 g13616 ( .a(n16879), .b(delay_add_ln22_unr11_stage5_stallmux_q_29_), .o(n17405) );
in01f01 g13617 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_29_), .o(n17406) );
no02f01 g13618 ( .a(n16882), .b(n17406), .o(n17407) );
no02f01 g13619 ( .a(n17407), .b(n17405), .o(n17408) );
in01f01 g13620 ( .a(n17408), .o(n17409) );
in01f01 g13621 ( .a(n17370), .o(n17410) );
no02f01 g13622 ( .a(n17377), .b(n17374), .o(n17411) );
oa12f01 g13623 ( .a(n17411), .b(n17378), .c(n17410), .o(n17412) );
no02f01 g13624 ( .a(n17412), .b(n17409), .o(n17413) );
na02f01 g13625 ( .a(n17412), .b(n17409), .o(n17414) );
in01f01 g13626 ( .a(n17414), .o(n17415) );
no02f01 g13627 ( .a(n17415), .b(n17413), .o(n17416) );
no02f01 g13628 ( .a(n17416), .b(n7550), .o(n17417) );
ao12f01 g13629 ( .a(n17417), .b(n17404), .c(n17396), .o(n17418) );
no02f01 g13630 ( .a(n17416), .b(n_17093), .o(n17419) );
no02f01 g13631 ( .a(n16879), .b(delay_add_ln22_unr11_stage5_stallmux_q_30_), .o(n17420) );
in01f01 g13632 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_30_), .o(n17421) );
no02f01 g13633 ( .a(n16882), .b(n17421), .o(n17422) );
no02f01 g13634 ( .a(n17422), .b(n17420), .o(n17423) );
in01f01 g13635 ( .a(n17423), .o(n17424) );
ao12f01 g13636 ( .a(n16882), .b(n17406), .c(n17376), .o(n17425) );
in01f01 g13637 ( .a(n17425), .o(n17426) );
no02f01 g13638 ( .a(n17405), .b(n17378), .o(n17427) );
in01f01 g13639 ( .a(n17427), .o(n17428) );
ao12f01 g13640 ( .a(n17428), .b(n17426), .c(n17375), .o(n17429) );
no02f01 g13641 ( .a(n17429), .b(n17424), .o(n17430) );
na02f01 g13642 ( .a(n17429), .b(n17424), .o(n17431) );
in01f01 g13643 ( .a(n17431), .o(n17432) );
no02f01 g13644 ( .a(n17432), .b(n17430), .o(n17433) );
no02f01 g13645 ( .a(n17433), .b(n_17093), .o(n17434) );
no02f01 g13646 ( .a(n17433), .b(n7550), .o(n17435) );
no02f01 g13647 ( .a(n17435), .b(n17434), .o(n17436) );
in01f01 g13648 ( .a(n17436), .o(n17437) );
oa12f01 g13649 ( .a(n17437), .b(n17419), .c(n17418), .o(n17438) );
no02f01 g13650 ( .a(n17332), .b(n7550), .o(n17439) );
no02f01 g13651 ( .a(n17255), .b(n17254), .o(n17440) );
ao12f01 g13652 ( .a(n_17093), .b(n17241), .c(n17240), .o(n17441) );
ao12f01 g13653 ( .a(n17441), .b(n17277), .c(n17276), .o(n17442) );
ao12f01 g13654 ( .a(n_17093), .b(n17442), .c(n17440), .o(n17443) );
na03f01 g13655 ( .a(n17194), .b(n17193), .c(n_17093), .o(n17444) );
oa12f01 g13656 ( .a(n7550), .b(n17255), .c(n17254), .o(n17445) );
ao12f01 g13657 ( .a(n17278), .b(n17445), .c(n17444), .o(n17446) );
no03f01 g13658 ( .a(n17446), .b(n17252), .c(n17443), .o(n17447) );
no02f01 g13659 ( .a(n17335), .b(n7550), .o(n17448) );
in01f01 g13660 ( .a(n17308), .o(n17449) );
ao12f01 g13661 ( .a(n7550), .b(n17449), .c(n17306), .o(n17450) );
no04f01 g13662 ( .a(n17450), .b(n17448), .c(n17447), .d(n17439), .o(n17451) );
na03f01 g13663 ( .a(n17320), .b(n17323), .c(n_17093), .o(n17452) );
oa12f01 g13664 ( .a(n7550), .b(n17321), .c(n17319), .o(n17453) );
oa12f01 g13665 ( .a(n7550), .b(n17308), .c(n17307), .o(n17454) );
na03f01 g13666 ( .a(n17454), .b(n17453), .c(n17452), .o(n17455) );
oa12f01 g13667 ( .a(n7550), .b(n17455), .c(n17451), .o(n17456) );
in01f01 g13668 ( .a(n17329), .o(n17457) );
ao12f01 g13669 ( .a(n17336), .b(n17457), .c(n17451), .o(n17458) );
no02f01 g13670 ( .a(n17398), .b(n7550), .o(n17459) );
ao12f01 g13671 ( .a(n17459), .b(n17458), .c(n17456), .o(n17460) );
in01f01 g13672 ( .a(n17361), .o(n17461) );
na02f01 g13673 ( .a(n17362), .b(n17461), .o(n17462) );
na02f01 g13674 ( .a(n17462), .b(n_17093), .o(n17463) );
na02f01 g13675 ( .a(n17463), .b(n17460), .o(n17464) );
no02f01 g13676 ( .a(n17401), .b(n7550), .o(n17465) );
no03f01 g13677 ( .a(n17394), .b(n17465), .c(n17464), .o(n17466) );
in01f01 g13678 ( .a(n17399), .o(n17467) );
na02f01 g13679 ( .a(n17383), .b(n7550), .o(n17468) );
in01f01 g13680 ( .a(n17403), .o(n17469) );
na03f01 g13681 ( .a(n17469), .b(n17468), .c(n17467), .o(n17470) );
in01f01 g13682 ( .a(n17413), .o(n17471) );
na02f01 g13683 ( .a(n17414), .b(n17471), .o(n17472) );
na02f01 g13684 ( .a(n17472), .b(n_17093), .o(n17473) );
oa12f01 g13685 ( .a(n17473), .b(n17470), .c(n17466), .o(n17474) );
na02f01 g13686 ( .a(n17472), .b(n7550), .o(n17475) );
na03f01 g13687 ( .a(n17436), .b(n17475), .c(n17474), .o(n17476) );
na03f01 g13688 ( .a(n17476), .b(n17438), .c(n16835), .o(n17477) );
na02f01 g13689 ( .a(n16772), .b(n16831), .o(n17478) );
ao22f01 g13690 ( .a(n16833), .b(n16831), .c(n16832), .d(n17478), .o(n17479) );
ao12f01 g13691 ( .a(n17436), .b(n17475), .c(n17474), .o(n17480) );
no03f01 g13692 ( .a(n17437), .b(n17419), .c(n17418), .o(n17481) );
oa12f01 g13693 ( .a(n17479), .b(n17481), .c(n17480), .o(n17482) );
na02f01 g13694 ( .a(n17482), .b(n17477), .o(n17483) );
in01f01 g13695 ( .a(n17483), .o(n17484) );
na03f01 g13696 ( .a(n17469), .b(n17467), .c(n17464), .o(n17485) );
no02f01 g13697 ( .a(n17402), .b(n17465), .o(n17486) );
in01f01 g13698 ( .a(n17486), .o(n17487) );
ao12f01 g13699 ( .a(n17487), .b(n17485), .c(n17395), .o(n17488) );
no03f01 g13700 ( .a(n17403), .b(n17399), .c(n17366), .o(n17489) );
no03f01 g13701 ( .a(n17486), .b(n17489), .c(n17394), .o(n17490) );
no02f01 g13702 ( .a(n16755), .b(n16595), .o(n17491) );
ao12f01 g13703 ( .a(n16757), .b(n16826), .c(n16789), .o(n17492) );
no03f01 g13704 ( .a(n17492), .b(n17491), .c(n16752), .o(n17493) );
in01f01 g13705 ( .a(n17491), .o(n17494) );
oa12f01 g13706 ( .a(n16756), .b(n16746), .c(n16606), .o(n17495) );
ao12f01 g13707 ( .a(n17494), .b(n17495), .c(n16827), .o(n17496) );
no02f01 g13708 ( .a(n17496), .b(n17493), .o(n17497) );
oa12f01 g13709 ( .a(n17497), .b(n17490), .c(n17488), .o(n17498) );
no02f01 g13710 ( .a(n17321), .b(n17319), .o(n17499) );
no03f01 g13711 ( .a(n17336), .b(n17326), .c(n17451), .o(n17500) );
no02f01 g13712 ( .a(n17500), .b(n17499), .o(n17501) );
in01f01 g13713 ( .a(n17501), .o(n17502) );
na02f01 g13714 ( .a(n17500), .b(n17499), .o(n17503) );
no02f01 g13715 ( .a(n16740), .b(n16625), .o(n17504) );
in01f01 g13716 ( .a(n17504), .o(n17505) );
no03f01 g13717 ( .a(n17505), .b(n16738), .c(n16637), .o(n17506) );
ao12f01 g13718 ( .a(n17504), .b(n16821), .c(n16792), .o(n17507) );
no02f01 g13719 ( .a(n17507), .b(n17506), .o(n17508) );
in01f01 g13720 ( .a(n17508), .o(n17509) );
ao12f01 g13721 ( .a(n17509), .b(n17503), .c(n17502), .o(n17510) );
no03f01 g13722 ( .a(n17448), .b(n17447), .c(n17439), .o(n17511) );
in01f01 g13723 ( .a(n17325), .o(n17512) );
oa12f01 g13724 ( .a(n17512), .b(n17336), .c(n17511), .o(n17513) );
in01f01 g13725 ( .a(n17513), .o(n17514) );
no03f01 g13726 ( .a(n17336), .b(n17512), .c(n17511), .o(n17515) );
no02f01 g13727 ( .a(n16736), .b(n16642), .o(n17516) );
in01f01 g13728 ( .a(n17516), .o(n17517) );
no02f01 g13729 ( .a(n16737), .b(n16637), .o(n17518) );
no02f01 g13730 ( .a(n17518), .b(n17517), .o(n17519) );
na02f01 g13731 ( .a(n17518), .b(n17517), .o(n17520) );
in01f01 g13732 ( .a(n17520), .o(n17521) );
no02f01 g13733 ( .a(n17521), .b(n17519), .o(n17522) );
no03f01 g13734 ( .a(n17522), .b(n17515), .c(n17514), .o(n17523) );
no02f01 g13735 ( .a(n17332), .b(n_17093), .o(n17524) );
ao12f01 g13736 ( .a(n17524), .b(n17281), .c(n17190), .o(n17525) );
no02f01 g13737 ( .a(n17335), .b(n_17093), .o(n17526) );
no02f01 g13738 ( .a(n17448), .b(n17526), .o(n17527) );
no02f01 g13739 ( .a(n17527), .b(n17525), .o(n17528) );
na02f01 g13740 ( .a(n17189), .b(n7550), .o(n17529) );
oa12f01 g13741 ( .a(n17529), .b(n17447), .c(n17439), .o(n17530) );
na02f01 g13742 ( .a(n17295), .b(n7550), .o(n17531) );
na02f01 g13743 ( .a(n17296), .b(n17531), .o(n17532) );
no02f01 g13744 ( .a(n17532), .b(n17530), .o(n17533) );
no02f01 g13745 ( .a(n16733), .b(n16650), .o(n17534) );
no02f01 g13746 ( .a(n16735), .b(n16642), .o(n17535) );
no02f01 g13747 ( .a(n17535), .b(n17534), .o(n17536) );
na02f01 g13748 ( .a(n17535), .b(n17534), .o(n17537) );
in01f01 g13749 ( .a(n17537), .o(n17538) );
no02f01 g13750 ( .a(n17538), .b(n17536), .o(n17539) );
no03f01 g13751 ( .a(n17539), .b(n17533), .c(n17528), .o(n17540) );
na02f01 g13752 ( .a(n17447), .b(n17332), .o(n17541) );
na02f01 g13753 ( .a(n17281), .b(n17189), .o(n17542) );
no02f01 g13754 ( .a(n16731), .b(n16656), .o(n17543) );
no02f01 g13755 ( .a(n16732), .b(n16650), .o(n17544) );
in01f01 g13756 ( .a(n17544), .o(n17545) );
no02f01 g13757 ( .a(n17545), .b(n17543), .o(n17546) );
na02f01 g13758 ( .a(n17545), .b(n17543), .o(n17547) );
in01f01 g13759 ( .a(n17547), .o(n17548) );
no02f01 g13760 ( .a(n17548), .b(n17546), .o(n17549) );
in01f01 g13761 ( .a(n17549), .o(n17550) );
na03f01 g13762 ( .a(n17550), .b(n17542), .c(n17541), .o(n17551) );
ao12f01 g13763 ( .a(n17550), .b(n17542), .c(n17541), .o(n17552) );
na02f01 g13764 ( .a(n17253), .b(n17442), .o(n17553) );
no02f01 g13765 ( .a(n17553), .b(n17195), .o(n17554) );
na02f01 g13766 ( .a(n17553), .b(n17195), .o(n17555) );
in01f01 g13767 ( .a(n17555), .o(n17556) );
no02f01 g13768 ( .a(n17556), .b(n17554), .o(n17557) );
no02f01 g13769 ( .a(n16730), .b(n16656), .o(n17558) );
in01f01 g13770 ( .a(n17558), .o(n17559) );
no03f01 g13771 ( .a(n17559), .b(n16728), .c(n16665), .o(n17560) );
ao12f01 g13772 ( .a(n17558), .b(n16815), .c(n16796), .o(n17561) );
no02f01 g13773 ( .a(n17561), .b(n17560), .o(n17562) );
in01f01 g13774 ( .a(n17562), .o(n17563) );
no02f01 g13775 ( .a(n16725), .b(n16672), .o(n17564) );
in01f01 g13776 ( .a(n17564), .o(n17565) );
no03f01 g13777 ( .a(n17565), .b(n16723), .c(n16686), .o(n17566) );
ao12f01 g13778 ( .a(n17564), .b(n16811), .c(n16685), .o(n17567) );
no02f01 g13779 ( .a(n17567), .b(n17566), .o(n17568) );
in01f01 g13780 ( .a(n17568), .o(n17569) );
in01f01 g13781 ( .a(n17236), .o(n17570) );
no02f01 g13782 ( .a(n17570), .b(n17229), .o(n17571) );
no02f01 g13783 ( .a(n17236), .b(n17272), .o(n17572) );
no02f01 g13784 ( .a(n17572), .b(n17571), .o(n17573) );
na02f01 g13785 ( .a(n17573), .b(n17569), .o(n17574) );
in01f01 g13786 ( .a(n17574), .o(n17575) );
no02f01 g13787 ( .a(n17228), .b(n17251), .o(n17576) );
no02f01 g13788 ( .a(n17271), .b(n17200), .o(n17577) );
no02f01 g13789 ( .a(n17577), .b(n17576), .o(n17578) );
no02f01 g13790 ( .a(n16721), .b(n16693), .o(n17579) );
in01f01 g13791 ( .a(n17579), .o(n17580) );
no02f01 g13792 ( .a(n16722), .b(n16686), .o(n17581) );
no02f01 g13793 ( .a(n17581), .b(n17580), .o(n17582) );
na02f01 g13794 ( .a(n17581), .b(n17580), .o(n17583) );
in01f01 g13795 ( .a(n17583), .o(n17584) );
no02f01 g13796 ( .a(n17584), .b(n17582), .o(n17585) );
in01f01 g13797 ( .a(n17585), .o(n17586) );
na02f01 g13798 ( .a(n17586), .b(n17578), .o(n17587) );
na02f01 g13799 ( .a(n17226), .b(n17263), .o(n17588) );
na02f01 g13800 ( .a(n17269), .b(n17214), .o(n17589) );
na02f01 g13801 ( .a(n17589), .b(n17588), .o(n17590) );
no03f01 g13802 ( .a(n16716), .b(n16805), .c(n16702), .o(n17591) );
ao12f01 g13803 ( .a(n16715), .b(n16806), .c(n16799), .o(n17592) );
no02f01 g13804 ( .a(n17592), .b(n17591), .o(n17593) );
no02f01 g13805 ( .a(n17593), .b(n17590), .o(n17594) );
in01f01 g13806 ( .a(n17594), .o(n17595) );
in01f01 g13807 ( .a(n17593), .o(n17596) );
ao12f01 g13808 ( .a(n17596), .b(n17589), .c(n17588), .o(n17597) );
in01f01 g13809 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_0_), .o(n17598) );
no02f01 g13810 ( .a(n16712), .b(n17598), .o(n17599) );
no02f01 g13811 ( .a(n16711), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_0_), .o(n17600) );
no02f01 g13812 ( .a(n17600), .b(n17599), .o(n17601) );
no02f01 g13813 ( .a(n17601), .b(n17225), .o(n17602) );
no03f01 g13814 ( .a(n16714), .b(n16804), .c(n16707), .o(n17603) );
ao12f01 g13815 ( .a(n16713), .b(n16708), .c(n16803), .o(n17604) );
no02f01 g13816 ( .a(n17604), .b(n17603), .o(n17605) );
no02f01 g13817 ( .a(n17605), .b(n17602), .o(n17606) );
no03f01 g13818 ( .a(n17225), .b(n17266), .c(n7550), .o(n17607) );
ao12f01 g13819 ( .a(n17219), .b(n17268), .c(n_17093), .o(n17608) );
no02f01 g13820 ( .a(n17608), .b(n17607), .o(n17609) );
na02f01 g13821 ( .a(n17605), .b(n17602), .o(n17610) );
ao12f01 g13822 ( .a(n17606), .b(n17610), .c(n17609), .o(n17611) );
oa12f01 g13823 ( .a(n17595), .b(n17611), .c(n17597), .o(n17612) );
na02f01 g13824 ( .a(n17227), .b(n17260), .o(n17613) );
na02f01 g13825 ( .a(n17270), .b(n17207), .o(n17614) );
na02f01 g13826 ( .a(n17614), .b(n17613), .o(n17615) );
no02f01 g13827 ( .a(n16717), .b(n16702), .o(n17616) );
no02f01 g13828 ( .a(n16720), .b(n16693), .o(n17617) );
no02f01 g13829 ( .a(n17617), .b(n17616), .o(n17618) );
na02f01 g13830 ( .a(n17617), .b(n17616), .o(n17619) );
in01f01 g13831 ( .a(n17619), .o(n17620) );
no02f01 g13832 ( .a(n17620), .b(n17618), .o(n17621) );
na02f01 g13833 ( .a(n17621), .b(n17615), .o(n17622) );
no02f01 g13834 ( .a(n17621), .b(n17615), .o(n17623) );
ao12f01 g13835 ( .a(n17623), .b(n17622), .c(n17612), .o(n17624) );
no02f01 g13836 ( .a(n17586), .b(n17578), .o(n17625) );
oa12f01 g13837 ( .a(n17587), .b(n17625), .c(n17624), .o(n17626) );
oa12f01 g13838 ( .a(n17568), .b(n17572), .c(n17571), .o(n17627) );
ao12f01 g13839 ( .a(n17575), .b(n17627), .c(n17626), .o(n17628) );
no02f01 g13840 ( .a(n17245), .b(n17243), .o(n17629) );
na02f01 g13841 ( .a(n17629), .b(n17237), .o(n17630) );
na02f01 g13842 ( .a(n17241), .b(n17240), .o(n17631) );
na02f01 g13843 ( .a(n17631), .b(n17276), .o(n17632) );
na02f01 g13844 ( .a(n17632), .b(n17630), .o(n17633) );
no02f01 g13845 ( .a(n16726), .b(n16672), .o(n17634) );
no02f01 g13846 ( .a(n16727), .b(n16665), .o(n17635) );
in01f01 g13847 ( .a(n17635), .o(n17636) );
no02f01 g13848 ( .a(n17636), .b(n17634), .o(n17637) );
na02f01 g13849 ( .a(n17636), .b(n17634), .o(n17638) );
in01f01 g13850 ( .a(n17638), .o(n17639) );
no02f01 g13851 ( .a(n17639), .b(n17637), .o(n17640) );
na02f01 g13852 ( .a(n17640), .b(n17633), .o(n17641) );
in01f01 g13853 ( .a(n17641), .o(n17642) );
in01f01 g13854 ( .a(n17640), .o(n17643) );
na03f01 g13855 ( .a(n17643), .b(n17632), .c(n17630), .o(n17644) );
na02f01 g13856 ( .a(n17644), .b(n17562), .o(n17645) );
in01f01 g13857 ( .a(n17645), .o(n17646) );
oa12f01 g13858 ( .a(n17646), .b(n17642), .c(n17628), .o(n17647) );
oa12f01 g13859 ( .a(n17644), .b(n17642), .c(n17628), .o(n17648) );
ao22f01 g13860 ( .a(n17648), .b(n17563), .c(n17647), .d(n17557), .o(n17649) );
oa12f01 g13861 ( .a(n17551), .b(n17649), .c(n17552), .o(n17650) );
oa12f01 g13862 ( .a(n17539), .b(n17533), .c(n17528), .o(n17651) );
oa12f01 g13863 ( .a(n17651), .b(n17650), .c(n17540), .o(n17652) );
in01f01 g13864 ( .a(n17515), .o(n17653) );
in01f01 g13865 ( .a(n17522), .o(n17654) );
ao12f01 g13866 ( .a(n17654), .b(n17653), .c(n17513), .o(n17655) );
no02f01 g13867 ( .a(n17655), .b(n17652), .o(n17656) );
in01f01 g13868 ( .a(n17503), .o(n17657) );
no03f01 g13869 ( .a(n17508), .b(n17657), .c(n17501), .o(n17658) );
no03f01 g13870 ( .a(n17658), .b(n17656), .c(n17523), .o(n17659) );
no02f01 g13871 ( .a(n17338), .b(n17328), .o(n17660) );
no02f01 g13872 ( .a(n17398), .b(n_17093), .o(n17661) );
no02f01 g13873 ( .a(n17661), .b(n17459), .o(n17662) );
na02f01 g13874 ( .a(n17662), .b(n17660), .o(n17663) );
no02f01 g13875 ( .a(n17662), .b(n17660), .o(n17664) );
in01f01 g13876 ( .a(n17664), .o(n17665) );
no02f01 g13877 ( .a(n16741), .b(n16625), .o(n17666) );
no02f01 g13878 ( .a(n16742), .b(n16616), .o(n17667) );
in01f01 g13879 ( .a(n17667), .o(n17668) );
no02f01 g13880 ( .a(n17668), .b(n17666), .o(n17669) );
na02f01 g13881 ( .a(n17668), .b(n17666), .o(n17670) );
in01f01 g13882 ( .a(n17670), .o(n17671) );
no02f01 g13883 ( .a(n17671), .b(n17669), .o(n17672) );
in01f01 g13884 ( .a(n17672), .o(n17673) );
ao12f01 g13885 ( .a(n17673), .b(n17665), .c(n17663), .o(n17674) );
no03f01 g13886 ( .a(n17674), .b(n17659), .c(n17510), .o(n17675) );
na03f01 g13887 ( .a(n17673), .b(n17665), .c(n17663), .o(n17676) );
in01f01 g13888 ( .a(n17661), .o(n17677) );
no02f01 g13889 ( .a(n17364), .b(n_17093), .o(n17678) );
no02f01 g13890 ( .a(n17678), .b(n17365), .o(n17679) );
na03f01 g13891 ( .a(n17679), .b(n17677), .c(n17351), .o(n17680) );
na02f01 g13892 ( .a(n17462), .b(n7550), .o(n17681) );
na02f01 g13893 ( .a(n17681), .b(n17463), .o(n17682) );
oa12f01 g13894 ( .a(n17682), .b(n17661), .c(n17460), .o(n17683) );
no02f01 g13895 ( .a(n16745), .b(n16606), .o(n17684) );
na03f01 g13896 ( .a(n17684), .b(n16825), .c(n16790), .o(n17685) );
in01f01 g13897 ( .a(n17684), .o(n17686) );
oa12f01 g13898 ( .a(n17686), .b(n16743), .c(n16616), .o(n17687) );
na02f01 g13899 ( .a(n17687), .b(n17685), .o(n17688) );
na03f01 g13900 ( .a(n17688), .b(n17683), .c(n17680), .o(n17689) );
na02f01 g13901 ( .a(n17689), .b(n17676), .o(n17690) );
ao12f01 g13902 ( .a(n17688), .b(n17683), .c(n17680), .o(n17691) );
in01f01 g13903 ( .a(n17691), .o(n17692) );
oa12f01 g13904 ( .a(n17692), .b(n17690), .c(n17675), .o(n17693) );
no02f01 g13905 ( .a(n17399), .b(n17366), .o(n17694) );
no02f01 g13906 ( .a(n17403), .b(n17394), .o(n17695) );
no02f01 g13907 ( .a(n17695), .b(n17694), .o(n17696) );
na02f01 g13908 ( .a(n17467), .b(n17464), .o(n17697) );
in01f01 g13909 ( .a(n17695), .o(n17698) );
no02f01 g13910 ( .a(n17698), .b(n17697), .o(n17699) );
no02f01 g13911 ( .a(n17699), .b(n17696), .o(n17700) );
no02f01 g13912 ( .a(n16757), .b(n16752), .o(n17701) );
oa12f01 g13913 ( .a(n17701), .b(n16746), .c(n16606), .o(n17702) );
in01f01 g13914 ( .a(n17701), .o(n17703) );
na03f01 g13915 ( .a(n17703), .b(n16826), .c(n16789), .o(n17704) );
na02f01 g13916 ( .a(n17704), .b(n17702), .o(n17705) );
no02f01 g13917 ( .a(n17705), .b(n17700), .o(n17706) );
na02f01 g13918 ( .a(n17698), .b(n17697), .o(n17707) );
na02f01 g13919 ( .a(n17695), .b(n17694), .o(n17708) );
na02f01 g13920 ( .a(n17708), .b(n17707), .o(n17709) );
ao12f01 g13921 ( .a(n17703), .b(n16826), .c(n16789), .o(n17710) );
no03f01 g13922 ( .a(n17701), .b(n16746), .c(n16606), .o(n17711) );
no02f01 g13923 ( .a(n17711), .b(n17710), .o(n17712) );
no02f01 g13924 ( .a(n17712), .b(n17709), .o(n17713) );
no03f01 g13925 ( .a(n17497), .b(n17490), .c(n17488), .o(n17714) );
no02f01 g13926 ( .a(n17714), .b(n17713), .o(n17715) );
oa12f01 g13927 ( .a(n17715), .b(n17706), .c(n17693), .o(n17716) );
na04f01 g13928 ( .a(n17475), .b(n17473), .c(n17404), .d(n17396), .o(n17717) );
oa22f01 g13929 ( .a(n17419), .b(n17417), .c(n17470), .d(n17466), .o(n17718) );
no02f01 g13930 ( .a(n16773), .b(n16770), .o(n17719) );
in01f01 g13931 ( .a(n17719), .o(n17720) );
na02f01 g13932 ( .a(n17720), .b(n16829), .o(n17721) );
na02f01 g13933 ( .a(n17719), .b(n16760), .o(n17722) );
na02f01 g13934 ( .a(n17722), .b(n17721), .o(n17723) );
ao12f01 g13935 ( .a(n17723), .b(n17718), .c(n17717), .o(n17724) );
in01f01 g13936 ( .a(n17724), .o(n17725) );
na03f01 g13937 ( .a(n17725), .b(n17716), .c(n17498), .o(n17726) );
na03f01 g13938 ( .a(n17723), .b(n17718), .c(n17717), .o(n17727) );
na03f01 g13939 ( .a(n17727), .b(n17726), .c(n17484), .o(n17728) );
oa12f01 g13940 ( .a(n17486), .b(n17489), .c(n17394), .o(n17729) );
na03f01 g13941 ( .a(n17487), .b(n17485), .c(n17395), .o(n17730) );
na03f01 g13942 ( .a(n17495), .b(n17494), .c(n16827), .o(n17731) );
oa12f01 g13943 ( .a(n17491), .b(n17492), .c(n16752), .o(n17732) );
na02f01 g13944 ( .a(n17732), .b(n17731), .o(n17733) );
ao12f01 g13945 ( .a(n17733), .b(n17730), .c(n17729), .o(n17734) );
in01f01 g13946 ( .a(n17510), .o(n17735) );
in01f01 g13947 ( .a(n17523), .o(n17736) );
na02f01 g13948 ( .a(n17532), .b(n17530), .o(n17737) );
na02f01 g13949 ( .a(n17527), .b(n17525), .o(n17738) );
in01f01 g13950 ( .a(n17539), .o(n17739) );
na03f01 g13951 ( .a(n17739), .b(n17738), .c(n17737), .o(n17740) );
no04f01 g13952 ( .a(n17446), .b(n17252), .c(n17443), .d(n17189), .o(n17741) );
no02f01 g13953 ( .a(n17447), .b(n17332), .o(n17742) );
no03f01 g13954 ( .a(n17549), .b(n17742), .c(n17741), .o(n17743) );
oa12f01 g13955 ( .a(n17549), .b(n17742), .c(n17741), .o(n17744) );
in01f01 g13956 ( .a(n17554), .o(n17745) );
na02f01 g13957 ( .a(n17555), .b(n17745), .o(n17746) );
na02f01 g13958 ( .a(n17271), .b(n17200), .o(n17747) );
na02f01 g13959 ( .a(n17228), .b(n17251), .o(n17748) );
na02f01 g13960 ( .a(n17748), .b(n17747), .o(n17749) );
no02f01 g13961 ( .a(n17585), .b(n17749), .o(n17750) );
no02f01 g13962 ( .a(n17611), .b(n17597), .o(n17751) );
no02f01 g13963 ( .a(n17751), .b(n17594), .o(n17752) );
no02f01 g13964 ( .a(n17270), .b(n17207), .o(n17753) );
no02f01 g13965 ( .a(n17227), .b(n17260), .o(n17754) );
no02f01 g13966 ( .a(n17754), .b(n17753), .o(n17755) );
in01f01 g13967 ( .a(n17621), .o(n17756) );
no02f01 g13968 ( .a(n17756), .b(n17755), .o(n17757) );
na02f01 g13969 ( .a(n17756), .b(n17755), .o(n17758) );
oa12f01 g13970 ( .a(n17758), .b(n17757), .c(n17752), .o(n17759) );
na02f01 g13971 ( .a(n17585), .b(n17749), .o(n17760) );
ao12f01 g13972 ( .a(n17750), .b(n17760), .c(n17759), .o(n17761) );
in01f01 g13973 ( .a(n17627), .o(n17762) );
oa12f01 g13974 ( .a(n17574), .b(n17762), .c(n17761), .o(n17763) );
ao12f01 g13975 ( .a(n17645), .b(n17641), .c(n17763), .o(n17764) );
in01f01 g13976 ( .a(n17644), .o(n17765) );
ao12f01 g13977 ( .a(n17765), .b(n17641), .c(n17763), .o(n17766) );
oa22f01 g13978 ( .a(n17766), .b(n17562), .c(n17764), .d(n17746), .o(n17767) );
ao12f01 g13979 ( .a(n17743), .b(n17767), .c(n17744), .o(n17768) );
ao12f01 g13980 ( .a(n17739), .b(n17738), .c(n17737), .o(n17769) );
ao12f01 g13981 ( .a(n17769), .b(n17768), .c(n17740), .o(n17770) );
oa12f01 g13982 ( .a(n17522), .b(n17515), .c(n17514), .o(n17771) );
na02f01 g13983 ( .a(n17771), .b(n17770), .o(n17772) );
na03f01 g13984 ( .a(n17509), .b(n17503), .c(n17502), .o(n17773) );
na03f01 g13985 ( .a(n17773), .b(n17772), .c(n17736), .o(n17774) );
in01f01 g13986 ( .a(n17663), .o(n17775) );
oa12f01 g13987 ( .a(n17672), .b(n17664), .c(n17775), .o(n17776) );
na03f01 g13988 ( .a(n17776), .b(n17774), .c(n17735), .o(n17777) );
no03f01 g13989 ( .a(n17672), .b(n17664), .c(n17775), .o(n17778) );
no03f01 g13990 ( .a(n17682), .b(n17661), .c(n17460), .o(n17779) );
ao12f01 g13991 ( .a(n17679), .b(n17677), .c(n17351), .o(n17780) );
no03f01 g13992 ( .a(n17686), .b(n16743), .c(n16616), .o(n17781) );
ao12f01 g13993 ( .a(n17684), .b(n16825), .c(n16790), .o(n17782) );
no02f01 g13994 ( .a(n17782), .b(n17781), .o(n17783) );
no03f01 g13995 ( .a(n17783), .b(n17780), .c(n17779), .o(n17784) );
no02f01 g13996 ( .a(n17784), .b(n17778), .o(n17785) );
ao12f01 g13997 ( .a(n17691), .b(n17785), .c(n17777), .o(n17786) );
na02f01 g13998 ( .a(n17712), .b(n17709), .o(n17787) );
na02f01 g13999 ( .a(n17705), .b(n17700), .o(n17788) );
na03f01 g14000 ( .a(n17733), .b(n17730), .c(n17729), .o(n17789) );
na02f01 g14001 ( .a(n17789), .b(n17788), .o(n17790) );
ao12f01 g14002 ( .a(n17790), .b(n17787), .c(n17786), .o(n17791) );
no03f01 g14003 ( .a(n17724), .b(n17791), .c(n17734), .o(n17792) );
in01f01 g14004 ( .a(n17727), .o(n17793) );
oa12f01 g14005 ( .a(n17483), .b(n17793), .c(n17792), .o(n17794) );
ao12f01 g14006 ( .a(n7682), .b(n17794), .c(n17728), .o(n17795) );
ao12f01 g14007 ( .a(n7712), .b(n17794), .c(n17728), .o(n17796) );
ao12f01 g14008 ( .a(n17523), .b(n17771), .c(n17770), .o(n17797) );
ao12f01 g14009 ( .a(n17510), .b(n17773), .c(n17797), .o(n17798) );
ao12f01 g14010 ( .a(n17690), .b(n17776), .c(n17798), .o(n17799) );
oa12f01 g14011 ( .a(n17788), .b(n17691), .c(n17799), .o(n17800) );
na02f01 g14012 ( .a(n17789), .b(n17498), .o(n17801) );
ao12f01 g14013 ( .a(n17801), .b(n17800), .c(n17787), .o(n17802) );
oa12f01 g14014 ( .a(n17736), .b(n17655), .c(n17652), .o(n17803) );
oa12f01 g14015 ( .a(n17735), .b(n17658), .c(n17803), .o(n17804) );
oa12f01 g14016 ( .a(n17785), .b(n17674), .c(n17804), .o(n17805) );
ao12f01 g14017 ( .a(n17713), .b(n17692), .c(n17805), .o(n17806) );
no02f01 g14018 ( .a(n17714), .b(n17734), .o(n17807) );
no03f01 g14019 ( .a(n17807), .b(n17806), .c(n17706), .o(n17808) );
no02f01 g14020 ( .a(n17808), .b(n17802), .o(n17809) );
no02f01 g14021 ( .a(n17713), .b(n17706), .o(n17810) );
no02f01 g14022 ( .a(n17810), .b(n17693), .o(n17811) );
na02f01 g14023 ( .a(n17788), .b(n17787), .o(n17812) );
no02f01 g14024 ( .a(n17812), .b(n17786), .o(n17813) );
no02f01 g14025 ( .a(n17813), .b(n17811), .o(n17814) );
ao12f01 g14026 ( .a(n7712), .b(n17814), .c(n17809), .o(n17815) );
no02f01 g14027 ( .a(n17793), .b(n17724), .o(n17816) );
oa12f01 g14028 ( .a(n17816), .b(n17791), .c(n17734), .o(n17817) );
na02f01 g14029 ( .a(n17727), .b(n17725), .o(n17818) );
na03f01 g14030 ( .a(n17818), .b(n17716), .c(n17498), .o(n17819) );
ao12f01 g14031 ( .a(n7712), .b(n17819), .c(n17817), .o(n17820) );
no02f01 g14032 ( .a(n17820), .b(n17815), .o(n17821) );
ao12f01 g14033 ( .a(n7682), .b(n17819), .c(n17817), .o(n17822) );
no04f01 g14034 ( .a(n17822), .b(n17821), .c(n17796), .d(n17795), .o(n17823) );
no03f01 g14035 ( .a(n17793), .b(n17792), .c(n17483), .o(n17824) );
ao12f01 g14036 ( .a(n17484), .b(n17727), .c(n17726), .o(n17825) );
oa12f01 g14037 ( .a(n7712), .b(n17825), .c(n17824), .o(n17826) );
oa12f01 g14038 ( .a(n7682), .b(n17825), .c(n17824), .o(n17827) );
oa12f01 g14039 ( .a(n17807), .b(n17806), .c(n17706), .o(n17828) );
na03f01 g14040 ( .a(n17801), .b(n17800), .c(n17787), .o(n17829) );
na02f01 g14041 ( .a(n17829), .b(n17828), .o(n17830) );
na02f01 g14042 ( .a(n17812), .b(n17786), .o(n17831) );
na02f01 g14043 ( .a(n17810), .b(n17693), .o(n17832) );
na02f01 g14044 ( .a(n17832), .b(n17831), .o(n17833) );
oa12f01 g14045 ( .a(n7682), .b(n17833), .c(n17830), .o(n17834) );
ao12f01 g14046 ( .a(n17818), .b(n17716), .c(n17498), .o(n17835) );
no03f01 g14047 ( .a(n17816), .b(n17791), .c(n17734), .o(n17836) );
oa12f01 g14048 ( .a(n7682), .b(n17836), .c(n17835), .o(n17837) );
na02f01 g14049 ( .a(n17837), .b(n17834), .o(n17838) );
oa12f01 g14050 ( .a(n7712), .b(n17836), .c(n17835), .o(n17839) );
ao22f01 g14051 ( .a(n17839), .b(n17838), .c(n17827), .d(n17826), .o(n17840) );
no02f01 g14052 ( .a(n17719), .b(n16760), .o(n17841) );
no02f01 g14053 ( .a(n17720), .b(n16829), .o(n17842) );
no02f01 g14054 ( .a(n17842), .b(n17841), .o(n17843) );
no02f01 g14055 ( .a(n17497), .b(n7550), .o(n17844) );
na02f01 g14056 ( .a(n17688), .b(n_17093), .o(n17845) );
oa12f01 g14057 ( .a(n17845), .b(n17712), .c(n7550), .o(n17846) );
oa12f01 g14058 ( .a(n17843), .b(n17846), .c(n17844), .o(n17847) );
na02f01 g14059 ( .a(n17733), .b(n_17093), .o(n17848) );
no02f01 g14060 ( .a(n17783), .b(n7550), .o(n17849) );
ao12f01 g14061 ( .a(n17849), .b(n17705), .c(n_17093), .o(n17850) );
na03f01 g14062 ( .a(n17850), .b(n17848), .c(n17723), .o(n17851) );
na02f01 g14063 ( .a(n17162), .b(n17153), .o(n17852) );
no02f01 g14064 ( .a(n17068), .b(n17034), .o(n17853) );
in01f01 g14065 ( .a(n17853), .o(n17854) );
no02f01 g14066 ( .a(n17854), .b(n17852), .o(n17855) );
na02f01 g14067 ( .a(n17854), .b(n17852), .o(n17856) );
in01f01 g14068 ( .a(n17856), .o(n17857) );
no02f01 g14069 ( .a(n17857), .b(n17855), .o(n17858) );
ao12f01 g14070 ( .a(n17858), .b(n17851), .c(n17847), .o(n17859) );
ao12f01 g14071 ( .a(n17723), .b(n17850), .c(n17848), .o(n17860) );
no03f01 g14072 ( .a(n17846), .b(n17844), .c(n17843), .o(n17861) );
in01f01 g14073 ( .a(n17858), .o(n17862) );
no03f01 g14074 ( .a(n17862), .b(n17861), .c(n17860), .o(n17863) );
no02f01 g14075 ( .a(n17863), .b(n17859), .o(n17864) );
no02f01 g14076 ( .a(n17062), .b(delay_add_ln22_unr11_stage5_stallmux_q_0_), .o(n17865) );
no02f01 g14077 ( .a(n17061), .b(n17057), .o(n17866) );
no02f01 g14078 ( .a(n17866), .b(n17865), .o(n17867) );
no02f01 g14079 ( .a(n17867), .b(n17783), .o(n17868) );
in01f01 g14080 ( .a(n17868), .o(n17869) );
no03f01 g14081 ( .a(n17063), .b(n17158), .c(n17055), .o(n17870) );
ao12f01 g14082 ( .a(n17159), .b(n17056), .c(n17157), .o(n17871) );
no02f01 g14083 ( .a(n17871), .b(n17870), .o(n17872) );
no02f01 g14084 ( .a(n17872), .b(n17869), .o(n17873) );
in01f01 g14085 ( .a(n17873), .o(n17874) );
in01f01 g14086 ( .a(n17872), .o(n17875) );
no02f01 g14087 ( .a(n17849), .b(n17712), .o(n17876) );
no02f01 g14088 ( .a(n17845), .b(n17705), .o(n17877) );
oa22f01 g14089 ( .a(n17877), .b(n17876), .c(n17875), .d(n17868), .o(n17878) );
no02f01 g14090 ( .a(n17065), .b(n17043), .o(n17879) );
no02f01 g14091 ( .a(n17879), .b(n17064), .o(n17880) );
na02f01 g14092 ( .a(n17879), .b(n17064), .o(n17881) );
in01f01 g14093 ( .a(n17881), .o(n17882) );
no02f01 g14094 ( .a(n17882), .b(n17880), .o(n17883) );
ao12f01 g14095 ( .a(n17883), .b(n17878), .c(n17874), .o(n17884) );
na03f01 g14096 ( .a(n17883), .b(n17878), .c(n17874), .o(n17885) );
na02f01 g14097 ( .a(n17846), .b(n17497), .o(n17886) );
na02f01 g14098 ( .a(n17850), .b(n17733), .o(n17887) );
na02f01 g14099 ( .a(n17887), .b(n17886), .o(n17888) );
ao12f01 g14100 ( .a(n17884), .b(n17888), .c(n17885), .o(n17889) );
no02f01 g14101 ( .a(n17889), .b(n17864), .o(n17890) );
na02f01 g14102 ( .a(n17889), .b(n17864), .o(n17891) );
in01f01 g14103 ( .a(n17891), .o(n17892) );
no02f01 g14104 ( .a(n17892), .b(n17890), .o(n17893) );
in01f01 g14105 ( .a(n17893), .o(n17894) );
oa12f01 g14106 ( .a(n17894), .b(n17840), .c(n17823), .o(n17895) );
na04f01 g14107 ( .a(n17839), .b(n17838), .c(n17827), .d(n17826), .o(n17896) );
oa22f01 g14108 ( .a(n17822), .b(n17821), .c(n17796), .d(n17795), .o(n17897) );
na03f01 g14109 ( .a(n17893), .b(n17897), .c(n17896), .o(n17898) );
oa12f01 g14110 ( .a(n17834), .b(n17822), .c(n17820), .o(n17899) );
na03f01 g14111 ( .a(n17839), .b(n17837), .c(n17815), .o(n17900) );
na02f01 g14112 ( .a(n17845), .b(n17705), .o(n17901) );
na02f01 g14113 ( .a(n17849), .b(n17712), .o(n17902) );
ao22f01 g14114 ( .a(n17902), .b(n17901), .c(n17872), .d(n17869), .o(n17903) );
no02f01 g14115 ( .a(n17903), .b(n17873), .o(n17904) );
no02f01 g14116 ( .a(n17850), .b(n17733), .o(n17905) );
no02f01 g14117 ( .a(n17846), .b(n17497), .o(n17906) );
no02f01 g14118 ( .a(n17906), .b(n17905), .o(n17907) );
no02f01 g14119 ( .a(n17907), .b(n17883), .o(n17908) );
in01f01 g14120 ( .a(n17883), .o(n17909) );
no02f01 g14121 ( .a(n17888), .b(n17909), .o(n17910) );
no02f01 g14122 ( .a(n17910), .b(n17908), .o(n17911) );
no02f01 g14123 ( .a(n17911), .b(n17904), .o(n17912) );
na02f01 g14124 ( .a(n17911), .b(n17904), .o(n17913) );
in01f01 g14125 ( .a(n17913), .o(n17914) );
no02f01 g14126 ( .a(n17914), .b(n17912), .o(n17915) );
na03f01 g14127 ( .a(n17915), .b(n17900), .c(n17899), .o(n17916) );
no02f01 g14128 ( .a(n17833), .b(n7712), .o(n17917) );
no02f01 g14129 ( .a(n17833), .b(n7682), .o(n17918) );
no02f01 g14130 ( .a(n17867), .b(n17688), .o(n17919) );
in01f01 g14131 ( .a(n17867), .o(n17920) );
no02f01 g14132 ( .a(n17920), .b(n17783), .o(n17921) );
no02f01 g14133 ( .a(n17921), .b(n17919), .o(n17922) );
no03f01 g14134 ( .a(n17922), .b(n17918), .c(n17917), .o(n17923) );
no03f01 g14135 ( .a(n17877), .b(n17876), .c(n17875), .o(n17924) );
ao12f01 g14136 ( .a(n17872), .b(n17902), .c(n17901), .o(n17925) );
no02f01 g14137 ( .a(n17925), .b(n17924), .o(n17926) );
no02f01 g14138 ( .a(n17926), .b(n17869), .o(n17927) );
na02f01 g14139 ( .a(n17926), .b(n17869), .o(n17928) );
in01f01 g14140 ( .a(n17928), .o(n17929) );
no02f01 g14141 ( .a(n17929), .b(n17927), .o(n17930) );
in01f01 g14142 ( .a(n17930), .o(n17931) );
no02f01 g14143 ( .a(n17931), .b(n17923), .o(n17932) );
no03f01 g14144 ( .a(n17814), .b(n17830), .c(n7712), .o(n17933) );
ao12f01 g14145 ( .a(n17809), .b(n17833), .c(n7682), .o(n17934) );
no02f01 g14146 ( .a(n17934), .b(n17933), .o(n17935) );
na02f01 g14147 ( .a(n17931), .b(n17923), .o(n17936) );
oa12f01 g14148 ( .a(n17936), .b(n17935), .c(n17932), .o(n17937) );
ao12f01 g14149 ( .a(n17915), .b(n17900), .c(n17899), .o(n17938) );
ao12f01 g14150 ( .a(n17938), .b(n17937), .c(n17916), .o(n17939) );
na03f01 g14151 ( .a(n17939), .b(n17898), .c(n17895), .o(n17940) );
ao12f01 g14152 ( .a(n17893), .b(n17897), .c(n17896), .o(n17941) );
no03f01 g14153 ( .a(n17894), .b(n17840), .c(n17823), .o(n17942) );
ao12f01 g14154 ( .a(n17815), .b(n17839), .c(n17837), .o(n17943) );
no03f01 g14155 ( .a(n17822), .b(n17820), .c(n17834), .o(n17944) );
in01f01 g14156 ( .a(n17915), .o(n17945) );
no03f01 g14157 ( .a(n17945), .b(n17944), .c(n17943), .o(n17946) );
na02f01 g14158 ( .a(n17814), .b(n7682), .o(n17947) );
na02f01 g14159 ( .a(n17814), .b(n7712), .o(n17948) );
in01f01 g14160 ( .a(n17922), .o(n17949) );
na03f01 g14161 ( .a(n17949), .b(n17948), .c(n17947), .o(n17950) );
na02f01 g14162 ( .a(n17930), .b(n17950), .o(n17951) );
na03f01 g14163 ( .a(n17833), .b(n17809), .c(n7682), .o(n17952) );
oa12f01 g14164 ( .a(n17830), .b(n17814), .c(n7712), .o(n17953) );
na02f01 g14165 ( .a(n17953), .b(n17952), .o(n17954) );
no02f01 g14166 ( .a(n17930), .b(n17950), .o(n17955) );
ao12f01 g14167 ( .a(n17955), .b(n17954), .c(n17951), .o(n17956) );
oa12f01 g14168 ( .a(n17945), .b(n17944), .c(n17943), .o(n17957) );
oa12f01 g14169 ( .a(n17957), .b(n17956), .c(n17946), .o(n17958) );
oa12f01 g14170 ( .a(n17958), .b(n17942), .c(n17941), .o(n17959) );
na02f01 g14171 ( .a(n17959), .b(n17940), .o(n263) );
na03f01 g14172 ( .a(n7546), .b(n7516), .c(n7466), .o(n17961) );
oa12f01 g14173 ( .a(n7545), .b(n7520), .c(n7465), .o(n17962) );
na02f01 g14174 ( .a(n17962), .b(n17961), .o(n268) );
na02f01 g14175 ( .a(delay_xor_ln23_unr6_stage3_stallmux_q), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(n17964) );
in01f01 g14176 ( .a(n17964), .o(n17965) );
in01f01 g14177 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(n17966) );
no02f01 g14178 ( .a(delay_xor_ln23_unr6_stage3_stallmux_q), .b(n17966), .o(n17967) );
in01f01 g14179 ( .a(n17967), .o(n17968) );
no02f01 g14180 ( .a(n17968), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_24_), .o(n17969) );
in01f01 g14181 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_8_), .o(n17970) );
in01f01 g14182 ( .a(delay_xor_ln23_unr6_stage3_stallmux_q), .o(n17971) );
no02f01 g14183 ( .a(n17971), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(n17972) );
in01f01 g14184 ( .a(n17972), .o(n17973) );
no02f01 g14185 ( .a(n17973), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_3_), .o(n17974) );
in01f01 g14186 ( .a(n17974), .o(n17975) );
in01f01 g14187 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_2_), .o(n17976) );
no02f01 g14188 ( .a(n17967), .b(n17976), .o(n17977) );
in01f01 g14189 ( .a(n17977), .o(n17978) );
no02f01 g14190 ( .a(delay_xor_ln23_unr6_stage3_stallmux_q), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(n17979) );
in01f01 g14191 ( .a(n17979), .o(n17980) );
na02f01 g14192 ( .a(n17980), .b(n17964), .o(n17981) );
no02f01 g14193 ( .a(n17981), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_1_), .o(n17982) );
no02f01 g14194 ( .a(n17968), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_2_), .o(n17983) );
oa12f01 g14195 ( .a(n17978), .b(n17983), .c(n17982), .o(n17984) );
na02f01 g14196 ( .a(n17984), .b(n17975), .o(n17985) );
in01f01 g14197 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_3_), .o(n17986) );
no02f01 g14198 ( .a(n17972), .b(n17986), .o(n17987) );
in01f01 g14199 ( .a(n17987), .o(n17988) );
na02f01 g14200 ( .a(n17988), .b(n17985), .o(n17989) );
in01f01 g14201 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_4_), .o(n17990) );
na02f01 g14202 ( .a(n17985), .b(n17990), .o(n17991) );
ao22f01 g14203 ( .a(n17991), .b(n17968), .c(n17989), .d(delay_sub_ln23_0_unr5_stage3_stallmux_q_4_), .o(n17992) );
no02f01 g14204 ( .a(n17973), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_5_), .o(n17993) );
no02f01 g14205 ( .a(n17993), .b(n17992), .o(n17994) );
in01f01 g14206 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_6_), .o(n17995) );
no02f01 g14207 ( .a(n17967), .b(n17995), .o(n17996) );
na02f01 g14208 ( .a(n17973), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_5_), .o(n17997) );
in01f01 g14209 ( .a(n17997), .o(n17998) );
no02f01 g14210 ( .a(n17998), .b(n17996), .o(n17999) );
in01f01 g14211 ( .a(n17999), .o(n18000) );
no02f01 g14212 ( .a(n17968), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_6_), .o(n18001) );
in01f01 g14213 ( .a(n18001), .o(n18002) );
oa12f01 g14214 ( .a(n18002), .b(n18000), .c(n17994), .o(n18003) );
no02f01 g14215 ( .a(n17973), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_7_), .o(n18004) );
no02f01 g14216 ( .a(n18004), .b(n18003), .o(n18005) );
na02f01 g14217 ( .a(n18005), .b(n17968), .o(n18006) );
na02f01 g14218 ( .a(n17973), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_7_), .o(n18007) );
in01f01 g14219 ( .a(n18007), .o(n18008) );
no02f01 g14220 ( .a(n18008), .b(n17968), .o(n18009) );
in01f01 g14221 ( .a(n18009), .o(n18010) );
no02f01 g14222 ( .a(n18010), .b(n18005), .o(n18011) );
oa12f01 g14223 ( .a(n18006), .b(n18011), .c(n17970), .o(n18012) );
no02f01 g14224 ( .a(n17968), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_10_), .o(n18013) );
no02f01 g14225 ( .a(n17973), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_9_), .o(n18014) );
no02f01 g14226 ( .a(n18014), .b(n18013), .o(n18015) );
na02f01 g14227 ( .a(n18015), .b(n18012), .o(n18016) );
na02f01 g14228 ( .a(n17968), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_10_), .o(n18017) );
na02f01 g14229 ( .a(n17973), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_9_), .o(n18018) );
ao12f01 g14230 ( .a(n18013), .b(n18018), .c(n18017), .o(n18019) );
in01f01 g14231 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_12_), .o(n18020) );
in01f01 g14232 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_11_), .o(n18021) );
ao12f01 g14233 ( .a(n17972), .b(n18021), .c(n18020), .o(n18022) );
no02f01 g14234 ( .a(n18022), .b(n18019), .o(n18023) );
no02f01 g14235 ( .a(n17973), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_12_), .o(n18024) );
no02f01 g14236 ( .a(n17973), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_11_), .o(n18025) );
no02f01 g14237 ( .a(n18025), .b(n18024), .o(n18026) );
in01f01 g14238 ( .a(n18026), .o(n18027) );
ao12f01 g14239 ( .a(n18027), .b(n18023), .c(n18016), .o(n18028) );
in01f01 g14240 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_16_), .o(n18029) );
in01f01 g14241 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_15_), .o(n18030) );
ao12f01 g14242 ( .a(n17972), .b(n18030), .c(n18029), .o(n18031) );
in01f01 g14243 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_14_), .o(n18032) );
in01f01 g14244 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_13_), .o(n18033) );
ao12f01 g14245 ( .a(n17972), .b(n18033), .c(n18032), .o(n18034) );
no02f01 g14246 ( .a(n18034), .b(n18031), .o(n18035) );
in01f01 g14247 ( .a(n18035), .o(n18036) );
no02f01 g14248 ( .a(n17973), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_15_), .o(n18037) );
ao12f01 g14249 ( .a(n17973), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_13_), .c(delay_sub_ln23_0_unr5_stage3_stallmux_q_14_), .o(n18038) );
no02f01 g14250 ( .a(n18038), .b(n18037), .o(n18039) );
in01f01 g14251 ( .a(n18039), .o(n18040) );
no02f01 g14252 ( .a(n17973), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_16_), .o(n18041) );
no02f01 g14253 ( .a(n18041), .b(n18040), .o(n18042) );
oa12f01 g14254 ( .a(n18042), .b(n18036), .c(n18028), .o(n18043) );
no02f01 g14255 ( .a(n17973), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_18_), .o(n18044) );
no02f01 g14256 ( .a(n17973), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_19_), .o(n18045) );
no02f01 g14257 ( .a(n17973), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_20_), .o(n18046) );
no02f01 g14258 ( .a(n17973), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_17_), .o(n18047) );
no04f01 g14259 ( .a(n18047), .b(n18046), .c(n18045), .d(n18044), .o(n18048) );
in01f01 g14260 ( .a(n18048), .o(n18049) );
in01f01 g14261 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_19_), .o(n18050) );
in01f01 g14262 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_20_), .o(n18051) );
ao12f01 g14263 ( .a(n17972), .b(n18051), .c(n18050), .o(n18052) );
in01f01 g14264 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_18_), .o(n18053) );
in01f01 g14265 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_17_), .o(n18054) );
ao12f01 g14266 ( .a(n17972), .b(n18054), .c(n18053), .o(n18055) );
no02f01 g14267 ( .a(n18055), .b(n18052), .o(n18056) );
oa12f01 g14268 ( .a(n18056), .b(n18049), .c(n18043), .o(n18057) );
no02f01 g14269 ( .a(n17973), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_21_), .o(n18058) );
no02f01 g14270 ( .a(n17973), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_22_), .o(n18059) );
no02f01 g14271 ( .a(n18059), .b(n18058), .o(n18060) );
in01f01 g14272 ( .a(n18060), .o(n18061) );
no02f01 g14273 ( .a(n17973), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_23_), .o(n18062) );
no02f01 g14274 ( .a(n18062), .b(n18061), .o(n18063) );
in01f01 g14275 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_21_), .o(n18064) );
in01f01 g14276 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_22_), .o(n18065) );
ao12f01 g14277 ( .a(n17972), .b(n18065), .c(n18064), .o(n18066) );
na02f01 g14278 ( .a(n17973), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_23_), .o(n18067) );
in01f01 g14279 ( .a(n18067), .o(n18068) );
no02f01 g14280 ( .a(n18068), .b(n18066), .o(n18069) );
in01f01 g14281 ( .a(n18069), .o(n18070) );
na02f01 g14282 ( .a(n17968), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_24_), .o(n18071) );
in01f01 g14283 ( .a(n18071), .o(n18072) );
no02f01 g14284 ( .a(n18072), .b(n18070), .o(n18073) );
in01f01 g14285 ( .a(n18073), .o(n18074) );
ao12f01 g14286 ( .a(n18074), .b(n18063), .c(n18057), .o(n18075) );
no02f01 g14287 ( .a(n17968), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_25_), .o(n18076) );
no02f01 g14288 ( .a(n17968), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_26_), .o(n18077) );
no02f01 g14289 ( .a(n18077), .b(n18076), .o(n18078) );
in01f01 g14290 ( .a(n18078), .o(n18079) );
no02f01 g14291 ( .a(n17968), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_27_), .o(n18080) );
no02f01 g14292 ( .a(n17968), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_28_), .o(n18081) );
no03f01 g14293 ( .a(n18081), .b(n18080), .c(n18079), .o(n18082) );
in01f01 g14294 ( .a(n18082), .o(n18083) );
no02f01 g14295 ( .a(n17968), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_29_), .o(n18084) );
no02f01 g14296 ( .a(n17968), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_30_), .o(n18085) );
no02f01 g14297 ( .a(n18085), .b(n18084), .o(n18086) );
in01f01 g14298 ( .a(n18086), .o(n18087) );
no04f01 g14299 ( .a(n18087), .b(n18083), .c(n18075), .d(n17969), .o(n18088) );
in01f01 g14300 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_28_), .o(n18089) );
in01f01 g14301 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_27_), .o(n18090) );
ao12f01 g14302 ( .a(n17967), .b(n18090), .c(n18089), .o(n18091) );
in01f01 g14303 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_26_), .o(n18092) );
in01f01 g14304 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_25_), .o(n18093) );
ao12f01 g14305 ( .a(n17967), .b(n18093), .c(n18092), .o(n18094) );
no02f01 g14306 ( .a(n18094), .b(n18091), .o(n18095) );
in01f01 g14307 ( .a(n18095), .o(n18096) );
in01f01 g14308 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_29_), .o(n18097) );
in01f01 g14309 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_30_), .o(n18098) );
ao12f01 g14310 ( .a(n17967), .b(n18098), .c(n18097), .o(n18099) );
no02f01 g14311 ( .a(n18099), .b(n18096), .o(n18100) );
in01f01 g14312 ( .a(n18100), .o(n18101) );
no02f01 g14313 ( .a(n18101), .b(n18088), .o(n18102) );
no02f01 g14314 ( .a(n18102), .b(n17965), .o(n18103) );
in01f01 g14315 ( .a(n18056), .o(n18104) );
no02f01 g14316 ( .a(n18049), .b(n18043), .o(n18105) );
in01f01 g14317 ( .a(n18105), .o(n18106) );
no02f01 g14318 ( .a(n18061), .b(n18106), .o(n18107) );
no03f01 g14319 ( .a(n18107), .b(n18066), .c(n18104), .o(n18108) );
in01f01 g14320 ( .a(n18108), .o(n18109) );
no02f01 g14321 ( .a(n18068), .b(n18062), .o(n18110) );
in01f01 g14322 ( .a(n18110), .o(n18111) );
no02f01 g14323 ( .a(n18111), .b(n18109), .o(n18112) );
no02f01 g14324 ( .a(n18110), .b(n18108), .o(n18113) );
no03f01 g14325 ( .a(n18113), .b(n18112), .c(n18103), .o(n18114) );
no02f01 g14326 ( .a(n17972), .b(n18050), .o(n18115) );
no03f01 g14327 ( .a(n18047), .b(n18044), .c(n18043), .o(n18116) );
in01f01 g14328 ( .a(n18116), .o(n18117) );
no02f01 g14329 ( .a(n18117), .b(n18045), .o(n18118) );
no03f01 g14330 ( .a(n18118), .b(n18055), .c(n18115), .o(n18119) );
in01f01 g14331 ( .a(n18119), .o(n18120) );
no02f01 g14332 ( .a(n17972), .b(n18051), .o(n18121) );
no02f01 g14333 ( .a(n18121), .b(n18046), .o(n18122) );
in01f01 g14334 ( .a(n18122), .o(n18123) );
no02f01 g14335 ( .a(n18123), .b(n18120), .o(n18124) );
no02f01 g14336 ( .a(n18122), .b(n18119), .o(n18125) );
no02f01 g14337 ( .a(n18125), .b(n18124), .o(n18126) );
in01f01 g14338 ( .a(n18057), .o(n18127) );
no02f01 g14339 ( .a(n17972), .b(n18064), .o(n18128) );
no02f01 g14340 ( .a(n18128), .b(n18058), .o(n18129) );
no02f01 g14341 ( .a(n18129), .b(n18127), .o(n18130) );
na02f01 g14342 ( .a(n18129), .b(n18127), .o(n18131) );
in01f01 g14343 ( .a(n18131), .o(n18132) );
no02f01 g14344 ( .a(n18132), .b(n18130), .o(n18133) );
ao12f01 g14345 ( .a(n18103), .b(n18133), .c(n18126), .o(n18134) );
no02f01 g14346 ( .a(n18058), .b(n18106), .o(n18135) );
no03f01 g14347 ( .a(n18135), .b(n18128), .c(n18104), .o(n18136) );
no02f01 g14348 ( .a(n17972), .b(n18065), .o(n18137) );
no02f01 g14349 ( .a(n18137), .b(n18059), .o(n18138) );
no02f01 g14350 ( .a(n18138), .b(n18136), .o(n18139) );
na02f01 g14351 ( .a(n18138), .b(n18136), .o(n18140) );
in01f01 g14352 ( .a(n18140), .o(n18141) );
no02f01 g14353 ( .a(n18141), .b(n18139), .o(n18142) );
no02f01 g14354 ( .a(n18142), .b(n18103), .o(n18143) );
no02f01 g14355 ( .a(n18143), .b(n18134), .o(n18144) );
oa12f01 g14356 ( .a(n17964), .b(n18101), .c(n18088), .o(n18145) );
no02f01 g14357 ( .a(n18113), .b(n18112), .o(n18146) );
no02f01 g14358 ( .a(n18146), .b(n18145), .o(n18147) );
in01f01 g14359 ( .a(n18147), .o(n18148) );
ao12f01 g14360 ( .a(n18114), .b(n18148), .c(n18144), .o(n18149) );
no02f01 g14361 ( .a(n18008), .b(n18004), .o(n18150) );
no02f01 g14362 ( .a(n18150), .b(n18003), .o(n18151) );
na02f01 g14363 ( .a(n18150), .b(n18003), .o(n18152) );
in01f01 g14364 ( .a(n18152), .o(n18153) );
no02f01 g14365 ( .a(n18153), .b(n18151), .o(n18154) );
in01f01 g14366 ( .a(n18154), .o(n18155) );
no02f01 g14367 ( .a(n18155), .b(n18103), .o(n18156) );
in01f01 g14368 ( .a(n18156), .o(n18157) );
in01f01 g14369 ( .a(n17992), .o(n18158) );
no02f01 g14370 ( .a(n17998), .b(n17993), .o(n18159) );
in01f01 g14371 ( .a(n18159), .o(n18160) );
no02f01 g14372 ( .a(n18160), .b(n18158), .o(n18161) );
no02f01 g14373 ( .a(n18159), .b(n17992), .o(n18162) );
no02f01 g14374 ( .a(n18162), .b(n18161), .o(n18163) );
in01f01 g14375 ( .a(n18163), .o(n18164) );
no02f01 g14376 ( .a(n18164), .b(n18103), .o(n18165) );
in01f01 g14377 ( .a(n18165), .o(n18166) );
no02f01 g14378 ( .a(n17987), .b(n17974), .o(n18167) );
in01f01 g14379 ( .a(n18167), .o(n18168) );
no02f01 g14380 ( .a(n18168), .b(n17984), .o(n18169) );
in01f01 g14381 ( .a(n17984), .o(n18170) );
no02f01 g14382 ( .a(n18167), .b(n18170), .o(n18171) );
no02f01 g14383 ( .a(n18171), .b(n18169), .o(n18172) );
no02f01 g14384 ( .a(n18172), .b(n18145), .o(n18173) );
no04f01 g14385 ( .a(n17983), .b(n17981), .c(n17977), .d(delay_sub_ln23_0_unr5_stage3_stallmux_q_1_), .o(n18174) );
no02f01 g14386 ( .a(n17983), .b(n17977), .o(n18175) );
no02f01 g14387 ( .a(n18175), .b(n17982), .o(n18176) );
no02f01 g14388 ( .a(n18176), .b(n18174), .o(n18177) );
no02f01 g14389 ( .a(n18177), .b(n18103), .o(n18178) );
in01f01 g14390 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_0_), .o(n4498) );
ao12f01 g14391 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_1_), .b(n17980), .c(n17964), .o(n18180) );
in01f01 g14392 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_1_), .o(n18181) );
no02f01 g14393 ( .a(n17981), .b(n18181), .o(n18182) );
no02f01 g14394 ( .a(n18182), .b(n18180), .o(n18183) );
no02f01 g14395 ( .a(n18183), .b(n18103), .o(n18184) );
na02f01 g14396 ( .a(n18183), .b(n18103), .o(n18185) );
oa12f01 g14397 ( .a(n18185), .b(n18184), .c(n4498), .o(n18186) );
in01f01 g14398 ( .a(n18177), .o(n18187) );
no02f01 g14399 ( .a(n18187), .b(n18145), .o(n18188) );
in01f01 g14400 ( .a(n18188), .o(n18189) );
ao12f01 g14401 ( .a(n18178), .b(n18189), .c(n18186), .o(n18190) );
na02f01 g14402 ( .a(n18172), .b(n18145), .o(n18191) );
in01f01 g14403 ( .a(n18191), .o(n18192) );
no02f01 g14404 ( .a(n18192), .b(n18190), .o(n18193) );
no02f01 g14405 ( .a(n18193), .b(n18173), .o(n18194) );
in01f01 g14406 ( .a(n17989), .o(n18195) );
no02f01 g14407 ( .a(n17968), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_4_), .o(n18196) );
no02f01 g14408 ( .a(n17967), .b(n17990), .o(n18197) );
no02f01 g14409 ( .a(n18197), .b(n18196), .o(n18198) );
no02f01 g14410 ( .a(n18198), .b(n18195), .o(n18199) );
na02f01 g14411 ( .a(n18198), .b(n18195), .o(n18200) );
in01f01 g14412 ( .a(n18200), .o(n18201) );
no02f01 g14413 ( .a(n18201), .b(n18199), .o(n18202) );
in01f01 g14414 ( .a(n18202), .o(n18203) );
no02f01 g14415 ( .a(n18203), .b(n18145), .o(n18204) );
no02f01 g14416 ( .a(n18204), .b(n18194), .o(n18205) );
no02f01 g14417 ( .a(n18202), .b(n18103), .o(n18206) );
no02f01 g14418 ( .a(n18163), .b(n18145), .o(n18207) );
no02f01 g14419 ( .a(n18207), .b(n18206), .o(n18208) );
in01f01 g14420 ( .a(n18208), .o(n18209) );
oa12f01 g14421 ( .a(n18166), .b(n18209), .c(n18205), .o(n18210) );
no02f01 g14422 ( .a(n18001), .b(n17996), .o(n18211) );
in01f01 g14423 ( .a(n18211), .o(n18212) );
no03f01 g14424 ( .a(n18212), .b(n17998), .c(n17994), .o(n18213) );
no02f01 g14425 ( .a(n17998), .b(n17994), .o(n18214) );
no02f01 g14426 ( .a(n18211), .b(n18214), .o(n18215) );
no02f01 g14427 ( .a(n18215), .b(n18213), .o(n18216) );
in01f01 g14428 ( .a(n18216), .o(n18217) );
no02f01 g14429 ( .a(n18217), .b(n18145), .o(n18218) );
ao12f01 g14430 ( .a(n18154), .b(n18216), .c(n18145), .o(n18219) );
in01f01 g14431 ( .a(n18219), .o(n18220) );
oa12f01 g14432 ( .a(n18220), .b(n18218), .c(n18210), .o(n18221) );
ao12f01 g14433 ( .a(n18004), .b(n18007), .c(n18003), .o(n18222) );
in01f01 g14434 ( .a(n18222), .o(n18223) );
no02f01 g14435 ( .a(n17968), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_8_), .o(n18224) );
no02f01 g14436 ( .a(n17967), .b(n17970), .o(n18225) );
no02f01 g14437 ( .a(n18225), .b(n18224), .o(n18226) );
no02f01 g14438 ( .a(n18226), .b(n18223), .o(n18227) );
na02f01 g14439 ( .a(n18226), .b(n18223), .o(n18228) );
in01f01 g14440 ( .a(n18228), .o(n18229) );
no02f01 g14441 ( .a(n18229), .b(n18227), .o(n18230) );
in01f01 g14442 ( .a(n18230), .o(n18231) );
no02f01 g14443 ( .a(n18231), .b(n18145), .o(n18232) );
in01f01 g14444 ( .a(n18012), .o(n18233) );
in01f01 g14445 ( .a(n18018), .o(n18234) );
no02f01 g14446 ( .a(n18234), .b(n18014), .o(n18235) );
no02f01 g14447 ( .a(n18235), .b(n18233), .o(n18236) );
na02f01 g14448 ( .a(n18235), .b(n18233), .o(n18237) );
in01f01 g14449 ( .a(n18237), .o(n18238) );
no02f01 g14450 ( .a(n18238), .b(n18236), .o(n18239) );
in01f01 g14451 ( .a(n18239), .o(n18240) );
no02f01 g14452 ( .a(n18240), .b(n18145), .o(n18241) );
no02f01 g14453 ( .a(n18241), .b(n18232), .o(n18242) );
in01f01 g14454 ( .a(n18013), .o(n18243) );
no02f01 g14455 ( .a(n18014), .b(n18233), .o(n18244) );
ao12f01 g14456 ( .a(n18019), .b(n18244), .c(n18243), .o(n18245) );
in01f01 g14457 ( .a(n18245), .o(n18246) );
no02f01 g14458 ( .a(n17972), .b(n18021), .o(n18247) );
no02f01 g14459 ( .a(n18025), .b(n18247), .o(n18248) );
in01f01 g14460 ( .a(n18248), .o(n18249) );
no02f01 g14461 ( .a(n18249), .b(n18246), .o(n18250) );
no02f01 g14462 ( .a(n18248), .b(n18245), .o(n18251) );
no02f01 g14463 ( .a(n18251), .b(n18250), .o(n18252) );
in01f01 g14464 ( .a(n18252), .o(n18253) );
no02f01 g14465 ( .a(n18253), .b(n18145), .o(n18254) );
no02f01 g14466 ( .a(n18244), .b(n18234), .o(n18255) );
in01f01 g14467 ( .a(n18255), .o(n18256) );
na02f01 g14468 ( .a(n18017), .b(n18243), .o(n18257) );
no02f01 g14469 ( .a(n18257), .b(n18256), .o(n18258) );
na02f01 g14470 ( .a(n18257), .b(n18256), .o(n18259) );
in01f01 g14471 ( .a(n18259), .o(n18260) );
no02f01 g14472 ( .a(n18260), .b(n18258), .o(n18261) );
in01f01 g14473 ( .a(n18261), .o(n18262) );
no02f01 g14474 ( .a(n18262), .b(n18145), .o(n18263) );
no02f01 g14475 ( .a(n18263), .b(n18254), .o(n18264) );
na04f01 g14476 ( .a(n18264), .b(n18242), .c(n18221), .d(n18157), .o(n18265) );
no02f01 g14477 ( .a(n17972), .b(n18033), .o(n18266) );
no02f01 g14478 ( .a(n17973), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_13_), .o(n18267) );
no02f01 g14479 ( .a(n18267), .b(n18266), .o(n18268) );
in01f01 g14480 ( .a(n18268), .o(n18269) );
no02f01 g14481 ( .a(n18269), .b(n18028), .o(n18270) );
in01f01 g14482 ( .a(n18028), .o(n18271) );
no02f01 g14483 ( .a(n18268), .b(n18271), .o(n18272) );
no02f01 g14484 ( .a(n18272), .b(n18270), .o(n18273) );
in01f01 g14485 ( .a(n18273), .o(n18274) );
no02f01 g14486 ( .a(n18274), .b(n18145), .o(n18275) );
no02f01 g14487 ( .a(n18245), .b(n18025), .o(n18276) );
no02f01 g14488 ( .a(n17972), .b(n18020), .o(n18277) );
no02f01 g14489 ( .a(n18277), .b(n18024), .o(n18278) );
in01f01 g14490 ( .a(n18278), .o(n18279) );
no03f01 g14491 ( .a(n18279), .b(n18276), .c(n18247), .o(n18280) );
no02f01 g14492 ( .a(n18276), .b(n18247), .o(n18281) );
no02f01 g14493 ( .a(n18278), .b(n18281), .o(n18282) );
no02f01 g14494 ( .a(n18282), .b(n18280), .o(n18283) );
in01f01 g14495 ( .a(n18283), .o(n18284) );
no02f01 g14496 ( .a(n18284), .b(n18145), .o(n18285) );
no02f01 g14497 ( .a(n18285), .b(n18275), .o(n18286) );
in01f01 g14498 ( .a(n18286), .o(n18287) );
in01f01 g14499 ( .a(n18267), .o(n18288) );
ao12f01 g14500 ( .a(n18266), .b(n18288), .c(n18028), .o(n18289) );
in01f01 g14501 ( .a(n18289), .o(n18290) );
no02f01 g14502 ( .a(n17972), .b(n18032), .o(n18291) );
no02f01 g14503 ( .a(n17973), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_14_), .o(n18292) );
no02f01 g14504 ( .a(n18292), .b(n18291), .o(n18293) );
in01f01 g14505 ( .a(n18293), .o(n18294) );
no02f01 g14506 ( .a(n18294), .b(n18290), .o(n18295) );
no02f01 g14507 ( .a(n18293), .b(n18289), .o(n18296) );
no02f01 g14508 ( .a(n18296), .b(n18295), .o(n18297) );
in01f01 g14509 ( .a(n18297), .o(n18298) );
no02f01 g14510 ( .a(n18298), .b(n18145), .o(n18299) );
no02f01 g14511 ( .a(n18034), .b(n18028), .o(n18300) );
no02f01 g14512 ( .a(n18300), .b(n18038), .o(n18301) );
in01f01 g14513 ( .a(n18301), .o(n18302) );
no02f01 g14514 ( .a(n17972), .b(n18030), .o(n18303) );
no02f01 g14515 ( .a(n18037), .b(n18303), .o(n18304) );
no02f01 g14516 ( .a(n18304), .b(n18302), .o(n18305) );
na02f01 g14517 ( .a(n18304), .b(n18302), .o(n18306) );
in01f01 g14518 ( .a(n18306), .o(n18307) );
no02f01 g14519 ( .a(n18307), .b(n18305), .o(n18308) );
in01f01 g14520 ( .a(n18308), .o(n18309) );
no02f01 g14521 ( .a(n18309), .b(n18145), .o(n18310) );
no02f01 g14522 ( .a(n18310), .b(n18299), .o(n18311) );
in01f01 g14523 ( .a(n18311), .o(n18312) );
no03f01 g14524 ( .a(n18312), .b(n18287), .c(n18265), .o(n18313) );
ao12f01 g14525 ( .a(n18103), .b(n18239), .c(n18230), .o(n18314) );
ao12f01 g14526 ( .a(n18103), .b(n18261), .c(n18252), .o(n18315) );
no02f01 g14527 ( .a(n18315), .b(n18314), .o(n18316) );
in01f01 g14528 ( .a(n18316), .o(n18317) );
ao12f01 g14529 ( .a(n18103), .b(n18283), .c(n18273), .o(n18318) );
no02f01 g14530 ( .a(n18318), .b(n18317), .o(n18319) );
in01f01 g14531 ( .a(n18319), .o(n18320) );
ao12f01 g14532 ( .a(n18103), .b(n18308), .c(n18297), .o(n18321) );
no02f01 g14533 ( .a(n18321), .b(n18320), .o(n18322) );
in01f01 g14534 ( .a(n18322), .o(n18323) );
no02f01 g14535 ( .a(n17972), .b(n18054), .o(n18324) );
no02f01 g14536 ( .a(n18324), .b(n18047), .o(n18325) );
no02f01 g14537 ( .a(n18325), .b(n18043), .o(n18326) );
na02f01 g14538 ( .a(n18325), .b(n18043), .o(n18327) );
in01f01 g14539 ( .a(n18327), .o(n18328) );
no02f01 g14540 ( .a(n18328), .b(n18326), .o(n18329) );
in01f01 g14541 ( .a(n18329), .o(n18330) );
no02f01 g14542 ( .a(n18330), .b(n18145), .o(n18331) );
no02f01 g14543 ( .a(n18040), .b(n18271), .o(n18332) );
no03f01 g14544 ( .a(n18332), .b(n18034), .c(n18303), .o(n18333) );
in01f01 g14545 ( .a(n18333), .o(n18334) );
no02f01 g14546 ( .a(n17972), .b(n18029), .o(n18335) );
no02f01 g14547 ( .a(n18335), .b(n18041), .o(n18336) );
in01f01 g14548 ( .a(n18336), .o(n18337) );
no02f01 g14549 ( .a(n18337), .b(n18334), .o(n18338) );
no02f01 g14550 ( .a(n18336), .b(n18333), .o(n18339) );
no02f01 g14551 ( .a(n18339), .b(n18338), .o(n18340) );
in01f01 g14552 ( .a(n18340), .o(n18341) );
no02f01 g14553 ( .a(n18341), .b(n18145), .o(n18342) );
no02f01 g14554 ( .a(n18342), .b(n18331), .o(n18343) );
in01f01 g14555 ( .a(n18343), .o(n18344) );
no02f01 g14556 ( .a(n18047), .b(n18043), .o(n18345) );
no02f01 g14557 ( .a(n17972), .b(n18053), .o(n18346) );
no02f01 g14558 ( .a(n18346), .b(n18044), .o(n18347) );
in01f01 g14559 ( .a(n18347), .o(n18348) );
no03f01 g14560 ( .a(n18348), .b(n18345), .c(n18324), .o(n18349) );
no02f01 g14561 ( .a(n18345), .b(n18324), .o(n18350) );
no02f01 g14562 ( .a(n18347), .b(n18350), .o(n18351) );
no02f01 g14563 ( .a(n18351), .b(n18349), .o(n18352) );
in01f01 g14564 ( .a(n18352), .o(n18353) );
no02f01 g14565 ( .a(n18353), .b(n18145), .o(n18354) );
no02f01 g14566 ( .a(n18115), .b(n18045), .o(n18355) );
in01f01 g14567 ( .a(n18355), .o(n18356) );
no03f01 g14568 ( .a(n18356), .b(n18116), .c(n18055), .o(n18357) );
no02f01 g14569 ( .a(n18116), .b(n18055), .o(n18358) );
no02f01 g14570 ( .a(n18355), .b(n18358), .o(n18359) );
no02f01 g14571 ( .a(n18359), .b(n18357), .o(n18360) );
in01f01 g14572 ( .a(n18360), .o(n18361) );
no02f01 g14573 ( .a(n18361), .b(n18145), .o(n18362) );
no03f01 g14574 ( .a(n18362), .b(n18354), .c(n18344), .o(n18363) );
oa12f01 g14575 ( .a(n18363), .b(n18323), .c(n18313), .o(n18364) );
ao12f01 g14576 ( .a(n18103), .b(n18340), .c(n18329), .o(n18365) );
ao12f01 g14577 ( .a(n18103), .b(n18360), .c(n18352), .o(n18366) );
no02f01 g14578 ( .a(n18366), .b(n18365), .o(n18367) );
in01f01 g14579 ( .a(n18133), .o(n18368) );
no02f01 g14580 ( .a(n18368), .b(n18145), .o(n18369) );
na02f01 g14581 ( .a(n18126), .b(n18103), .o(n18370) );
in01f01 g14582 ( .a(n18370), .o(n18371) );
no02f01 g14583 ( .a(n18371), .b(n18369), .o(n18372) );
in01f01 g14584 ( .a(n18372), .o(n18373) );
na02f01 g14585 ( .a(n18142), .b(n18103), .o(n18374) );
in01f01 g14586 ( .a(n18374), .o(n18375) );
no03f01 g14587 ( .a(n18375), .b(n18373), .c(n18114), .o(n18376) );
in01f01 g14588 ( .a(n18376), .o(n18377) );
ao12f01 g14589 ( .a(n18377), .b(n18367), .c(n18364), .o(n18378) );
no02f01 g14590 ( .a(n18075), .b(n17969), .o(n18379) );
no02f01 g14591 ( .a(n17967), .b(n18093), .o(n18380) );
no02f01 g14592 ( .a(n18380), .b(n18076), .o(n18381) );
in01f01 g14593 ( .a(n18381), .o(n18382) );
no02f01 g14594 ( .a(n18382), .b(n18379), .o(n18383) );
in01f01 g14595 ( .a(n18379), .o(n18384) );
no02f01 g14596 ( .a(n18381), .b(n18384), .o(n18385) );
no03f01 g14597 ( .a(n18385), .b(n18383), .c(n18103), .o(n18386) );
no03f01 g14598 ( .a(n18062), .b(n18061), .c(n18106), .o(n18387) );
no03f01 g14599 ( .a(n18387), .b(n18070), .c(n18104), .o(n18388) );
no02f01 g14600 ( .a(n18072), .b(n17969), .o(n18389) );
no02f01 g14601 ( .a(n18389), .b(n18388), .o(n18390) );
na02f01 g14602 ( .a(n18389), .b(n18388), .o(n18391) );
in01f01 g14603 ( .a(n18391), .o(n18392) );
no03f01 g14604 ( .a(n18392), .b(n18390), .c(n18103), .o(n18393) );
no02f01 g14605 ( .a(n18393), .b(n18386), .o(n18394) );
in01f01 g14606 ( .a(n18394), .o(n18395) );
no02f01 g14607 ( .a(n18079), .b(n18384), .o(n18396) );
no02f01 g14608 ( .a(n17967), .b(n18090), .o(n18397) );
no02f01 g14609 ( .a(n18397), .b(n18080), .o(n18398) );
in01f01 g14610 ( .a(n18398), .o(n18399) );
no03f01 g14611 ( .a(n18399), .b(n18396), .c(n18094), .o(n18400) );
no02f01 g14612 ( .a(n18396), .b(n18094), .o(n18401) );
no02f01 g14613 ( .a(n18398), .b(n18401), .o(n18402) );
no03f01 g14614 ( .a(n18402), .b(n18400), .c(n18103), .o(n18403) );
in01f01 g14615 ( .a(n18076), .o(n18404) );
ao12f01 g14616 ( .a(n18380), .b(n18404), .c(n18379), .o(n18405) );
in01f01 g14617 ( .a(n18405), .o(n18406) );
no02f01 g14618 ( .a(n17967), .b(n18092), .o(n18407) );
no02f01 g14619 ( .a(n18407), .b(n18077), .o(n18408) );
in01f01 g14620 ( .a(n18408), .o(n18409) );
no02f01 g14621 ( .a(n18409), .b(n18406), .o(n18410) );
no02f01 g14622 ( .a(n18408), .b(n18405), .o(n18411) );
no03f01 g14623 ( .a(n18411), .b(n18410), .c(n18103), .o(n18412) );
no03f01 g14624 ( .a(n18412), .b(n18403), .c(n18395), .o(n18413) );
oa12f01 g14625 ( .a(n18413), .b(n18378), .c(n18149), .o(n18414) );
ao12f01 g14626 ( .a(n18096), .b(n18082), .c(n18379), .o(n18415) );
no02f01 g14627 ( .a(n17967), .b(n18097), .o(n18416) );
no02f01 g14628 ( .a(n18416), .b(n18084), .o(n18417) );
no02f01 g14629 ( .a(n18417), .b(n18415), .o(n18418) );
na02f01 g14630 ( .a(n18417), .b(n18415), .o(n18419) );
in01f01 g14631 ( .a(n18419), .o(n18420) );
no03f01 g14632 ( .a(n18420), .b(n18418), .c(n18103), .o(n18421) );
no03f01 g14633 ( .a(n18080), .b(n18079), .c(n18384), .o(n18422) );
no03f01 g14634 ( .a(n18422), .b(n18094), .c(n18397), .o(n18423) );
in01f01 g14635 ( .a(n18423), .o(n18424) );
no02f01 g14636 ( .a(n17967), .b(n18089), .o(n18425) );
no02f01 g14637 ( .a(n18425), .b(n18081), .o(n18426) );
in01f01 g14638 ( .a(n18426), .o(n18427) );
no02f01 g14639 ( .a(n18427), .b(n18424), .o(n18428) );
no02f01 g14640 ( .a(n18426), .b(n18423), .o(n18429) );
no03f01 g14641 ( .a(n18429), .b(n18428), .c(n18103), .o(n18430) );
no02f01 g14642 ( .a(n18430), .b(n18421), .o(n18431) );
in01f01 g14643 ( .a(n18431), .o(n18432) );
no03f01 g14644 ( .a(n18084), .b(n18083), .c(n18384), .o(n18433) );
no03f01 g14645 ( .a(n18433), .b(n18416), .c(n18096), .o(n18434) );
in01f01 g14646 ( .a(n18434), .o(n18435) );
no02f01 g14647 ( .a(n17967), .b(n18098), .o(n18436) );
no02f01 g14648 ( .a(n18436), .b(n18085), .o(n18437) );
in01f01 g14649 ( .a(n18437), .o(n18438) );
no02f01 g14650 ( .a(n18438), .b(n18435), .o(n18439) );
no02f01 g14651 ( .a(n18437), .b(n18434), .o(n18440) );
no03f01 g14652 ( .a(n18440), .b(n18439), .c(n18103), .o(n18441) );
no02f01 g14653 ( .a(n18441), .b(n18432), .o(n18442) );
in01f01 g14654 ( .a(n18442), .o(n18443) );
no02f01 g14655 ( .a(n18440), .b(n18439), .o(n18444) );
no02f01 g14656 ( .a(n18420), .b(n18418), .o(n18445) );
no02f01 g14657 ( .a(n18429), .b(n18428), .o(n18446) );
ao12f01 g14658 ( .a(n18145), .b(n18446), .c(n18445), .o(n18447) );
in01f01 g14659 ( .a(n18447), .o(n18448) );
ao12f01 g14660 ( .a(n18145), .b(n18448), .c(n18444), .o(n18449) );
no02f01 g14661 ( .a(n18385), .b(n18383), .o(n18450) );
no02f01 g14662 ( .a(n18392), .b(n18390), .o(n18451) );
ao12f01 g14663 ( .a(n18145), .b(n18451), .c(n18450), .o(n18452) );
no02f01 g14664 ( .a(n18402), .b(n18400), .o(n18453) );
no02f01 g14665 ( .a(n18411), .b(n18410), .o(n18454) );
ao12f01 g14666 ( .a(n18145), .b(n18454), .c(n18453), .o(n18455) );
no02f01 g14667 ( .a(n18455), .b(n18452), .o(n18456) );
in01f01 g14668 ( .a(n18456), .o(n18457) );
no02f01 g14669 ( .a(n18457), .b(n18449), .o(n18458) );
oa12f01 g14670 ( .a(n18458), .b(n18443), .c(n18414), .o(n18459) );
in01f01 g14671 ( .a(n18459), .o(n18460) );
in01f01 g14672 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_25_), .o(n18461) );
no02f01 g14673 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .b(n18461), .o(n18462) );
no02f01 g14674 ( .a(n17966), .b(delay_xor_ln21_unr6_stage3_stallmux_q_4_), .o(n18463) );
no02f01 g14675 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_3_), .b(n17966), .o(n18464) );
no02f01 g14676 ( .a(n17966), .b(delay_xor_ln21_unr6_stage3_stallmux_q_2_), .o(n18465) );
in01f01 g14677 ( .a(n18465), .o(n18466) );
no02f01 g14678 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_1_), .b(n17966), .o(n18467) );
no02f01 g14679 ( .a(n17966), .b(delay_xor_ln21_unr6_stage3_stallmux_q_0_), .o(n18468) );
no02f01 g14680 ( .a(n18468), .b(n18467), .o(n18469) );
na02f01 g14681 ( .a(n18469), .b(n18466), .o(n18470) );
no03f01 g14682 ( .a(n18470), .b(n18464), .c(n18463), .o(n18471) );
in01f01 g14683 ( .a(n18471), .o(n18472) );
no02f01 g14684 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_5_), .b(n17966), .o(n18473) );
no02f01 g14685 ( .a(n18473), .b(n18472), .o(n18474) );
no02f01 g14686 ( .a(n17966), .b(delay_xor_ln21_unr6_stage3_stallmux_q_7_), .o(n18475) );
no02f01 g14687 ( .a(n17966), .b(delay_xor_ln21_unr6_stage3_stallmux_q_8_), .o(n18476) );
no02f01 g14688 ( .a(n17966), .b(delay_xor_ln21_unr6_stage3_stallmux_q_6_), .o(n18477) );
no03f01 g14689 ( .a(n18477), .b(n18476), .c(n18475), .o(n18478) );
na02f01 g14690 ( .a(n18478), .b(n18474), .o(n18479) );
no02f01 g14691 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_9_), .b(n17966), .o(n18480) );
no02f01 g14692 ( .a(n18480), .b(n18479), .o(n18481) );
in01f01 g14693 ( .a(n18481), .o(n18482) );
no02f01 g14694 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_10_), .b(n17966), .o(n18483) );
no02f01 g14695 ( .a(n18483), .b(n18482), .o(n18484) );
in01f01 g14696 ( .a(n18484), .o(n18485) );
no02f01 g14697 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_11_), .b(n17966), .o(n18486) );
no02f01 g14698 ( .a(n18486), .b(n18485), .o(n18487) );
in01f01 g14699 ( .a(n18487), .o(n18488) );
no02f01 g14700 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_12_), .b(n17966), .o(n18489) );
no02f01 g14701 ( .a(n18489), .b(n18488), .o(n18490) );
in01f01 g14702 ( .a(n18490), .o(n18491) );
no02f01 g14703 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_13_), .b(n17966), .o(n18492) );
no02f01 g14704 ( .a(n18492), .b(n18491), .o(n18493) );
in01f01 g14705 ( .a(n18493), .o(n18494) );
no02f01 g14706 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_14_), .b(n17966), .o(n18495) );
no02f01 g14707 ( .a(n18495), .b(n18494), .o(n18496) );
in01f01 g14708 ( .a(n18496), .o(n18497) );
no02f01 g14709 ( .a(n17966), .b(delay_xor_ln21_unr6_stage3_stallmux_q_15_), .o(n18498) );
no02f01 g14710 ( .a(n18498), .b(n18497), .o(n18499) );
in01f01 g14711 ( .a(n18499), .o(n18500) );
no02f01 g14712 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_16_), .b(n17966), .o(n18501) );
no02f01 g14713 ( .a(n18501), .b(n18500), .o(n18502) );
in01f01 g14714 ( .a(n18502), .o(n18503) );
no02f01 g14715 ( .a(n17966), .b(delay_xor_ln21_unr6_stage3_stallmux_q_17_), .o(n18504) );
no02f01 g14716 ( .a(n18504), .b(n18503), .o(n18505) );
in01f01 g14717 ( .a(n18505), .o(n18506) );
no02f01 g14718 ( .a(n17966), .b(delay_xor_ln21_unr6_stage3_stallmux_q_18_), .o(n18507) );
no02f01 g14719 ( .a(n18507), .b(n18506), .o(n18508) );
in01f01 g14720 ( .a(n18508), .o(n18509) );
no02f01 g14721 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_19_), .b(n17966), .o(n18510) );
no02f01 g14722 ( .a(n18510), .b(n18509), .o(n18511) );
in01f01 g14723 ( .a(n18511), .o(n18512) );
no02f01 g14724 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_20_), .b(n17966), .o(n18513) );
no02f01 g14725 ( .a(n18513), .b(n18512), .o(n18514) );
in01f01 g14726 ( .a(n18514), .o(n18515) );
no02f01 g14727 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_21_), .b(n17966), .o(n18516) );
no02f01 g14728 ( .a(n18516), .b(n18515), .o(n18517) );
in01f01 g14729 ( .a(n18517), .o(n18518) );
no02f01 g14730 ( .a(n17966), .b(delay_xor_ln21_unr6_stage3_stallmux_q_22_), .o(n18519) );
no02f01 g14731 ( .a(n18519), .b(n18518), .o(n18520) );
in01f01 g14732 ( .a(n18520), .o(n18521) );
no02f01 g14733 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_23_), .b(n17966), .o(n18522) );
no02f01 g14734 ( .a(n18522), .b(n18521), .o(n18523) );
in01f01 g14735 ( .a(n18523), .o(n18524) );
no02f01 g14736 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_24_), .b(n17966), .o(n18525) );
no02f01 g14737 ( .a(n18525), .b(n18524), .o(n18526) );
no02f01 g14738 ( .a(n17966), .b(delay_xor_ln21_unr6_stage3_stallmux_q_25_), .o(n18527) );
no02f01 g14739 ( .a(n18527), .b(n18462), .o(n18528) );
in01f01 g14740 ( .a(n18528), .o(n18529) );
no02f01 g14741 ( .a(n18529), .b(n18526), .o(n18530) );
no02f01 g14742 ( .a(n18530), .b(n18462), .o(n18531) );
in01f01 g14743 ( .a(n18531), .o(n18532) );
na02f01 g14744 ( .a(n18529), .b(n18526), .o(n18533) );
in01f01 g14745 ( .a(n18533), .o(n18534) );
no02f01 g14746 ( .a(n18534), .b(n18530), .o(n18535) );
no02f01 g14747 ( .a(n18535), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_25_), .o(n18536) );
in01f01 g14748 ( .a(n18536), .o(n18537) );
in01f01 g14749 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_24_), .o(n18538) );
na02f01 g14750 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_24_), .b(n17966), .o(n18539) );
in01f01 g14751 ( .a(n18539), .o(n18540) );
no02f01 g14752 ( .a(n18540), .b(n18525), .o(n18541) );
no02f01 g14753 ( .a(n18541), .b(n18524), .o(n18542) );
na02f01 g14754 ( .a(n18541), .b(n18524), .o(n18543) );
in01f01 g14755 ( .a(n18543), .o(n18544) );
no02f01 g14756 ( .a(n18544), .b(n18542), .o(n18545) );
in01f01 g14757 ( .a(n18545), .o(n18546) );
no02f01 g14758 ( .a(n18546), .b(n18538), .o(n18547) );
in01f01 g14759 ( .a(n18547), .o(n18548) );
in01f01 g14760 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_23_), .o(n18549) );
na02f01 g14761 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_23_), .b(n17966), .o(n18550) );
in01f01 g14762 ( .a(n18550), .o(n18551) );
no02f01 g14763 ( .a(n18551), .b(n18522), .o(n18552) );
no02f01 g14764 ( .a(n18552), .b(n18521), .o(n18553) );
in01f01 g14765 ( .a(n18553), .o(n18554) );
na02f01 g14766 ( .a(n18552), .b(n18521), .o(n18555) );
na02f01 g14767 ( .a(n18555), .b(n18554), .o(n18556) );
no02f01 g14768 ( .a(n18556), .b(n18549), .o(n18557) );
ao12f01 g14769 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_23_), .b(n18555), .c(n18554), .o(n18558) );
na02f01 g14770 ( .a(n17966), .b(delay_xor_ln21_unr6_stage3_stallmux_q_22_), .o(n18559) );
in01f01 g14771 ( .a(n18559), .o(n18560) );
no02f01 g14772 ( .a(n18560), .b(n18519), .o(n18561) );
no02f01 g14773 ( .a(n18561), .b(n18518), .o(n18562) );
na02f01 g14774 ( .a(n18561), .b(n18518), .o(n18563) );
in01f01 g14775 ( .a(n18563), .o(n18564) );
no02f01 g14776 ( .a(n18564), .b(n18562), .o(n18565) );
no02f01 g14777 ( .a(n18565), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_22_), .o(n18566) );
in01f01 g14778 ( .a(n18566), .o(n18567) );
na02f01 g14779 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_21_), .b(n17966), .o(n18568) );
in01f01 g14780 ( .a(n18568), .o(n18569) );
no02f01 g14781 ( .a(n18569), .b(n18516), .o(n18570) );
no02f01 g14782 ( .a(n18570), .b(n18515), .o(n18571) );
na02f01 g14783 ( .a(n18570), .b(n18515), .o(n18572) );
in01f01 g14784 ( .a(n18572), .o(n18573) );
no02f01 g14785 ( .a(n18573), .b(n18571), .o(n18574) );
na02f01 g14786 ( .a(n18574), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_21_), .o(n18575) );
in01f01 g14787 ( .a(n18575), .o(n18576) );
in01f01 g14788 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_20_), .o(n18577) );
na02f01 g14789 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_20_), .b(n17966), .o(n18578) );
in01f01 g14790 ( .a(n18578), .o(n18579) );
no02f01 g14791 ( .a(n18579), .b(n18513), .o(n18580) );
in01f01 g14792 ( .a(n18580), .o(n18581) );
no02f01 g14793 ( .a(n18581), .b(n18511), .o(n18582) );
no02f01 g14794 ( .a(n18580), .b(n18512), .o(n18583) );
no02f01 g14795 ( .a(n18583), .b(n18582), .o(n18584) );
in01f01 g14796 ( .a(n18584), .o(n18585) );
no02f01 g14797 ( .a(n18585), .b(n18577), .o(n18586) );
in01f01 g14798 ( .a(n18586), .o(n18587) );
in01f01 g14799 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_19_), .o(n18588) );
na02f01 g14800 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_19_), .b(n17966), .o(n18589) );
in01f01 g14801 ( .a(n18589), .o(n18590) );
no02f01 g14802 ( .a(n18590), .b(n18510), .o(n18591) );
no02f01 g14803 ( .a(n18591), .b(n18509), .o(n18592) );
na02f01 g14804 ( .a(n18591), .b(n18509), .o(n18593) );
in01f01 g14805 ( .a(n18593), .o(n18594) );
no02f01 g14806 ( .a(n18594), .b(n18592), .o(n18595) );
in01f01 g14807 ( .a(n18595), .o(n18596) );
no02f01 g14808 ( .a(n18596), .b(n18588), .o(n18597) );
in01f01 g14809 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_18_), .o(n18598) );
na02f01 g14810 ( .a(n17966), .b(delay_xor_ln21_unr6_stage3_stallmux_q_18_), .o(n18599) );
in01f01 g14811 ( .a(n18599), .o(n18600) );
no02f01 g14812 ( .a(n18600), .b(n18507), .o(n18601) );
in01f01 g14813 ( .a(n18601), .o(n18602) );
no02f01 g14814 ( .a(n18602), .b(n18505), .o(n18603) );
no02f01 g14815 ( .a(n18601), .b(n18506), .o(n18604) );
no02f01 g14816 ( .a(n18604), .b(n18603), .o(n18605) );
in01f01 g14817 ( .a(n18605), .o(n18606) );
no02f01 g14818 ( .a(n18606), .b(n18598), .o(n18607) );
in01f01 g14819 ( .a(n18607), .o(n18608) );
in01f01 g14820 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_17_), .o(n18609) );
na02f01 g14821 ( .a(n17966), .b(delay_xor_ln21_unr6_stage3_stallmux_q_17_), .o(n18610) );
in01f01 g14822 ( .a(n18610), .o(n18611) );
no02f01 g14823 ( .a(n18611), .b(n18504), .o(n18612) );
in01f01 g14824 ( .a(n18612), .o(n18613) );
no02f01 g14825 ( .a(n18613), .b(n18502), .o(n18614) );
no02f01 g14826 ( .a(n18612), .b(n18503), .o(n18615) );
no02f01 g14827 ( .a(n18615), .b(n18614), .o(n18616) );
in01f01 g14828 ( .a(n18616), .o(n18617) );
no02f01 g14829 ( .a(n18617), .b(n18609), .o(n18618) );
in01f01 g14830 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_16_), .o(n18619) );
na02f01 g14831 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_16_), .b(n17966), .o(n18620) );
in01f01 g14832 ( .a(n18620), .o(n18621) );
no02f01 g14833 ( .a(n18621), .b(n18501), .o(n18622) );
in01f01 g14834 ( .a(n18622), .o(n18623) );
no02f01 g14835 ( .a(n18623), .b(n18499), .o(n18624) );
no02f01 g14836 ( .a(n18622), .b(n18500), .o(n18625) );
no02f01 g14837 ( .a(n18625), .b(n18624), .o(n18626) );
in01f01 g14838 ( .a(n18626), .o(n18627) );
no02f01 g14839 ( .a(n18627), .b(n18619), .o(n18628) );
in01f01 g14840 ( .a(n18628), .o(n18629) );
in01f01 g14841 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_15_), .o(n18630) );
na02f01 g14842 ( .a(n17966), .b(delay_xor_ln21_unr6_stage3_stallmux_q_15_), .o(n18631) );
in01f01 g14843 ( .a(n18631), .o(n18632) );
no02f01 g14844 ( .a(n18632), .b(n18498), .o(n18633) );
no02f01 g14845 ( .a(n18633), .b(n18497), .o(n18634) );
na02f01 g14846 ( .a(n18633), .b(n18497), .o(n18635) );
in01f01 g14847 ( .a(n18635), .o(n18636) );
no02f01 g14848 ( .a(n18636), .b(n18634), .o(n18637) );
in01f01 g14849 ( .a(n18637), .o(n18638) );
no02f01 g14850 ( .a(n18638), .b(n18630), .o(n18639) );
in01f01 g14851 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_14_), .o(n18640) );
na02f01 g14852 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_14_), .b(n17966), .o(n18641) );
in01f01 g14853 ( .a(n18641), .o(n18642) );
no02f01 g14854 ( .a(n18642), .b(n18495), .o(n18643) );
no02f01 g14855 ( .a(n18643), .b(n18494), .o(n18644) );
na02f01 g14856 ( .a(n18643), .b(n18494), .o(n18645) );
in01f01 g14857 ( .a(n18645), .o(n18646) );
no02f01 g14858 ( .a(n18646), .b(n18644), .o(n18647) );
in01f01 g14859 ( .a(n18647), .o(n18648) );
no02f01 g14860 ( .a(n18648), .b(n18640), .o(n18649) );
in01f01 g14861 ( .a(n18649), .o(n18650) );
in01f01 g14862 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_13_), .o(n18651) );
na02f01 g14863 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_13_), .b(n17966), .o(n18652) );
in01f01 g14864 ( .a(n18652), .o(n18653) );
no02f01 g14865 ( .a(n18653), .b(n18492), .o(n18654) );
no02f01 g14866 ( .a(n18654), .b(n18491), .o(n18655) );
na02f01 g14867 ( .a(n18654), .b(n18491), .o(n18656) );
in01f01 g14868 ( .a(n18656), .o(n18657) );
no02f01 g14869 ( .a(n18657), .b(n18655), .o(n18658) );
in01f01 g14870 ( .a(n18658), .o(n18659) );
no02f01 g14871 ( .a(n18659), .b(n18651), .o(n18660) );
na02f01 g14872 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_12_), .b(n17966), .o(n18661) );
in01f01 g14873 ( .a(n18661), .o(n18662) );
no02f01 g14874 ( .a(n18662), .b(n18489), .o(n18663) );
no02f01 g14875 ( .a(n18663), .b(n18488), .o(n18664) );
na02f01 g14876 ( .a(n18663), .b(n18488), .o(n18665) );
in01f01 g14877 ( .a(n18665), .o(n18666) );
no02f01 g14878 ( .a(n18666), .b(n18664), .o(n18667) );
no02f01 g14879 ( .a(n18667), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_12_), .o(n18668) );
in01f01 g14880 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_11_), .o(n18669) );
na02f01 g14881 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_11_), .b(n17966), .o(n18670) );
in01f01 g14882 ( .a(n18670), .o(n18671) );
no02f01 g14883 ( .a(n18671), .b(n18486), .o(n18672) );
no02f01 g14884 ( .a(n18672), .b(n18485), .o(n18673) );
na02f01 g14885 ( .a(n18672), .b(n18485), .o(n18674) );
in01f01 g14886 ( .a(n18674), .o(n18675) );
no03f01 g14887 ( .a(n18675), .b(n18673), .c(n18669), .o(n18676) );
in01f01 g14888 ( .a(n18673), .o(n18677) );
ao12f01 g14889 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_11_), .b(n18674), .c(n18677), .o(n18678) );
in01f01 g14890 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_10_), .o(n18679) );
na02f01 g14891 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_10_), .b(n17966), .o(n18680) );
in01f01 g14892 ( .a(n18680), .o(n18681) );
no02f01 g14893 ( .a(n18681), .b(n18483), .o(n18682) );
no02f01 g14894 ( .a(n18682), .b(n18482), .o(n18683) );
na02f01 g14895 ( .a(n18682), .b(n18482), .o(n18684) );
in01f01 g14896 ( .a(n18684), .o(n18685) );
no02f01 g14897 ( .a(n18685), .b(n18683), .o(n18686) );
in01f01 g14898 ( .a(n18686), .o(n18687) );
no02f01 g14899 ( .a(n18687), .b(n18679), .o(n18688) );
in01f01 g14900 ( .a(n18688), .o(n18689) );
no02f01 g14901 ( .a(n18686), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_10_), .o(n18690) );
in01f01 g14902 ( .a(n18690), .o(n18691) );
in01f01 g14903 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_9_), .o(n18692) );
na02f01 g14904 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_9_), .b(n17966), .o(n18693) );
in01f01 g14905 ( .a(n18693), .o(n18694) );
no02f01 g14906 ( .a(n18694), .b(n18480), .o(n18695) );
no02f01 g14907 ( .a(n18695), .b(n18479), .o(n18696) );
na02f01 g14908 ( .a(n18695), .b(n18479), .o(n18697) );
in01f01 g14909 ( .a(n18697), .o(n18698) );
no03f01 g14910 ( .a(n18698), .b(n18696), .c(n18692), .o(n18699) );
in01f01 g14911 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_4_), .o(n18700) );
no02f01 g14912 ( .a(n18470), .b(n18464), .o(n18701) );
na02f01 g14913 ( .a(n17966), .b(delay_xor_ln21_unr6_stage3_stallmux_q_4_), .o(n18702) );
in01f01 g14914 ( .a(n18702), .o(n18703) );
no02f01 g14915 ( .a(n18703), .b(n18463), .o(n18704) );
in01f01 g14916 ( .a(n18704), .o(n18705) );
no02f01 g14917 ( .a(n18705), .b(n18701), .o(n18706) );
in01f01 g14918 ( .a(n18706), .o(n18707) );
na02f01 g14919 ( .a(n18705), .b(n18701), .o(n18708) );
na02f01 g14920 ( .a(n18708), .b(n18707), .o(n18709) );
no02f01 g14921 ( .a(n18709), .b(n18700), .o(n18710) );
in01f01 g14922 ( .a(n18710), .o(n18711) );
in01f01 g14923 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_3_), .o(n18712) );
na02f01 g14924 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_3_), .b(n17966), .o(n18713) );
in01f01 g14925 ( .a(n18713), .o(n18714) );
no02f01 g14926 ( .a(n18714), .b(n18464), .o(n18715) );
in01f01 g14927 ( .a(n18715), .o(n18716) );
na03f01 g14928 ( .a(n18716), .b(n18469), .c(n18466), .o(n18717) );
na02f01 g14929 ( .a(n18715), .b(n18470), .o(n18718) );
na02f01 g14930 ( .a(n18718), .b(n18717), .o(n18719) );
no02f01 g14931 ( .a(n18719), .b(n18712), .o(n18720) );
na02f01 g14932 ( .a(n17966), .b(delay_xor_ln21_unr6_stage3_stallmux_q_2_), .o(n18721) );
na02f01 g14933 ( .a(n18721), .b(n18466), .o(n18722) );
no02f01 g14934 ( .a(n18722), .b(n18469), .o(n18723) );
in01f01 g14935 ( .a(n18469), .o(n18724) );
ao12f01 g14936 ( .a(n18724), .b(n18721), .c(n18466), .o(n18725) );
no02f01 g14937 ( .a(n18725), .b(n18723), .o(n18726) );
na02f01 g14938 ( .a(n18726), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_2_), .o(n18727) );
no02f01 g14939 ( .a(n18726), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_2_), .o(n18728) );
in01f01 g14940 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_1_), .o(n18729) );
no02f01 g14941 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .b(delay_xor_ln21_unr6_stage3_stallmux_q_0_), .o(n18730) );
in01f01 g14942 ( .a(n18730), .o(n18731) );
na02f01 g14943 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .b(delay_xor_ln21_unr6_stage3_stallmux_q_0_), .o(n18732) );
na02f01 g14944 ( .a(n18732), .b(n18731), .o(n18733) );
no02f01 g14945 ( .a(n18733), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_0_), .o(n18734) );
no02f01 g14946 ( .a(n18734), .b(n18729), .o(n18735) );
na02f01 g14947 ( .a(n18734), .b(n18729), .o(n18736) );
in01f01 g14948 ( .a(n18468), .o(n18737) );
in01f01 g14949 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_1_), .o(n18738) );
na02f01 g14950 ( .a(n18738), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(n18739) );
na02f01 g14951 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_1_), .b(n17966), .o(n18740) );
na02f01 g14952 ( .a(n18740), .b(n18739), .o(n18741) );
no02f01 g14953 ( .a(n18741), .b(n18737), .o(n18742) );
ao12f01 g14954 ( .a(n18468), .b(n18740), .c(n18739), .o(n18743) );
no02f01 g14955 ( .a(n18743), .b(n18742), .o(n18744) );
ao12f01 g14956 ( .a(n18735), .b(n18744), .c(n18736), .o(n18745) );
oa12f01 g14957 ( .a(n18727), .b(n18745), .c(n18728), .o(n18746) );
ao12f01 g14958 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_3_), .b(n18718), .c(n18717), .o(n18747) );
in01f01 g14959 ( .a(n18747), .o(n18748) );
ao12f01 g14960 ( .a(n18720), .b(n18748), .c(n18746), .o(n18749) );
ao12f01 g14961 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_4_), .b(n18708), .c(n18707), .o(n18750) );
oa12f01 g14962 ( .a(n18711), .b(n18750), .c(n18749), .o(n18751) );
in01f01 g14963 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_5_), .o(n18752) );
na02f01 g14964 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_5_), .b(n17966), .o(n18753) );
in01f01 g14965 ( .a(n18753), .o(n18754) );
no02f01 g14966 ( .a(n18754), .b(n18473), .o(n18755) );
no02f01 g14967 ( .a(n18755), .b(n18472), .o(n18756) );
in01f01 g14968 ( .a(n18756), .o(n18757) );
na02f01 g14969 ( .a(n18755), .b(n18472), .o(n18758) );
na02f01 g14970 ( .a(n18758), .b(n18757), .o(n18759) );
na02f01 g14971 ( .a(n18759), .b(n18752), .o(n18760) );
no02f01 g14972 ( .a(n18759), .b(n18752), .o(n18761) );
ao12f01 g14973 ( .a(n18761), .b(n18760), .c(n18751), .o(n18762) );
in01f01 g14974 ( .a(n18477), .o(n18763) );
na02f01 g14975 ( .a(n17966), .b(delay_xor_ln21_unr6_stage3_stallmux_q_6_), .o(n18764) );
na02f01 g14976 ( .a(n18764), .b(n18763), .o(n18765) );
no02f01 g14977 ( .a(n18765), .b(n18474), .o(n18766) );
na02f01 g14978 ( .a(n18765), .b(n18474), .o(n18767) );
in01f01 g14979 ( .a(n18767), .o(n18768) );
no02f01 g14980 ( .a(n18768), .b(n18766), .o(n18769) );
no02f01 g14981 ( .a(n18769), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_6_), .o(n18770) );
no02f01 g14982 ( .a(n18770), .b(n18762), .o(n18771) );
na02f01 g14983 ( .a(n18769), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_6_), .o(n18772) );
in01f01 g14984 ( .a(n18772), .o(n18773) );
no02f01 g14985 ( .a(n18773), .b(n18771), .o(n18774) );
in01f01 g14986 ( .a(n18475), .o(n18775) );
na02f01 g14987 ( .a(n17966), .b(delay_xor_ln21_unr6_stage3_stallmux_q_7_), .o(n18776) );
na02f01 g14988 ( .a(n18776), .b(n18775), .o(n18777) );
in01f01 g14989 ( .a(n18777), .o(n18778) );
na02f01 g14990 ( .a(n18763), .b(n18474), .o(n18779) );
no02f01 g14991 ( .a(n18779), .b(n18778), .o(n18780) );
ao12f01 g14992 ( .a(n18777), .b(n18763), .c(n18474), .o(n18781) );
no02f01 g14993 ( .a(n18781), .b(n18780), .o(n18782) );
no02f01 g14994 ( .a(n18782), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_7_), .o(n18783) );
no02f01 g14995 ( .a(n18783), .b(n18774), .o(n18784) );
na02f01 g14996 ( .a(n18782), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_7_), .o(n18785) );
in01f01 g14997 ( .a(n18785), .o(n18786) );
no02f01 g14998 ( .a(n18786), .b(n18784), .o(n18787) );
na02f01 g14999 ( .a(n17966), .b(delay_xor_ln21_unr6_stage3_stallmux_q_8_), .o(n18788) );
in01f01 g15000 ( .a(n18788), .o(n18789) );
no02f01 g15001 ( .a(n18789), .b(n18476), .o(n18790) );
in01f01 g15002 ( .a(n18790), .o(n18791) );
no02f01 g15003 ( .a(n18779), .b(n18475), .o(n18792) );
no02f01 g15004 ( .a(n18792), .b(n18791), .o(n18793) );
na02f01 g15005 ( .a(n18792), .b(n18791), .o(n18794) );
in01f01 g15006 ( .a(n18794), .o(n18795) );
no02f01 g15007 ( .a(n18795), .b(n18793), .o(n18796) );
no02f01 g15008 ( .a(n18796), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_8_), .o(n18797) );
no02f01 g15009 ( .a(n18797), .b(n18787), .o(n18798) );
na02f01 g15010 ( .a(n18796), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_8_), .o(n18799) );
in01f01 g15011 ( .a(n18799), .o(n18800) );
no02f01 g15012 ( .a(n18800), .b(n18798), .o(n18801) );
in01f01 g15013 ( .a(n18696), .o(n18802) );
ao12f01 g15014 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_9_), .b(n18697), .c(n18802), .o(n18803) );
no02f01 g15015 ( .a(n18803), .b(n18801), .o(n18804) );
oa12f01 g15016 ( .a(n18691), .b(n18804), .c(n18699), .o(n18805) );
ao12f01 g15017 ( .a(n18678), .b(n18805), .c(n18689), .o(n18806) );
na02f01 g15018 ( .a(n18667), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_12_), .o(n18807) );
in01f01 g15019 ( .a(n18807), .o(n18808) );
no03f01 g15020 ( .a(n18808), .b(n18806), .c(n18676), .o(n18809) );
no02f01 g15021 ( .a(n18658), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_13_), .o(n18810) );
no03f01 g15022 ( .a(n18810), .b(n18809), .c(n18668), .o(n18811) );
no02f01 g15023 ( .a(n18647), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_14_), .o(n18812) );
in01f01 g15024 ( .a(n18812), .o(n18813) );
oa12f01 g15025 ( .a(n18813), .b(n18811), .c(n18660), .o(n18814) );
no02f01 g15026 ( .a(n18637), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_15_), .o(n18815) );
ao12f01 g15027 ( .a(n18815), .b(n18814), .c(n18650), .o(n18816) );
no02f01 g15028 ( .a(n18626), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_16_), .o(n18817) );
in01f01 g15029 ( .a(n18817), .o(n18818) );
oa12f01 g15030 ( .a(n18818), .b(n18816), .c(n18639), .o(n18819) );
no02f01 g15031 ( .a(n18616), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_17_), .o(n18820) );
ao12f01 g15032 ( .a(n18820), .b(n18819), .c(n18629), .o(n18821) );
no02f01 g15033 ( .a(n18605), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_18_), .o(n18822) );
in01f01 g15034 ( .a(n18822), .o(n18823) );
oa12f01 g15035 ( .a(n18823), .b(n18821), .c(n18618), .o(n18824) );
no02f01 g15036 ( .a(n18595), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_19_), .o(n18825) );
ao12f01 g15037 ( .a(n18825), .b(n18824), .c(n18608), .o(n18826) );
no02f01 g15038 ( .a(n18584), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_20_), .o(n18827) );
in01f01 g15039 ( .a(n18827), .o(n18828) );
oa12f01 g15040 ( .a(n18828), .b(n18826), .c(n18597), .o(n18829) );
no02f01 g15041 ( .a(n18574), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_21_), .o(n18830) );
ao12f01 g15042 ( .a(n18830), .b(n18829), .c(n18587), .o(n18831) );
oa12f01 g15043 ( .a(n18567), .b(n18831), .c(n18576), .o(n18832) );
na02f01 g15044 ( .a(n18565), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_22_), .o(n18833) );
ao12f01 g15045 ( .a(n18558), .b(n18833), .c(n18832), .o(n18834) );
no02f01 g15046 ( .a(n18545), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_24_), .o(n18835) );
in01f01 g15047 ( .a(n18835), .o(n18836) );
oa12f01 g15048 ( .a(n18836), .b(n18834), .c(n18557), .o(n18837) );
in01f01 g15049 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_25_), .o(n18838) );
no03f01 g15050 ( .a(n18534), .b(n18530), .c(n18838), .o(n18839) );
in01f01 g15051 ( .a(n18839), .o(n18840) );
na03f01 g15052 ( .a(n18840), .b(n18837), .c(n18548), .o(n18841) );
in01f01 g15053 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_26_), .o(n18842) );
no02f01 g15054 ( .a(n18532), .b(n18842), .o(n18843) );
ao12f01 g15055 ( .a(n18843), .b(n18841), .c(n18537), .o(n18844) );
in01f01 g15056 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_27_), .o(n18845) );
no02f01 g15057 ( .a(n18531), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_26_), .o(n18846) );
no02f01 g15058 ( .a(n18846), .b(n18845), .o(n18847) );
in01f01 g15059 ( .a(n18847), .o(n18848) );
ao12f01 g15060 ( .a(n18532), .b(n18848), .c(n18844), .o(n18849) );
na02f01 g15061 ( .a(n18841), .b(n18537), .o(n18850) );
no02f01 g15062 ( .a(n18848), .b(n18850), .o(n18851) );
no02f01 g15063 ( .a(n18851), .b(n18849), .o(n18852) );
no02f01 g15064 ( .a(n18531), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_30_), .o(n18853) );
ao12f01 g15065 ( .a(n18531), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_29_), .c(delay_sub_ln21_0_unr5_stage3_stallmux_q_28_), .o(n18854) );
no03f01 g15066 ( .a(n18854), .b(n18853), .c(n18852), .o(n18855) );
in01f01 g15067 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_30_), .o(n18856) );
no02f01 g15068 ( .a(n18532), .b(n18856), .o(n18857) );
no02f01 g15069 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_29_), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_28_), .o(n18858) );
no02f01 g15070 ( .a(n18858), .b(n18532), .o(n18859) );
no03f01 g15071 ( .a(n18859), .b(n18857), .c(n18855), .o(n18860) );
in01f01 g15072 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_31_), .o(n18861) );
no02f01 g15073 ( .a(n18532), .b(n18861), .o(n18862) );
no02f01 g15074 ( .a(n18531), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_31_), .o(n18863) );
no02f01 g15075 ( .a(n18863), .b(n18862), .o(n18864) );
na02f01 g15076 ( .a(n18864), .b(n18860), .o(n18865) );
in01f01 g15077 ( .a(n18865), .o(n18866) );
no02f01 g15078 ( .a(n18864), .b(n18860), .o(n18867) );
no02f01 g15079 ( .a(n18867), .b(n18866), .o(n18868) );
in01f01 g15080 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_29_), .o(n18869) );
no02f01 g15081 ( .a(n18532), .b(n18869), .o(n18870) );
no02f01 g15082 ( .a(n18531), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_29_), .o(n18871) );
no02f01 g15083 ( .a(n18871), .b(n18870), .o(n18872) );
in01f01 g15084 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_28_), .o(n18873) );
no02f01 g15085 ( .a(n18532), .b(n18873), .o(n18874) );
in01f01 g15086 ( .a(n18874), .o(n18875) );
no02f01 g15087 ( .a(n18531), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_28_), .o(n18876) );
in01f01 g15088 ( .a(n18876), .o(n18877) );
oa12f01 g15089 ( .a(n18877), .b(n18851), .c(n18849), .o(n18878) );
na03f01 g15090 ( .a(n18878), .b(n18875), .c(n18872), .o(n18879) );
in01f01 g15091 ( .a(n18879), .o(n18880) );
ao12f01 g15092 ( .a(n18872), .b(n18878), .c(n18875), .o(n18881) );
no02f01 g15093 ( .a(n18881), .b(n18880), .o(n18882) );
no02f01 g15094 ( .a(n18882), .b(n18103), .o(n18883) );
in01f01 g15095 ( .a(n18854), .o(n18884) );
no02f01 g15096 ( .a(n18857), .b(n18853), .o(n18885) );
in01f01 g15097 ( .a(n18885), .o(n18886) );
in01f01 g15098 ( .a(n18859), .o(n18887) );
na02f01 g15099 ( .a(n18887), .b(n18852), .o(n18888) );
ao12f01 g15100 ( .a(n18886), .b(n18888), .c(n18884), .o(n18889) );
in01f01 g15101 ( .a(n18850), .o(n18890) );
no03f01 g15102 ( .a(n18847), .b(n18843), .c(n18890), .o(n18891) );
in01f01 g15103 ( .a(n18851), .o(n18892) );
oa12f01 g15104 ( .a(n18892), .b(n18891), .c(n18532), .o(n18893) );
no02f01 g15105 ( .a(n18859), .b(n18893), .o(n18894) );
no03f01 g15106 ( .a(n18894), .b(n18885), .c(n18854), .o(n18895) );
no02f01 g15107 ( .a(n18895), .b(n18889), .o(n18896) );
no02f01 g15108 ( .a(n18896), .b(n18103), .o(n18897) );
no02f01 g15109 ( .a(n18831), .b(n18576), .o(n18898) );
in01f01 g15110 ( .a(n18898), .o(n18899) );
in01f01 g15111 ( .a(n18833), .o(n18900) );
no02f01 g15112 ( .a(n18900), .b(n18566), .o(n18901) );
in01f01 g15113 ( .a(n18901), .o(n18902) );
no02f01 g15114 ( .a(n18902), .b(n18899), .o(n18903) );
no02f01 g15115 ( .a(n18901), .b(n18898), .o(n18904) );
no02f01 g15116 ( .a(n18904), .b(n18903), .o(n18905) );
in01f01 g15117 ( .a(n18905), .o(n18906) );
na02f01 g15118 ( .a(n18906), .b(n18145), .o(n18907) );
no02f01 g15119 ( .a(n18803), .b(n18699), .o(n18908) );
in01f01 g15120 ( .a(n18908), .o(n18909) );
no03f01 g15121 ( .a(n18909), .b(n18800), .c(n18798), .o(n18910) );
no02f01 g15122 ( .a(n18908), .b(n18801), .o(n18911) );
no02f01 g15123 ( .a(n18911), .b(n18910), .o(n18912) );
in01f01 g15124 ( .a(n18912), .o(n18913) );
no02f01 g15125 ( .a(n18786), .b(n18783), .o(n18914) );
no02f01 g15126 ( .a(n18914), .b(n18774), .o(n18915) );
na02f01 g15127 ( .a(n18914), .b(n18774), .o(n18916) );
in01f01 g15128 ( .a(n18916), .o(n18917) );
no02f01 g15129 ( .a(n18917), .b(n18915), .o(n18918) );
in01f01 g15130 ( .a(n18918), .o(n18919) );
no02f01 g15131 ( .a(n18800), .b(n18797), .o(n18920) );
no02f01 g15132 ( .a(n18920), .b(n18787), .o(n18921) );
na02f01 g15133 ( .a(n18920), .b(n18787), .o(n18922) );
in01f01 g15134 ( .a(n18922), .o(n18923) );
no02f01 g15135 ( .a(n18923), .b(n18921), .o(n18924) );
in01f01 g15136 ( .a(n18924), .o(n18925) );
oa12f01 g15137 ( .a(n18145), .b(n18925), .c(n18919), .o(n18926) );
in01f01 g15138 ( .a(n18926), .o(n18927) );
ao12f01 g15139 ( .a(n18927), .b(n18913), .c(n18145), .o(n18928) );
no02f01 g15140 ( .a(n18804), .b(n18699), .o(n18929) );
no02f01 g15141 ( .a(n18690), .b(n18688), .o(n18930) );
no02f01 g15142 ( .a(n18930), .b(n18929), .o(n18931) );
na02f01 g15143 ( .a(n18930), .b(n18929), .o(n18932) );
in01f01 g15144 ( .a(n18932), .o(n18933) );
no02f01 g15145 ( .a(n18933), .b(n18931), .o(n18934) );
in01f01 g15146 ( .a(n18934), .o(n18935) );
na02f01 g15147 ( .a(n18935), .b(n18145), .o(n18936) );
na02f01 g15148 ( .a(n18936), .b(n18928), .o(n18937) );
na02f01 g15149 ( .a(n18805), .b(n18689), .o(n18938) );
no02f01 g15150 ( .a(n18678), .b(n18676), .o(n18939) );
in01f01 g15151 ( .a(n18939), .o(n18940) );
no02f01 g15152 ( .a(n18940), .b(n18938), .o(n18941) );
na02f01 g15153 ( .a(n18940), .b(n18938), .o(n18942) );
in01f01 g15154 ( .a(n18942), .o(n18943) );
no02f01 g15155 ( .a(n18943), .b(n18941), .o(n18944) );
no02f01 g15156 ( .a(n18944), .b(n18103), .o(n18945) );
no02f01 g15157 ( .a(n18945), .b(n18937), .o(n18946) );
no02f01 g15158 ( .a(n18806), .b(n18676), .o(n18947) );
no02f01 g15159 ( .a(n18808), .b(n18668), .o(n18948) );
no02f01 g15160 ( .a(n18948), .b(n18947), .o(n18949) );
na02f01 g15161 ( .a(n18948), .b(n18947), .o(n18950) );
in01f01 g15162 ( .a(n18950), .o(n18951) );
no02f01 g15163 ( .a(n18951), .b(n18949), .o(n18952) );
no02f01 g15164 ( .a(n18952), .b(n18103), .o(n18953) );
in01f01 g15165 ( .a(n18953), .o(n18954) );
na02f01 g15166 ( .a(n18954), .b(n18946), .o(n18955) );
no02f01 g15167 ( .a(n18809), .b(n18668), .o(n18956) );
in01f01 g15168 ( .a(n18956), .o(n18957) );
no02f01 g15169 ( .a(n18810), .b(n18660), .o(n18958) );
no02f01 g15170 ( .a(n18958), .b(n18957), .o(n18959) );
na02f01 g15171 ( .a(n18958), .b(n18957), .o(n18960) );
in01f01 g15172 ( .a(n18960), .o(n18961) );
no02f01 g15173 ( .a(n18961), .b(n18959), .o(n18962) );
in01f01 g15174 ( .a(n18962), .o(n18963) );
ao12f01 g15175 ( .a(n18955), .b(n18963), .c(n18145), .o(n18964) );
no02f01 g15176 ( .a(n18812), .b(n18649), .o(n18965) );
in01f01 g15177 ( .a(n18965), .o(n18966) );
no03f01 g15178 ( .a(n18966), .b(n18811), .c(n18660), .o(n18967) );
no02f01 g15179 ( .a(n18811), .b(n18660), .o(n18968) );
no02f01 g15180 ( .a(n18965), .b(n18968), .o(n18969) );
no02f01 g15181 ( .a(n18969), .b(n18967), .o(n18970) );
ao12f01 g15182 ( .a(n18103), .b(n18970), .c(n18964), .o(n18971) );
na02f01 g15183 ( .a(n18814), .b(n18650), .o(n18972) );
no02f01 g15184 ( .a(n18815), .b(n18639), .o(n18973) );
in01f01 g15185 ( .a(n18973), .o(n18974) );
no02f01 g15186 ( .a(n18974), .b(n18972), .o(n18975) );
na02f01 g15187 ( .a(n18974), .b(n18972), .o(n18976) );
in01f01 g15188 ( .a(n18976), .o(n18977) );
no02f01 g15189 ( .a(n18977), .b(n18975), .o(n18978) );
in01f01 g15190 ( .a(n18978), .o(n18979) );
ao12f01 g15191 ( .a(n18971), .b(n18979), .c(n18145), .o(n18980) );
no02f01 g15192 ( .a(n18817), .b(n18628), .o(n18981) );
in01f01 g15193 ( .a(n18981), .o(n18982) );
no03f01 g15194 ( .a(n18982), .b(n18816), .c(n18639), .o(n18983) );
no02f01 g15195 ( .a(n18816), .b(n18639), .o(n18984) );
no02f01 g15196 ( .a(n18981), .b(n18984), .o(n18985) );
no02f01 g15197 ( .a(n18985), .b(n18983), .o(n18986) );
oa12f01 g15198 ( .a(n18980), .b(n18986), .c(n18103), .o(n18987) );
na02f01 g15199 ( .a(n18819), .b(n18629), .o(n18988) );
in01f01 g15200 ( .a(n18988), .o(n18989) );
no02f01 g15201 ( .a(n18820), .b(n18618), .o(n18990) );
no02f01 g15202 ( .a(n18990), .b(n18989), .o(n18991) );
na02f01 g15203 ( .a(n18990), .b(n18989), .o(n18992) );
in01f01 g15204 ( .a(n18992), .o(n18993) );
no02f01 g15205 ( .a(n18993), .b(n18991), .o(n18994) );
in01f01 g15206 ( .a(n18994), .o(n18995) );
ao12f01 g15207 ( .a(n18987), .b(n18995), .c(n18145), .o(n18996) );
no02f01 g15208 ( .a(n18822), .b(n18607), .o(n18997) );
in01f01 g15209 ( .a(n18997), .o(n18998) );
no03f01 g15210 ( .a(n18998), .b(n18821), .c(n18618), .o(n18999) );
no02f01 g15211 ( .a(n18821), .b(n18618), .o(n19000) );
no02f01 g15212 ( .a(n18997), .b(n19000), .o(n19001) );
no02f01 g15213 ( .a(n19001), .b(n18999), .o(n19002) );
oa12f01 g15214 ( .a(n18996), .b(n19002), .c(n18103), .o(n19003) );
in01f01 g15215 ( .a(n19002), .o(n19004) );
in01f01 g15216 ( .a(n18986), .o(n19005) );
no02f01 g15217 ( .a(n18978), .b(n18145), .o(n19006) );
ao12f01 g15218 ( .a(n19006), .b(n19005), .c(n18103), .o(n19007) );
oa12f01 g15219 ( .a(n19007), .b(n18994), .c(n18145), .o(n19008) );
ao12f01 g15220 ( .a(n19008), .b(n19004), .c(n18103), .o(n19009) );
na02f01 g15221 ( .a(n19009), .b(n19003), .o(n19010) );
in01f01 g15222 ( .a(n19010), .o(n19011) );
no02f01 g15223 ( .a(n18826), .b(n18597), .o(n19012) );
no02f01 g15224 ( .a(n18827), .b(n18586), .o(n19013) );
na02f01 g15225 ( .a(n19013), .b(n19012), .o(n19014) );
no02f01 g15226 ( .a(n19013), .b(n19012), .o(n19015) );
in01f01 g15227 ( .a(n19015), .o(n19016) );
na02f01 g15228 ( .a(n19016), .b(n19014), .o(n19017) );
na02f01 g15229 ( .a(n18824), .b(n18608), .o(n19018) );
no02f01 g15230 ( .a(n18825), .b(n18597), .o(n19019) );
in01f01 g15231 ( .a(n19019), .o(n19020) );
no02f01 g15232 ( .a(n19020), .b(n19018), .o(n19021) );
na02f01 g15233 ( .a(n19020), .b(n19018), .o(n19022) );
in01f01 g15234 ( .a(n19022), .o(n19023) );
no02f01 g15235 ( .a(n19023), .b(n19021), .o(n19024) );
no02f01 g15236 ( .a(n19024), .b(n18103), .o(n19025) );
ao12f01 g15237 ( .a(n19025), .b(n19017), .c(n18145), .o(n19026) );
na02f01 g15238 ( .a(n18829), .b(n18587), .o(n19027) );
no02f01 g15239 ( .a(n18830), .b(n18576), .o(n19028) );
in01f01 g15240 ( .a(n19028), .o(n19029) );
no02f01 g15241 ( .a(n19029), .b(n19027), .o(n19030) );
no02f01 g15242 ( .a(n18827), .b(n19012), .o(n19031) );
no02f01 g15243 ( .a(n19031), .b(n18586), .o(n19032) );
no02f01 g15244 ( .a(n19028), .b(n19032), .o(n19033) );
no02f01 g15245 ( .a(n19033), .b(n19030), .o(n19034) );
oa12f01 g15246 ( .a(n19026), .b(n19034), .c(n18103), .o(n19035) );
no02f01 g15247 ( .a(n19035), .b(n19011), .o(n19036) );
no02f01 g15248 ( .a(n19034), .b(n18145), .o(n19037) );
no02f01 g15249 ( .a(n19024), .b(n18145), .o(n19038) );
ao12f01 g15250 ( .a(n19038), .b(n19017), .c(n18103), .o(n19039) );
in01f01 g15251 ( .a(n19039), .o(n19040) );
no02f01 g15252 ( .a(n19040), .b(n19037), .o(n19041) );
oa12f01 g15253 ( .a(n19041), .b(n18905), .c(n18145), .o(n19042) );
ao12f01 g15254 ( .a(n19042), .b(n19036), .c(n18907), .o(n19043) );
ao12f01 g15255 ( .a(n18566), .b(n18833), .c(n18898), .o(n19044) );
in01f01 g15256 ( .a(n19044), .o(n19045) );
no02f01 g15257 ( .a(n18558), .b(n18557), .o(n19046) );
no02f01 g15258 ( .a(n19046), .b(n19045), .o(n19047) );
na02f01 g15259 ( .a(n19046), .b(n19045), .o(n19048) );
in01f01 g15260 ( .a(n19048), .o(n19049) );
no02f01 g15261 ( .a(n19049), .b(n19047), .o(n19050) );
in01f01 g15262 ( .a(n19050), .o(n19051) );
ao12f01 g15263 ( .a(n19043), .b(n19051), .c(n18145), .o(n19052) );
no02f01 g15264 ( .a(n18834), .b(n18557), .o(n19053) );
in01f01 g15265 ( .a(n19053), .o(n19054) );
no02f01 g15266 ( .a(n18835), .b(n18547), .o(n19055) );
in01f01 g15267 ( .a(n19055), .o(n19056) );
no02f01 g15268 ( .a(n19056), .b(n19054), .o(n19057) );
no02f01 g15269 ( .a(n19055), .b(n19053), .o(n19058) );
no02f01 g15270 ( .a(n19058), .b(n19057), .o(n19059) );
oa12f01 g15271 ( .a(n19052), .b(n19059), .c(n18103), .o(n19060) );
na02f01 g15272 ( .a(n18837), .b(n18548), .o(n19061) );
no02f01 g15273 ( .a(n18839), .b(n18536), .o(n19062) );
in01f01 g15274 ( .a(n19062), .o(n19063) );
no02f01 g15275 ( .a(n19063), .b(n19061), .o(n19064) );
na02f01 g15276 ( .a(n19063), .b(n19061), .o(n19065) );
in01f01 g15277 ( .a(n19065), .o(n19066) );
no02f01 g15278 ( .a(n19066), .b(n19064), .o(n19067) );
in01f01 g15279 ( .a(n19067), .o(n19068) );
ao12f01 g15280 ( .a(n19060), .b(n19068), .c(n18145), .o(n19069) );
no02f01 g15281 ( .a(n18846), .b(n18843), .o(n19070) );
na02f01 g15282 ( .a(n19070), .b(n18850), .o(n19071) );
in01f01 g15283 ( .a(n19071), .o(n19072) );
no02f01 g15284 ( .a(n19070), .b(n18850), .o(n19073) );
no02f01 g15285 ( .a(n19073), .b(n19072), .o(n19074) );
oa12f01 g15286 ( .a(n19069), .b(n19074), .c(n18103), .o(n19075) );
in01f01 g15287 ( .a(n19073), .o(n19076) );
na02f01 g15288 ( .a(n19076), .b(n19071), .o(n19077) );
ao12f01 g15289 ( .a(n18145), .b(n19059), .c(n19050), .o(n19078) );
in01f01 g15290 ( .a(n19078), .o(n19079) );
oa12f01 g15291 ( .a(n19079), .b(n19067), .c(n18145), .o(n19080) );
ao12f01 g15292 ( .a(n19080), .b(n19077), .c(n18103), .o(n19081) );
no02f01 g15293 ( .a(n18532), .b(n18845), .o(n19082) );
no02f01 g15294 ( .a(n18531), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_27_), .o(n19083) );
no02f01 g15295 ( .a(n19083), .b(n19082), .o(n19084) );
in01f01 g15296 ( .a(n19084), .o(n19085) );
no02f01 g15297 ( .a(n18846), .b(n18844), .o(n19086) );
na02f01 g15298 ( .a(n19086), .b(n19085), .o(n19087) );
no02f01 g15299 ( .a(n19086), .b(n19085), .o(n19088) );
in01f01 g15300 ( .a(n19088), .o(n19089) );
na02f01 g15301 ( .a(n19089), .b(n19087), .o(n19090) );
ao22f01 g15302 ( .a(n19090), .b(n18145), .c(n19081), .d(n19075), .o(n19091) );
no02f01 g15303 ( .a(n18876), .b(n18874), .o(n19092) );
no02f01 g15304 ( .a(n19092), .b(n18852), .o(n19093) );
na02f01 g15305 ( .a(n19092), .b(n18852), .o(n19094) );
in01f01 g15306 ( .a(n19094), .o(n19095) );
no02f01 g15307 ( .a(n19095), .b(n19093), .o(n19096) );
oa12f01 g15308 ( .a(n19091), .b(n19096), .c(n18103), .o(n19097) );
no03f01 g15309 ( .a(n19097), .b(n18897), .c(n18883), .o(n19098) );
in01f01 g15310 ( .a(n18872), .o(n19099) );
na02f01 g15311 ( .a(n18878), .b(n18875), .o(n19100) );
na02f01 g15312 ( .a(n19100), .b(n19099), .o(n19101) );
na02f01 g15313 ( .a(n19101), .b(n18879), .o(n19102) );
na02f01 g15314 ( .a(n19102), .b(n18103), .o(n19103) );
oa12f01 g15315 ( .a(n18103), .b(n18895), .c(n18889), .o(n19104) );
in01f01 g15316 ( .a(n19093), .o(n19105) );
na02f01 g15317 ( .a(n19094), .b(n19105), .o(n19106) );
in01f01 g15318 ( .a(n19087), .o(n19107) );
no02f01 g15319 ( .a(n19088), .b(n19107), .o(n19108) );
no02f01 g15320 ( .a(n19108), .b(n18145), .o(n19109) );
ao12f01 g15321 ( .a(n19109), .b(n19106), .c(n18103), .o(n19110) );
na03f01 g15322 ( .a(n19110), .b(n19104), .c(n19103), .o(n19111) );
no02f01 g15323 ( .a(n19111), .b(n19098), .o(n19112) );
no02f01 g15324 ( .a(n18868), .b(n18145), .o(n19113) );
in01f01 g15325 ( .a(n18868), .o(n19114) );
no02f01 g15326 ( .a(n18868), .b(n18145), .o(n19115) );
ao12f01 g15327 ( .a(n19112), .b(n19114), .c(n18145), .o(n19116) );
no03f01 g15328 ( .a(n19116), .b(n19115), .c(n19114), .o(n19117) );
no02f01 g15329 ( .a(n19117), .b(n19113), .o(n19118) );
in01f01 g15330 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_25_), .o(n19119) );
no02f01 g15331 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_2_), .b(n17966), .o(n19120) );
in01f01 g15332 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_1_), .o(n19121) );
na02f01 g15333 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .b(n19121), .o(n19122) );
in01f01 g15334 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_0_), .o(n19123) );
na02f01 g15335 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .b(n19123), .o(n19124) );
na02f01 g15336 ( .a(n19124), .b(n19122), .o(n19125) );
no02f01 g15337 ( .a(n19125), .b(n19120), .o(n19126) );
no02f01 g15338 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_4_), .b(n17966), .o(n19127) );
no02f01 g15339 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_5_), .b(n17966), .o(n19128) );
no02f01 g15340 ( .a(n17966), .b(delay_xor_ln22_unr6_stage3_stallmux_q_3_), .o(n19129) );
no03f01 g15341 ( .a(n19129), .b(n19128), .c(n19127), .o(n19130) );
na02f01 g15342 ( .a(n19130), .b(n19126), .o(n19131) );
in01f01 g15343 ( .a(n19131), .o(n19132) );
no02f01 g15344 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_6_), .b(n17966), .o(n19133) );
no02f01 g15345 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_8_), .b(n17966), .o(n19134) );
no02f01 g15346 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_7_), .b(n17966), .o(n19135) );
no03f01 g15347 ( .a(n19135), .b(n19134), .c(n19133), .o(n19136) );
na02f01 g15348 ( .a(n19136), .b(n19132), .o(n19137) );
no02f01 g15349 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_9_), .b(n17966), .o(n19138) );
no02f01 g15350 ( .a(n19138), .b(n19137), .o(n19139) );
in01f01 g15351 ( .a(n19139), .o(n19140) );
no02f01 g15352 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_10_), .b(n17966), .o(n19141) );
no02f01 g15353 ( .a(n19141), .b(n19140), .o(n19142) );
in01f01 g15354 ( .a(n19142), .o(n19143) );
no02f01 g15355 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_11_), .b(n17966), .o(n19144) );
no02f01 g15356 ( .a(n19144), .b(n19143), .o(n19145) );
in01f01 g15357 ( .a(n19145), .o(n19146) );
no02f01 g15358 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_12_), .b(n17966), .o(n19147) );
no02f01 g15359 ( .a(n19147), .b(n19146), .o(n19148) );
in01f01 g15360 ( .a(n19148), .o(n19149) );
no02f01 g15361 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_13_), .b(n17966), .o(n19150) );
no02f01 g15362 ( .a(n19150), .b(n19149), .o(n19151) );
in01f01 g15363 ( .a(n19151), .o(n19152) );
no02f01 g15364 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_14_), .b(n17966), .o(n19153) );
no02f01 g15365 ( .a(n19153), .b(n19152), .o(n19154) );
in01f01 g15366 ( .a(n19154), .o(n19155) );
no02f01 g15367 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_15_), .b(n17966), .o(n19156) );
no02f01 g15368 ( .a(n19156), .b(n19155), .o(n19157) );
in01f01 g15369 ( .a(n19157), .o(n19158) );
no02f01 g15370 ( .a(n17966), .b(delay_xor_ln22_unr6_stage3_stallmux_q_16_), .o(n19159) );
no02f01 g15371 ( .a(n19159), .b(n19158), .o(n19160) );
in01f01 g15372 ( .a(n19160), .o(n19161) );
no02f01 g15373 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_17_), .b(n17966), .o(n19162) );
no02f01 g15374 ( .a(n19162), .b(n19161), .o(n19163) );
in01f01 g15375 ( .a(n19163), .o(n19164) );
no02f01 g15376 ( .a(n17966), .b(delay_xor_ln22_unr6_stage3_stallmux_q_18_), .o(n19165) );
no02f01 g15377 ( .a(n19165), .b(n19164), .o(n19166) );
in01f01 g15378 ( .a(n19166), .o(n19167) );
no02f01 g15379 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_19_), .b(n17966), .o(n19168) );
no02f01 g15380 ( .a(n19168), .b(n19167), .o(n19169) );
in01f01 g15381 ( .a(n19169), .o(n19170) );
no02f01 g15382 ( .a(n17966), .b(delay_xor_ln22_unr6_stage3_stallmux_q_20_), .o(n19171) );
no02f01 g15383 ( .a(n19171), .b(n19170), .o(n19172) );
in01f01 g15384 ( .a(n19172), .o(n19173) );
no02f01 g15385 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_21_), .b(n17966), .o(n19174) );
no02f01 g15386 ( .a(n19174), .b(n19173), .o(n19175) );
in01f01 g15387 ( .a(n19175), .o(n19176) );
no02f01 g15388 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_22_), .b(n17966), .o(n19177) );
no02f01 g15389 ( .a(n19177), .b(n19176), .o(n19178) );
in01f01 g15390 ( .a(n19178), .o(n19179) );
no02f01 g15391 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_23_), .b(n17966), .o(n19180) );
no02f01 g15392 ( .a(n19180), .b(n19179), .o(n19181) );
in01f01 g15393 ( .a(n19181), .o(n19182) );
no02f01 g15394 ( .a(n17966), .b(delay_xor_ln22_unr6_stage3_stallmux_q_24_), .o(n19183) );
no02f01 g15395 ( .a(n19183), .b(n19182), .o(n19184) );
in01f01 g15396 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_25_), .o(n19185) );
no02f01 g15397 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .b(n19185), .o(n19186) );
no02f01 g15398 ( .a(n17966), .b(delay_xor_ln22_unr6_stage3_stallmux_q_25_), .o(n19187) );
no02f01 g15399 ( .a(n19187), .b(n19186), .o(n19188) );
in01f01 g15400 ( .a(n19188), .o(n19189) );
no02f01 g15401 ( .a(n19189), .b(n19184), .o(n19190) );
in01f01 g15402 ( .a(n19190), .o(n19191) );
na02f01 g15403 ( .a(n19189), .b(n19184), .o(n19192) );
na02f01 g15404 ( .a(n19192), .b(n19191), .o(n19193) );
in01f01 g15405 ( .a(n19193), .o(n19194) );
no02f01 g15406 ( .a(n19194), .b(n19119), .o(n19195) );
in01f01 g15407 ( .a(n19195), .o(n19196) );
in01f01 g15408 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_24_), .o(n19197) );
na02f01 g15409 ( .a(n17966), .b(delay_xor_ln22_unr6_stage3_stallmux_q_24_), .o(n19198) );
in01f01 g15410 ( .a(n19198), .o(n19199) );
no02f01 g15411 ( .a(n19199), .b(n19183), .o(n19200) );
in01f01 g15412 ( .a(n19200), .o(n19201) );
no02f01 g15413 ( .a(n19201), .b(n19181), .o(n19202) );
no02f01 g15414 ( .a(n19200), .b(n19182), .o(n19203) );
no02f01 g15415 ( .a(n19203), .b(n19202), .o(n19204) );
no02f01 g15416 ( .a(n19204), .b(n19197), .o(n19205) );
in01f01 g15417 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_23_), .o(n19206) );
na02f01 g15418 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_23_), .b(n17966), .o(n19207) );
in01f01 g15419 ( .a(n19207), .o(n19208) );
no02f01 g15420 ( .a(n19208), .b(n19180), .o(n19209) );
in01f01 g15421 ( .a(n19209), .o(n19210) );
no02f01 g15422 ( .a(n19210), .b(n19178), .o(n19211) );
no02f01 g15423 ( .a(n19209), .b(n19179), .o(n19212) );
no02f01 g15424 ( .a(n19212), .b(n19211), .o(n19213) );
no02f01 g15425 ( .a(n19213), .b(n19206), .o(n19214) );
in01f01 g15426 ( .a(n19214), .o(n19215) );
in01f01 g15427 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_22_), .o(n19216) );
na02f01 g15428 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_22_), .b(n17966), .o(n19217) );
in01f01 g15429 ( .a(n19217), .o(n19218) );
no02f01 g15430 ( .a(n19218), .b(n19177), .o(n19219) );
in01f01 g15431 ( .a(n19219), .o(n19220) );
no02f01 g15432 ( .a(n19220), .b(n19175), .o(n19221) );
no02f01 g15433 ( .a(n19219), .b(n19176), .o(n19222) );
no02f01 g15434 ( .a(n19222), .b(n19221), .o(n19223) );
no02f01 g15435 ( .a(n19223), .b(n19216), .o(n19224) );
in01f01 g15436 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_21_), .o(n19225) );
na02f01 g15437 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_21_), .b(n17966), .o(n19226) );
in01f01 g15438 ( .a(n19226), .o(n19227) );
no02f01 g15439 ( .a(n19227), .b(n19174), .o(n19228) );
no02f01 g15440 ( .a(n19228), .b(n19173), .o(n19229) );
na02f01 g15441 ( .a(n19228), .b(n19173), .o(n19230) );
in01f01 g15442 ( .a(n19230), .o(n19231) );
no02f01 g15443 ( .a(n19231), .b(n19229), .o(n19232) );
no02f01 g15444 ( .a(n19232), .b(n19225), .o(n19233) );
in01f01 g15445 ( .a(n19233), .o(n19234) );
in01f01 g15446 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_20_), .o(n19235) );
na02f01 g15447 ( .a(n17966), .b(delay_xor_ln22_unr6_stage3_stallmux_q_20_), .o(n19236) );
in01f01 g15448 ( .a(n19236), .o(n19237) );
no02f01 g15449 ( .a(n19237), .b(n19171), .o(n19238) );
in01f01 g15450 ( .a(n19238), .o(n19239) );
no02f01 g15451 ( .a(n19239), .b(n19169), .o(n19240) );
no02f01 g15452 ( .a(n19238), .b(n19170), .o(n19241) );
no02f01 g15453 ( .a(n19241), .b(n19240), .o(n19242) );
no02f01 g15454 ( .a(n19242), .b(n19235), .o(n19243) );
in01f01 g15455 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_19_), .o(n19244) );
na02f01 g15456 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_19_), .b(n17966), .o(n19245) );
in01f01 g15457 ( .a(n19245), .o(n19246) );
no02f01 g15458 ( .a(n19246), .b(n19168), .o(n19247) );
no02f01 g15459 ( .a(n19247), .b(n19167), .o(n19248) );
na02f01 g15460 ( .a(n19247), .b(n19167), .o(n19249) );
in01f01 g15461 ( .a(n19249), .o(n19250) );
no02f01 g15462 ( .a(n19250), .b(n19248), .o(n19251) );
no02f01 g15463 ( .a(n19251), .b(n19244), .o(n19252) );
in01f01 g15464 ( .a(n19252), .o(n19253) );
in01f01 g15465 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_18_), .o(n19254) );
na02f01 g15466 ( .a(n17966), .b(delay_xor_ln22_unr6_stage3_stallmux_q_18_), .o(n19255) );
in01f01 g15467 ( .a(n19255), .o(n19256) );
no02f01 g15468 ( .a(n19256), .b(n19165), .o(n19257) );
no02f01 g15469 ( .a(n19257), .b(n19164), .o(n19258) );
na02f01 g15470 ( .a(n19257), .b(n19164), .o(n19259) );
in01f01 g15471 ( .a(n19259), .o(n19260) );
no02f01 g15472 ( .a(n19260), .b(n19258), .o(n19261) );
no02f01 g15473 ( .a(n19261), .b(n19254), .o(n19262) );
in01f01 g15474 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_17_), .o(n19263) );
na02f01 g15475 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_17_), .b(n17966), .o(n19264) );
in01f01 g15476 ( .a(n19264), .o(n19265) );
no02f01 g15477 ( .a(n19265), .b(n19162), .o(n19266) );
no02f01 g15478 ( .a(n19266), .b(n19161), .o(n19267) );
na02f01 g15479 ( .a(n19266), .b(n19161), .o(n19268) );
in01f01 g15480 ( .a(n19268), .o(n19269) );
no02f01 g15481 ( .a(n19269), .b(n19267), .o(n19270) );
no02f01 g15482 ( .a(n19270), .b(n19263), .o(n19271) );
in01f01 g15483 ( .a(n19271), .o(n19272) );
in01f01 g15484 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_16_), .o(n19273) );
na02f01 g15485 ( .a(n17966), .b(delay_xor_ln22_unr6_stage3_stallmux_q_16_), .o(n19274) );
in01f01 g15486 ( .a(n19274), .o(n19275) );
no02f01 g15487 ( .a(n19275), .b(n19159), .o(n19276) );
in01f01 g15488 ( .a(n19276), .o(n19277) );
no02f01 g15489 ( .a(n19277), .b(n19157), .o(n19278) );
no02f01 g15490 ( .a(n19276), .b(n19158), .o(n19279) );
no02f01 g15491 ( .a(n19279), .b(n19278), .o(n19280) );
no02f01 g15492 ( .a(n19280), .b(n19273), .o(n19281) );
in01f01 g15493 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_15_), .o(n19282) );
na02f01 g15494 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_15_), .b(n17966), .o(n19283) );
in01f01 g15495 ( .a(n19283), .o(n19284) );
no02f01 g15496 ( .a(n19284), .b(n19156), .o(n19285) );
no02f01 g15497 ( .a(n19285), .b(n19155), .o(n19286) );
na02f01 g15498 ( .a(n19285), .b(n19155), .o(n19287) );
in01f01 g15499 ( .a(n19287), .o(n19288) );
no02f01 g15500 ( .a(n19288), .b(n19286), .o(n19289) );
no02f01 g15501 ( .a(n19289), .b(n19282), .o(n19290) );
in01f01 g15502 ( .a(n19290), .o(n19291) );
na02f01 g15503 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_14_), .b(n17966), .o(n19292) );
in01f01 g15504 ( .a(n19292), .o(n19293) );
no02f01 g15505 ( .a(n19293), .b(n19153), .o(n19294) );
no02f01 g15506 ( .a(n19294), .b(n19152), .o(n19295) );
na02f01 g15507 ( .a(n19294), .b(n19152), .o(n19296) );
in01f01 g15508 ( .a(n19296), .o(n19297) );
no02f01 g15509 ( .a(n19297), .b(n19295), .o(n19298) );
in01f01 g15510 ( .a(n19298), .o(n19299) );
no02f01 g15511 ( .a(n19299), .b(delay_add_ln22_unr5_stage3_stallmux_q_14_), .o(n19300) );
in01f01 g15512 ( .a(n19300), .o(n19301) );
in01f01 g15513 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_13_), .o(n19302) );
na02f01 g15514 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_13_), .b(n17966), .o(n19303) );
in01f01 g15515 ( .a(n19303), .o(n19304) );
no02f01 g15516 ( .a(n19304), .b(n19150), .o(n19305) );
no02f01 g15517 ( .a(n19305), .b(n19149), .o(n19306) );
na02f01 g15518 ( .a(n19305), .b(n19149), .o(n19307) );
in01f01 g15519 ( .a(n19307), .o(n19308) );
no02f01 g15520 ( .a(n19308), .b(n19306), .o(n19309) );
no02f01 g15521 ( .a(n19309), .b(n19302), .o(n19310) );
in01f01 g15522 ( .a(n19310), .o(n19311) );
in01f01 g15523 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_6_), .o(n19312) );
in01f01 g15524 ( .a(n19133), .o(n19313) );
na02f01 g15525 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_6_), .b(n17966), .o(n19314) );
na02f01 g15526 ( .a(n19314), .b(n19313), .o(n19315) );
no02f01 g15527 ( .a(n19315), .b(n19132), .o(n19316) );
na02f01 g15528 ( .a(n19315), .b(n19132), .o(n19317) );
in01f01 g15529 ( .a(n19317), .o(n19318) );
no02f01 g15530 ( .a(n19318), .b(n19316), .o(n19319) );
no02f01 g15531 ( .a(n19319), .b(n19312), .o(n19320) );
in01f01 g15532 ( .a(n19320), .o(n19321) );
na02f01 g15533 ( .a(n19319), .b(n19312), .o(n19322) );
in01f01 g15534 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_2_), .o(n19323) );
in01f01 g15535 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_2_), .o(n19324) );
no02f01 g15536 ( .a(n19324), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(n19325) );
no02f01 g15537 ( .a(n19325), .b(n19120), .o(n19326) );
no02f01 g15538 ( .a(n19326), .b(n19125), .o(n19327) );
no02f01 g15539 ( .a(n17966), .b(delay_xor_ln22_unr6_stage3_stallmux_q_1_), .o(n19328) );
no02f01 g15540 ( .a(n17966), .b(delay_xor_ln22_unr6_stage3_stallmux_q_0_), .o(n19329) );
no02f01 g15541 ( .a(n19329), .b(n19328), .o(n19330) );
no03f01 g15542 ( .a(n19325), .b(n19330), .c(n19120), .o(n19331) );
no02f01 g15543 ( .a(n19331), .b(n19327), .o(n19332) );
no02f01 g15544 ( .a(n19332), .b(n19323), .o(n19333) );
na02f01 g15545 ( .a(n17966), .b(delay_xor_ln22_unr6_stage3_stallmux_q_1_), .o(n19334) );
na02f01 g15546 ( .a(n19334), .b(n19122), .o(n19335) );
no02f01 g15547 ( .a(n19335), .b(n19124), .o(n19336) );
ao12f01 g15548 ( .a(n19329), .b(n19334), .c(n19122), .o(n19337) );
no02f01 g15549 ( .a(n19337), .b(n19336), .o(n19338) );
in01f01 g15550 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_0_), .o(n19339) );
no02f01 g15551 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .b(delay_xor_ln22_unr6_stage3_stallmux_q_0_), .o(n19340) );
in01f01 g15552 ( .a(n19340), .o(n19341) );
na02f01 g15553 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .b(delay_xor_ln22_unr6_stage3_stallmux_q_0_), .o(n19342) );
na02f01 g15554 ( .a(n19342), .b(n19341), .o(n19343) );
no02f01 g15555 ( .a(n19343), .b(n19339), .o(n19344) );
no02f01 g15556 ( .a(n19344), .b(delay_add_ln22_unr5_stage3_stallmux_q_1_), .o(n19345) );
na02f01 g15557 ( .a(n19344), .b(delay_add_ln22_unr5_stage3_stallmux_q_1_), .o(n19346) );
oa12f01 g15558 ( .a(n19346), .b(n19345), .c(n19338), .o(n19347) );
na02f01 g15559 ( .a(n19332), .b(n19323), .o(n19348) );
ao12f01 g15560 ( .a(n19333), .b(n19348), .c(n19347), .o(n19349) );
na02f01 g15561 ( .a(n19324), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(n19350) );
na02f01 g15562 ( .a(n19330), .b(n19350), .o(n19351) );
na02f01 g15563 ( .a(n17966), .b(delay_xor_ln22_unr6_stage3_stallmux_q_3_), .o(n19352) );
in01f01 g15564 ( .a(n19352), .o(n19353) );
no02f01 g15565 ( .a(n19353), .b(n19129), .o(n19354) );
no02f01 g15566 ( .a(n19354), .b(n19351), .o(n19355) );
no03f01 g15567 ( .a(n19353), .b(n19129), .c(n19126), .o(n19356) );
no03f01 g15568 ( .a(n19356), .b(n19355), .c(delay_add_ln22_unr5_stage3_stallmux_q_3_), .o(n19357) );
in01f01 g15569 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_3_), .o(n19358) );
no02f01 g15570 ( .a(n19356), .b(n19355), .o(n19359) );
no02f01 g15571 ( .a(n19359), .b(n19358), .o(n19360) );
in01f01 g15572 ( .a(n19360), .o(n19361) );
oa12f01 g15573 ( .a(n19361), .b(n19357), .c(n19349), .o(n19362) );
in01f01 g15574 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_4_), .o(n19363) );
in01f01 g15575 ( .a(n19127), .o(n19364) );
na02f01 g15576 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_4_), .b(n17966), .o(n19365) );
na02f01 g15577 ( .a(n19365), .b(n19364), .o(n19366) );
no02f01 g15578 ( .a(n19129), .b(n19351), .o(n19367) );
na02f01 g15579 ( .a(n19367), .b(n19366), .o(n19368) );
in01f01 g15580 ( .a(n19368), .o(n19369) );
no02f01 g15581 ( .a(n19367), .b(n19366), .o(n19370) );
no02f01 g15582 ( .a(n19370), .b(n19369), .o(n19371) );
na02f01 g15583 ( .a(n19371), .b(n19363), .o(n19372) );
no02f01 g15584 ( .a(n19371), .b(n19363), .o(n19373) );
ao12f01 g15585 ( .a(n19373), .b(n19372), .c(n19362), .o(n19374) );
na02f01 g15586 ( .a(n19367), .b(n19364), .o(n19375) );
na02f01 g15587 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_5_), .b(n17966), .o(n19376) );
in01f01 g15588 ( .a(n19376), .o(n19377) );
no02f01 g15589 ( .a(n19377), .b(n19128), .o(n19378) );
no02f01 g15590 ( .a(n19378), .b(n19375), .o(n19379) );
na02f01 g15591 ( .a(n19378), .b(n19375), .o(n19380) );
in01f01 g15592 ( .a(n19380), .o(n19381) );
no02f01 g15593 ( .a(n19381), .b(n19379), .o(n19382) );
in01f01 g15594 ( .a(n19382), .o(n19383) );
no02f01 g15595 ( .a(n19383), .b(delay_add_ln22_unr5_stage3_stallmux_q_5_), .o(n19384) );
na02f01 g15596 ( .a(n19383), .b(delay_add_ln22_unr5_stage3_stallmux_q_5_), .o(n19385) );
oa12f01 g15597 ( .a(n19385), .b(n19384), .c(n19374), .o(n19386) );
na02f01 g15598 ( .a(n19386), .b(n19322), .o(n19387) );
na02f01 g15599 ( .a(n19387), .b(n19321), .o(n19388) );
no02f01 g15600 ( .a(n19133), .b(n19131), .o(n19389) );
in01f01 g15601 ( .a(n19135), .o(n19390) );
na02f01 g15602 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_7_), .b(n17966), .o(n19391) );
na02f01 g15603 ( .a(n19391), .b(n19390), .o(n19392) );
no02f01 g15604 ( .a(n19392), .b(n19389), .o(n19393) );
na02f01 g15605 ( .a(n19392), .b(n19389), .o(n19394) );
in01f01 g15606 ( .a(n19394), .o(n19395) );
no02f01 g15607 ( .a(n19395), .b(n19393), .o(n19396) );
in01f01 g15608 ( .a(n19396), .o(n19397) );
no02f01 g15609 ( .a(n19397), .b(delay_add_ln22_unr5_stage3_stallmux_q_7_), .o(n19398) );
in01f01 g15610 ( .a(n19398), .o(n19399) );
na02f01 g15611 ( .a(n19399), .b(n19388), .o(n19400) );
na02f01 g15612 ( .a(n19397), .b(delay_add_ln22_unr5_stage3_stallmux_q_7_), .o(n19401) );
na02f01 g15613 ( .a(n19401), .b(n19400), .o(n19402) );
na02f01 g15614 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_8_), .b(n17966), .o(n19403) );
in01f01 g15615 ( .a(n19403), .o(n19404) );
no02f01 g15616 ( .a(n19404), .b(n19134), .o(n19405) );
in01f01 g15617 ( .a(n19405), .o(n19406) );
ao12f01 g15618 ( .a(n19406), .b(n19389), .c(n19390), .o(n19407) );
no04f01 g15619 ( .a(n19405), .b(n19135), .c(n19133), .d(n19131), .o(n19408) );
no02f01 g15620 ( .a(n19408), .b(n19407), .o(n19409) );
in01f01 g15621 ( .a(n19409), .o(n19410) );
no02f01 g15622 ( .a(n19410), .b(delay_add_ln22_unr5_stage3_stallmux_q_8_), .o(n19411) );
in01f01 g15623 ( .a(n19411), .o(n19412) );
na02f01 g15624 ( .a(n19412), .b(n19402), .o(n19413) );
na02f01 g15625 ( .a(n19410), .b(delay_add_ln22_unr5_stage3_stallmux_q_8_), .o(n19414) );
na02f01 g15626 ( .a(n19414), .b(n19413), .o(n19415) );
na02f01 g15627 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_9_), .b(n17966), .o(n19416) );
in01f01 g15628 ( .a(n19416), .o(n19417) );
no02f01 g15629 ( .a(n19417), .b(n19138), .o(n19418) );
no02f01 g15630 ( .a(n19418), .b(n19137), .o(n19419) );
na02f01 g15631 ( .a(n19418), .b(n19137), .o(n19420) );
in01f01 g15632 ( .a(n19420), .o(n19421) );
no02f01 g15633 ( .a(n19421), .b(n19419), .o(n19422) );
in01f01 g15634 ( .a(n19422), .o(n19423) );
no02f01 g15635 ( .a(n19423), .b(delay_add_ln22_unr5_stage3_stallmux_q_9_), .o(n19424) );
in01f01 g15636 ( .a(n19424), .o(n19425) );
na02f01 g15637 ( .a(n19425), .b(n19415), .o(n19426) );
na02f01 g15638 ( .a(n19423), .b(delay_add_ln22_unr5_stage3_stallmux_q_9_), .o(n19427) );
na02f01 g15639 ( .a(n19427), .b(n19426), .o(n19428) );
na02f01 g15640 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_10_), .b(n17966), .o(n19429) );
in01f01 g15641 ( .a(n19429), .o(n19430) );
no02f01 g15642 ( .a(n19430), .b(n19141), .o(n19431) );
in01f01 g15643 ( .a(n19431), .o(n19432) );
no02f01 g15644 ( .a(n19432), .b(n19139), .o(n19433) );
no02f01 g15645 ( .a(n19431), .b(n19140), .o(n19434) );
no02f01 g15646 ( .a(n19434), .b(n19433), .o(n19435) );
in01f01 g15647 ( .a(n19435), .o(n19436) );
no02f01 g15648 ( .a(n19436), .b(delay_add_ln22_unr5_stage3_stallmux_q_10_), .o(n19437) );
in01f01 g15649 ( .a(n19437), .o(n19438) );
na02f01 g15650 ( .a(n19438), .b(n19428), .o(n19439) );
na02f01 g15651 ( .a(n19436), .b(delay_add_ln22_unr5_stage3_stallmux_q_10_), .o(n19440) );
na02f01 g15652 ( .a(n19440), .b(n19439), .o(n19441) );
na02f01 g15653 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_11_), .b(n17966), .o(n19442) );
in01f01 g15654 ( .a(n19442), .o(n19443) );
no02f01 g15655 ( .a(n19443), .b(n19144), .o(n19444) );
no02f01 g15656 ( .a(n19444), .b(n19143), .o(n19445) );
na02f01 g15657 ( .a(n19444), .b(n19143), .o(n19446) );
in01f01 g15658 ( .a(n19446), .o(n19447) );
no02f01 g15659 ( .a(n19447), .b(n19445), .o(n19448) );
in01f01 g15660 ( .a(n19448), .o(n19449) );
no02f01 g15661 ( .a(n19449), .b(delay_add_ln22_unr5_stage3_stallmux_q_11_), .o(n19450) );
in01f01 g15662 ( .a(n19450), .o(n19451) );
na02f01 g15663 ( .a(n19451), .b(n19441), .o(n19452) );
na02f01 g15664 ( .a(n19449), .b(delay_add_ln22_unr5_stage3_stallmux_q_11_), .o(n19453) );
na02f01 g15665 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_12_), .b(n17966), .o(n19454) );
in01f01 g15666 ( .a(n19454), .o(n19455) );
no02f01 g15667 ( .a(n19455), .b(n19147), .o(n19456) );
no02f01 g15668 ( .a(n19456), .b(n19146), .o(n19457) );
na02f01 g15669 ( .a(n19456), .b(n19146), .o(n19458) );
in01f01 g15670 ( .a(n19458), .o(n19459) );
no02f01 g15671 ( .a(n19459), .b(n19457), .o(n19460) );
in01f01 g15672 ( .a(n19460), .o(n19461) );
no02f01 g15673 ( .a(n19461), .b(delay_add_ln22_unr5_stage3_stallmux_q_12_), .o(n19462) );
ao12f01 g15674 ( .a(n19462), .b(n19453), .c(n19452), .o(n19463) );
na02f01 g15675 ( .a(n19461), .b(delay_add_ln22_unr5_stage3_stallmux_q_12_), .o(n19464) );
in01f01 g15676 ( .a(n19464), .o(n19465) );
na02f01 g15677 ( .a(n19309), .b(n19302), .o(n19466) );
oa12f01 g15678 ( .a(n19466), .b(n19465), .c(n19463), .o(n19467) );
na02f01 g15679 ( .a(n19299), .b(delay_add_ln22_unr5_stage3_stallmux_q_14_), .o(n19468) );
na03f01 g15680 ( .a(n19468), .b(n19467), .c(n19311), .o(n19469) );
na02f01 g15681 ( .a(n19289), .b(n19282), .o(n19470) );
na03f01 g15682 ( .a(n19470), .b(n19469), .c(n19301), .o(n19471) );
na02f01 g15683 ( .a(n19280), .b(n19273), .o(n19472) );
in01f01 g15684 ( .a(n19472), .o(n19473) );
ao12f01 g15685 ( .a(n19473), .b(n19471), .c(n19291), .o(n19474) );
na02f01 g15686 ( .a(n19270), .b(n19263), .o(n19475) );
oa12f01 g15687 ( .a(n19475), .b(n19474), .c(n19281), .o(n19476) );
na02f01 g15688 ( .a(n19261), .b(n19254), .o(n19477) );
in01f01 g15689 ( .a(n19477), .o(n19478) );
ao12f01 g15690 ( .a(n19478), .b(n19476), .c(n19272), .o(n19479) );
na02f01 g15691 ( .a(n19251), .b(n19244), .o(n19480) );
oa12f01 g15692 ( .a(n19480), .b(n19479), .c(n19262), .o(n19481) );
na02f01 g15693 ( .a(n19242), .b(n19235), .o(n19482) );
in01f01 g15694 ( .a(n19482), .o(n19483) );
ao12f01 g15695 ( .a(n19483), .b(n19481), .c(n19253), .o(n19484) );
na02f01 g15696 ( .a(n19232), .b(n19225), .o(n19485) );
oa12f01 g15697 ( .a(n19485), .b(n19484), .c(n19243), .o(n19486) );
na02f01 g15698 ( .a(n19223), .b(n19216), .o(n19487) );
in01f01 g15699 ( .a(n19487), .o(n19488) );
ao12f01 g15700 ( .a(n19488), .b(n19486), .c(n19234), .o(n19489) );
na02f01 g15701 ( .a(n19213), .b(n19206), .o(n19490) );
oa12f01 g15702 ( .a(n19490), .b(n19489), .c(n19224), .o(n19491) );
na02f01 g15703 ( .a(n19204), .b(n19197), .o(n19492) );
in01f01 g15704 ( .a(n19492), .o(n19493) );
ao12f01 g15705 ( .a(n19493), .b(n19491), .c(n19215), .o(n19494) );
no02f01 g15706 ( .a(n19193), .b(delay_add_ln22_unr5_stage3_stallmux_q_25_), .o(n19495) );
in01f01 g15707 ( .a(n19495), .o(n19496) );
oa12f01 g15708 ( .a(n19496), .b(n19494), .c(n19205), .o(n19497) );
na02f01 g15709 ( .a(n19497), .b(n19196), .o(n19498) );
no02f01 g15710 ( .a(n19190), .b(n19186), .o(n19499) );
in01f01 g15711 ( .a(n19499), .o(n19500) );
in01f01 g15712 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_27_), .o(n19501) );
in01f01 g15713 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_26_), .o(n19502) );
no02f01 g15714 ( .a(n19502), .b(n19501), .o(n19503) );
no02f01 g15715 ( .a(n19503), .b(n19500), .o(n19504) );
in01f01 g15716 ( .a(n19504), .o(n19505) );
na02f01 g15717 ( .a(n19505), .b(n19498), .o(n19506) );
no02f01 g15718 ( .a(n19499), .b(n19502), .o(n19507) );
no02f01 g15719 ( .a(n19499), .b(n19501), .o(n19508) );
no02f01 g15720 ( .a(n19508), .b(n19507), .o(n19509) );
na02f01 g15721 ( .a(n19509), .b(n19506), .o(n19510) );
no02f01 g15722 ( .a(n19500), .b(delay_add_ln22_unr5_stage3_stallmux_q_29_), .o(n19511) );
no02f01 g15723 ( .a(n19500), .b(delay_add_ln22_unr5_stage3_stallmux_q_28_), .o(n19512) );
no02f01 g15724 ( .a(n19512), .b(n19511), .o(n19513) );
na02f01 g15725 ( .a(n19513), .b(n19510), .o(n19514) );
no02f01 g15726 ( .a(n19500), .b(delay_add_ln22_unr5_stage3_stallmux_q_30_), .o(n19515) );
in01f01 g15727 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_30_), .o(n19516) );
no02f01 g15728 ( .a(n19499), .b(n19516), .o(n19517) );
no02f01 g15729 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_29_), .b(delay_add_ln22_unr5_stage3_stallmux_q_28_), .o(n19518) );
no02f01 g15730 ( .a(n19518), .b(n19499), .o(n19519) );
no02f01 g15731 ( .a(n19519), .b(n19517), .o(n19520) );
oa12f01 g15732 ( .a(n19520), .b(n19515), .c(n19514), .o(n19521) );
in01f01 g15733 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_31_), .o(n19522) );
no02f01 g15734 ( .a(n19499), .b(n19522), .o(n19523) );
no02f01 g15735 ( .a(n19500), .b(delay_add_ln22_unr5_stage3_stallmux_q_31_), .o(n19524) );
no02f01 g15736 ( .a(n19524), .b(n19523), .o(n19525) );
in01f01 g15737 ( .a(n19525), .o(n19526) );
no02f01 g15738 ( .a(n19526), .b(n19521), .o(n19527) );
na02f01 g15739 ( .a(n19526), .b(n19521), .o(n19528) );
in01f01 g15740 ( .a(n19528), .o(n19529) );
no02f01 g15741 ( .a(n19529), .b(n19527), .o(n19530) );
no02f01 g15742 ( .a(n19530), .b(n19118), .o(n19531) );
in01f01 g15743 ( .a(n19118), .o(n19532) );
in01f01 g15744 ( .a(n19527), .o(n19533) );
na02f01 g15745 ( .a(n19528), .b(n19533), .o(n19534) );
no02f01 g15746 ( .a(n19534), .b(n19532), .o(n19535) );
no02f01 g15747 ( .a(n19535), .b(n19531), .o(n19536) );
no02f01 g15748 ( .a(n19500), .b(delay_add_ln22_unr5_stage3_stallmux_q_27_), .o(n19537) );
no02f01 g15749 ( .a(n19537), .b(n19508), .o(n19538) );
in01f01 g15750 ( .a(n19538), .o(n19539) );
no02f01 g15751 ( .a(n19500), .b(delay_add_ln22_unr5_stage3_stallmux_q_26_), .o(n19540) );
ao12f01 g15752 ( .a(n19540), .b(n19497), .c(n19196), .o(n19541) );
no03f01 g15753 ( .a(n19541), .b(n19539), .c(n19507), .o(n19542) );
in01f01 g15754 ( .a(n19542), .o(n19543) );
oa12f01 g15755 ( .a(n19539), .b(n19541), .c(n19507), .o(n19544) );
na02f01 g15756 ( .a(n19544), .b(n19543), .o(n19545) );
no02f01 g15757 ( .a(n19495), .b(n19195), .o(n19546) );
in01f01 g15758 ( .a(n19546), .o(n19547) );
oa12f01 g15759 ( .a(n19547), .b(n19494), .c(n19205), .o(n19548) );
no03f01 g15760 ( .a(n19547), .b(n19494), .c(n19205), .o(n19549) );
in01f01 g15761 ( .a(n19549), .o(n19550) );
na02f01 g15762 ( .a(n19550), .b(n19548), .o(n19551) );
no03f01 g15763 ( .a(n19551), .b(n19117), .c(n19113), .o(n19552) );
na02f01 g15764 ( .a(n19112), .b(n18868), .o(n19553) );
na02f01 g15765 ( .a(n19102), .b(n18145), .o(n19554) );
oa12f01 g15766 ( .a(n18145), .b(n18895), .c(n18889), .o(n19555) );
oa12f01 g15767 ( .a(n19036), .b(n18905), .c(n18103), .o(n19556) );
na02f01 g15768 ( .a(n19028), .b(n19032), .o(n19557) );
na02f01 g15769 ( .a(n19029), .b(n19027), .o(n19558) );
na02f01 g15770 ( .a(n19558), .b(n19557), .o(n19559) );
na02f01 g15771 ( .a(n19559), .b(n18103), .o(n19560) );
na02f01 g15772 ( .a(n19039), .b(n19560), .o(n19561) );
ao12f01 g15773 ( .a(n19561), .b(n18906), .c(n18103), .o(n19562) );
na02f01 g15774 ( .a(n19562), .b(n19556), .o(n19563) );
oa12f01 g15775 ( .a(n19563), .b(n19050), .c(n18103), .o(n19564) );
in01f01 g15776 ( .a(n19059), .o(n19565) );
ao12f01 g15777 ( .a(n19564), .b(n19565), .c(n18145), .o(n19566) );
oa12f01 g15778 ( .a(n19566), .b(n19067), .c(n18103), .o(n19567) );
ao12f01 g15779 ( .a(n19567), .b(n19077), .c(n18145), .o(n19568) );
ao12f01 g15780 ( .a(n19078), .b(n19068), .c(n18103), .o(n19569) );
oa12f01 g15781 ( .a(n19569), .b(n19074), .c(n18145), .o(n19570) );
oa22f01 g15782 ( .a(n19108), .b(n18103), .c(n19570), .d(n19568), .o(n19571) );
ao12f01 g15783 ( .a(n19571), .b(n19106), .c(n18145), .o(n19572) );
na03f01 g15784 ( .a(n19572), .b(n19555), .c(n19554), .o(n19573) );
in01f01 g15785 ( .a(n19111), .o(n19574) );
na02f01 g15786 ( .a(n19574), .b(n19573), .o(n19575) );
na02f01 g15787 ( .a(n19575), .b(n19114), .o(n19576) );
na02f01 g15788 ( .a(n19491), .b(n19215), .o(n19577) );
no02f01 g15789 ( .a(n19493), .b(n19205), .o(n19578) );
in01f01 g15790 ( .a(n19578), .o(n19579) );
no02f01 g15791 ( .a(n19579), .b(n19577), .o(n19580) );
na02f01 g15792 ( .a(n19579), .b(n19577), .o(n19581) );
in01f01 g15793 ( .a(n19581), .o(n19582) );
no02f01 g15794 ( .a(n19582), .b(n19580), .o(n19583) );
ao12f01 g15795 ( .a(n19583), .b(n19576), .c(n19553), .o(n19584) );
na02f01 g15796 ( .a(n19090), .b(n18103), .o(n19585) );
ao12f01 g15797 ( .a(n19096), .b(n19585), .c(n19571), .o(n19586) );
no03f01 g15798 ( .a(n19109), .b(n19106), .c(n19091), .o(n19587) );
no02f01 g15799 ( .a(n19484), .b(n19243), .o(n19588) );
in01f01 g15800 ( .a(n19485), .o(n19589) );
no02f01 g15801 ( .a(n19589), .b(n19233), .o(n19590) );
na02f01 g15802 ( .a(n19590), .b(n19588), .o(n19591) );
no02f01 g15803 ( .a(n19590), .b(n19588), .o(n19592) );
in01f01 g15804 ( .a(n19592), .o(n19593) );
na02f01 g15805 ( .a(n19593), .b(n19591), .o(n19594) );
no03f01 g15806 ( .a(n19594), .b(n19587), .c(n19586), .o(n19595) );
no02f01 g15807 ( .a(n19570), .b(n19568), .o(n19596) );
no02f01 g15808 ( .a(n19108), .b(n18103), .o(n19597) );
no02f01 g15809 ( .a(n19109), .b(n19597), .o(n19598) );
no02f01 g15810 ( .a(n19598), .b(n19596), .o(n19599) );
na02f01 g15811 ( .a(n19081), .b(n19075), .o(n19600) );
na02f01 g15812 ( .a(n19090), .b(n18145), .o(n19601) );
na02f01 g15813 ( .a(n19585), .b(n19601), .o(n19602) );
no02f01 g15814 ( .a(n19602), .b(n19600), .o(n19603) );
na02f01 g15815 ( .a(n19481), .b(n19253), .o(n19604) );
no02f01 g15816 ( .a(n19483), .b(n19243), .o(n19605) );
in01f01 g15817 ( .a(n19605), .o(n19606) );
no02f01 g15818 ( .a(n19606), .b(n19604), .o(n19607) );
in01f01 g15819 ( .a(n19607), .o(n19608) );
na02f01 g15820 ( .a(n19606), .b(n19604), .o(n19609) );
na02f01 g15821 ( .a(n19609), .b(n19608), .o(n19610) );
oa12f01 g15822 ( .a(n19610), .b(n19603), .c(n19599), .o(n19611) );
oa12f01 g15823 ( .a(n19594), .b(n19587), .c(n19586), .o(n19612) );
ao12f01 g15824 ( .a(n19595), .b(n19612), .c(n19611), .o(n19613) );
na02f01 g15825 ( .a(n19569), .b(n19567), .o(n19614) );
na02f01 g15826 ( .a(n19614), .b(n19077), .o(n19615) );
no02f01 g15827 ( .a(n19080), .b(n19069), .o(n19616) );
na02f01 g15828 ( .a(n19616), .b(n19074), .o(n19617) );
na02f01 g15829 ( .a(n19617), .b(n19615), .o(n19618) );
no02f01 g15830 ( .a(n19479), .b(n19262), .o(n19619) );
in01f01 g15831 ( .a(n19480), .o(n19620) );
no02f01 g15832 ( .a(n19620), .b(n19252), .o(n19621) );
na02f01 g15833 ( .a(n19621), .b(n19619), .o(n19622) );
no02f01 g15834 ( .a(n19621), .b(n19619), .o(n19623) );
in01f01 g15835 ( .a(n19623), .o(n19624) );
na02f01 g15836 ( .a(n19624), .b(n19622), .o(n19625) );
no02f01 g15837 ( .a(n19625), .b(n19618), .o(n19626) );
no02f01 g15838 ( .a(n19078), .b(n19566), .o(n19627) );
no02f01 g15839 ( .a(n19627), .b(n19067), .o(n19628) );
na02f01 g15840 ( .a(n19079), .b(n19060), .o(n19629) );
no02f01 g15841 ( .a(n19629), .b(n19068), .o(n19630) );
no02f01 g15842 ( .a(n19630), .b(n19628), .o(n19631) );
na02f01 g15843 ( .a(n19476), .b(n19272), .o(n19632) );
no02f01 g15844 ( .a(n19478), .b(n19262), .o(n19633) );
in01f01 g15845 ( .a(n19633), .o(n19634) );
no02f01 g15846 ( .a(n19634), .b(n19632), .o(n19635) );
na02f01 g15847 ( .a(n19634), .b(n19632), .o(n19636) );
in01f01 g15848 ( .a(n19636), .o(n19637) );
no02f01 g15849 ( .a(n19637), .b(n19635), .o(n19638) );
no02f01 g15850 ( .a(n19638), .b(n19631), .o(n19639) );
na02f01 g15851 ( .a(n19039), .b(n19009), .o(n19640) );
no02f01 g15852 ( .a(n19640), .b(n19037), .o(n19641) );
oa12f01 g15853 ( .a(n19641), .b(n19035), .c(n19003), .o(n19642) );
no02f01 g15854 ( .a(n19642), .b(n18906), .o(n19643) );
in01f01 g15855 ( .a(n19642), .o(n19644) );
no02f01 g15856 ( .a(n19644), .b(n18905), .o(n19645) );
na02f01 g15857 ( .a(n19469), .b(n19301), .o(n19646) );
in01f01 g15858 ( .a(n19470), .o(n19647) );
no02f01 g15859 ( .a(n19647), .b(n19290), .o(n19648) );
no02f01 g15860 ( .a(n19648), .b(n19646), .o(n19649) );
na02f01 g15861 ( .a(n19648), .b(n19646), .o(n19650) );
in01f01 g15862 ( .a(n19650), .o(n19651) );
no02f01 g15863 ( .a(n19651), .b(n19649), .o(n19652) );
in01f01 g15864 ( .a(n19652), .o(n19653) );
no03f01 g15865 ( .a(n19653), .b(n19645), .c(n19643), .o(n19654) );
in01f01 g15866 ( .a(n19654), .o(n19655) );
in01f01 g15867 ( .a(n19003), .o(n19656) );
in01f01 g15868 ( .a(n19025), .o(n19657) );
in01f01 g15869 ( .a(n19038), .o(n19658) );
na02f01 g15870 ( .a(n19658), .b(n19009), .o(n19659) );
ao12f01 g15871 ( .a(n19659), .b(n19657), .c(n19656), .o(n19660) );
in01f01 g15872 ( .a(n19660), .o(n19661) );
no02f01 g15873 ( .a(n19661), .b(n19017), .o(n19662) );
in01f01 g15874 ( .a(n19014), .o(n19663) );
no02f01 g15875 ( .a(n19015), .b(n19663), .o(n19664) );
no02f01 g15876 ( .a(n19660), .b(n19664), .o(n19665) );
no02f01 g15877 ( .a(n19465), .b(n19463), .o(n19666) );
in01f01 g15878 ( .a(n19666), .o(n19667) );
in01f01 g15879 ( .a(n19466), .o(n19668) );
no02f01 g15880 ( .a(n19668), .b(n19310), .o(n19669) );
in01f01 g15881 ( .a(n19669), .o(n19670) );
no02f01 g15882 ( .a(n19670), .b(n19667), .o(n19671) );
no02f01 g15883 ( .a(n19669), .b(n19666), .o(n19672) );
no02f01 g15884 ( .a(n19672), .b(n19671), .o(n19673) );
in01f01 g15885 ( .a(n19673), .o(n19674) );
no03f01 g15886 ( .a(n19674), .b(n19665), .c(n19662), .o(n19675) );
in01f01 g15887 ( .a(n19675), .o(n19676) );
no02f01 g15888 ( .a(n19008), .b(n18996), .o(n19677) );
no02f01 g15889 ( .a(n19677), .b(n19002), .o(n19678) );
na02f01 g15890 ( .a(n19677), .b(n19002), .o(n19679) );
in01f01 g15891 ( .a(n19679), .o(n19680) );
no02f01 g15892 ( .a(n19680), .b(n19678), .o(n19681) );
in01f01 g15893 ( .a(n19441), .o(n19682) );
in01f01 g15894 ( .a(n19453), .o(n19683) );
no02f01 g15895 ( .a(n19683), .b(n19450), .o(n19684) );
no02f01 g15896 ( .a(n19684), .b(n19682), .o(n19685) );
na02f01 g15897 ( .a(n19684), .b(n19682), .o(n19686) );
in01f01 g15898 ( .a(n19686), .o(n19687) );
no02f01 g15899 ( .a(n19687), .b(n19685), .o(n19688) );
no02f01 g15900 ( .a(n19688), .b(n19681), .o(n19689) );
in01f01 g15901 ( .a(n19689), .o(n19690) );
na02f01 g15902 ( .a(n19007), .b(n18987), .o(n19691) );
na02f01 g15903 ( .a(n19691), .b(n18995), .o(n19692) );
in01f01 g15904 ( .a(n19692), .o(n19693) );
no02f01 g15905 ( .a(n19691), .b(n18995), .o(n19694) );
no02f01 g15906 ( .a(n19694), .b(n19693), .o(n19695) );
in01f01 g15907 ( .a(n19440), .o(n19696) );
no02f01 g15908 ( .a(n19696), .b(n19437), .o(n19697) );
in01f01 g15909 ( .a(n19697), .o(n19698) );
no02f01 g15910 ( .a(n19698), .b(n19428), .o(n19699) );
ao12f01 g15911 ( .a(n19697), .b(n19427), .c(n19426), .o(n19700) );
no02f01 g15912 ( .a(n19700), .b(n19699), .o(n19701) );
no02f01 g15913 ( .a(n19701), .b(n19695), .o(n19702) );
no03f01 g15914 ( .a(n19006), .b(n19005), .c(n18980), .o(n19703) );
no02f01 g15915 ( .a(n19006), .b(n18980), .o(n19704) );
no02f01 g15916 ( .a(n19704), .b(n18986), .o(n19705) );
no02f01 g15917 ( .a(n19705), .b(n19703), .o(n19706) );
in01f01 g15918 ( .a(n19415), .o(n19707) );
in01f01 g15919 ( .a(n19427), .o(n19708) );
no02f01 g15920 ( .a(n19708), .b(n19424), .o(n19709) );
no02f01 g15921 ( .a(n19709), .b(n19707), .o(n19710) );
na02f01 g15922 ( .a(n19709), .b(n19707), .o(n19711) );
in01f01 g15923 ( .a(n19711), .o(n19712) );
no02f01 g15924 ( .a(n19712), .b(n19710), .o(n19713) );
na02f01 g15925 ( .a(n19713), .b(n19706), .o(n19714) );
in01f01 g15926 ( .a(n19714), .o(n19715) );
no02f01 g15927 ( .a(n19713), .b(n19706), .o(n19716) );
in01f01 g15928 ( .a(n18971), .o(n19717) );
no02f01 g15929 ( .a(n18979), .b(n19717), .o(n19718) );
na02f01 g15930 ( .a(n18979), .b(n19717), .o(n19719) );
in01f01 g15931 ( .a(n19719), .o(n19720) );
no02f01 g15932 ( .a(n19720), .b(n19718), .o(n19721) );
in01f01 g15933 ( .a(n19414), .o(n19722) );
no02f01 g15934 ( .a(n19722), .b(n19411), .o(n19723) );
in01f01 g15935 ( .a(n19723), .o(n19724) );
no02f01 g15936 ( .a(n19724), .b(n19402), .o(n19725) );
ao12f01 g15937 ( .a(n19723), .b(n19401), .c(n19400), .o(n19726) );
no02f01 g15938 ( .a(n19726), .b(n19725), .o(n19727) );
no02f01 g15939 ( .a(n19727), .b(n19721), .o(n19728) );
in01f01 g15940 ( .a(n18964), .o(n19729) );
no02f01 g15941 ( .a(n18970), .b(n19729), .o(n19730) );
na02f01 g15942 ( .a(n18970), .b(n19729), .o(n19731) );
in01f01 g15943 ( .a(n19731), .o(n19732) );
no02f01 g15944 ( .a(n19732), .b(n19730), .o(n19733) );
na02f01 g15945 ( .a(n19401), .b(n19399), .o(n19734) );
in01f01 g15946 ( .a(n19734), .o(n19735) );
ao12f01 g15947 ( .a(n19735), .b(n19387), .c(n19321), .o(n19736) );
no02f01 g15948 ( .a(n19734), .b(n19388), .o(n19737) );
no02f01 g15949 ( .a(n19737), .b(n19736), .o(n19738) );
no02f01 g15950 ( .a(n19738), .b(n19733), .o(n19739) );
in01f01 g15951 ( .a(n19739), .o(n19740) );
in01f01 g15952 ( .a(n18955), .o(n19741) );
no02f01 g15953 ( .a(n18963), .b(n19741), .o(n19742) );
na02f01 g15954 ( .a(n18963), .b(n19741), .o(n19743) );
in01f01 g15955 ( .a(n19743), .o(n19744) );
no02f01 g15956 ( .a(n19744), .b(n19742), .o(n19745) );
in01f01 g15957 ( .a(n19386), .o(n19746) );
na02f01 g15958 ( .a(n19322), .b(n19321), .o(n19747) );
in01f01 g15959 ( .a(n19747), .o(n19748) );
no02f01 g15960 ( .a(n19748), .b(n19746), .o(n19749) );
no02f01 g15961 ( .a(n19747), .b(n19386), .o(n19750) );
no02f01 g15962 ( .a(n19750), .b(n19749), .o(n19751) );
no02f01 g15963 ( .a(n19751), .b(n19745), .o(n19752) );
no03f01 g15964 ( .a(n18952), .b(n18945), .c(n18937), .o(n19753) );
in01f01 g15965 ( .a(n18952), .o(n19754) );
no02f01 g15966 ( .a(n19754), .b(n18946), .o(n19755) );
no02f01 g15967 ( .a(n19755), .b(n19753), .o(n19756) );
in01f01 g15968 ( .a(n19374), .o(n19757) );
in01f01 g15969 ( .a(n19385), .o(n19758) );
no03f01 g15970 ( .a(n19758), .b(n19384), .c(n19757), .o(n19759) );
in01f01 g15971 ( .a(n19384), .o(n19760) );
ao12f01 g15972 ( .a(n19374), .b(n19385), .c(n19760), .o(n19761) );
no02f01 g15973 ( .a(n19761), .b(n19759), .o(n19762) );
no02f01 g15974 ( .a(n19762), .b(n19756), .o(n19763) );
in01f01 g15975 ( .a(n19763), .o(n19764) );
na02f01 g15976 ( .a(n18944), .b(n18937), .o(n19765) );
in01f01 g15977 ( .a(n19765), .o(n19766) );
no02f01 g15978 ( .a(n18944), .b(n18937), .o(n19767) );
no02f01 g15979 ( .a(n19767), .b(n19766), .o(n19768) );
in01f01 g15980 ( .a(n19362), .o(n19769) );
in01f01 g15981 ( .a(n19372), .o(n19770) );
no02f01 g15982 ( .a(n19373), .b(n19770), .o(n19771) );
no02f01 g15983 ( .a(n19771), .b(n19769), .o(n19772) );
na02f01 g15984 ( .a(n19771), .b(n19769), .o(n19773) );
in01f01 g15985 ( .a(n19773), .o(n19774) );
no02f01 g15986 ( .a(n19774), .b(n19772), .o(n19775) );
no02f01 g15987 ( .a(n19775), .b(n19768), .o(n19776) );
in01f01 g15988 ( .a(n19775), .o(n19777) );
no03f01 g15989 ( .a(n19777), .b(n19767), .c(n19766), .o(n19778) );
no02f01 g15990 ( .a(n18935), .b(n18928), .o(n19779) );
in01f01 g15991 ( .a(n19779), .o(n19780) );
na02f01 g15992 ( .a(n18935), .b(n18928), .o(n19781) );
in01f01 g15993 ( .a(n19349), .o(n19782) );
no03f01 g15994 ( .a(n19360), .b(n19357), .c(n19782), .o(n19783) );
no02f01 g15995 ( .a(n19360), .b(n19357), .o(n19784) );
no02f01 g15996 ( .a(n19784), .b(n19349), .o(n19785) );
no02f01 g15997 ( .a(n19785), .b(n19783), .o(n19786) );
ao12f01 g15998 ( .a(n19786), .b(n19781), .c(n19780), .o(n19787) );
in01f01 g15999 ( .a(n19787), .o(n19788) );
no02f01 g16000 ( .a(n18926), .b(n18913), .o(n19789) );
in01f01 g16001 ( .a(n19789), .o(n19790) );
na02f01 g16002 ( .a(n18926), .b(n18913), .o(n19791) );
na02f01 g16003 ( .a(n19791), .b(n19790), .o(n19792) );
in01f01 g16004 ( .a(n19348), .o(n19793) );
no03f01 g16005 ( .a(n19793), .b(n19347), .c(n19333), .o(n19794) );
in01f01 g16006 ( .a(n19333), .o(n19795) );
in01f01 g16007 ( .a(n19347), .o(n19796) );
ao12f01 g16008 ( .a(n19796), .b(n19348), .c(n19795), .o(n19797) );
no02f01 g16009 ( .a(n19797), .b(n19794), .o(n19798) );
in01f01 g16010 ( .a(n19798), .o(n19799) );
na02f01 g16011 ( .a(n19799), .b(n19792), .o(n19800) );
in01f01 g16012 ( .a(n19800), .o(n19801) );
no02f01 g16013 ( .a(n19799), .b(n19792), .o(n19802) );
ao12f01 g16014 ( .a(n19339), .b(n19342), .c(n19341), .o(n19803) );
no02f01 g16015 ( .a(n19343), .b(delay_add_ln22_unr5_stage3_stallmux_q_0_), .o(n19804) );
no02f01 g16016 ( .a(n19804), .b(n19803), .o(n19805) );
no02f01 g16017 ( .a(n19805), .b(n18918), .o(n19806) );
in01f01 g16018 ( .a(n19806), .o(n19807) );
in01f01 g16019 ( .a(n19344), .o(n19808) );
no03f01 g16020 ( .a(n19337), .b(n19336), .c(delay_add_ln22_unr5_stage3_stallmux_q_1_), .o(n19809) );
in01f01 g16021 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_1_), .o(n19810) );
no02f01 g16022 ( .a(n19338), .b(n19810), .o(n19811) );
no02f01 g16023 ( .a(n19811), .b(n19809), .o(n19812) );
no02f01 g16024 ( .a(n19812), .b(n19808), .o(n19813) );
na02f01 g16025 ( .a(n19812), .b(n19808), .o(n19814) );
in01f01 g16026 ( .a(n19814), .o(n19815) );
no02f01 g16027 ( .a(n19815), .b(n19813), .o(n19816) );
no02f01 g16028 ( .a(n19816), .b(n19807), .o(n19817) );
in01f01 g16029 ( .a(n19817), .o(n19818) );
in01f01 g16030 ( .a(n19816), .o(n19819) );
na02f01 g16031 ( .a(n18919), .b(n18145), .o(n19820) );
na02f01 g16032 ( .a(n18925), .b(n19820), .o(n19821) );
no02f01 g16033 ( .a(n18925), .b(n19820), .o(n19822) );
in01f01 g16034 ( .a(n19822), .o(n19823) );
na02f01 g16035 ( .a(n19823), .b(n19821), .o(n19824) );
oa12f01 g16036 ( .a(n19824), .b(n19819), .c(n19806), .o(n19825) );
ao12f01 g16037 ( .a(n19802), .b(n19825), .c(n19818), .o(n19826) );
na03f01 g16038 ( .a(n19786), .b(n19781), .c(n19780), .o(n19827) );
oa12f01 g16039 ( .a(n19827), .b(n19826), .c(n19801), .o(n19828) );
ao12f01 g16040 ( .a(n19778), .b(n19828), .c(n19788), .o(n19829) );
na02f01 g16041 ( .a(n19762), .b(n19756), .o(n19830) );
oa12f01 g16042 ( .a(n19830), .b(n19829), .c(n19776), .o(n19831) );
in01f01 g16043 ( .a(n19751), .o(n19832) );
no03f01 g16044 ( .a(n19832), .b(n19744), .c(n19742), .o(n19833) );
ao12f01 g16045 ( .a(n19833), .b(n19831), .c(n19764), .o(n19834) );
in01f01 g16046 ( .a(n19738), .o(n19835) );
no03f01 g16047 ( .a(n19835), .b(n19732), .c(n19730), .o(n19836) );
in01f01 g16048 ( .a(n19836), .o(n19837) );
oa12f01 g16049 ( .a(n19837), .b(n19834), .c(n19752), .o(n19838) );
in01f01 g16050 ( .a(n19727), .o(n19839) );
no03f01 g16051 ( .a(n19839), .b(n19720), .c(n19718), .o(n19840) );
ao12f01 g16052 ( .a(n19840), .b(n19838), .c(n19740), .o(n19841) );
no03f01 g16053 ( .a(n19841), .b(n19728), .c(n19716), .o(n19842) );
in01f01 g16054 ( .a(n19701), .o(n19843) );
no03f01 g16055 ( .a(n19843), .b(n19694), .c(n19693), .o(n19844) );
no03f01 g16056 ( .a(n19844), .b(n19842), .c(n19715), .o(n19845) );
na02f01 g16057 ( .a(n19688), .b(n19681), .o(n19846) );
oa12f01 g16058 ( .a(n19846), .b(n19845), .c(n19702), .o(n19847) );
in01f01 g16059 ( .a(n19024), .o(n19848) );
no02f01 g16060 ( .a(n19848), .b(n19010), .o(n19849) );
na02f01 g16061 ( .a(n19848), .b(n19010), .o(n19850) );
in01f01 g16062 ( .a(n19850), .o(n19851) );
no02f01 g16063 ( .a(n19851), .b(n19849), .o(n19852) );
na02f01 g16064 ( .a(n19453), .b(n19452), .o(n19853) );
in01f01 g16065 ( .a(n19853), .o(n19854) );
no02f01 g16066 ( .a(n19465), .b(n19462), .o(n19855) );
no02f01 g16067 ( .a(n19855), .b(n19854), .o(n19856) );
na02f01 g16068 ( .a(n19855), .b(n19854), .o(n19857) );
in01f01 g16069 ( .a(n19857), .o(n19858) );
no02f01 g16070 ( .a(n19858), .b(n19856), .o(n19859) );
na02f01 g16071 ( .a(n19859), .b(n19852), .o(n19860) );
in01f01 g16072 ( .a(n19860), .o(n19861) );
ao12f01 g16073 ( .a(n19861), .b(n19847), .c(n19690), .o(n19862) );
oa12f01 g16074 ( .a(n19674), .b(n19665), .c(n19662), .o(n19863) );
in01f01 g16075 ( .a(n19859), .o(n19864) );
oa12f01 g16076 ( .a(n19864), .b(n19851), .c(n19849), .o(n19865) );
na02f01 g16077 ( .a(n19865), .b(n19863), .o(n19866) );
oa12f01 g16078 ( .a(n19676), .b(n19866), .c(n19862), .o(n19867) );
ao12f01 g16079 ( .a(n19640), .b(n19026), .c(n19656), .o(n19868) );
in01f01 g16080 ( .a(n19868), .o(n19869) );
no02f01 g16081 ( .a(n19869), .b(n19559), .o(n19870) );
no02f01 g16082 ( .a(n19868), .b(n19034), .o(n19871) );
no02f01 g16083 ( .a(n19871), .b(n19870), .o(n19872) );
na02f01 g16084 ( .a(n19467), .b(n19311), .o(n19873) );
in01f01 g16085 ( .a(n19873), .o(n19874) );
in01f01 g16086 ( .a(n19468), .o(n19875) );
no02f01 g16087 ( .a(n19875), .b(n19300), .o(n19876) );
no02f01 g16088 ( .a(n19876), .b(n19874), .o(n19877) );
in01f01 g16089 ( .a(n19877), .o(n19878) );
na02f01 g16090 ( .a(n19876), .b(n19874), .o(n19879) );
na02f01 g16091 ( .a(n19879), .b(n19878), .o(n19880) );
in01f01 g16092 ( .a(n19880), .o(n19881) );
na02f01 g16093 ( .a(n19881), .b(n19872), .o(n19882) );
in01f01 g16094 ( .a(n19882), .o(n19883) );
oa12f01 g16095 ( .a(n19653), .b(n19645), .c(n19643), .o(n19884) );
in01f01 g16096 ( .a(n19884), .o(n19885) );
no02f01 g16097 ( .a(n19881), .b(n19872), .o(n19886) );
no02f01 g16098 ( .a(n19886), .b(n19885), .o(n19887) );
oa12f01 g16099 ( .a(n19887), .b(n19883), .c(n19867), .o(n19888) );
no02f01 g16100 ( .a(n19051), .b(n19563), .o(n19889) );
no02f01 g16101 ( .a(n19050), .b(n19043), .o(n19890) );
no02f01 g16102 ( .a(n19890), .b(n19889), .o(n19891) );
in01f01 g16103 ( .a(n19891), .o(n19892) );
na02f01 g16104 ( .a(n19471), .b(n19291), .o(n19893) );
no02f01 g16105 ( .a(n19473), .b(n19281), .o(n19894) );
in01f01 g16106 ( .a(n19894), .o(n19895) );
no02f01 g16107 ( .a(n19895), .b(n19893), .o(n19896) );
na02f01 g16108 ( .a(n19895), .b(n19893), .o(n19897) );
in01f01 g16109 ( .a(n19897), .o(n19898) );
no02f01 g16110 ( .a(n19898), .b(n19896), .o(n19899) );
in01f01 g16111 ( .a(n19899), .o(n19900) );
no02f01 g16112 ( .a(n19900), .b(n19892), .o(n19901) );
in01f01 g16113 ( .a(n19901), .o(n19902) );
no02f01 g16114 ( .a(n19050), .b(n18145), .o(n19903) );
no02f01 g16115 ( .a(n19903), .b(n19052), .o(n19904) );
na02f01 g16116 ( .a(n19904), .b(n19059), .o(n19905) );
in01f01 g16117 ( .a(n19903), .o(n19906) );
na02f01 g16118 ( .a(n19906), .b(n19564), .o(n19907) );
na02f01 g16119 ( .a(n19907), .b(n19565), .o(n19908) );
no02f01 g16120 ( .a(n19474), .b(n19281), .o(n19909) );
in01f01 g16121 ( .a(n19475), .o(n19910) );
no02f01 g16122 ( .a(n19910), .b(n19271), .o(n19911) );
no02f01 g16123 ( .a(n19911), .b(n19909), .o(n19912) );
na02f01 g16124 ( .a(n19911), .b(n19909), .o(n19913) );
in01f01 g16125 ( .a(n19913), .o(n19914) );
no02f01 g16126 ( .a(n19914), .b(n19912), .o(n19915) );
na03f01 g16127 ( .a(n19915), .b(n19908), .c(n19905), .o(n19916) );
na04f01 g16128 ( .a(n19916), .b(n19902), .c(n19888), .d(n19655), .o(n19917) );
ao12f01 g16129 ( .a(n19915), .b(n19908), .c(n19905), .o(n19918) );
no02f01 g16130 ( .a(n19899), .b(n19891), .o(n19919) );
oa12f01 g16131 ( .a(n19916), .b(n19919), .c(n19918), .o(n19920) );
na02f01 g16132 ( .a(n19629), .b(n19068), .o(n19921) );
na02f01 g16133 ( .a(n19627), .b(n19067), .o(n19922) );
na02f01 g16134 ( .a(n19922), .b(n19921), .o(n19923) );
in01f01 g16135 ( .a(n19638), .o(n19924) );
no02f01 g16136 ( .a(n19924), .b(n19923), .o(n19925) );
ao12f01 g16137 ( .a(n19925), .b(n19920), .c(n19917), .o(n19926) );
no02f01 g16138 ( .a(n19616), .b(n19074), .o(n19927) );
no02f01 g16139 ( .a(n19614), .b(n19077), .o(n19928) );
no02f01 g16140 ( .a(n19928), .b(n19927), .o(n19929) );
in01f01 g16141 ( .a(n19622), .o(n19930) );
no02f01 g16142 ( .a(n19623), .b(n19930), .o(n19931) );
no02f01 g16143 ( .a(n19931), .b(n19929), .o(n19932) );
no03f01 g16144 ( .a(n19932), .b(n19926), .c(n19639), .o(n19933) );
no03f01 g16145 ( .a(n19610), .b(n19603), .c(n19599), .o(n19934) );
no04f01 g16146 ( .a(n19934), .b(n19933), .c(n19626), .d(n19595), .o(n19935) );
oa12f01 g16147 ( .a(n19585), .b(n19096), .c(n18145), .o(n19936) );
no02f01 g16148 ( .a(n19936), .b(n19572), .o(n19937) );
no02f01 g16149 ( .a(n18882), .b(n18145), .o(n19938) );
no02f01 g16150 ( .a(n19938), .b(n18883), .o(n19939) );
na02f01 g16151 ( .a(n19939), .b(n19937), .o(n19940) );
na02f01 g16152 ( .a(n19110), .b(n19097), .o(n19941) );
na02f01 g16153 ( .a(n19103), .b(n19554), .o(n19942) );
na02f01 g16154 ( .a(n19942), .b(n19941), .o(n19943) );
na02f01 g16155 ( .a(n19486), .b(n19234), .o(n19944) );
no02f01 g16156 ( .a(n19488), .b(n19224), .o(n19945) );
in01f01 g16157 ( .a(n19945), .o(n19946) );
no02f01 g16158 ( .a(n19946), .b(n19944), .o(n19947) );
in01f01 g16159 ( .a(n19944), .o(n19948) );
no02f01 g16160 ( .a(n19945), .b(n19948), .o(n19949) );
no02f01 g16161 ( .a(n19949), .b(n19947), .o(n19950) );
na03f01 g16162 ( .a(n19950), .b(n19943), .c(n19940), .o(n19951) );
oa12f01 g16163 ( .a(n19951), .b(n19935), .c(n19613), .o(n19952) );
na02f01 g16164 ( .a(n19104), .b(n19555), .o(n19953) );
na03f01 g16165 ( .a(n19110), .b(n19103), .c(n19097), .o(n19954) );
na03f01 g16166 ( .a(n19954), .b(n19953), .c(n19554), .o(n19955) );
no02f01 g16167 ( .a(n18896), .b(n18145), .o(n19956) );
no02f01 g16168 ( .a(n19956), .b(n18897), .o(n19957) );
no03f01 g16169 ( .a(n19936), .b(n19938), .c(n19572), .o(n19958) );
oa12f01 g16170 ( .a(n19957), .b(n19958), .c(n18883), .o(n19959) );
in01f01 g16171 ( .a(n19490), .o(n19960) );
no02f01 g16172 ( .a(n19960), .b(n19214), .o(n19961) );
no02f01 g16173 ( .a(n19944), .b(n19224), .o(n19962) );
no03f01 g16174 ( .a(n19962), .b(n19961), .c(n19488), .o(n19963) );
oa12f01 g16175 ( .a(n19961), .b(n19962), .c(n19488), .o(n19964) );
in01f01 g16176 ( .a(n19964), .o(n19965) );
no02f01 g16177 ( .a(n19965), .b(n19963), .o(n19966) );
ao12f01 g16178 ( .a(n19966), .b(n19959), .c(n19955), .o(n19967) );
ao12f01 g16179 ( .a(n19950), .b(n19943), .c(n19940), .o(n19968) );
no02f01 g16180 ( .a(n19968), .b(n19967), .o(n19969) );
no03f01 g16181 ( .a(n19958), .b(n19957), .c(n18883), .o(n19970) );
ao12f01 g16182 ( .a(n19953), .b(n19954), .c(n19554), .o(n19971) );
in01f01 g16183 ( .a(n19966), .o(n19972) );
no03f01 g16184 ( .a(n19972), .b(n19971), .c(n19970), .o(n19973) );
ao12f01 g16185 ( .a(n19973), .b(n19969), .c(n19952), .o(n19974) );
na03f01 g16186 ( .a(n19583), .b(n19576), .c(n19553), .o(n19975) );
ao12f01 g16187 ( .a(n19584), .b(n19975), .c(n19974), .o(n19976) );
oa12f01 g16188 ( .a(n19551), .b(n19117), .c(n19113), .o(n19977) );
ao12f01 g16189 ( .a(n19552), .b(n19977), .c(n19976), .o(n19978) );
ao12f01 g16190 ( .a(n19532), .b(n19978), .c(n19545), .o(n19979) );
no02f01 g16191 ( .a(n19540), .b(n19507), .o(n19980) );
ao12f01 g16192 ( .a(n19980), .b(n19497), .c(n19196), .o(n19981) );
na03f01 g16193 ( .a(n19980), .b(n19497), .c(n19196), .o(n19982) );
in01f01 g16194 ( .a(n19982), .o(n19983) );
no02f01 g16195 ( .a(n19983), .b(n19981), .o(n19984) );
no02f01 g16196 ( .a(n19984), .b(n19118), .o(n19985) );
no03f01 g16197 ( .a(n19985), .b(n19978), .c(n19545), .o(n19986) );
na02f01 g16198 ( .a(n19984), .b(n19118), .o(n19987) );
in01f01 g16199 ( .a(n19987), .o(n19988) );
na02f01 g16200 ( .a(n19500), .b(delay_add_ln22_unr5_stage3_stallmux_q_29_), .o(n19989) );
in01f01 g16201 ( .a(n19989), .o(n19990) );
no02f01 g16202 ( .a(n19990), .b(n19511), .o(n19991) );
in01f01 g16203 ( .a(n19991), .o(n19992) );
ao12f01 g16204 ( .a(n19504), .b(n19497), .c(n19196), .o(n19993) );
in01f01 g16205 ( .a(n19509), .o(n19994) );
no02f01 g16206 ( .a(n19994), .b(n19993), .o(n19995) );
no02f01 g16207 ( .a(n19512), .b(n19995), .o(n19996) );
na02f01 g16208 ( .a(n19500), .b(delay_add_ln22_unr5_stage3_stallmux_q_28_), .o(n19997) );
in01f01 g16209 ( .a(n19997), .o(n19998) );
no03f01 g16210 ( .a(n19998), .b(n19996), .c(n19992), .o(n19999) );
in01f01 g16211 ( .a(n19999), .o(n20000) );
oa12f01 g16212 ( .a(n19992), .b(n19998), .c(n19996), .o(n20001) );
na02f01 g16213 ( .a(n20001), .b(n20000), .o(n20002) );
no02f01 g16214 ( .a(n19998), .b(n19512), .o(n20003) );
in01f01 g16215 ( .a(n20003), .o(n20004) );
no03f01 g16216 ( .a(n20004), .b(n19994), .c(n19993), .o(n20005) );
in01f01 g16217 ( .a(n20005), .o(n20006) );
oa12f01 g16218 ( .a(n20004), .b(n19994), .c(n19993), .o(n20007) );
na02f01 g16219 ( .a(n20007), .b(n20006), .o(n20008) );
ao12f01 g16220 ( .a(n19532), .b(n20008), .c(n20002), .o(n20009) );
no04f01 g16221 ( .a(n20009), .b(n19988), .c(n19986), .d(n19979), .o(n20010) );
in01f01 g16222 ( .a(n19513), .o(n20011) );
no02f01 g16223 ( .a(n20011), .b(n19995), .o(n20012) );
no02f01 g16224 ( .a(n19517), .b(n19515), .o(n20013) );
in01f01 g16225 ( .a(n20013), .o(n20014) );
no03f01 g16226 ( .a(n20014), .b(n19519), .c(n20012), .o(n20015) );
in01f01 g16227 ( .a(n20015), .o(n20016) );
oa12f01 g16228 ( .a(n20014), .b(n19519), .c(n20012), .o(n20017) );
na02f01 g16229 ( .a(n20017), .b(n20016), .o(n20018) );
in01f01 g16230 ( .a(n19544), .o(n20019) );
no02f01 g16231 ( .a(n20019), .b(n19542), .o(n20020) );
in01f01 g16232 ( .a(n19552), .o(n20021) );
no02f01 g16233 ( .a(n19575), .b(n19114), .o(n20022) );
no02f01 g16234 ( .a(n19112), .b(n18868), .o(n20023) );
in01f01 g16235 ( .a(n19580), .o(n20024) );
na02f01 g16236 ( .a(n19581), .b(n20024), .o(n20025) );
oa12f01 g16237 ( .a(n20025), .b(n20023), .c(n20022), .o(n20026) );
oa12f01 g16238 ( .a(n19106), .b(n19109), .c(n19091), .o(n20027) );
na03f01 g16239 ( .a(n19585), .b(n19096), .c(n19571), .o(n20028) );
in01f01 g16240 ( .a(n19591), .o(n20029) );
no02f01 g16241 ( .a(n19592), .b(n20029), .o(n20030) );
na03f01 g16242 ( .a(n20030), .b(n20028), .c(n20027), .o(n20031) );
na02f01 g16243 ( .a(n19602), .b(n19600), .o(n20032) );
na02f01 g16244 ( .a(n19598), .b(n19596), .o(n20033) );
in01f01 g16245 ( .a(n19609), .o(n20034) );
no02f01 g16246 ( .a(n20034), .b(n19607), .o(n20035) );
ao12f01 g16247 ( .a(n20035), .b(n20033), .c(n20032), .o(n20036) );
ao12f01 g16248 ( .a(n20030), .b(n20028), .c(n20027), .o(n20037) );
oa12f01 g16249 ( .a(n20031), .b(n20037), .c(n20036), .o(n20038) );
na02f01 g16250 ( .a(n19931), .b(n19929), .o(n20039) );
na02f01 g16251 ( .a(n19924), .b(n19923), .o(n20040) );
in01f01 g16252 ( .a(n19702), .o(n20041) );
in01f01 g16253 ( .a(n19716), .o(n20042) );
in01f01 g16254 ( .a(n19728), .o(n20043) );
in01f01 g16255 ( .a(n19752), .o(n20044) );
in01f01 g16256 ( .a(n19776), .o(n20045) );
in01f01 g16257 ( .a(n19778), .o(n20046) );
in01f01 g16258 ( .a(n19821), .o(n20047) );
no02f01 g16259 ( .a(n19822), .b(n20047), .o(n20048) );
ao12f01 g16260 ( .a(n20048), .b(n19816), .c(n19807), .o(n20049) );
oa22f01 g16261 ( .a(n20049), .b(n19817), .c(n19799), .d(n19792), .o(n20050) );
in01f01 g16262 ( .a(n19827), .o(n20051) );
ao12f01 g16263 ( .a(n20051), .b(n20050), .c(n19800), .o(n20052) );
oa12f01 g16264 ( .a(n20046), .b(n20052), .c(n19787), .o(n20053) );
in01f01 g16265 ( .a(n19830), .o(n20054) );
ao12f01 g16266 ( .a(n20054), .b(n20053), .c(n20045), .o(n20055) );
in01f01 g16267 ( .a(n19833), .o(n20056) );
oa12f01 g16268 ( .a(n20056), .b(n20055), .c(n19763), .o(n20057) );
ao12f01 g16269 ( .a(n19836), .b(n20057), .c(n20044), .o(n20058) );
in01f01 g16270 ( .a(n19840), .o(n20059) );
oa12f01 g16271 ( .a(n20059), .b(n20058), .c(n19739), .o(n20060) );
na03f01 g16272 ( .a(n20060), .b(n20043), .c(n20042), .o(n20061) );
in01f01 g16273 ( .a(n19844), .o(n20062) );
na03f01 g16274 ( .a(n20062), .b(n20061), .c(n19714), .o(n20063) );
in01f01 g16275 ( .a(n19846), .o(n20064) );
ao12f01 g16276 ( .a(n20064), .b(n20063), .c(n20041), .o(n20065) );
oa12f01 g16277 ( .a(n19860), .b(n20065), .c(n19689), .o(n20066) );
in01f01 g16278 ( .a(n19866), .o(n20067) );
ao12f01 g16279 ( .a(n19675), .b(n20067), .c(n20066), .o(n20068) );
in01f01 g16280 ( .a(n19886), .o(n20069) );
na02f01 g16281 ( .a(n20069), .b(n19884), .o(n20070) );
ao12f01 g16282 ( .a(n20070), .b(n19882), .c(n20068), .o(n20071) );
no02f01 g16283 ( .a(n19907), .b(n19565), .o(n20072) );
no02f01 g16284 ( .a(n19904), .b(n19059), .o(n20073) );
in01f01 g16285 ( .a(n19915), .o(n20074) );
no03f01 g16286 ( .a(n20074), .b(n20073), .c(n20072), .o(n20075) );
no04f01 g16287 ( .a(n20075), .b(n19901), .c(n20071), .d(n19654), .o(n20076) );
oa12f01 g16288 ( .a(n20074), .b(n20073), .c(n20072), .o(n20077) );
in01f01 g16289 ( .a(n19919), .o(n20078) );
ao12f01 g16290 ( .a(n20075), .b(n20078), .c(n20077), .o(n20079) );
na02f01 g16291 ( .a(n19638), .b(n19631), .o(n20080) );
oa12f01 g16292 ( .a(n20080), .b(n20079), .c(n20076), .o(n20081) );
na02f01 g16293 ( .a(n19625), .b(n19618), .o(n20082) );
na03f01 g16294 ( .a(n20082), .b(n20081), .c(n20040), .o(n20083) );
na03f01 g16295 ( .a(n20035), .b(n20033), .c(n20032), .o(n20084) );
na04f01 g16296 ( .a(n20084), .b(n20083), .c(n20039), .d(n20031), .o(n20085) );
no02f01 g16297 ( .a(n19942), .b(n19941), .o(n20086) );
no02f01 g16298 ( .a(n19939), .b(n19937), .o(n20087) );
in01f01 g16299 ( .a(n19950), .o(n20088) );
no03f01 g16300 ( .a(n20088), .b(n20087), .c(n20086), .o(n20089) );
ao12f01 g16301 ( .a(n20089), .b(n20085), .c(n20038), .o(n20090) );
oa12f01 g16302 ( .a(n19972), .b(n19971), .c(n19970), .o(n20091) );
oa12f01 g16303 ( .a(n20088), .b(n20087), .c(n20086), .o(n20092) );
na02f01 g16304 ( .a(n20092), .b(n20091), .o(n20093) );
na03f01 g16305 ( .a(n19966), .b(n19959), .c(n19955), .o(n20094) );
oa12f01 g16306 ( .a(n20094), .b(n20093), .c(n20090), .o(n20095) );
no03f01 g16307 ( .a(n20025), .b(n20023), .c(n20022), .o(n20096) );
oa12f01 g16308 ( .a(n20026), .b(n20096), .c(n20095), .o(n20097) );
in01f01 g16309 ( .a(n19977), .o(n20098) );
oa12f01 g16310 ( .a(n20021), .b(n20098), .c(n20097), .o(n20099) );
oa12f01 g16311 ( .a(n19118), .b(n20099), .c(n20020), .o(n20100) );
in01f01 g16312 ( .a(n19985), .o(n20101) );
na03f01 g16313 ( .a(n20101), .b(n20099), .c(n20020), .o(n20102) );
in01f01 g16314 ( .a(n20009), .o(n20103) );
na04f01 g16315 ( .a(n20103), .b(n19987), .c(n20102), .d(n20100), .o(n20104) );
no02f01 g16316 ( .a(n19519), .b(n20012), .o(n20105) );
no02f01 g16317 ( .a(n20013), .b(n20105), .o(n20106) );
no02f01 g16318 ( .a(n20106), .b(n20015), .o(n20107) );
no02f01 g16319 ( .a(n19998), .b(n19996), .o(n20108) );
no02f01 g16320 ( .a(n20108), .b(n19991), .o(n20109) );
no02f01 g16321 ( .a(n20109), .b(n19999), .o(n20110) );
in01f01 g16322 ( .a(n20007), .o(n20111) );
no02f01 g16323 ( .a(n20111), .b(n20005), .o(n20112) );
ao12f01 g16324 ( .a(n19118), .b(n20112), .c(n20110), .o(n20113) );
in01f01 g16325 ( .a(n20113), .o(n20114) );
na03f01 g16326 ( .a(n20114), .b(n20107), .c(n20104), .o(n20115) );
ao22f01 g16327 ( .a(n20115), .b(n19532), .c(n20018), .d(n20010), .o(n20116) );
na02f01 g16328 ( .a(n20116), .b(n19536), .o(n20117) );
in01f01 g16329 ( .a(n19536), .o(n20118) );
no03f01 g16330 ( .a(n20113), .b(n20018), .c(n20010), .o(n20119) );
oa22f01 g16331 ( .a(n20119), .b(n19118), .c(n20107), .d(n20104), .o(n20120) );
na02f01 g16332 ( .a(n20120), .b(n20118), .o(n20121) );
ao12f01 g16333 ( .a(n18460), .b(n20121), .c(n20117), .o(n20122) );
ao12f01 g16334 ( .a(n18459), .b(n20121), .c(n20117), .o(n20123) );
no02f01 g16335 ( .a(n20123), .b(n20122), .o(n20124) );
no02f01 g16336 ( .a(n20110), .b(n19118), .o(n20125) );
no02f01 g16337 ( .a(n20002), .b(n19532), .o(n20126) );
no02f01 g16338 ( .a(n20126), .b(n20125), .o(n20127) );
in01f01 g16339 ( .a(n20127), .o(n20128) );
no02f01 g16340 ( .a(n20112), .b(n19118), .o(n20129) );
na02f01 g16341 ( .a(n20112), .b(n19118), .o(n20130) );
in01f01 g16342 ( .a(n20130), .o(n20131) );
no04f01 g16343 ( .a(n20131), .b(n19988), .c(n19986), .d(n19979), .o(n20132) );
no03f01 g16344 ( .a(n20132), .b(n20129), .c(n20128), .o(n20133) );
in01f01 g16345 ( .a(n20129), .o(n20134) );
na04f01 g16346 ( .a(n20130), .b(n19987), .c(n20102), .d(n20100), .o(n20135) );
ao12f01 g16347 ( .a(n20127), .b(n20135), .c(n20134), .o(n20136) );
oa12f01 g16348 ( .a(n18460), .b(n20136), .c(n20133), .o(n20137) );
no02f01 g16349 ( .a(n20093), .b(n20090), .o(n20138) );
no03f01 g16350 ( .a(n20096), .b(n19973), .c(n20138), .o(n20139) );
no03f01 g16351 ( .a(n20098), .b(n20139), .c(n19584), .o(n20140) );
oa12f01 g16352 ( .a(n20101), .b(n20140), .c(n19552), .o(n20141) );
oa12f01 g16353 ( .a(n19987), .b(n20141), .c(n19545), .o(n20142) );
no02f01 g16354 ( .a(n20131), .b(n20129), .o(n20143) );
oa12f01 g16355 ( .a(n20143), .b(n20142), .c(n19979), .o(n20144) );
na02f01 g16356 ( .a(n19969), .b(n19952), .o(n20145) );
na03f01 g16357 ( .a(n19975), .b(n20094), .c(n20145), .o(n20146) );
na03f01 g16358 ( .a(n19977), .b(n20146), .c(n20026), .o(n20147) );
ao12f01 g16359 ( .a(n19985), .b(n20147), .c(n20021), .o(n20148) );
ao12f01 g16360 ( .a(n19988), .b(n20148), .c(n20020), .o(n20149) );
in01f01 g16361 ( .a(n20143), .o(n20150) );
na03f01 g16362 ( .a(n20150), .b(n20149), .c(n20100), .o(n20151) );
na02f01 g16363 ( .a(n20151), .b(n20144), .o(n20152) );
no02f01 g16364 ( .a(n19545), .b(n19532), .o(n20153) );
no02f01 g16365 ( .a(n20020), .b(n19118), .o(n20154) );
no02f01 g16366 ( .a(n20154), .b(n20153), .o(n20155) );
in01f01 g16367 ( .a(n20155), .o(n20156) );
ao12f01 g16368 ( .a(n20156), .b(n19987), .c(n20141), .o(n20157) );
no03f01 g16369 ( .a(n20155), .b(n19988), .c(n20148), .o(n20158) );
no02f01 g16370 ( .a(n20158), .b(n20157), .o(n20159) );
no02f01 g16371 ( .a(n20096), .b(n19584), .o(n20160) );
no02f01 g16372 ( .a(n20160), .b(n20095), .o(n20161) );
na02f01 g16373 ( .a(n19975), .b(n20026), .o(n20162) );
no02f01 g16374 ( .a(n20162), .b(n19974), .o(n20163) );
no02f01 g16375 ( .a(n20163), .b(n20161), .o(n20164) );
no02f01 g16376 ( .a(n20164), .b(n18459), .o(n20165) );
no02f01 g16377 ( .a(n19973), .b(n19967), .o(n20166) );
no03f01 g16378 ( .a(n19968), .b(n19935), .c(n19613), .o(n20167) );
no03f01 g16379 ( .a(n20167), .b(n20166), .c(n20089), .o(n20168) );
na02f01 g16380 ( .a(n20094), .b(n20091), .o(n20169) );
in01f01 g16381 ( .a(n20167), .o(n20170) );
ao12f01 g16382 ( .a(n20169), .b(n20170), .c(n19951), .o(n20171) );
no02f01 g16383 ( .a(n20171), .b(n20168), .o(n20172) );
na03f01 g16384 ( .a(n20084), .b(n20083), .c(n20039), .o(n20173) );
no02f01 g16385 ( .a(n20037), .b(n19595), .o(n20174) );
ao12f01 g16386 ( .a(n20174), .b(n20173), .c(n19611), .o(n20175) );
no03f01 g16387 ( .a(n19934), .b(n19933), .c(n19626), .o(n20176) );
in01f01 g16388 ( .a(n20174), .o(n20177) );
no03f01 g16389 ( .a(n20177), .b(n20176), .c(n20036), .o(n20178) );
no02f01 g16390 ( .a(n20178), .b(n20175), .o(n20179) );
no02f01 g16391 ( .a(n20179), .b(n18459), .o(n20180) );
na02f01 g16392 ( .a(n20082), .b(n20039), .o(n20181) );
no03f01 g16393 ( .a(n20181), .b(n19926), .c(n19639), .o(n20182) );
no02f01 g16394 ( .a(n19932), .b(n19626), .o(n20183) );
ao12f01 g16395 ( .a(n20183), .b(n20081), .c(n20040), .o(n20184) );
no02f01 g16396 ( .a(n20184), .b(n20182), .o(n20185) );
no02f01 g16397 ( .a(n20185), .b(n18459), .o(n20186) );
in01f01 g16398 ( .a(n20186), .o(n20187) );
na02f01 g16399 ( .a(n20080), .b(n20040), .o(n20188) );
no03f01 g16400 ( .a(n20188), .b(n20079), .c(n20076), .o(n20189) );
no02f01 g16401 ( .a(n19925), .b(n19639), .o(n20190) );
ao12f01 g16402 ( .a(n20190), .b(n19920), .c(n19917), .o(n20191) );
oa12f01 g16403 ( .a(n18460), .b(n20191), .c(n20189), .o(n20192) );
ao12f01 g16404 ( .a(n19883), .b(n20069), .c(n19867), .o(n20193) );
no02f01 g16405 ( .a(n19885), .b(n19654), .o(n20194) );
in01f01 g16406 ( .a(n20194), .o(n20195) );
no02f01 g16407 ( .a(n20195), .b(n20193), .o(n20196) );
oa12f01 g16408 ( .a(n19882), .b(n19886), .c(n20068), .o(n20197) );
no02f01 g16409 ( .a(n20194), .b(n20197), .o(n20198) );
no02f01 g16410 ( .a(n20198), .b(n20196), .o(n20199) );
no02f01 g16411 ( .a(n20199), .b(n18459), .o(n20200) );
no02f01 g16412 ( .a(n20199), .b(n18460), .o(n20201) );
no02f01 g16413 ( .a(n20058), .b(n19739), .o(n20202) );
no02f01 g16414 ( .a(n19840), .b(n19728), .o(n20203) );
no02f01 g16415 ( .a(n20203), .b(n20202), .o(n20204) );
na02f01 g16416 ( .a(n20203), .b(n20202), .o(n20205) );
in01f01 g16417 ( .a(n20205), .o(n20206) );
no02f01 g16418 ( .a(n20206), .b(n20204), .o(n20207) );
no02f01 g16419 ( .a(n19841), .b(n19728), .o(n20208) );
in01f01 g16420 ( .a(n20208), .o(n20209) );
na02f01 g16421 ( .a(n20042), .b(n19714), .o(n20210) );
no02f01 g16422 ( .a(n20210), .b(n20209), .o(n20211) );
na02f01 g16423 ( .a(n20210), .b(n20209), .o(n20212) );
in01f01 g16424 ( .a(n20212), .o(n20213) );
no02f01 g16425 ( .a(n20213), .b(n20211), .o(n20214) );
ao12f01 g16426 ( .a(n18459), .b(n20214), .c(n20207), .o(n20215) );
no02f01 g16427 ( .a(n19842), .b(n19715), .o(n20216) );
no02f01 g16428 ( .a(n19844), .b(n19702), .o(n20217) );
in01f01 g16429 ( .a(n20217), .o(n20218) );
no02f01 g16430 ( .a(n20218), .b(n20216), .o(n20219) );
no03f01 g16431 ( .a(n20217), .b(n19842), .c(n19715), .o(n20220) );
no02f01 g16432 ( .a(n20220), .b(n20219), .o(n20221) );
no02f01 g16433 ( .a(n20221), .b(n18459), .o(n20222) );
no02f01 g16434 ( .a(n20222), .b(n20215), .o(n20223) );
na02f01 g16435 ( .a(n20063), .b(n20041), .o(n20224) );
na02f01 g16436 ( .a(n19846), .b(n19690), .o(n20225) );
no02f01 g16437 ( .a(n20225), .b(n20224), .o(n20226) );
no02f01 g16438 ( .a(n19845), .b(n19702), .o(n20227) );
no02f01 g16439 ( .a(n20064), .b(n19689), .o(n20228) );
no02f01 g16440 ( .a(n20228), .b(n20227), .o(n20229) );
oa12f01 g16441 ( .a(n18460), .b(n20229), .c(n20226), .o(n20230) );
na02f01 g16442 ( .a(n20230), .b(n20223), .o(n20231) );
na02f01 g16443 ( .a(n19865), .b(n19860), .o(n20232) );
no03f01 g16444 ( .a(n20232), .b(n20065), .c(n19689), .o(n20233) );
in01f01 g16445 ( .a(n20232), .o(n20234) );
ao12f01 g16446 ( .a(n20234), .b(n19847), .c(n19690), .o(n20235) );
no02f01 g16447 ( .a(n20235), .b(n20233), .o(n20236) );
no02f01 g16448 ( .a(n20236), .b(n18459), .o(n20237) );
no02f01 g16449 ( .a(n20237), .b(n20231), .o(n20238) );
in01f01 g16450 ( .a(n19863), .o(n20239) );
no02f01 g16451 ( .a(n20239), .b(n19675), .o(n20240) );
in01f01 g16452 ( .a(n19865), .o(n20241) );
no03f01 g16453 ( .a(n20241), .b(n20065), .c(n19689), .o(n20242) );
no03f01 g16454 ( .a(n20242), .b(n20240), .c(n19861), .o(n20243) );
na02f01 g16455 ( .a(n19863), .b(n19676), .o(n20244) );
na03f01 g16456 ( .a(n19865), .b(n19847), .c(n19690), .o(n20245) );
ao12f01 g16457 ( .a(n20244), .b(n20245), .c(n19860), .o(n20246) );
no02f01 g16458 ( .a(n20246), .b(n20243), .o(n20247) );
oa12f01 g16459 ( .a(n20238), .b(n20247), .c(n18459), .o(n20248) );
ao12f01 g16460 ( .a(n18460), .b(n20247), .c(n20236), .o(n20249) );
in01f01 g16461 ( .a(n20249), .o(n20250) );
na02f01 g16462 ( .a(n20069), .b(n19882), .o(n20251) );
no02f01 g16463 ( .a(n20251), .b(n20068), .o(n20252) );
no02f01 g16464 ( .a(n19886), .b(n19883), .o(n20253) );
no02f01 g16465 ( .a(n20253), .b(n19867), .o(n20254) );
no02f01 g16466 ( .a(n20254), .b(n20252), .o(n20255) );
no02f01 g16467 ( .a(n20255), .b(n18459), .o(n20256) );
ao12f01 g16468 ( .a(n20256), .b(n20250), .c(n20248), .o(n20257) );
no02f01 g16469 ( .a(n20255), .b(n18460), .o(n20258) );
no03f01 g16470 ( .a(n20258), .b(n20257), .c(n20201), .o(n20259) );
na02f01 g16471 ( .a(n19888), .b(n19655), .o(n20260) );
no02f01 g16472 ( .a(n19919), .b(n19901), .o(n20261) );
no02f01 g16473 ( .a(n20261), .b(n20260), .o(n20262) );
no02f01 g16474 ( .a(n20071), .b(n19654), .o(n20263) );
in01f01 g16475 ( .a(n20261), .o(n20264) );
no02f01 g16476 ( .a(n20264), .b(n20263), .o(n20265) );
no02f01 g16477 ( .a(n20265), .b(n20262), .o(n20266) );
no02f01 g16478 ( .a(n20266), .b(n18459), .o(n20267) );
no03f01 g16479 ( .a(n20267), .b(n20259), .c(n20200), .o(n20268) );
no02f01 g16480 ( .a(n19901), .b(n20260), .o(n20269) );
no02f01 g16481 ( .a(n19918), .b(n20075), .o(n20270) );
in01f01 g16482 ( .a(n20270), .o(n20271) );
no03f01 g16483 ( .a(n20271), .b(n19919), .c(n20269), .o(n20272) );
ao12f01 g16484 ( .a(n19919), .b(n19902), .c(n20263), .o(n20273) );
no02f01 g16485 ( .a(n20273), .b(n20270), .o(n20274) );
oa12f01 g16486 ( .a(n18460), .b(n20274), .c(n20272), .o(n20275) );
na03f01 g16487 ( .a(n20275), .b(n20268), .c(n20192), .o(n20276) );
oa12f01 g16488 ( .a(n18459), .b(n20274), .c(n20272), .o(n20277) );
in01f01 g16489 ( .a(n20277), .o(n20278) );
no02f01 g16490 ( .a(n20266), .b(n18460), .o(n20279) );
na03f01 g16491 ( .a(n20190), .b(n19920), .c(n19917), .o(n20280) );
oa12f01 g16492 ( .a(n20188), .b(n20079), .c(n20076), .o(n20281) );
ao12f01 g16493 ( .a(n18460), .b(n20281), .c(n20280), .o(n20282) );
no03f01 g16494 ( .a(n20282), .b(n20279), .c(n20278), .o(n20283) );
oa12f01 g16495 ( .a(n18459), .b(n20184), .c(n20182), .o(n20284) );
na03f01 g16496 ( .a(n20284), .b(n20283), .c(n20276), .o(n20285) );
no02f01 g16497 ( .a(n19934), .b(n20036), .o(n20286) );
oa12f01 g16498 ( .a(n20286), .b(n19933), .c(n19626), .o(n20287) );
na02f01 g16499 ( .a(n20084), .b(n19611), .o(n20288) );
na03f01 g16500 ( .a(n20288), .b(n20083), .c(n20039), .o(n20289) );
na02f01 g16501 ( .a(n20289), .b(n20287), .o(n20290) );
na02f01 g16502 ( .a(n20290), .b(n18460), .o(n20291) );
na03f01 g16503 ( .a(n20291), .b(n20285), .c(n20187), .o(n20292) );
na04f01 g16504 ( .a(n20092), .b(n19951), .c(n20085), .d(n20038), .o(n20293) );
oa22f01 g16505 ( .a(n19968), .b(n20089), .c(n19935), .d(n19613), .o(n20294) );
ao12f01 g16506 ( .a(n18459), .b(n20294), .c(n20293), .o(n20295) );
no03f01 g16507 ( .a(n20295), .b(n20292), .c(n20180), .o(n20296) );
oa12f01 g16508 ( .a(n20296), .b(n20172), .c(n18459), .o(n20297) );
na03f01 g16509 ( .a(n20170), .b(n20169), .c(n19951), .o(n20298) );
oa12f01 g16510 ( .a(n20166), .b(n20167), .c(n20089), .o(n20299) );
na02f01 g16511 ( .a(n20299), .b(n20298), .o(n20300) );
oa12f01 g16512 ( .a(n20177), .b(n20176), .c(n20036), .o(n20301) );
na03f01 g16513 ( .a(n20174), .b(n20173), .c(n19611), .o(n20302) );
na02f01 g16514 ( .a(n20302), .b(n20301), .o(n20303) );
na02f01 g16515 ( .a(n20303), .b(n18459), .o(n20304) );
ao12f01 g16516 ( .a(n20288), .b(n20083), .c(n20039), .o(n20305) );
no03f01 g16517 ( .a(n20286), .b(n19933), .c(n19626), .o(n20306) );
no02f01 g16518 ( .a(n20306), .b(n20305), .o(n20307) );
no02f01 g16519 ( .a(n20307), .b(n18460), .o(n20308) );
in01f01 g16520 ( .a(n20308), .o(n20309) );
no04f01 g16521 ( .a(n19968), .b(n20089), .c(n19935), .d(n19613), .o(n20310) );
ao22f01 g16522 ( .a(n20092), .b(n19951), .c(n20085), .d(n20038), .o(n20311) );
oa12f01 g16523 ( .a(n18459), .b(n20311), .c(n20310), .o(n20312) );
na03f01 g16524 ( .a(n20312), .b(n20309), .c(n20304), .o(n20313) );
ao12f01 g16525 ( .a(n20313), .b(n20300), .c(n18459), .o(n20314) );
ao12f01 g16526 ( .a(n20165), .b(n20314), .c(n20297), .o(n20315) );
na02f01 g16527 ( .a(n19977), .b(n20021), .o(n20316) );
no02f01 g16528 ( .a(n20316), .b(n20097), .o(n20317) );
no02f01 g16529 ( .a(n20098), .b(n19552), .o(n20318) );
no02f01 g16530 ( .a(n20318), .b(n19976), .o(n20319) );
oa12f01 g16531 ( .a(n18460), .b(n20319), .c(n20317), .o(n20320) );
na02f01 g16532 ( .a(n20320), .b(n20315), .o(n20321) );
na02f01 g16533 ( .a(n19987), .b(n20101), .o(n20322) );
na02f01 g16534 ( .a(n20322), .b(n19978), .o(n20323) );
no02f01 g16535 ( .a(n19988), .b(n19985), .o(n20324) );
na02f01 g16536 ( .a(n20324), .b(n20099), .o(n20325) );
na02f01 g16537 ( .a(n20325), .b(n20323), .o(n20326) );
ao12f01 g16538 ( .a(n20321), .b(n20326), .c(n18460), .o(n20327) );
oa12f01 g16539 ( .a(n20327), .b(n20159), .c(n18459), .o(n20328) );
oa12f01 g16540 ( .a(n20155), .b(n19988), .c(n20148), .o(n20329) );
na03f01 g16541 ( .a(n20156), .b(n19987), .c(n20141), .o(n20330) );
na02f01 g16542 ( .a(n20330), .b(n20329), .o(n20331) );
no02f01 g16543 ( .a(n20324), .b(n20099), .o(n20332) );
no02f01 g16544 ( .a(n20322), .b(n19978), .o(n20333) );
no02f01 g16545 ( .a(n20333), .b(n20332), .o(n20334) );
na02f01 g16546 ( .a(n20318), .b(n19976), .o(n20335) );
na02f01 g16547 ( .a(n20316), .b(n20097), .o(n20336) );
na02f01 g16548 ( .a(n20336), .b(n20335), .o(n20337) );
no02f01 g16549 ( .a(n20164), .b(n18460), .o(n20338) );
ao12f01 g16550 ( .a(n20338), .b(n20337), .c(n18459), .o(n20339) );
oa12f01 g16551 ( .a(n20339), .b(n20334), .c(n18460), .o(n20340) );
ao12f01 g16552 ( .a(n20340), .b(n20331), .c(n18459), .o(n20341) );
ao22f01 g16553 ( .a(n20341), .b(n20328), .c(n20152), .d(n18460), .o(n20342) );
na02f01 g16554 ( .a(n20342), .b(n20137), .o(n20343) );
na03f01 g16555 ( .a(n20135), .b(n20134), .c(n20127), .o(n20344) );
oa12f01 g16556 ( .a(n20128), .b(n20132), .c(n20129), .o(n20345) );
na02f01 g16557 ( .a(n20345), .b(n20344), .o(n20346) );
ao12f01 g16558 ( .a(n20150), .b(n20149), .c(n20100), .o(n20347) );
no03f01 g16559 ( .a(n20143), .b(n20142), .c(n19979), .o(n20348) );
no02f01 g16560 ( .a(n20348), .b(n20347), .o(n20349) );
no02f01 g16561 ( .a(n20349), .b(n18460), .o(n20350) );
ao12f01 g16562 ( .a(n20350), .b(n20346), .c(n18459), .o(n20351) );
no02f01 g16563 ( .a(n20113), .b(n20010), .o(n20352) );
no02f01 g16564 ( .a(n20018), .b(n19532), .o(n20353) );
no02f01 g16565 ( .a(n20107), .b(n19118), .o(n20354) );
no02f01 g16566 ( .a(n20354), .b(n20353), .o(n20355) );
na02f01 g16567 ( .a(n20355), .b(n20352), .o(n20356) );
na02f01 g16568 ( .a(n20114), .b(n20104), .o(n20357) );
in01f01 g16569 ( .a(n20355), .o(n20358) );
na02f01 g16570 ( .a(n20358), .b(n20357), .o(n20359) );
na02f01 g16571 ( .a(n20359), .b(n20356), .o(n20360) );
na02f01 g16572 ( .a(n20360), .b(n18459), .o(n20361) );
na03f01 g16573 ( .a(n20361), .b(n20351), .c(n20343), .o(n20362) );
na02f01 g16574 ( .a(n20360), .b(n18460), .o(n20363) );
na02f01 g16575 ( .a(n20363), .b(n20362), .o(n20364) );
na02f01 g16576 ( .a(n20364), .b(n20124), .o(n20365) );
no02f01 g16577 ( .a(n20120), .b(n20118), .o(n20366) );
no02f01 g16578 ( .a(n20116), .b(n19536), .o(n20367) );
oa12f01 g16579 ( .a(n18459), .b(n20367), .c(n20366), .o(n20368) );
oa12f01 g16580 ( .a(n18460), .b(n20367), .c(n20366), .o(n20369) );
na02f01 g16581 ( .a(n20369), .b(n20368), .o(n20370) );
ao12f01 g16582 ( .a(n18459), .b(n20345), .c(n20344), .o(n20371) );
na02f01 g16583 ( .a(n20303), .b(n18460), .o(n20372) );
ao12f01 g16584 ( .a(n18459), .b(n20281), .c(n20280), .o(n20373) );
in01f01 g16585 ( .a(n20200), .o(n20374) );
na02f01 g16586 ( .a(n20194), .b(n20197), .o(n20375) );
na02f01 g16587 ( .a(n20195), .b(n20193), .o(n20376) );
na02f01 g16588 ( .a(n20376), .b(n20375), .o(n20377) );
na02f01 g16589 ( .a(n20377), .b(n18459), .o(n20378) );
no02f01 g16590 ( .a(n20229), .b(n20226), .o(n20379) );
no02f01 g16591 ( .a(n20379), .b(n18459), .o(n20380) );
no03f01 g16592 ( .a(n20380), .b(n20222), .c(n20215), .o(n20381) );
na03f01 g16593 ( .a(n20234), .b(n19847), .c(n19690), .o(n20382) );
oa12f01 g16594 ( .a(n20232), .b(n20065), .c(n19689), .o(n20383) );
na02f01 g16595 ( .a(n20383), .b(n20382), .o(n20384) );
na02f01 g16596 ( .a(n20384), .b(n18460), .o(n20385) );
na02f01 g16597 ( .a(n20385), .b(n20381), .o(n20386) );
no02f01 g16598 ( .a(n20247), .b(n18459), .o(n20387) );
no02f01 g16599 ( .a(n20387), .b(n20386), .o(n20388) );
na02f01 g16600 ( .a(n20253), .b(n19867), .o(n20389) );
na02f01 g16601 ( .a(n20251), .b(n20068), .o(n20390) );
na02f01 g16602 ( .a(n20390), .b(n20389), .o(n20391) );
na02f01 g16603 ( .a(n20391), .b(n18460), .o(n20392) );
oa12f01 g16604 ( .a(n20392), .b(n20249), .c(n20388), .o(n20393) );
in01f01 g16605 ( .a(n20258), .o(n20394) );
na03f01 g16606 ( .a(n20394), .b(n20393), .c(n20378), .o(n20395) );
na02f01 g16607 ( .a(n20264), .b(n20263), .o(n20396) );
na02f01 g16608 ( .a(n20261), .b(n20260), .o(n20397) );
na02f01 g16609 ( .a(n20397), .b(n20396), .o(n20398) );
na02f01 g16610 ( .a(n20398), .b(n18460), .o(n20399) );
na03f01 g16611 ( .a(n20399), .b(n20395), .c(n20374), .o(n20400) );
in01f01 g16612 ( .a(n20275), .o(n20401) );
no03f01 g16613 ( .a(n20401), .b(n20400), .c(n20373), .o(n20402) );
in01f01 g16614 ( .a(n20279), .o(n20403) );
oa12f01 g16615 ( .a(n18459), .b(n20191), .c(n20189), .o(n20404) );
na03f01 g16616 ( .a(n20404), .b(n20403), .c(n20277), .o(n20405) );
na03f01 g16617 ( .a(n20183), .b(n20081), .c(n20040), .o(n20406) );
oa12f01 g16618 ( .a(n20181), .b(n19926), .c(n19639), .o(n20407) );
ao12f01 g16619 ( .a(n18460), .b(n20407), .c(n20406), .o(n20408) );
no03f01 g16620 ( .a(n20408), .b(n20405), .c(n20402), .o(n20409) );
no02f01 g16621 ( .a(n20307), .b(n18459), .o(n20410) );
no03f01 g16622 ( .a(n20410), .b(n20409), .c(n20186), .o(n20411) );
oa12f01 g16623 ( .a(n18460), .b(n20311), .c(n20310), .o(n20412) );
na03f01 g16624 ( .a(n20412), .b(n20411), .c(n20372), .o(n20413) );
ao12f01 g16625 ( .a(n20413), .b(n20300), .c(n18460), .o(n20414) );
no02f01 g16626 ( .a(n20179), .b(n18460), .o(n20415) );
ao12f01 g16627 ( .a(n18460), .b(n20294), .c(n20293), .o(n20416) );
no03f01 g16628 ( .a(n20416), .b(n20308), .c(n20415), .o(n20417) );
oa12f01 g16629 ( .a(n20417), .b(n20172), .c(n18460), .o(n20418) );
oa22f01 g16630 ( .a(n20418), .b(n20414), .c(n20164), .d(n18459), .o(n20419) );
ao12f01 g16631 ( .a(n18459), .b(n20336), .c(n20335), .o(n20420) );
no02f01 g16632 ( .a(n20420), .b(n20419), .o(n20421) );
oa12f01 g16633 ( .a(n20421), .b(n20334), .c(n18459), .o(n20422) );
ao12f01 g16634 ( .a(n20422), .b(n20331), .c(n18460), .o(n20423) );
no02f01 g16635 ( .a(n20319), .b(n20317), .o(n20424) );
in01f01 g16636 ( .a(n20338), .o(n20425) );
oa12f01 g16637 ( .a(n20425), .b(n20424), .c(n18460), .o(n20426) );
ao12f01 g16638 ( .a(n20426), .b(n20326), .c(n18459), .o(n20427) );
oa12f01 g16639 ( .a(n20427), .b(n20159), .c(n18460), .o(n20428) );
oa22f01 g16640 ( .a(n20428), .b(n20423), .c(n20349), .d(n18459), .o(n20429) );
no02f01 g16641 ( .a(n20429), .b(n20371), .o(n20430) );
no02f01 g16642 ( .a(n20136), .b(n20133), .o(n20431) );
na02f01 g16643 ( .a(n20152), .b(n18459), .o(n20432) );
oa12f01 g16644 ( .a(n20432), .b(n20431), .c(n18460), .o(n20433) );
no02f01 g16645 ( .a(n20358), .b(n20357), .o(n20434) );
no02f01 g16646 ( .a(n20355), .b(n20352), .o(n20435) );
no02f01 g16647 ( .a(n20435), .b(n20434), .o(n20436) );
no02f01 g16648 ( .a(n20436), .b(n18460), .o(n20437) );
no03f01 g16649 ( .a(n20437), .b(n20433), .c(n20430), .o(n20438) );
no02f01 g16650 ( .a(n20436), .b(n18459), .o(n20439) );
no02f01 g16651 ( .a(n20439), .b(n20438), .o(n20440) );
na02f01 g16652 ( .a(n20440), .b(n20370), .o(n20441) );
no02f01 g16653 ( .a(n20107), .b(n18145), .o(n20442) );
no02f01 g16654 ( .a(n20107), .b(n18103), .o(n20443) );
no02f01 g16655 ( .a(n20443), .b(n20442), .o(n20444) );
no02f01 g16656 ( .a(n19984), .b(n18103), .o(n20445) );
in01f01 g16657 ( .a(n20445), .o(n20446) );
oa12f01 g16658 ( .a(n18103), .b(n19983), .c(n19981), .o(n20447) );
na02f01 g16659 ( .a(n19594), .b(n18145), .o(n20448) );
in01f01 g16660 ( .a(n19688), .o(n20449) );
in01f01 g16661 ( .a(n19713), .o(n20450) );
ao12f01 g16662 ( .a(n18103), .b(n19738), .c(n19727), .o(n20451) );
ao12f01 g16663 ( .a(n20451), .b(n20450), .c(n18145), .o(n20452) );
oa12f01 g16664 ( .a(n20452), .b(n19701), .c(n18103), .o(n20453) );
ao12f01 g16665 ( .a(n20453), .b(n20449), .c(n18145), .o(n20454) );
oa12f01 g16666 ( .a(n20454), .b(n19859), .c(n18103), .o(n20455) );
no02f01 g16667 ( .a(n19673), .b(n18103), .o(n20456) );
no02f01 g16668 ( .a(n20456), .b(n20455), .o(n20457) );
na02f01 g16669 ( .a(n19880), .b(n18145), .o(n20458) );
na02f01 g16670 ( .a(n20458), .b(n20457), .o(n20459) );
ao12f01 g16671 ( .a(n20459), .b(n19653), .c(n18145), .o(n20460) );
oa12f01 g16672 ( .a(n20460), .b(n19899), .c(n18103), .o(n20461) );
ao12f01 g16673 ( .a(n20461), .b(n20074), .c(n18145), .o(n20462) );
oa12f01 g16674 ( .a(n20462), .b(n19638), .c(n18103), .o(n20463) );
ao12f01 g16675 ( .a(n18145), .b(n19899), .c(n19652), .o(n20464) );
in01f01 g16676 ( .a(n20464), .o(n20465) );
oa12f01 g16677 ( .a(n20465), .b(n19915), .c(n18145), .o(n20466) );
ao12f01 g16678 ( .a(n20466), .b(n19924), .c(n18103), .o(n20467) );
na02f01 g16679 ( .a(n20467), .b(n20463), .o(n20468) );
oa12f01 g16680 ( .a(n18145), .b(n19625), .c(n19610), .o(n20469) );
na03f01 g16681 ( .a(n20469), .b(n20468), .c(n20448), .o(n20470) );
ao12f01 g16682 ( .a(n20470), .b(n20088), .c(n18145), .o(n20471) );
no02f01 g16683 ( .a(n20030), .b(n18145), .o(n20472) );
no02f01 g16684 ( .a(n19931), .b(n18145), .o(n20473) );
ao12f01 g16685 ( .a(n20473), .b(n19610), .c(n18103), .o(n20474) );
in01f01 g16686 ( .a(n20474), .o(n20475) );
no02f01 g16687 ( .a(n20475), .b(n20472), .o(n20476) );
oa12f01 g16688 ( .a(n20476), .b(n19950), .c(n18145), .o(n20477) );
oa22f01 g16689 ( .a(n20477), .b(n20471), .c(n19966), .d(n18103), .o(n20478) );
ao12f01 g16690 ( .a(n20478), .b(n20025), .c(n18145), .o(n20479) );
na02f01 g16691 ( .a(n19551), .b(n18145), .o(n20480) );
na02f01 g16692 ( .a(n20480), .b(n20479), .o(n20481) );
in01f01 g16693 ( .a(n19548), .o(n20482) );
no02f01 g16694 ( .a(n19549), .b(n20482), .o(n20483) );
no02f01 g16695 ( .a(n20483), .b(n18145), .o(n20484) );
no02f01 g16696 ( .a(n19966), .b(n18145), .o(n20485) );
in01f01 g16697 ( .a(n20485), .o(n20486) );
oa12f01 g16698 ( .a(n20486), .b(n19583), .c(n18145), .o(n20487) );
no02f01 g16699 ( .a(n20487), .b(n20484), .o(n20488) );
na03f01 g16700 ( .a(n20488), .b(n20481), .c(n20447), .o(n20489) );
oa12f01 g16701 ( .a(n18145), .b(n20019), .c(n19542), .o(n20490) );
na03f01 g16702 ( .a(n20490), .b(n20489), .c(n20446), .o(n20491) );
no02f01 g16703 ( .a(n20112), .b(n18103), .o(n20492) );
no02f01 g16704 ( .a(n20492), .b(n20491), .o(n20493) );
no02f01 g16705 ( .a(n20112), .b(n18145), .o(n20494) );
no02f01 g16706 ( .a(n20020), .b(n18145), .o(n20495) );
no02f01 g16707 ( .a(n20495), .b(n20494), .o(n20496) );
in01f01 g16708 ( .a(n20496), .o(n20497) );
ao12f01 g16709 ( .a(n18145), .b(n20001), .c(n20000), .o(n20498) );
no03f01 g16710 ( .a(n20498), .b(n20497), .c(n20493), .o(n20499) );
no02f01 g16711 ( .a(n20110), .b(n18103), .o(n20500) );
oa12f01 g16712 ( .a(n20444), .b(n20500), .c(n20499), .o(n20501) );
na02f01 g16713 ( .a(n20018), .b(n18103), .o(n20502) );
na02f01 g16714 ( .a(n20018), .b(n18145), .o(n20503) );
na02f01 g16715 ( .a(n20503), .b(n20502), .o(n20504) );
in01f01 g16716 ( .a(n19981), .o(n20505) );
ao12f01 g16717 ( .a(n18145), .b(n19982), .c(n20505), .o(n20506) );
no02f01 g16718 ( .a(n20030), .b(n18103), .o(n20507) );
oa12f01 g16719 ( .a(n18145), .b(n19835), .c(n19839), .o(n20508) );
oa12f01 g16720 ( .a(n20508), .b(n19713), .c(n18103), .o(n20509) );
ao12f01 g16721 ( .a(n20509), .b(n19843), .c(n18145), .o(n20510) );
oa12f01 g16722 ( .a(n20510), .b(n19688), .c(n18103), .o(n20511) );
ao12f01 g16723 ( .a(n20511), .b(n19864), .c(n18145), .o(n20512) );
oa12f01 g16724 ( .a(n20512), .b(n19673), .c(n18103), .o(n20513) );
ao12f01 g16725 ( .a(n20513), .b(n19880), .c(n18145), .o(n20514) );
oa12f01 g16726 ( .a(n20514), .b(n19652), .c(n18103), .o(n20515) );
ao12f01 g16727 ( .a(n20515), .b(n19900), .c(n18145), .o(n20516) );
oa12f01 g16728 ( .a(n20516), .b(n19915), .c(n18103), .o(n20517) );
ao12f01 g16729 ( .a(n20517), .b(n19924), .c(n18145), .o(n20518) );
in01f01 g16730 ( .a(n20466), .o(n20519) );
oa12f01 g16731 ( .a(n20519), .b(n19638), .c(n18145), .o(n20520) );
no02f01 g16732 ( .a(n20520), .b(n20518), .o(n20521) );
in01f01 g16733 ( .a(n20469), .o(n20522) );
no03f01 g16734 ( .a(n20522), .b(n20521), .c(n20507), .o(n20523) );
oa12f01 g16735 ( .a(n20523), .b(n19950), .c(n18103), .o(n20524) );
na02f01 g16736 ( .a(n19594), .b(n18103), .o(n20525) );
na02f01 g16737 ( .a(n20474), .b(n20525), .o(n20526) );
ao12f01 g16738 ( .a(n20526), .b(n20088), .c(n18103), .o(n20527) );
ao22f01 g16739 ( .a(n20527), .b(n20524), .c(n19972), .d(n18145), .o(n20528) );
oa12f01 g16740 ( .a(n20528), .b(n19583), .c(n18103), .o(n20529) );
no02f01 g16741 ( .a(n20483), .b(n18103), .o(n20530) );
no02f01 g16742 ( .a(n20530), .b(n20529), .o(n20531) );
na02f01 g16743 ( .a(n19551), .b(n18103), .o(n20532) );
ao12f01 g16744 ( .a(n20485), .b(n20025), .c(n18103), .o(n20533) );
na02f01 g16745 ( .a(n20533), .b(n20532), .o(n20534) );
no03f01 g16746 ( .a(n20534), .b(n20531), .c(n20506), .o(n20535) );
ao12f01 g16747 ( .a(n18103), .b(n19544), .c(n19543), .o(n20536) );
no03f01 g16748 ( .a(n20536), .b(n20535), .c(n20445), .o(n20537) );
na02f01 g16749 ( .a(n20008), .b(n18145), .o(n20538) );
na02f01 g16750 ( .a(n20538), .b(n20537), .o(n20539) );
oa12f01 g16751 ( .a(n18103), .b(n20109), .c(n19999), .o(n20540) );
na03f01 g16752 ( .a(n20540), .b(n20496), .c(n20539), .o(n20541) );
na02f01 g16753 ( .a(n20002), .b(n18145), .o(n20542) );
na03f01 g16754 ( .a(n20542), .b(n20541), .c(n20504), .o(n20543) );
na03f01 g16755 ( .a(n20543), .b(n20501), .c(n19051), .o(n20544) );
ao12f01 g16756 ( .a(n20504), .b(n20542), .c(n20541), .o(n20545) );
no03f01 g16757 ( .a(n20500), .b(n20499), .c(n20444), .o(n20546) );
oa12f01 g16758 ( .a(n19050), .b(n20546), .c(n20545), .o(n20547) );
na02f01 g16759 ( .a(n20547), .b(n20544), .o(n20548) );
na02f01 g16760 ( .a(n20496), .b(n20539), .o(n20549) );
no03f01 g16761 ( .a(n20500), .b(n20498), .c(n20549), .o(n20550) );
no02f01 g16762 ( .a(n20497), .b(n20493), .o(n20551) );
ao12f01 g16763 ( .a(n20551), .b(n20542), .c(n20540), .o(n20552) );
oa12f01 g16764 ( .a(n18905), .b(n20552), .c(n20550), .o(n20553) );
na03f01 g16765 ( .a(n20542), .b(n20540), .c(n20551), .o(n20554) );
oa12f01 g16766 ( .a(n20549), .b(n20500), .c(n20498), .o(n20555) );
na03f01 g16767 ( .a(n20555), .b(n20554), .c(n18906), .o(n20556) );
no02f01 g16768 ( .a(n20534), .b(n20531), .o(n20557) );
no02f01 g16769 ( .a(n20506), .b(n20445), .o(n20558) );
no02f01 g16770 ( .a(n20558), .b(n20557), .o(n20559) );
na02f01 g16771 ( .a(n20558), .b(n20557), .o(n20560) );
in01f01 g16772 ( .a(n20560), .o(n20561) );
oa12f01 g16773 ( .a(n19024), .b(n20561), .c(n20559), .o(n20562) );
no02f01 g16774 ( .a(n20484), .b(n20530), .o(n20563) );
no02f01 g16775 ( .a(n20487), .b(n20479), .o(n20564) );
no02f01 g16776 ( .a(n20564), .b(n20563), .o(n20565) );
na02f01 g16777 ( .a(n20532), .b(n20480), .o(n20566) );
na02f01 g16778 ( .a(n20533), .b(n20529), .o(n20567) );
no02f01 g16779 ( .a(n20567), .b(n20566), .o(n20568) );
no02f01 g16780 ( .a(n20568), .b(n20565), .o(n20569) );
na02f01 g16781 ( .a(n20569), .b(n19004), .o(n20570) );
na02f01 g16782 ( .a(n20469), .b(n20518), .o(n20571) );
na02f01 g16783 ( .a(n20474), .b(n20467), .o(n20572) );
no02f01 g16784 ( .a(n20572), .b(n20472), .o(n20573) );
oa12f01 g16785 ( .a(n20573), .b(n20571), .c(n20507), .o(n20574) );
no02f01 g16786 ( .a(n20574), .b(n20088), .o(n20575) );
in01f01 g16787 ( .a(n20575), .o(n20576) );
na02f01 g16788 ( .a(n20574), .b(n20088), .o(n20577) );
na02f01 g16789 ( .a(n20577), .b(n20576), .o(n20578) );
no02f01 g16790 ( .a(n20578), .b(n18978), .o(n20579) );
in01f01 g16791 ( .a(n18970), .o(n20580) );
ao12f01 g16792 ( .a(n20572), .b(n20469), .c(n20518), .o(n20581) );
na02f01 g16793 ( .a(n20581), .b(n20030), .o(n20582) );
in01f01 g16794 ( .a(n20582), .o(n20583) );
no02f01 g16795 ( .a(n20581), .b(n20030), .o(n20584) );
no02f01 g16796 ( .a(n20584), .b(n20583), .o(n20585) );
na02f01 g16797 ( .a(n20585), .b(n20580), .o(n20586) );
no02f01 g16798 ( .a(n19931), .b(n18103), .o(n20587) );
no02f01 g16799 ( .a(n20587), .b(n20463), .o(n20588) );
no03f01 g16800 ( .a(n20588), .b(n20473), .c(n20520), .o(n20589) );
na02f01 g16801 ( .a(n20589), .b(n20035), .o(n20590) );
no02f01 g16802 ( .a(n20473), .b(n20520), .o(n20591) );
oa12f01 g16803 ( .a(n20591), .b(n20587), .c(n20463), .o(n20592) );
na02f01 g16804 ( .a(n20592), .b(n19610), .o(n20593) );
na02f01 g16805 ( .a(n20593), .b(n20590), .o(n20594) );
no02f01 g16806 ( .a(n20594), .b(n18962), .o(n20595) );
na02f01 g16807 ( .a(n20521), .b(n19931), .o(n20596) );
na02f01 g16808 ( .a(n20468), .b(n19625), .o(n20597) );
na02f01 g16809 ( .a(n20597), .b(n20596), .o(n20598) );
no02f01 g16810 ( .a(n20598), .b(n18952), .o(n20599) );
in01f01 g16811 ( .a(n20599), .o(n20600) );
in01f01 g16812 ( .a(n18944), .o(n20601) );
na02f01 g16813 ( .a(n20519), .b(n20517), .o(n20602) );
no02f01 g16814 ( .a(n20602), .b(n19924), .o(n20603) );
no02f01 g16815 ( .a(n20466), .b(n20462), .o(n20604) );
no02f01 g16816 ( .a(n20604), .b(n19638), .o(n20605) );
no02f01 g16817 ( .a(n20605), .b(n20603), .o(n20606) );
no02f01 g16818 ( .a(n20606), .b(n20601), .o(n20607) );
in01f01 g16819 ( .a(n20607), .o(n20608) );
na02f01 g16820 ( .a(n20465), .b(n20461), .o(n20609) );
na02f01 g16821 ( .a(n20609), .b(n20074), .o(n20610) );
no02f01 g16822 ( .a(n20464), .b(n20516), .o(n20611) );
na02f01 g16823 ( .a(n20611), .b(n19915), .o(n20612) );
na02f01 g16824 ( .a(n20612), .b(n20610), .o(n20613) );
no02f01 g16825 ( .a(n20613), .b(n18934), .o(n20614) );
in01f01 g16826 ( .a(n20614), .o(n20615) );
no02f01 g16827 ( .a(n19652), .b(n18145), .o(n20616) );
oa12f01 g16828 ( .a(n19900), .b(n20616), .c(n20460), .o(n20617) );
in01f01 g16829 ( .a(n20616), .o(n20618) );
na03f01 g16830 ( .a(n20618), .b(n20515), .c(n19899), .o(n20619) );
ao12f01 g16831 ( .a(n18913), .b(n20619), .c(n20617), .o(n20620) );
in01f01 g16832 ( .a(n20620), .o(n20621) );
no02f01 g16833 ( .a(n20513), .b(n19881), .o(n20622) );
no02f01 g16834 ( .a(n20457), .b(n19880), .o(n20623) );
no02f01 g16835 ( .a(n20623), .b(n20622), .o(n20624) );
in01f01 g16836 ( .a(n20624), .o(n20625) );
no02f01 g16837 ( .a(n20625), .b(n18918), .o(n20626) );
no02f01 g16838 ( .a(n20512), .b(n19674), .o(n20627) );
no02f01 g16839 ( .a(n20455), .b(n19673), .o(n20628) );
no02f01 g16840 ( .a(n20628), .b(n20627), .o(n20629) );
no02f01 g16841 ( .a(n18773), .b(n18770), .o(n20630) );
no02f01 g16842 ( .a(n20630), .b(n18762), .o(n20631) );
na02f01 g16843 ( .a(n20630), .b(n18762), .o(n20632) );
in01f01 g16844 ( .a(n20632), .o(n20633) );
no02f01 g16845 ( .a(n20633), .b(n20631), .o(n20634) );
in01f01 g16846 ( .a(n20634), .o(n20635) );
na02f01 g16847 ( .a(n20635), .b(n20629), .o(n20636) );
no02f01 g16848 ( .a(n20454), .b(n19864), .o(n20637) );
no02f01 g16849 ( .a(n20511), .b(n19859), .o(n20638) );
no02f01 g16850 ( .a(n20638), .b(n20637), .o(n20639) );
in01f01 g16851 ( .a(n18761), .o(n20640) );
na02f01 g16852 ( .a(n20640), .b(n18760), .o(n20641) );
no02f01 g16853 ( .a(n20641), .b(n18751), .o(n20642) );
na02f01 g16854 ( .a(n20641), .b(n18751), .o(n20643) );
in01f01 g16855 ( .a(n20643), .o(n20644) );
no02f01 g16856 ( .a(n20644), .b(n20642), .o(n20645) );
in01f01 g16857 ( .a(n20645), .o(n20646) );
na02f01 g16858 ( .a(n20646), .b(n20639), .o(n20647) );
in01f01 g16859 ( .a(n20647), .o(n20648) );
no02f01 g16860 ( .a(n20510), .b(n20449), .o(n20649) );
na02f01 g16861 ( .a(n20510), .b(n20449), .o(n20650) );
in01f01 g16862 ( .a(n20650), .o(n20651) );
no02f01 g16863 ( .a(n20651), .b(n20649), .o(n20652) );
in01f01 g16864 ( .a(n18749), .o(n20653) );
no02f01 g16865 ( .a(n18750), .b(n18710), .o(n20654) );
in01f01 g16866 ( .a(n20654), .o(n20655) );
no02f01 g16867 ( .a(n20655), .b(n20653), .o(n20656) );
no02f01 g16868 ( .a(n20654), .b(n18749), .o(n20657) );
no02f01 g16869 ( .a(n20657), .b(n20656), .o(n20658) );
in01f01 g16870 ( .a(n20658), .o(n20659) );
na02f01 g16871 ( .a(n20659), .b(n20652), .o(n20660) );
na02f01 g16872 ( .a(n20509), .b(n19701), .o(n20661) );
no02f01 g16873 ( .a(n20509), .b(n19701), .o(n20662) );
in01f01 g16874 ( .a(n20662), .o(n20663) );
na02f01 g16875 ( .a(n20663), .b(n20661), .o(n20664) );
no03f01 g16876 ( .a(n18747), .b(n18746), .c(n18720), .o(n20665) );
in01f01 g16877 ( .a(n18746), .o(n20666) );
no02f01 g16878 ( .a(n18747), .b(n18720), .o(n20667) );
no02f01 g16879 ( .a(n20667), .b(n20666), .o(n20668) );
no02f01 g16880 ( .a(n20668), .b(n20665), .o(n20669) );
no02f01 g16881 ( .a(n20669), .b(n20664), .o(n20670) );
in01f01 g16882 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_0_), .o(n20671) );
no02f01 g16883 ( .a(n18733), .b(n20671), .o(n20672) );
ao12f01 g16884 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_0_), .b(n18732), .c(n18731), .o(n20673) );
no02f01 g16885 ( .a(n20673), .b(n20672), .o(n20674) );
no02f01 g16886 ( .a(n20674), .b(n19738), .o(n20675) );
in01f01 g16887 ( .a(n18734), .o(n20676) );
no02f01 g16888 ( .a(n18744), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_1_), .o(n20677) );
no03f01 g16889 ( .a(n18743), .b(n18742), .c(n18729), .o(n20678) );
no03f01 g16890 ( .a(n20678), .b(n20677), .c(n20676), .o(n20679) );
no02f01 g16891 ( .a(n20678), .b(n20677), .o(n20680) );
no02f01 g16892 ( .a(n20680), .b(n18734), .o(n20681) );
no02f01 g16893 ( .a(n20681), .b(n20679), .o(n20682) );
no02f01 g16894 ( .a(n20682), .b(n20675), .o(n20683) );
ao12f01 g16895 ( .a(n19727), .b(n19835), .c(n18145), .o(n20684) );
na03f01 g16896 ( .a(n19835), .b(n19727), .c(n18145), .o(n20685) );
in01f01 g16897 ( .a(n20685), .o(n20686) );
no02f01 g16898 ( .a(n20686), .b(n20684), .o(n20687) );
in01f01 g16899 ( .a(n20682), .o(n20688) );
no03f01 g16900 ( .a(n20688), .b(n20674), .c(n19738), .o(n20689) );
in01f01 g16901 ( .a(n20689), .o(n20690) );
ao12f01 g16902 ( .a(n20683), .b(n20690), .c(n20687), .o(n20691) );
no02f01 g16903 ( .a(n20508), .b(n20450), .o(n20692) );
in01f01 g16904 ( .a(n20692), .o(n20693) );
na02f01 g16905 ( .a(n20508), .b(n20450), .o(n20694) );
in01f01 g16906 ( .a(n18727), .o(n20695) );
no02f01 g16907 ( .a(n18728), .b(n20695), .o(n20696) );
no02f01 g16908 ( .a(n20696), .b(n18745), .o(n20697) );
na02f01 g16909 ( .a(n20696), .b(n18745), .o(n20698) );
in01f01 g16910 ( .a(n20698), .o(n20699) );
no02f01 g16911 ( .a(n20699), .b(n20697), .o(n20700) );
in01f01 g16912 ( .a(n20700), .o(n20701) );
ao12f01 g16913 ( .a(n20701), .b(n20694), .c(n20693), .o(n20702) );
in01f01 g16914 ( .a(n20694), .o(n20703) );
no03f01 g16915 ( .a(n20700), .b(n20703), .c(n20692), .o(n20704) );
in01f01 g16916 ( .a(n20704), .o(n20705) );
oa12f01 g16917 ( .a(n20705), .b(n20702), .c(n20691), .o(n20706) );
na02f01 g16918 ( .a(n20669), .b(n20664), .o(n20707) );
ao12f01 g16919 ( .a(n20670), .b(n20707), .c(n20706), .o(n20708) );
no02f01 g16920 ( .a(n20659), .b(n20652), .o(n20709) );
oa12f01 g16921 ( .a(n20660), .b(n20709), .c(n20708), .o(n20710) );
no02f01 g16922 ( .a(n20646), .b(n20639), .o(n20711) );
in01f01 g16923 ( .a(n20711), .o(n20712) );
ao12f01 g16924 ( .a(n20648), .b(n20712), .c(n20710), .o(n20713) );
no02f01 g16925 ( .a(n20635), .b(n20629), .o(n20714) );
oa12f01 g16926 ( .a(n20636), .b(n20714), .c(n20713), .o(n20715) );
no02f01 g16927 ( .a(n20624), .b(n18919), .o(n20716) );
in01f01 g16928 ( .a(n20716), .o(n20717) );
ao12f01 g16929 ( .a(n20626), .b(n20717), .c(n20715), .o(n20718) );
no02f01 g16930 ( .a(n20459), .b(n19652), .o(n20719) );
no02f01 g16931 ( .a(n20514), .b(n19653), .o(n20720) );
no02f01 g16932 ( .a(n20720), .b(n20719), .o(n20721) );
no02f01 g16933 ( .a(n20721), .b(n18925), .o(n20722) );
na02f01 g16934 ( .a(n20721), .b(n18925), .o(n20723) );
in01f01 g16935 ( .a(n20723), .o(n20724) );
ao12f01 g16936 ( .a(n19899), .b(n20618), .c(n20515), .o(n20725) );
in01f01 g16937 ( .a(n20619), .o(n20726) );
no03f01 g16938 ( .a(n20726), .b(n20725), .c(n18912), .o(n20727) );
no02f01 g16939 ( .a(n20727), .b(n20724), .o(n20728) );
oa12f01 g16940 ( .a(n20728), .b(n20722), .c(n20718), .o(n20729) );
na02f01 g16941 ( .a(n20613), .b(n18934), .o(n20730) );
na03f01 g16942 ( .a(n20730), .b(n20729), .c(n20621), .o(n20731) );
no03f01 g16943 ( .a(n20605), .b(n20603), .c(n18944), .o(n20732) );
in01f01 g16944 ( .a(n20732), .o(n20733) );
na03f01 g16945 ( .a(n20733), .b(n20731), .c(n20615), .o(n20734) );
ao12f01 g16946 ( .a(n19754), .b(n20597), .c(n20596), .o(n20735) );
in01f01 g16947 ( .a(n20735), .o(n20736) );
na03f01 g16948 ( .a(n20736), .b(n20734), .c(n20608), .o(n20737) );
ao12f01 g16949 ( .a(n18963), .b(n20593), .c(n20590), .o(n20738) );
ao12f01 g16950 ( .a(n20738), .b(n20737), .c(n20600), .o(n20739) );
no02f01 g16951 ( .a(n20739), .b(n20595), .o(n20740) );
no02f01 g16952 ( .a(n20585), .b(n20580), .o(n20741) );
oa12f01 g16953 ( .a(n20586), .b(n20741), .c(n20740), .o(n20742) );
na02f01 g16954 ( .a(n20578), .b(n18978), .o(n20743) );
ao12f01 g16955 ( .a(n20579), .b(n20743), .c(n20742), .o(n20744) );
na02f01 g16956 ( .a(n20527), .b(n20524), .o(n20745) );
no02f01 g16957 ( .a(n20745), .b(n19972), .o(n20746) );
no02f01 g16958 ( .a(n20477), .b(n20471), .o(n20747) );
no02f01 g16959 ( .a(n20747), .b(n19966), .o(n20748) );
no02f01 g16960 ( .a(n20748), .b(n20746), .o(n20749) );
no02f01 g16961 ( .a(n20749), .b(n19005), .o(n20750) );
no02f01 g16962 ( .a(n20485), .b(n20528), .o(n20751) );
na02f01 g16963 ( .a(n20751), .b(n19583), .o(n20752) );
na02f01 g16964 ( .a(n20486), .b(n20478), .o(n20753) );
na02f01 g16965 ( .a(n20753), .b(n20025), .o(n20754) );
ao12f01 g16966 ( .a(n18995), .b(n20754), .c(n20752), .o(n20755) );
no03f01 g16967 ( .a(n20755), .b(n20750), .c(n20744), .o(n20756) );
na03f01 g16968 ( .a(n20754), .b(n20752), .c(n18995), .o(n20757) );
na02f01 g16969 ( .a(n20749), .b(n19005), .o(n20758) );
ao12f01 g16970 ( .a(n20755), .b(n20758), .c(n20757), .o(n20759) );
na02f01 g16971 ( .a(n20567), .b(n20566), .o(n20760) );
na02f01 g16972 ( .a(n20564), .b(n20563), .o(n20761) );
na02f01 g16973 ( .a(n20761), .b(n20760), .o(n20762) );
na02f01 g16974 ( .a(n20762), .b(n19002), .o(n20763) );
oa12f01 g16975 ( .a(n20763), .b(n20759), .c(n20756), .o(n20764) );
in01f01 g16976 ( .a(n20559), .o(n20765) );
na03f01 g16977 ( .a(n20560), .b(n20765), .c(n19848), .o(n20766) );
na03f01 g16978 ( .a(n20766), .b(n20764), .c(n20570), .o(n20767) );
no02f01 g16979 ( .a(n20535), .b(n20445), .o(n20768) );
in01f01 g16980 ( .a(n20768), .o(n20769) );
no02f01 g16981 ( .a(n20495), .b(n20536), .o(n20770) );
no02f01 g16982 ( .a(n20770), .b(n20769), .o(n20771) );
na02f01 g16983 ( .a(n19545), .b(n18103), .o(n20772) );
na02f01 g16984 ( .a(n20772), .b(n20490), .o(n20773) );
no02f01 g16985 ( .a(n20773), .b(n20768), .o(n20774) );
oa12f01 g16986 ( .a(n19664), .b(n20774), .c(n20771), .o(n20775) );
na02f01 g16987 ( .a(n20008), .b(n18103), .o(n20776) );
na02f01 g16988 ( .a(n20776), .b(n20538), .o(n20777) );
no03f01 g16989 ( .a(n20777), .b(n20495), .c(n20537), .o(n20778) );
no02f01 g16990 ( .a(n20494), .b(n20492), .o(n20779) );
ao12f01 g16991 ( .a(n20779), .b(n20772), .c(n20491), .o(n20780) );
oa12f01 g16992 ( .a(n19034), .b(n20780), .c(n20778), .o(n20781) );
na04f01 g16993 ( .a(n20781), .b(n20775), .c(n20767), .d(n20562), .o(n20782) );
no03f01 g16994 ( .a(n20780), .b(n20778), .c(n19034), .o(n20783) );
no03f01 g16995 ( .a(n20774), .b(n20771), .c(n19664), .o(n20784) );
oa12f01 g16996 ( .a(n20781), .b(n20784), .c(n20783), .o(n20785) );
na03f01 g16997 ( .a(n20785), .b(n20782), .c(n20556), .o(n20786) );
ao12f01 g16998 ( .a(n20548), .b(n20786), .c(n20553), .o(n20787) );
no03f01 g16999 ( .a(n20546), .b(n20545), .c(n19050), .o(n20788) );
ao12f01 g17000 ( .a(n19051), .b(n20543), .c(n20501), .o(n20789) );
no02f01 g17001 ( .a(n20789), .b(n20788), .o(n20790) );
ao12f01 g17002 ( .a(n18906), .b(n20555), .c(n20554), .o(n20791) );
no03f01 g17003 ( .a(n20552), .b(n20550), .c(n18905), .o(n20792) );
ao12f01 g17004 ( .a(n19848), .b(n20560), .c(n20765), .o(n20793) );
no02f01 g17005 ( .a(n20762), .b(n19002), .o(n20794) );
in01f01 g17006 ( .a(n20577), .o(n20795) );
no02f01 g17007 ( .a(n20795), .b(n20575), .o(n20796) );
na02f01 g17008 ( .a(n20796), .b(n18979), .o(n20797) );
in01f01 g17009 ( .a(n20584), .o(n20798) );
na02f01 g17010 ( .a(n20798), .b(n20582), .o(n20799) );
no02f01 g17011 ( .a(n20799), .b(n18970), .o(n20800) );
in01f01 g17012 ( .a(n20595), .o(n20801) );
in01f01 g17013 ( .a(n20626), .o(n20802) );
in01f01 g17014 ( .a(n20636), .o(n20803) );
in01f01 g17015 ( .a(n20649), .o(n20804) );
na02f01 g17016 ( .a(n20650), .b(n20804), .o(n20805) );
no02f01 g17017 ( .a(n20658), .b(n20805), .o(n20806) );
in01f01 g17018 ( .a(n20661), .o(n20807) );
no02f01 g17019 ( .a(n20662), .b(n20807), .o(n20808) );
in01f01 g17020 ( .a(n20669), .o(n20809) );
na02f01 g17021 ( .a(n20809), .b(n20808), .o(n20810) );
in01f01 g17022 ( .a(n20683), .o(n20811) );
in01f01 g17023 ( .a(n20684), .o(n20812) );
na03f01 g17024 ( .a(n20690), .b(n20685), .c(n20812), .o(n20813) );
na02f01 g17025 ( .a(n20813), .b(n20811), .o(n20814) );
oa12f01 g17026 ( .a(n20700), .b(n20703), .c(n20692), .o(n20815) );
ao12f01 g17027 ( .a(n20704), .b(n20815), .c(n20814), .o(n20816) );
no02f01 g17028 ( .a(n20809), .b(n20808), .o(n20817) );
oa12f01 g17029 ( .a(n20810), .b(n20817), .c(n20816), .o(n20818) );
na02f01 g17030 ( .a(n20658), .b(n20805), .o(n20819) );
ao12f01 g17031 ( .a(n20806), .b(n20819), .c(n20818), .o(n20820) );
oa12f01 g17032 ( .a(n20647), .b(n20711), .c(n20820), .o(n20821) );
in01f01 g17033 ( .a(n20714), .o(n20822) );
ao12f01 g17034 ( .a(n20803), .b(n20822), .c(n20821), .o(n20823) );
oa12f01 g17035 ( .a(n20802), .b(n20716), .c(n20823), .o(n20824) );
in01f01 g17036 ( .a(n20722), .o(n20825) );
na03f01 g17037 ( .a(n20619), .b(n20617), .c(n18913), .o(n20826) );
na02f01 g17038 ( .a(n20826), .b(n20723), .o(n20827) );
ao12f01 g17039 ( .a(n20827), .b(n20825), .c(n20824), .o(n20828) );
ao12f01 g17040 ( .a(n18935), .b(n20612), .c(n20610), .o(n20829) );
no03f01 g17041 ( .a(n20829), .b(n20828), .c(n20620), .o(n20830) );
no03f01 g17042 ( .a(n20732), .b(n20830), .c(n20614), .o(n20831) );
no03f01 g17043 ( .a(n20735), .b(n20831), .c(n20607), .o(n20832) );
in01f01 g17044 ( .a(n20738), .o(n20833) );
oa12f01 g17045 ( .a(n20833), .b(n20832), .c(n20599), .o(n20834) );
na02f01 g17046 ( .a(n20834), .b(n20801), .o(n20835) );
na02f01 g17047 ( .a(n20799), .b(n18970), .o(n20836) );
ao12f01 g17048 ( .a(n20800), .b(n20836), .c(n20835), .o(n20837) );
no02f01 g17049 ( .a(n20796), .b(n18979), .o(n20838) );
oa12f01 g17050 ( .a(n20797), .b(n20838), .c(n20837), .o(n20839) );
na02f01 g17051 ( .a(n20747), .b(n19966), .o(n20840) );
na02f01 g17052 ( .a(n20745), .b(n19972), .o(n20841) );
na02f01 g17053 ( .a(n20841), .b(n20840), .o(n20842) );
na02f01 g17054 ( .a(n20842), .b(n18986), .o(n20843) );
no02f01 g17055 ( .a(n20753), .b(n20025), .o(n20844) );
no02f01 g17056 ( .a(n20751), .b(n19583), .o(n20845) );
oa12f01 g17057 ( .a(n18994), .b(n20845), .c(n20844), .o(n20846) );
na03f01 g17058 ( .a(n20846), .b(n20843), .c(n20839), .o(n20847) );
no03f01 g17059 ( .a(n20845), .b(n20844), .c(n18994), .o(n20848) );
no02f01 g17060 ( .a(n20842), .b(n18986), .o(n20849) );
oa12f01 g17061 ( .a(n20846), .b(n20849), .c(n20848), .o(n20850) );
no02f01 g17062 ( .a(n20569), .b(n19004), .o(n20851) );
ao12f01 g17063 ( .a(n20851), .b(n20850), .c(n20847), .o(n20852) );
no03f01 g17064 ( .a(n20561), .b(n20559), .c(n19024), .o(n20853) );
no03f01 g17065 ( .a(n20853), .b(n20852), .c(n20794), .o(n20854) );
na02f01 g17066 ( .a(n20773), .b(n20768), .o(n20855) );
na02f01 g17067 ( .a(n20770), .b(n20769), .o(n20856) );
ao12f01 g17068 ( .a(n19017), .b(n20856), .c(n20855), .o(n20857) );
na03f01 g17069 ( .a(n20779), .b(n20772), .c(n20491), .o(n20858) );
oa12f01 g17070 ( .a(n20777), .b(n20495), .c(n20537), .o(n20859) );
ao12f01 g17071 ( .a(n19559), .b(n20859), .c(n20858), .o(n20860) );
no04f01 g17072 ( .a(n20860), .b(n20857), .c(n20854), .d(n20793), .o(n20861) );
na03f01 g17073 ( .a(n20859), .b(n20858), .c(n19559), .o(n20862) );
na03f01 g17074 ( .a(n20856), .b(n20855), .c(n19017), .o(n20863) );
ao12f01 g17075 ( .a(n20860), .b(n20863), .c(n20862), .o(n20864) );
no03f01 g17076 ( .a(n20864), .b(n20861), .c(n20792), .o(n20865) );
no03f01 g17077 ( .a(n20865), .b(n20791), .c(n20790), .o(n20866) );
no02f01 g17078 ( .a(n20866), .b(n20787), .o(n20867) );
in01f01 g17079 ( .a(n20867), .o(n20868) );
ao12f01 g17080 ( .a(n20868), .b(n20441), .c(n20365), .o(n20869) );
no02f01 g17081 ( .a(n20440), .b(n20370), .o(n20870) );
no02f01 g17082 ( .a(n20364), .b(n20124), .o(n20871) );
no03f01 g17083 ( .a(n20867), .b(n20871), .c(n20870), .o(n20872) );
in01f01 g17084 ( .a(n20872), .o(n20873) );
no02f01 g17085 ( .a(n20433), .b(n20430), .o(n20874) );
no02f01 g17086 ( .a(n20439), .b(n20437), .o(n20875) );
no02f01 g17087 ( .a(n20875), .b(n20874), .o(n20876) );
na02f01 g17088 ( .a(n20351), .b(n20343), .o(n20877) );
na02f01 g17089 ( .a(n20363), .b(n20361), .o(n20878) );
no02f01 g17090 ( .a(n20878), .b(n20877), .o(n20879) );
na02f01 g17091 ( .a(n20785), .b(n20782), .o(n20880) );
na02f01 g17092 ( .a(n20556), .b(n20553), .o(n20881) );
no02f01 g17093 ( .a(n20881), .b(n20880), .o(n20882) );
no02f01 g17094 ( .a(n20864), .b(n20861), .o(n20883) );
no02f01 g17095 ( .a(n20792), .b(n20791), .o(n20884) );
no02f01 g17096 ( .a(n20884), .b(n20883), .o(n20885) );
no02f01 g17097 ( .a(n20885), .b(n20882), .o(n20886) );
no03f01 g17098 ( .a(n20886), .b(n20879), .c(n20876), .o(n20887) );
oa12f01 g17099 ( .a(n20886), .b(n20879), .c(n20876), .o(n20888) );
no02f01 g17100 ( .a(n20431), .b(n18460), .o(n20889) );
na02f01 g17101 ( .a(n20432), .b(n20429), .o(n20890) );
oa12f01 g17102 ( .a(n20890), .b(n20889), .c(n20371), .o(n20891) );
na02f01 g17103 ( .a(n20346), .b(n18459), .o(n20892) );
no02f01 g17104 ( .a(n20350), .b(n20342), .o(n20893) );
na03f01 g17105 ( .a(n20893), .b(n20892), .c(n20137), .o(n20894) );
no02f01 g17106 ( .a(n20854), .b(n20793), .o(n20895) );
na02f01 g17107 ( .a(n20775), .b(n20895), .o(n20896) );
no02f01 g17108 ( .a(n20783), .b(n20860), .o(n20897) );
na03f01 g17109 ( .a(n20897), .b(n20863), .c(n20896), .o(n20898) );
na02f01 g17110 ( .a(n20767), .b(n20562), .o(n20899) );
no02f01 g17111 ( .a(n20857), .b(n20899), .o(n20900) );
in01f01 g17112 ( .a(n20897), .o(n20901) );
oa12f01 g17113 ( .a(n20901), .b(n20784), .c(n20900), .o(n20902) );
na02f01 g17114 ( .a(n20902), .b(n20898), .o(n20903) );
ao12f01 g17115 ( .a(n20903), .b(n20894), .c(n20891), .o(n20904) );
na03f01 g17116 ( .a(n20903), .b(n20894), .c(n20891), .o(n20905) );
no02f01 g17117 ( .a(n20428), .b(n20423), .o(n20906) );
no02f01 g17118 ( .a(n20349), .b(n18459), .o(n20907) );
no02f01 g17119 ( .a(n20350), .b(n20907), .o(n20908) );
no02f01 g17120 ( .a(n20908), .b(n20906), .o(n20909) );
in01f01 g17121 ( .a(n20906), .o(n20910) );
na02f01 g17122 ( .a(n20152), .b(n18460), .o(n20911) );
na02f01 g17123 ( .a(n20432), .b(n20911), .o(n20912) );
no02f01 g17124 ( .a(n20912), .b(n20910), .o(n20913) );
no02f01 g17125 ( .a(n20913), .b(n20909), .o(n20914) );
no02f01 g17126 ( .a(n20784), .b(n20857), .o(n20915) );
in01f01 g17127 ( .a(n20915), .o(n20916) );
na02f01 g17128 ( .a(n20916), .b(n20895), .o(n20917) );
na02f01 g17129 ( .a(n20915), .b(n20899), .o(n20918) );
na02f01 g17130 ( .a(n20918), .b(n20917), .o(n20919) );
na02f01 g17131 ( .a(n20919), .b(n20914), .o(n20920) );
ao12f01 g17132 ( .a(n20904), .b(n20920), .c(n20905), .o(n20921) );
ao12f01 g17133 ( .a(n20887), .b(n20921), .c(n20888), .o(n20922) );
ao12f01 g17134 ( .a(n20869), .b(n20922), .c(n20873), .o(n20923) );
oa12f01 g17135 ( .a(n20867), .b(n20871), .c(n20870), .o(n20924) );
na02f01 g17136 ( .a(n20878), .b(n20877), .o(n20925) );
na02f01 g17137 ( .a(n20875), .b(n20874), .o(n20926) );
na02f01 g17138 ( .a(n20884), .b(n20883), .o(n20927) );
na02f01 g17139 ( .a(n20881), .b(n20880), .o(n20928) );
na02f01 g17140 ( .a(n20928), .b(n20927), .o(n20929) );
ao12f01 g17141 ( .a(n20929), .b(n20926), .c(n20925), .o(n20930) );
no02f01 g17142 ( .a(n20919), .b(n20914), .o(n20931) );
no03f01 g17143 ( .a(n20931), .b(n20904), .c(n20930), .o(n20932) );
na02f01 g17144 ( .a(n20932), .b(n20924), .o(n20933) );
no02f01 g17145 ( .a(n20159), .b(n18459), .o(n20934) );
no02f01 g17146 ( .a(n20159), .b(n18460), .o(n20935) );
no02f01 g17147 ( .a(n20935), .b(n20934), .o(n20936) );
in01f01 g17148 ( .a(n20936), .o(n20937) );
no02f01 g17149 ( .a(n20340), .b(n20327), .o(n20938) );
in01f01 g17150 ( .a(n20938), .o(n20939) );
no02f01 g17151 ( .a(n20939), .b(n20937), .o(n20940) );
no02f01 g17152 ( .a(n20938), .b(n20936), .o(n20941) );
no02f01 g17153 ( .a(n20941), .b(n20940), .o(n20942) );
no02f01 g17154 ( .a(n20852), .b(n20794), .o(n20943) );
no02f01 g17155 ( .a(n20853), .b(n20793), .o(n20944) );
na02f01 g17156 ( .a(n20944), .b(n20943), .o(n20945) );
in01f01 g17157 ( .a(n20945), .o(n20946) );
oa22f01 g17158 ( .a(n20853), .b(n20793), .c(n20852), .d(n20794), .o(n20947) );
in01f01 g17159 ( .a(n20947), .o(n20948) );
no02f01 g17160 ( .a(n20948), .b(n20946), .o(n20949) );
in01f01 g17161 ( .a(n20949), .o(n20950) );
no02f01 g17162 ( .a(n20950), .b(n20942), .o(n20951) );
in01f01 g17163 ( .a(n20942), .o(n20952) );
no02f01 g17164 ( .a(n20949), .b(n20952), .o(n20953) );
in01f01 g17165 ( .a(n20953), .o(n20954) );
no02f01 g17166 ( .a(n20426), .b(n20421), .o(n20955) );
no02f01 g17167 ( .a(n20334), .b(n18459), .o(n20956) );
no02f01 g17168 ( .a(n20334), .b(n18460), .o(n20957) );
no02f01 g17169 ( .a(n20957), .b(n20956), .o(n20958) );
no02f01 g17170 ( .a(n20958), .b(n20955), .o(n20959) );
no04f01 g17171 ( .a(n20957), .b(n20426), .c(n20956), .d(n20421), .o(n20960) );
no02f01 g17172 ( .a(n20960), .b(n20959), .o(n20961) );
no02f01 g17173 ( .a(n20759), .b(n20756), .o(n20962) );
no02f01 g17174 ( .a(n20851), .b(n20794), .o(n20963) );
na02f01 g17175 ( .a(n20963), .b(n20962), .o(n20964) );
na02f01 g17176 ( .a(n20850), .b(n20847), .o(n20965) );
na02f01 g17177 ( .a(n20763), .b(n20570), .o(n20966) );
na02f01 g17178 ( .a(n20966), .b(n20965), .o(n20967) );
na02f01 g17179 ( .a(n20967), .b(n20964), .o(n20968) );
na02f01 g17180 ( .a(n20968), .b(n20961), .o(n20969) );
in01f01 g17181 ( .a(n20969), .o(n20970) );
no02f01 g17182 ( .a(n20966), .b(n20965), .o(n20971) );
no02f01 g17183 ( .a(n20963), .b(n20962), .o(n20972) );
no02f01 g17184 ( .a(n20972), .b(n20971), .o(n20973) );
oa12f01 g17185 ( .a(n20973), .b(n20960), .c(n20959), .o(n20974) );
no02f01 g17186 ( .a(n20424), .b(n18460), .o(n20975) );
no02f01 g17187 ( .a(n20975), .b(n20420), .o(n20976) );
no02f01 g17188 ( .a(n20338), .b(n20315), .o(n20977) );
na02f01 g17189 ( .a(n20977), .b(n20976), .o(n20978) );
oa22f01 g17190 ( .a(n20338), .b(n20315), .c(n20975), .d(n20420), .o(n20979) );
na02f01 g17191 ( .a(n20979), .b(n20978), .o(n20980) );
oa12f01 g17192 ( .a(n20758), .b(n20750), .c(n20744), .o(n20981) );
no02f01 g17193 ( .a(n20848), .b(n20755), .o(n20982) );
in01f01 g17194 ( .a(n20982), .o(n20983) );
no02f01 g17195 ( .a(n20983), .b(n20981), .o(n20984) );
ao12f01 g17196 ( .a(n20849), .b(n20843), .c(n20839), .o(n20985) );
no02f01 g17197 ( .a(n20982), .b(n20985), .o(n20986) );
no02f01 g17198 ( .a(n20986), .b(n20984), .o(n20987) );
na02f01 g17199 ( .a(n20987), .b(n20980), .o(n20988) );
in01f01 g17200 ( .a(n20988), .o(n20989) );
na02f01 g17201 ( .a(n20982), .b(n20985), .o(n20990) );
na02f01 g17202 ( .a(n20983), .b(n20981), .o(n20991) );
na02f01 g17203 ( .a(n20991), .b(n20990), .o(n20992) );
na03f01 g17204 ( .a(n20992), .b(n20979), .c(n20978), .o(n20993) );
no04f01 g17205 ( .a(n20338), .b(n20418), .c(n20414), .d(n20165), .o(n20994) );
in01f01 g17206 ( .a(n20165), .o(n20995) );
ao22f01 g17207 ( .a(n20425), .b(n20995), .c(n20314), .d(n20297), .o(n20996) );
no02f01 g17208 ( .a(n20996), .b(n20994), .o(n20997) );
na02f01 g17209 ( .a(n20758), .b(n20843), .o(n20998) );
no02f01 g17210 ( .a(n20998), .b(n20839), .o(n20999) );
ao12f01 g17211 ( .a(n20744), .b(n20758), .c(n20843), .o(n21000) );
no02f01 g17212 ( .a(n21000), .b(n20999), .o(n21001) );
in01f01 g17213 ( .a(n21001), .o(n21002) );
na02f01 g17214 ( .a(n21002), .b(n20997), .o(n21003) );
ao12f01 g17215 ( .a(n20989), .b(n21003), .c(n20993), .o(n21004) );
ao12f01 g17216 ( .a(n20970), .b(n21004), .c(n20974), .o(n21005) );
ao12f01 g17217 ( .a(n20951), .b(n21005), .c(n20954), .o(n21006) );
in01f01 g17218 ( .a(n21006), .o(n21007) );
in01f01 g17219 ( .a(n20951), .o(n21008) );
no02f01 g17220 ( .a(n20172), .b(n18459), .o(n21009) );
no02f01 g17221 ( .a(n20172), .b(n18460), .o(n21010) );
no02f01 g17222 ( .a(n21010), .b(n21009), .o(n21011) );
no02f01 g17223 ( .a(n20308), .b(n20415), .o(n21012) );
oa12f01 g17224 ( .a(n21012), .b(n20292), .c(n20180), .o(n21013) );
in01f01 g17225 ( .a(n21013), .o(n21014) );
ao12f01 g17226 ( .a(n20295), .b(n21014), .c(n20312), .o(n21015) );
in01f01 g17227 ( .a(n21015), .o(n21016) );
no02f01 g17228 ( .a(n21016), .b(n21011), .o(n21017) );
in01f01 g17229 ( .a(n21011), .o(n21018) );
no02f01 g17230 ( .a(n21015), .b(n21018), .o(n21019) );
no02f01 g17231 ( .a(n21019), .b(n21017), .o(n21020) );
ao12f01 g17232 ( .a(n20741), .b(n20740), .c(n20586), .o(n21021) );
in01f01 g17233 ( .a(n21021), .o(n21022) );
na03f01 g17234 ( .a(n21022), .b(n20743), .c(n20797), .o(n21023) );
oa12f01 g17235 ( .a(n21021), .b(n20838), .c(n20579), .o(n21024) );
na02f01 g17236 ( .a(n21024), .b(n21023), .o(n21025) );
no02f01 g17237 ( .a(n21025), .b(n21020), .o(n21026) );
no02f01 g17238 ( .a(n20738), .b(n20595), .o(n21027) );
no02f01 g17239 ( .a(n20831), .b(n20607), .o(n21028) );
oa12f01 g17240 ( .a(n20736), .b(n21028), .c(n20599), .o(n21029) );
no02f01 g17241 ( .a(n21029), .b(n21027), .o(n21030) );
in01f01 g17242 ( .a(n21030), .o(n21031) );
na02f01 g17243 ( .a(n21029), .b(n21027), .o(n21032) );
na02f01 g17244 ( .a(n21032), .b(n21031), .o(n21033) );
in01f01 g17245 ( .a(n21033), .o(n21034) );
no02f01 g17246 ( .a(n20405), .b(n20402), .o(n21035) );
no02f01 g17247 ( .a(n20408), .b(n20186), .o(n21036) );
no02f01 g17248 ( .a(n21036), .b(n21035), .o(n21037) );
na02f01 g17249 ( .a(n21036), .b(n21035), .o(n21038) );
in01f01 g17250 ( .a(n21038), .o(n21039) );
no02f01 g17251 ( .a(n21039), .b(n21037), .o(n21040) );
in01f01 g17252 ( .a(n21040), .o(n21041) );
no02f01 g17253 ( .a(n20830), .b(n20614), .o(n21042) );
no02f01 g17254 ( .a(n20732), .b(n20607), .o(n21043) );
na02f01 g17255 ( .a(n21043), .b(n21042), .o(n21044) );
no02f01 g17256 ( .a(n21043), .b(n21042), .o(n21045) );
in01f01 g17257 ( .a(n21045), .o(n21046) );
na02f01 g17258 ( .a(n21046), .b(n21044), .o(n21047) );
in01f01 g17259 ( .a(n21047), .o(n21048) );
no02f01 g17260 ( .a(n21048), .b(n21041), .o(n21049) );
in01f01 g17261 ( .a(n21049), .o(n21050) );
no02f01 g17262 ( .a(n20279), .b(n20278), .o(n21051) );
oa12f01 g17263 ( .a(n21051), .b(n20401), .c(n20400), .o(n21052) );
in01f01 g17264 ( .a(n21052), .o(n21053) );
no02f01 g17265 ( .a(n20282), .b(n20373), .o(n21054) );
no02f01 g17266 ( .a(n21054), .b(n21053), .o(n21055) );
in01f01 g17267 ( .a(n21055), .o(n21056) );
na02f01 g17268 ( .a(n21054), .b(n21053), .o(n21057) );
na02f01 g17269 ( .a(n21057), .b(n21056), .o(n21058) );
no02f01 g17270 ( .a(n20828), .b(n20620), .o(n21059) );
no02f01 g17271 ( .a(n20829), .b(n20614), .o(n21060) );
in01f01 g17272 ( .a(n21060), .o(n21061) );
no02f01 g17273 ( .a(n21061), .b(n21059), .o(n21062) );
na02f01 g17274 ( .a(n21061), .b(n21059), .o(n21063) );
in01f01 g17275 ( .a(n21063), .o(n21064) );
no02f01 g17276 ( .a(n21064), .b(n21062), .o(n21065) );
no02f01 g17277 ( .a(n21065), .b(n21058), .o(n21066) );
no02f01 g17278 ( .a(n20279), .b(n20268), .o(n21067) );
no02f01 g17279 ( .a(n20278), .b(n20401), .o(n21068) );
no02f01 g17280 ( .a(n21068), .b(n21067), .o(n21069) );
na02f01 g17281 ( .a(n21068), .b(n21067), .o(n21070) );
in01f01 g17282 ( .a(n21070), .o(n21071) );
no02f01 g17283 ( .a(n21071), .b(n21069), .o(n21072) );
ao12f01 g17284 ( .a(n20724), .b(n20825), .c(n20824), .o(n21073) );
no02f01 g17285 ( .a(n20727), .b(n20620), .o(n21074) );
na02f01 g17286 ( .a(n21074), .b(n21073), .o(n21075) );
in01f01 g17287 ( .a(n21075), .o(n21076) );
no02f01 g17288 ( .a(n21074), .b(n21073), .o(n21077) );
no02f01 g17289 ( .a(n21077), .b(n21076), .o(n21078) );
in01f01 g17290 ( .a(n21078), .o(n21079) );
na02f01 g17291 ( .a(n21079), .b(n21072), .o(n21080) );
no02f01 g17292 ( .a(n20259), .b(n20200), .o(n21081) );
no02f01 g17293 ( .a(n20279), .b(n20267), .o(n21082) );
in01f01 g17294 ( .a(n21082), .o(n21083) );
no02f01 g17295 ( .a(n21083), .b(n21081), .o(n21084) );
in01f01 g17296 ( .a(n21084), .o(n21085) );
na02f01 g17297 ( .a(n21083), .b(n21081), .o(n21086) );
na02f01 g17298 ( .a(n21086), .b(n21085), .o(n21087) );
no02f01 g17299 ( .a(n20724), .b(n20722), .o(n21088) );
no02f01 g17300 ( .a(n21088), .b(n20718), .o(n21089) );
na02f01 g17301 ( .a(n21088), .b(n20718), .o(n21090) );
in01f01 g17302 ( .a(n21090), .o(n21091) );
no02f01 g17303 ( .a(n21091), .b(n21089), .o(n21092) );
no02f01 g17304 ( .a(n21092), .b(n21087), .o(n21093) );
no02f01 g17305 ( .a(n20249), .b(n20388), .o(n21094) );
ao12f01 g17306 ( .a(n20256), .b(n20394), .c(n21094), .o(n21095) );
in01f01 g17307 ( .a(n21095), .o(n21096) );
na03f01 g17308 ( .a(n21096), .b(n20378), .c(n20374), .o(n21097) );
oa12f01 g17309 ( .a(n21095), .b(n20201), .c(n20200), .o(n21098) );
ao12f01 g17310 ( .a(n20714), .b(n20713), .c(n20636), .o(n21099) );
no02f01 g17311 ( .a(n20716), .b(n20626), .o(n21100) );
in01f01 g17312 ( .a(n21100), .o(n21101) );
no02f01 g17313 ( .a(n21101), .b(n21099), .o(n21102) );
na02f01 g17314 ( .a(n21101), .b(n21099), .o(n21103) );
in01f01 g17315 ( .a(n21103), .o(n21104) );
no02f01 g17316 ( .a(n21104), .b(n21102), .o(n21105) );
in01f01 g17317 ( .a(n21105), .o(n21106) );
ao12f01 g17318 ( .a(n21106), .b(n21098), .c(n21097), .o(n21107) );
no02f01 g17319 ( .a(n20247), .b(n18460), .o(n21108) );
no02f01 g17320 ( .a(n20236), .b(n18460), .o(n21109) );
no04f01 g17321 ( .a(n21109), .b(n21108), .c(n20387), .d(n20238), .o(n21110) );
no02f01 g17322 ( .a(n21109), .b(n20238), .o(n21111) );
no02f01 g17323 ( .a(n21108), .b(n20387), .o(n21112) );
no02f01 g17324 ( .a(n21112), .b(n21111), .o(n21113) );
no02f01 g17325 ( .a(n20711), .b(n20648), .o(n21114) );
no02f01 g17326 ( .a(n21114), .b(n20820), .o(n21115) );
na02f01 g17327 ( .a(n21114), .b(n20820), .o(n21116) );
in01f01 g17328 ( .a(n21116), .o(n21117) );
no02f01 g17329 ( .a(n21117), .b(n21115), .o(n21118) );
no03f01 g17330 ( .a(n21118), .b(n21113), .c(n21110), .o(n21119) );
no02f01 g17331 ( .a(n21109), .b(n20237), .o(n21120) );
no02f01 g17332 ( .a(n21120), .b(n20231), .o(n21121) );
in01f01 g17333 ( .a(n21121), .o(n21122) );
na02f01 g17334 ( .a(n21120), .b(n20231), .o(n21123) );
na02f01 g17335 ( .a(n21123), .b(n21122), .o(n21124) );
no02f01 g17336 ( .a(n20709), .b(n20806), .o(n21125) );
no02f01 g17337 ( .a(n21125), .b(n20708), .o(n21126) );
na02f01 g17338 ( .a(n21125), .b(n20708), .o(n21127) );
in01f01 g17339 ( .a(n21127), .o(n21128) );
no02f01 g17340 ( .a(n21128), .b(n21126), .o(n21129) );
no02f01 g17341 ( .a(n21129), .b(n21124), .o(n21130) );
in01f01 g17342 ( .a(n21130), .o(n21131) );
in01f01 g17343 ( .a(n20223), .o(n21132) );
no02f01 g17344 ( .a(n20379), .b(n18460), .o(n21133) );
no02f01 g17345 ( .a(n21133), .b(n20380), .o(n21134) );
na02f01 g17346 ( .a(n21134), .b(n21132), .o(n21135) );
oa12f01 g17347 ( .a(n20223), .b(n21133), .c(n20380), .o(n21136) );
na02f01 g17348 ( .a(n21136), .b(n21135), .o(n21137) );
no03f01 g17349 ( .a(n20817), .b(n20706), .c(n20670), .o(n21138) );
ao12f01 g17350 ( .a(n20816), .b(n20707), .c(n20810), .o(n21139) );
no02f01 g17351 ( .a(n21139), .b(n21138), .o(n21140) );
no02f01 g17352 ( .a(n21140), .b(n21137), .o(n21141) );
in01f01 g17353 ( .a(n21141), .o(n21142) );
in01f01 g17354 ( .a(n20215), .o(n21143) );
oa12f01 g17355 ( .a(n18459), .b(n20220), .c(n20219), .o(n21144) );
in01f01 g17356 ( .a(n21144), .o(n21145) );
oa12f01 g17357 ( .a(n21143), .b(n21145), .c(n20222), .o(n21146) );
in01f01 g17358 ( .a(n20222), .o(n21147) );
na03f01 g17359 ( .a(n21144), .b(n21147), .c(n20215), .o(n21148) );
na02f01 g17360 ( .a(n21148), .b(n21146), .o(n21149) );
no03f01 g17361 ( .a(n20704), .b(n20702), .c(n20814), .o(n21150) );
ao12f01 g17362 ( .a(n20691), .b(n20705), .c(n20815), .o(n21151) );
no02f01 g17363 ( .a(n21151), .b(n21150), .o(n21152) );
na02f01 g17364 ( .a(n21152), .b(n21149), .o(n21153) );
in01f01 g17365 ( .a(n20207), .o(n21154) );
no02f01 g17366 ( .a(n21154), .b(n18460), .o(n21155) );
no02f01 g17367 ( .a(n21154), .b(n18459), .o(n21156) );
no02f01 g17368 ( .a(n21156), .b(n21155), .o(n21157) );
no02f01 g17369 ( .a(n20674), .b(n19835), .o(n21158) );
na02f01 g17370 ( .a(n20674), .b(n19835), .o(n21159) );
in01f01 g17371 ( .a(n21159), .o(n21160) );
no02f01 g17372 ( .a(n21160), .b(n21158), .o(n21161) );
in01f01 g17373 ( .a(n21161), .o(n21162) );
na02f01 g17374 ( .a(n21162), .b(n21157), .o(n21163) );
no03f01 g17375 ( .a(n20686), .b(n20684), .c(n20682), .o(n21164) );
no02f01 g17376 ( .a(n20687), .b(n20688), .o(n21165) );
no02f01 g17377 ( .a(n21165), .b(n21164), .o(n21166) );
no02f01 g17378 ( .a(n21166), .b(n20675), .o(n21167) );
na02f01 g17379 ( .a(n21166), .b(n20675), .o(n21168) );
in01f01 g17380 ( .a(n21168), .o(n21169) );
no02f01 g17381 ( .a(n21169), .b(n21167), .o(n21170) );
in01f01 g17382 ( .a(n21170), .o(n21171) );
na02f01 g17383 ( .a(n21171), .b(n21163), .o(n21172) );
no04f01 g17384 ( .a(n20213), .b(n20211), .c(n20207), .d(n18459), .o(n21173) );
ao12f01 g17385 ( .a(n20214), .b(n21154), .c(n18460), .o(n21174) );
no02f01 g17386 ( .a(n21174), .b(n21173), .o(n21175) );
oa12f01 g17387 ( .a(n21175), .b(n21171), .c(n21163), .o(n21176) );
na02f01 g17388 ( .a(n21176), .b(n21172), .o(n21177) );
na02f01 g17389 ( .a(n21177), .b(n21153), .o(n21178) );
in01f01 g17390 ( .a(n21152), .o(n21179) );
na03f01 g17391 ( .a(n21179), .b(n21148), .c(n21146), .o(n21180) );
na02f01 g17392 ( .a(n21180), .b(n21178), .o(n21181) );
na02f01 g17393 ( .a(n21140), .b(n21137), .o(n21182) );
na02f01 g17394 ( .a(n21182), .b(n21181), .o(n21183) );
na02f01 g17395 ( .a(n21183), .b(n21142), .o(n21184) );
na02f01 g17396 ( .a(n21129), .b(n21124), .o(n21185) );
na02f01 g17397 ( .a(n21185), .b(n21184), .o(n21186) );
no02f01 g17398 ( .a(n21113), .b(n21110), .o(n21187) );
in01f01 g17399 ( .a(n21118), .o(n21188) );
no02f01 g17400 ( .a(n21188), .b(n21187), .o(n21189) );
ao12f01 g17401 ( .a(n21189), .b(n21186), .c(n21131), .o(n21190) );
no02f01 g17402 ( .a(n20258), .b(n20256), .o(n21191) );
no02f01 g17403 ( .a(n21191), .b(n21094), .o(n21192) );
in01f01 g17404 ( .a(n21192), .o(n21193) );
na02f01 g17405 ( .a(n21191), .b(n21094), .o(n21194) );
na02f01 g17406 ( .a(n21194), .b(n21193), .o(n21195) );
no03f01 g17407 ( .a(n20714), .b(n20821), .c(n20803), .o(n21196) );
ao12f01 g17408 ( .a(n20713), .b(n20822), .c(n20636), .o(n21197) );
no02f01 g17409 ( .a(n21197), .b(n21196), .o(n21198) );
na02f01 g17410 ( .a(n21198), .b(n21195), .o(n21199) );
oa12f01 g17411 ( .a(n21199), .b(n21190), .c(n21119), .o(n21200) );
na02f01 g17412 ( .a(n21098), .b(n21097), .o(n21201) );
no02f01 g17413 ( .a(n21105), .b(n21201), .o(n21202) );
no02f01 g17414 ( .a(n21198), .b(n21195), .o(n21203) );
no02f01 g17415 ( .a(n21203), .b(n21202), .o(n21204) );
ao12f01 g17416 ( .a(n21107), .b(n21204), .c(n21200), .o(n21205) );
na02f01 g17417 ( .a(n21092), .b(n21087), .o(n21206) );
ao12f01 g17418 ( .a(n21093), .b(n21206), .c(n21205), .o(n21207) );
no02f01 g17419 ( .a(n21079), .b(n21072), .o(n21208) );
oa12f01 g17420 ( .a(n21080), .b(n21208), .c(n21207), .o(n21209) );
na02f01 g17421 ( .a(n21065), .b(n21058), .o(n21210) );
ao12f01 g17422 ( .a(n21066), .b(n21210), .c(n21209), .o(n21211) );
no02f01 g17423 ( .a(n21047), .b(n21040), .o(n21212) );
oa12f01 g17424 ( .a(n21050), .b(n21212), .c(n21211), .o(n21213) );
na02f01 g17425 ( .a(n20285), .b(n20187), .o(n21214) );
no02f01 g17426 ( .a(n20308), .b(n20410), .o(n21215) );
no02f01 g17427 ( .a(n21215), .b(n21214), .o(n21216) );
na02f01 g17428 ( .a(n21215), .b(n21214), .o(n21217) );
in01f01 g17429 ( .a(n21217), .o(n21218) );
no02f01 g17430 ( .a(n21218), .b(n21216), .o(n21219) );
no02f01 g17431 ( .a(n20735), .b(n20599), .o(n21220) );
in01f01 g17432 ( .a(n21220), .o(n21221) );
no02f01 g17433 ( .a(n21221), .b(n21028), .o(n21222) );
na02f01 g17434 ( .a(n21221), .b(n21028), .o(n21223) );
in01f01 g17435 ( .a(n21223), .o(n21224) );
no02f01 g17436 ( .a(n21224), .b(n21222), .o(n21225) );
in01f01 g17437 ( .a(n21225), .o(n21226) );
no02f01 g17438 ( .a(n21226), .b(n21219), .o(n21227) );
in01f01 g17439 ( .a(n21227), .o(n21228) );
na02f01 g17440 ( .a(n21226), .b(n21219), .o(n21229) );
in01f01 g17441 ( .a(n21229), .o(n21230) );
ao12f01 g17442 ( .a(n21230), .b(n21228), .c(n21213), .o(n21231) );
na02f01 g17443 ( .a(n20309), .b(n21214), .o(n21232) );
na02f01 g17444 ( .a(n21232), .b(n20291), .o(n21233) );
no02f01 g17445 ( .a(n20415), .b(n20180), .o(n21234) );
no02f01 g17446 ( .a(n21234), .b(n21233), .o(n21235) );
na02f01 g17447 ( .a(n21234), .b(n21233), .o(n21236) );
in01f01 g17448 ( .a(n21236), .o(n21237) );
no02f01 g17449 ( .a(n21237), .b(n21235), .o(n21238) );
in01f01 g17450 ( .a(n21238), .o(n21239) );
no02f01 g17451 ( .a(n21230), .b(n21033), .o(n21240) );
in01f01 g17452 ( .a(n21240), .o(n21241) );
ao12f01 g17453 ( .a(n21241), .b(n21228), .c(n21213), .o(n21242) );
oa22f01 g17454 ( .a(n21242), .b(n21239), .c(n21231), .d(n21034), .o(n21243) );
no02f01 g17455 ( .a(n20416), .b(n20295), .o(n21244) );
in01f01 g17456 ( .a(n21244), .o(n21245) );
no02f01 g17457 ( .a(n21245), .b(n21013), .o(n21246) );
no02f01 g17458 ( .a(n21244), .b(n21014), .o(n21247) );
no02f01 g17459 ( .a(n21247), .b(n21246), .o(n21248) );
na02f01 g17460 ( .a(n20836), .b(n20586), .o(n21249) );
no02f01 g17461 ( .a(n21249), .b(n20835), .o(n21250) );
ao12f01 g17462 ( .a(n20740), .b(n20836), .c(n20586), .o(n21251) );
no02f01 g17463 ( .a(n21251), .b(n21250), .o(n21252) );
in01f01 g17464 ( .a(n21252), .o(n21253) );
no02f01 g17465 ( .a(n21253), .b(n21248), .o(n21254) );
in01f01 g17466 ( .a(n21254), .o(n21255) );
na02f01 g17467 ( .a(n21025), .b(n21020), .o(n21256) );
na02f01 g17468 ( .a(n21253), .b(n21248), .o(n21257) );
na02f01 g17469 ( .a(n21257), .b(n21256), .o(n21258) );
ao12f01 g17470 ( .a(n21258), .b(n21255), .c(n21243), .o(n21259) );
no02f01 g17471 ( .a(n21002), .b(n20997), .o(n21260) );
no04f01 g17472 ( .a(n21260), .b(n21259), .c(n21026), .d(n20989), .o(n21261) );
na03f01 g17473 ( .a(n21261), .b(n20974), .c(n21008), .o(n21262) );
ao12f01 g17474 ( .a(n20933), .b(n21262), .c(n21007), .o(n21263) );
no02f01 g17475 ( .a(n21263), .b(n20923), .o(n21264) );
no02f01 g17476 ( .a(n20367), .b(n20366), .o(n21265) );
no02f01 g17477 ( .a(n21265), .b(n18460), .o(n21266) );
in01f01 g17478 ( .a(n21266), .o(n21267) );
na02f01 g17479 ( .a(n20363), .b(n20877), .o(n21268) );
na04f01 g17480 ( .a(n21268), .b(n20361), .c(n20369), .d(n20368), .o(n21269) );
na02f01 g17481 ( .a(n21269), .b(n21267), .o(n21270) );
na03f01 g17482 ( .a(n20542), .b(n20493), .c(n20503), .o(n21271) );
na04f01 g17483 ( .a(n21271), .b(n20540), .c(n20496), .d(n20502), .o(n21272) );
na02f01 g17484 ( .a(n19534), .b(n18103), .o(n21273) );
na02f01 g17485 ( .a(n19534), .b(n18145), .o(n21274) );
na02f01 g17486 ( .a(n21274), .b(n21273), .o(n21275) );
no02f01 g17487 ( .a(n21275), .b(n21272), .o(n21276) );
no03f01 g17488 ( .a(n20500), .b(n20539), .c(n20443), .o(n21277) );
no04f01 g17489 ( .a(n21277), .b(n20498), .c(n20497), .d(n20442), .o(n21278) );
no02f01 g17490 ( .a(n19530), .b(n18145), .o(n21279) );
no02f01 g17491 ( .a(n19530), .b(n18103), .o(n21280) );
no02f01 g17492 ( .a(n21280), .b(n21279), .o(n21281) );
no02f01 g17493 ( .a(n21281), .b(n21278), .o(n21282) );
no02f01 g17494 ( .a(n21282), .b(n21276), .o(n21283) );
no02f01 g17495 ( .a(n21283), .b(n19565), .o(n21284) );
na02f01 g17496 ( .a(n21281), .b(n21278), .o(n21285) );
na02f01 g17497 ( .a(n21275), .b(n21272), .o(n21286) );
na02f01 g17498 ( .a(n21286), .b(n21285), .o(n21287) );
no02f01 g17499 ( .a(n21287), .b(n19059), .o(n21288) );
no02f01 g17500 ( .a(n21288), .b(n21284), .o(n21289) );
ao12f01 g17501 ( .a(n20791), .b(n20785), .c(n20782), .o(n21290) );
na02f01 g17502 ( .a(n20556), .b(n20544), .o(n21291) );
oa12f01 g17503 ( .a(n20547), .b(n21291), .c(n21290), .o(n21292) );
no02f01 g17504 ( .a(n21292), .b(n21289), .o(n21293) );
na02f01 g17505 ( .a(n21287), .b(n19059), .o(n21294) );
na02f01 g17506 ( .a(n21283), .b(n19565), .o(n21295) );
na02f01 g17507 ( .a(n21295), .b(n21294), .o(n21296) );
oa12f01 g17508 ( .a(n20553), .b(n20864), .c(n20861), .o(n21297) );
no02f01 g17509 ( .a(n20792), .b(n20788), .o(n21298) );
ao12f01 g17510 ( .a(n20789), .b(n21298), .c(n21297), .o(n21299) );
no02f01 g17511 ( .a(n21299), .b(n21296), .o(n21300) );
no02f01 g17512 ( .a(n21300), .b(n21293), .o(n21301) );
no02f01 g17513 ( .a(n21301), .b(n21270), .o(n21302) );
no02f01 g17514 ( .a(n20439), .b(n20874), .o(n21303) );
no04f01 g17515 ( .a(n21303), .b(n20437), .c(n20123), .d(n20122), .o(n21304) );
no02f01 g17516 ( .a(n21304), .b(n21266), .o(n21305) );
na02f01 g17517 ( .a(n21299), .b(n21296), .o(n21306) );
na02f01 g17518 ( .a(n21292), .b(n21289), .o(n21307) );
na02f01 g17519 ( .a(n21307), .b(n21306), .o(n21308) );
no02f01 g17520 ( .a(n21308), .b(n21305), .o(n21309) );
no02f01 g17521 ( .a(n21309), .b(n21302), .o(n21310) );
na02f01 g17522 ( .a(n21310), .b(n21264), .o(n21311) );
in01f01 g17523 ( .a(n20887), .o(n21312) );
ao12f01 g17524 ( .a(n20893), .b(n20892), .c(n20137), .o(n21313) );
no03f01 g17525 ( .a(n20890), .b(n20889), .c(n20371), .o(n21314) );
no03f01 g17526 ( .a(n20901), .b(n20784), .c(n20900), .o(n21315) );
ao12f01 g17527 ( .a(n20897), .b(n20863), .c(n20896), .o(n21316) );
no02f01 g17528 ( .a(n21316), .b(n21315), .o(n21317) );
oa12f01 g17529 ( .a(n21317), .b(n21314), .c(n21313), .o(n21318) );
no03f01 g17530 ( .a(n21317), .b(n21314), .c(n21313), .o(n21319) );
na02f01 g17531 ( .a(n20912), .b(n20910), .o(n21320) );
na02f01 g17532 ( .a(n20908), .b(n20906), .o(n21321) );
na02f01 g17533 ( .a(n21321), .b(n21320), .o(n21322) );
in01f01 g17534 ( .a(n20919), .o(n21323) );
no02f01 g17535 ( .a(n21323), .b(n21322), .o(n21324) );
oa12f01 g17536 ( .a(n21318), .b(n21324), .c(n21319), .o(n21325) );
oa12f01 g17537 ( .a(n21312), .b(n21325), .c(n20930), .o(n21326) );
oa12f01 g17538 ( .a(n20924), .b(n21326), .c(n20872), .o(n21327) );
in01f01 g17539 ( .a(n20931), .o(n21328) );
na03f01 g17540 ( .a(n21328), .b(n21318), .c(n20888), .o(n21329) );
no02f01 g17541 ( .a(n21329), .b(n20869), .o(n21330) );
in01f01 g17542 ( .a(n21261), .o(n21331) );
na02f01 g17543 ( .a(n20974), .b(n21008), .o(n21332) );
no02f01 g17544 ( .a(n21332), .b(n21331), .o(n21333) );
oa12f01 g17545 ( .a(n21330), .b(n21333), .c(n21006), .o(n21334) );
na02f01 g17546 ( .a(n21334), .b(n21327), .o(n21335) );
in01f01 g17547 ( .a(n21310), .o(n21336) );
na02f01 g17548 ( .a(n21336), .b(n21335), .o(n21337) );
na02f01 g17549 ( .a(n21337), .b(n21311), .o(n273) );
no02f01 g17550 ( .a(n16326), .b(n16236), .o(n21339) );
no02f01 g17551 ( .a(n16435), .b(n21339), .o(n21340) );
no02f01 g17552 ( .a(n16354), .b(n16329), .o(n21341) );
no02f01 g17553 ( .a(n21341), .b(n16356), .o(n21342) );
na02f01 g17554 ( .a(n21342), .b(n21340), .o(n21343) );
in01f01 g17555 ( .a(n21342), .o(n21344) );
oa12f01 g17556 ( .a(n21344), .b(n16435), .c(n21339), .o(n21345) );
na02f01 g17557 ( .a(n21345), .b(n21343), .o(n278) );
na02f01 g17558 ( .a(n15993), .b(n15989), .o(n21347) );
na02f01 g17559 ( .a(n15977), .b(n15948), .o(n21348) );
in01f01 g17560 ( .a(n16055), .o(n21349) );
na03f01 g17561 ( .a(n21349), .b(n21348), .c(n21347), .o(n21350) );
ao12f01 g17562 ( .a(n15988), .b(n16059), .c(n15924), .o(n21351) );
no03f01 g17563 ( .a(n16057), .b(n15947), .c(n15981), .o(n21352) );
no03f01 g17564 ( .a(n16067), .b(n21352), .c(n21351), .o(n21353) );
oa12f01 g17565 ( .a(n16067), .b(n21352), .c(n21351), .o(n21354) );
oa12f01 g17566 ( .a(n15946), .b(n15984), .c(n15949), .o(n21355) );
na03f01 g17567 ( .a(n15987), .b(n15941), .c(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .o(n21356) );
in01f01 g17568 ( .a(n16075), .o(n21357) );
ao12f01 g17569 ( .a(n21357), .b(n21356), .c(n21355), .o(n21358) );
no02f01 g17570 ( .a(n15941), .b(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .o(n21359) );
no02f01 g17571 ( .a(n15941), .b(n15949), .o(n21360) );
no03f01 g17572 ( .a(n16082), .b(n21360), .c(n21359), .o(n21361) );
na03f01 g17573 ( .a(n21357), .b(n21356), .c(n21355), .o(n21362) );
oa12f01 g17574 ( .a(n21362), .b(n21361), .c(n21358), .o(n21363) );
ao12f01 g17575 ( .a(n21353), .b(n21363), .c(n21354), .o(n21364) );
ao12f01 g17576 ( .a(n21349), .b(n21348), .c(n21347), .o(n21365) );
oa12f01 g17577 ( .a(n21350), .b(n21365), .c(n21364), .o(n21366) );
na02f01 g17578 ( .a(n16182), .b(n16329), .o(n21367) );
oa12f01 g17579 ( .a(n16329), .b(n16227), .c(n16208), .o(n21368) );
na04f01 g17580 ( .a(n21368), .b(n21367), .c(n16149), .d(n21366), .o(n21369) );
in01f01 g17581 ( .a(n16235), .o(n21370) );
na02f01 g17582 ( .a(n21370), .b(n21369), .o(n21371) );
na04f01 g17583 ( .a(n16426), .b(n16380), .c(n16325), .d(n21371), .o(n21372) );
in01f01 g17584 ( .a(n16440), .o(n21373) );
na02f01 g17585 ( .a(n21373), .b(n21372), .o(n21374) );
in01f01 g17586 ( .a(n16488), .o(n21375) );
no02f01 g17587 ( .a(n16542), .b(n16512), .o(n21376) );
no03f01 g17588 ( .a(n16532), .b(n16504), .c(n16491), .o(n21377) );
in01f01 g17589 ( .a(n21377), .o(n21378) );
no02f01 g17590 ( .a(n21378), .b(n16481), .o(n21379) );
ao12f01 g17591 ( .a(n16193), .b(n16530), .c(n16502), .o(n21380) );
no02f01 g17592 ( .a(n21380), .b(n16493), .o(n21381) );
in01f01 g17593 ( .a(n21381), .o(n21382) );
no02f01 g17594 ( .a(n14732), .b(n14714), .o(n21383) );
na02f01 g17595 ( .a(n14992), .b(n15099), .o(n21384) );
na02f01 g17596 ( .a(n21384), .b(n21383), .o(n21385) );
no02f01 g17597 ( .a(n14772), .b(n14553), .o(n21386) );
no02f01 g17598 ( .a(n14771), .b(n14552), .o(n21387) );
no02f01 g17599 ( .a(n21387), .b(n21386), .o(n21388) );
in01f01 g17600 ( .a(n21388), .o(n21389) );
no02f01 g17601 ( .a(n21389), .b(n21385), .o(n21390) );
ao12f01 g17602 ( .a(n21388), .b(n21384), .c(n21383), .o(n21391) );
no02f01 g17603 ( .a(n21391), .b(n21390), .o(n21392) );
no02f01 g17604 ( .a(n21392), .b(n16193), .o(n21393) );
na02f01 g17605 ( .a(n21392), .b(n16193), .o(n21394) );
in01f01 g17606 ( .a(n21394), .o(n21395) );
no02f01 g17607 ( .a(n21395), .b(n21393), .o(n21396) );
in01f01 g17608 ( .a(n21396), .o(n21397) );
no03f01 g17609 ( .a(n21397), .b(n21382), .c(n21379), .o(n21398) );
no02f01 g17610 ( .a(n21382), .b(n21379), .o(n21399) );
no02f01 g17611 ( .a(n21396), .b(n21399), .o(n21400) );
no02f01 g17612 ( .a(n21400), .b(n21398), .o(n21401) );
in01f01 g17613 ( .a(n21401), .o(n21402) );
no02f01 g17614 ( .a(n21402), .b(n16155), .o(n21403) );
na02f01 g17615 ( .a(n21394), .b(n21379), .o(n21404) );
no02f01 g17616 ( .a(n21393), .b(n21382), .o(n21405) );
na02f01 g17617 ( .a(n21405), .b(n21404), .o(n21406) );
in01f01 g17618 ( .a(n21386), .o(n21407) );
ao12f01 g17619 ( .a(n21387), .b(n21407), .c(n21385), .o(n21408) );
no02f01 g17620 ( .a(n14765), .b(n14553), .o(n21409) );
no02f01 g17621 ( .a(n14764), .b(n14552), .o(n21410) );
no02f01 g17622 ( .a(n21410), .b(n21409), .o(n21411) );
no02f01 g17623 ( .a(n21411), .b(n21408), .o(n21412) );
na02f01 g17624 ( .a(n21411), .b(n21408), .o(n21413) );
in01f01 g17625 ( .a(n21413), .o(n21414) );
no02f01 g17626 ( .a(n21414), .b(n21412), .o(n21415) );
in01f01 g17627 ( .a(n21415), .o(n21416) );
no02f01 g17628 ( .a(n21416), .b(n16194), .o(n21417) );
no02f01 g17629 ( .a(n21415), .b(n16193), .o(n21418) );
no02f01 g17630 ( .a(n21418), .b(n21417), .o(n21419) );
in01f01 g17631 ( .a(n21419), .o(n21420) );
no02f01 g17632 ( .a(n21420), .b(n21406), .o(n21421) );
na02f01 g17633 ( .a(n21420), .b(n21406), .o(n21422) );
in01f01 g17634 ( .a(n21422), .o(n21423) );
no02f01 g17635 ( .a(n21423), .b(n21421), .o(n21424) );
in01f01 g17636 ( .a(n21424), .o(n21425) );
no02f01 g17637 ( .a(n21425), .b(n16155), .o(n21426) );
no02f01 g17638 ( .a(n21426), .b(n21403), .o(n21427) );
na04f01 g17639 ( .a(n21427), .b(n21376), .c(n21375), .d(n21374), .o(n21428) );
in01f01 g17640 ( .a(n14996), .o(n21429) );
ao12f01 g17641 ( .a(n14552), .b(n14771), .c(n14764), .o(n21430) );
ao12f01 g17642 ( .a(n21430), .b(n21385), .c(n21429), .o(n21431) );
no02f01 g17643 ( .a(n14742), .b(n14552), .o(n21432) );
no02f01 g17644 ( .a(n14994), .b(n21432), .o(n21433) );
no02f01 g17645 ( .a(n21433), .b(n21431), .o(n21434) );
na02f01 g17646 ( .a(n21433), .b(n21431), .o(n21435) );
in01f01 g17647 ( .a(n21435), .o(n21436) );
no02f01 g17648 ( .a(n21436), .b(n21434), .o(n21437) );
in01f01 g17649 ( .a(n21437), .o(n21438) );
no02f01 g17650 ( .a(n21438), .b(n16194), .o(n21439) );
ao12f01 g17651 ( .a(n16193), .b(n21415), .c(n21392), .o(n21440) );
no02f01 g17652 ( .a(n21440), .b(n21382), .o(n21441) );
oa12f01 g17653 ( .a(n21441), .b(n21417), .c(n21404), .o(n21442) );
no02f01 g17654 ( .a(n21437), .b(n16193), .o(n21443) );
no02f01 g17655 ( .a(n21443), .b(n21442), .o(n21444) );
no02f01 g17656 ( .a(n21444), .b(n21439), .o(n21445) );
in01f01 g17657 ( .a(n21445), .o(n21446) );
in01f01 g17658 ( .a(n21431), .o(n21447) );
oa12f01 g17659 ( .a(n14993), .b(n21447), .c(n21432), .o(n21448) );
in01f01 g17660 ( .a(n21448), .o(n21449) );
no02f01 g17661 ( .a(n14752), .b(n14552), .o(n21450) );
no02f01 g17662 ( .a(n21450), .b(n14997), .o(n21451) );
in01f01 g17663 ( .a(n21451), .o(n21452) );
no02f01 g17664 ( .a(n21452), .b(n21449), .o(n21453) );
no02f01 g17665 ( .a(n21451), .b(n21448), .o(n21454) );
no02f01 g17666 ( .a(n21454), .b(n21453), .o(n21455) );
in01f01 g17667 ( .a(n21455), .o(n21456) );
no02f01 g17668 ( .a(n21456), .b(n16194), .o(n21457) );
no02f01 g17669 ( .a(n21455), .b(n16193), .o(n21458) );
no02f01 g17670 ( .a(n21458), .b(n21457), .o(n21459) );
no02f01 g17671 ( .a(n21459), .b(n21446), .o(n21460) );
na02f01 g17672 ( .a(n21459), .b(n21446), .o(n21461) );
in01f01 g17673 ( .a(n21461), .o(n21462) );
no02f01 g17674 ( .a(n21462), .b(n21460), .o(n21463) );
in01f01 g17675 ( .a(n21463), .o(n21464) );
no02f01 g17676 ( .a(n21464), .b(n16155), .o(n21465) );
in01f01 g17677 ( .a(n21442), .o(n21466) );
no02f01 g17678 ( .a(n21443), .b(n21439), .o(n21467) );
no02f01 g17679 ( .a(n21467), .b(n21466), .o(n21468) );
na02f01 g17680 ( .a(n21467), .b(n21466), .o(n21469) );
in01f01 g17681 ( .a(n21469), .o(n21470) );
no02f01 g17682 ( .a(n21470), .b(n21468), .o(n21471) );
in01f01 g17683 ( .a(n21471), .o(n21472) );
no02f01 g17684 ( .a(n21472), .b(n16155), .o(n21473) );
no02f01 g17685 ( .a(n21473), .b(n21465), .o(n21474) );
in01f01 g17686 ( .a(n21474), .o(n21475) );
no04f01 g17687 ( .a(n21457), .b(n21439), .c(n21417), .d(n21395), .o(n21476) );
na02f01 g17688 ( .a(n21476), .b(n21377), .o(n21477) );
in01f01 g17689 ( .a(n21477), .o(n21478) );
na02f01 g17690 ( .a(n21476), .b(n21382), .o(n21479) );
ao12f01 g17691 ( .a(n16193), .b(n21455), .c(n21437), .o(n21480) );
no02f01 g17692 ( .a(n21480), .b(n21440), .o(n21481) );
na02f01 g17693 ( .a(n21481), .b(n21479), .o(n21482) );
ao12f01 g17694 ( .a(n21482), .b(n21478), .c(n16456), .o(n21483) );
in01f01 g17695 ( .a(n21483), .o(n21484) );
no02f01 g17696 ( .a(n15010), .b(n14553), .o(n21485) );
no02f01 g17697 ( .a(n15009), .b(n14552), .o(n21486) );
no02f01 g17698 ( .a(n21486), .b(n21485), .o(n21487) );
in01f01 g17699 ( .a(n21487), .o(n21488) );
no03f01 g17700 ( .a(n21488), .b(n15000), .c(n14776), .o(n21489) );
no02f01 g17701 ( .a(n15000), .b(n14776), .o(n21490) );
no02f01 g17702 ( .a(n21487), .b(n21490), .o(n21491) );
no02f01 g17703 ( .a(n21491), .b(n21489), .o(n21492) );
in01f01 g17704 ( .a(n21492), .o(n21493) );
no02f01 g17705 ( .a(n21493), .b(n16194), .o(n21494) );
no02f01 g17706 ( .a(n21492), .b(n16193), .o(n21495) );
no02f01 g17707 ( .a(n21495), .b(n21494), .o(n21496) );
in01f01 g17708 ( .a(n21496), .o(n21497) );
no02f01 g17709 ( .a(n21497), .b(n21484), .o(n21498) );
no02f01 g17710 ( .a(n21496), .b(n21483), .o(n21499) );
no02f01 g17711 ( .a(n21499), .b(n21498), .o(n21500) );
in01f01 g17712 ( .a(n21500), .o(n21501) );
no02f01 g17713 ( .a(n21501), .b(n16155), .o(n21502) );
in01f01 g17714 ( .a(n21495), .o(n21503) );
oa12f01 g17715 ( .a(n21503), .b(n21494), .c(n21483), .o(n21504) );
in01f01 g17716 ( .a(n21504), .o(n21505) );
no02f01 g17717 ( .a(n21485), .b(n21490), .o(n21506) );
no02f01 g17718 ( .a(n21506), .b(n21486), .o(n21507) );
no02f01 g17719 ( .a(n15021), .b(n14553), .o(n21508) );
no02f01 g17720 ( .a(n15020), .b(n14552), .o(n21509) );
no02f01 g17721 ( .a(n21509), .b(n21508), .o(n21510) );
no02f01 g17722 ( .a(n21510), .b(n21507), .o(n21511) );
na02f01 g17723 ( .a(n21510), .b(n21507), .o(n21512) );
in01f01 g17724 ( .a(n21512), .o(n21513) );
no02f01 g17725 ( .a(n21513), .b(n21511), .o(n21514) );
in01f01 g17726 ( .a(n21514), .o(n21515) );
no02f01 g17727 ( .a(n21515), .b(n16194), .o(n21516) );
no02f01 g17728 ( .a(n21514), .b(n16193), .o(n21517) );
no02f01 g17729 ( .a(n21517), .b(n21516), .o(n21518) );
no02f01 g17730 ( .a(n21518), .b(n21505), .o(n21519) );
na02f01 g17731 ( .a(n21518), .b(n21505), .o(n21520) );
in01f01 g17732 ( .a(n21520), .o(n21521) );
no02f01 g17733 ( .a(n21521), .b(n21519), .o(n21522) );
in01f01 g17734 ( .a(n21522), .o(n21523) );
no02f01 g17735 ( .a(n21523), .b(n16155), .o(n21524) );
no02f01 g17736 ( .a(n21524), .b(n21502), .o(n21525) );
in01f01 g17737 ( .a(n21525), .o(n21526) );
no02f01 g17738 ( .a(n16194), .b(n15160), .o(n21527) );
no02f01 g17739 ( .a(n16193), .b(n15107), .o(n21528) );
no02f01 g17740 ( .a(n21528), .b(n21527), .o(n21529) );
in01f01 g17741 ( .a(n21529), .o(n21530) );
no02f01 g17742 ( .a(n16194), .b(n15162), .o(n21531) );
in01f01 g17743 ( .a(n21531), .o(n21532) );
in01f01 g17744 ( .a(n21482), .o(n21533) );
no02f01 g17745 ( .a(n21514), .b(n21492), .o(n21534) );
no02f01 g17746 ( .a(n21534), .b(n16194), .o(n21535) );
no02f01 g17747 ( .a(n21535), .b(n21477), .o(n21536) );
na02f01 g17748 ( .a(n21536), .b(n16456), .o(n21537) );
ao12f01 g17749 ( .a(n16193), .b(n21514), .c(n21492), .o(n21538) );
in01f01 g17750 ( .a(n21538), .o(n21539) );
no02f01 g17751 ( .a(n16193), .b(n15114), .o(n21540) );
in01f01 g17752 ( .a(n21540), .o(n21541) );
na04f01 g17753 ( .a(n21541), .b(n21539), .c(n21537), .d(n21533), .o(n21542) );
na03f01 g17754 ( .a(n21542), .b(n21532), .c(n21530), .o(n21543) );
in01f01 g17755 ( .a(n21537), .o(n21544) );
na02f01 g17756 ( .a(n21539), .b(n21533), .o(n21545) );
no03f01 g17757 ( .a(n21540), .b(n21545), .c(n21544), .o(n21546) );
oa12f01 g17758 ( .a(n21529), .b(n21546), .c(n21531), .o(n21547) );
na02f01 g17759 ( .a(n21547), .b(n21543), .o(n21548) );
no02f01 g17760 ( .a(n21548), .b(n16155), .o(n21549) );
no02f01 g17761 ( .a(n21540), .b(n21531), .o(n21550) );
in01f01 g17762 ( .a(n21550), .o(n21551) );
no03f01 g17763 ( .a(n21551), .b(n21545), .c(n21544), .o(n21552) );
no02f01 g17764 ( .a(n21545), .b(n21544), .o(n21553) );
no02f01 g17765 ( .a(n21550), .b(n21553), .o(n21554) );
no02f01 g17766 ( .a(n21554), .b(n21552), .o(n21555) );
in01f01 g17767 ( .a(n21555), .o(n21556) );
no02f01 g17768 ( .a(n21556), .b(n16155), .o(n21557) );
no03f01 g17769 ( .a(n21557), .b(n21549), .c(n21526), .o(n21558) );
in01f01 g17770 ( .a(n21558), .o(n21559) );
no03f01 g17771 ( .a(n21535), .b(n21531), .c(n21527), .o(n21560) );
na03f01 g17772 ( .a(n21560), .b(n21478), .c(n16456), .o(n21561) );
ao12f01 g17773 ( .a(n16193), .b(n15114), .c(n15107), .o(n21562) );
no02f01 g17774 ( .a(n21562), .b(n21538), .o(n21563) );
in01f01 g17775 ( .a(n21563), .o(n21564) );
no02f01 g17776 ( .a(n21564), .b(n21482), .o(n21565) );
na02f01 g17777 ( .a(n21565), .b(n21561), .o(n21566) );
no02f01 g17778 ( .a(n16194), .b(n15123), .o(n21567) );
in01f01 g17779 ( .a(n15123), .o(n21568) );
no02f01 g17780 ( .a(n16193), .b(n21568), .o(n21569) );
no02f01 g17781 ( .a(n21569), .b(n21567), .o(n21570) );
in01f01 g17782 ( .a(n21570), .o(n21571) );
no02f01 g17783 ( .a(n21571), .b(n21566), .o(n21572) );
in01f01 g17784 ( .a(n21572), .o(n21573) );
na02f01 g17785 ( .a(n21571), .b(n21566), .o(n21574) );
na02f01 g17786 ( .a(n21574), .b(n21573), .o(n21575) );
no02f01 g17787 ( .a(n21575), .b(n16155), .o(n21576) );
no04f01 g17788 ( .a(n21576), .b(n21559), .c(n21475), .d(n21428), .o(n21577) );
ao12f01 g17789 ( .a(n16329), .b(n16539), .c(n16510), .o(n21578) );
no02f01 g17790 ( .a(n21578), .b(n16515), .o(n21579) );
in01f01 g17791 ( .a(n21579), .o(n21580) );
ao12f01 g17792 ( .a(n16329), .b(n21424), .c(n21401), .o(n21581) );
no02f01 g17793 ( .a(n21581), .b(n21580), .o(n21582) );
ao12f01 g17794 ( .a(n16329), .b(n21471), .c(n21463), .o(n21583) );
in01f01 g17795 ( .a(n21583), .o(n21584) );
na02f01 g17796 ( .a(n21584), .b(n21582), .o(n21585) );
ao12f01 g17797 ( .a(n16329), .b(n21522), .c(n21500), .o(n21586) );
in01f01 g17798 ( .a(n21543), .o(n21587) );
ao12f01 g17799 ( .a(n21530), .b(n21542), .c(n21532), .o(n21588) );
no02f01 g17800 ( .a(n21588), .b(n21587), .o(n21589) );
ao12f01 g17801 ( .a(n16329), .b(n21555), .c(n21589), .o(n21590) );
no02f01 g17802 ( .a(n21590), .b(n21586), .o(n21591) );
in01f01 g17803 ( .a(n21591), .o(n21592) );
no02f01 g17804 ( .a(n21592), .b(n21585), .o(n21593) );
in01f01 g17805 ( .a(n21574), .o(n21594) );
no02f01 g17806 ( .a(n21594), .b(n21572), .o(n21595) );
no02f01 g17807 ( .a(n21595), .b(n16329), .o(n21596) );
in01f01 g17808 ( .a(n21596), .o(n21597) );
na02f01 g17809 ( .a(n21597), .b(n21593), .o(n21598) );
no02f01 g17810 ( .a(n21569), .b(n21566), .o(n21599) );
no02f01 g17811 ( .a(n16194), .b(n15140), .o(n21600) );
no02f01 g17812 ( .a(n16193), .b(n15136), .o(n21601) );
no02f01 g17813 ( .a(n21601), .b(n21600), .o(n21602) );
oa12f01 g17814 ( .a(n21602), .b(n21599), .c(n21567), .o(n21603) );
in01f01 g17815 ( .a(n21603), .o(n21604) );
no03f01 g17816 ( .a(n21602), .b(n21599), .c(n21567), .o(n21605) );
no02f01 g17817 ( .a(n21605), .b(n21604), .o(n21606) );
in01f01 g17818 ( .a(n21606), .o(n21607) );
no02f01 g17819 ( .a(n21607), .b(n16155), .o(n21608) );
no02f01 g17820 ( .a(n21606), .b(n16329), .o(n21609) );
no02f01 g17821 ( .a(n21609), .b(n21608), .o(n21610) );
in01f01 g17822 ( .a(n21610), .o(n21611) );
oa12f01 g17823 ( .a(n21611), .b(n21598), .c(n21577), .o(n21612) );
in01f01 g17824 ( .a(n21376), .o(n21613) );
in01f01 g17825 ( .a(n21427), .o(n21614) );
no04f01 g17826 ( .a(n21614), .b(n21613), .c(n16488), .d(n16441), .o(n21615) );
in01f01 g17827 ( .a(n21576), .o(n21616) );
na04f01 g17828 ( .a(n21616), .b(n21558), .c(n21474), .d(n21615), .o(n21617) );
in01f01 g17829 ( .a(n21598), .o(n21618) );
na03f01 g17830 ( .a(n21610), .b(n21618), .c(n21617), .o(n21619) );
na03f01 g17831 ( .a(n21619), .b(n21612), .c(delay_sub_ln23_0_unr27_stage10_stallmux_z), .o(n21620) );
in01f01 g17832 ( .a(delay_sub_ln23_0_unr27_stage10_stallmux_z), .o(n21621) );
ao12f01 g17833 ( .a(n21610), .b(n21618), .c(n21617), .o(n21622) );
no03f01 g17834 ( .a(n21611), .b(n21598), .c(n21577), .o(n21623) );
oa12f01 g17835 ( .a(n21621), .b(n21623), .c(n21622), .o(n21624) );
na02f01 g17836 ( .a(n21624), .b(n21620), .o(n283) );
in01f01 g17837 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_28_), .o(n21626) );
no02f01 g17838 ( .a(n21626), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(n21627) );
na02f01 g17839 ( .a(n14281), .b(n14279), .o(n21628) );
no02f01 g17840 ( .a(n11021), .b(delay_xor_ln21_unr3_stage2_stallmux_q_27_), .o(n21629) );
no02f01 g17841 ( .a(n21629), .b(n21628), .o(n21630) );
no02f01 g17842 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_28_), .b(n11021), .o(n21631) );
no02f01 g17843 ( .a(n21631), .b(n21627), .o(n21632) );
in01f01 g17844 ( .a(n21632), .o(n21633) );
no02f01 g17845 ( .a(n21633), .b(n21630), .o(n21634) );
no02f01 g17846 ( .a(n21634), .b(n21627), .o(n21635) );
in01f01 g17847 ( .a(n21635), .o(n21636) );
in01f01 g17848 ( .a(delay_sub_ln21_0_unr2_stage2_stallmux_q_28_), .o(n21637) );
na02f01 g17849 ( .a(n21633), .b(n21630), .o(n21638) );
in01f01 g17850 ( .a(n21638), .o(n21639) );
no03f01 g17851 ( .a(n21639), .b(n21634), .c(n21637), .o(n21640) );
oa12f01 g17852 ( .a(n21635), .b(n21640), .c(delay_sub_ln21_0_unr2_stage2_stallmux_q_29_), .o(n21641) );
na02f01 g17853 ( .a(n11021), .b(delay_xor_ln21_unr3_stage2_stallmux_q_27_), .o(n21642) );
in01f01 g17854 ( .a(n21642), .o(n21643) );
no02f01 g17855 ( .a(n21643), .b(n21629), .o(n21644) );
no02f01 g17856 ( .a(n21644), .b(n21628), .o(n21645) );
na02f01 g17857 ( .a(n21644), .b(n21628), .o(n21646) );
in01f01 g17858 ( .a(n21646), .o(n21647) );
no02f01 g17859 ( .a(n21647), .b(n21645), .o(n21648) );
no02f01 g17860 ( .a(n21648), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_27_), .o(n21649) );
in01f01 g17861 ( .a(n21649), .o(n21650) );
oa12f01 g17862 ( .a(n14289), .b(n14288), .c(n14294), .o(n21651) );
na02f01 g17863 ( .a(n21651), .b(n21650), .o(n21652) );
na02f01 g17864 ( .a(n21648), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_27_), .o(n21653) );
na02f01 g17865 ( .a(n21653), .b(n21652), .o(n21654) );
no02f01 g17866 ( .a(n21635), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_29_), .o(n21655) );
no02f01 g17867 ( .a(n21639), .b(n21634), .o(n21656) );
no02f01 g17868 ( .a(n21656), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_28_), .o(n21657) );
no02f01 g17869 ( .a(n21657), .b(n21655), .o(n21658) );
na02f01 g17870 ( .a(n21658), .b(n21654), .o(n21659) );
na02f01 g17871 ( .a(n21659), .b(n21641), .o(n21660) );
no02f01 g17872 ( .a(n21660), .b(n21636), .o(n21661) );
in01f01 g17873 ( .a(n21661), .o(n21662) );
na02f01 g17874 ( .a(n21660), .b(n21636), .o(n21663) );
in01f01 g17875 ( .a(n21663), .o(n21664) );
no02f01 g17876 ( .a(n21664), .b(n21661), .o(n21665) );
in01f01 g17877 ( .a(n21665), .o(n21666) );
na02f01 g17878 ( .a(n21666), .b(n11158), .o(n21667) );
no02f01 g17879 ( .a(n21654), .b(n21640), .o(n21668) );
in01f01 g17880 ( .a(n21655), .o(n21669) );
na02f01 g17881 ( .a(n21635), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_29_), .o(n21670) );
na02f01 g17882 ( .a(n21670), .b(n21669), .o(n21671) );
in01f01 g17883 ( .a(n21671), .o(n21672) );
no03f01 g17884 ( .a(n21672), .b(n21668), .c(n21657), .o(n21673) );
oa12f01 g17885 ( .a(n21672), .b(n21668), .c(n21657), .o(n21674) );
in01f01 g17886 ( .a(n21674), .o(n21675) );
no02f01 g17887 ( .a(n21675), .b(n21673), .o(n21676) );
no02f01 g17888 ( .a(n21676), .b(n11179), .o(n21677) );
ao12f01 g17889 ( .a(n14288), .b(n14289), .c(n14294), .o(n21678) );
na02f01 g17890 ( .a(n21653), .b(n21650), .o(n21679) );
no02f01 g17891 ( .a(n21679), .b(n21678), .o(n21680) );
na02f01 g17892 ( .a(n21679), .b(n21678), .o(n21681) );
in01f01 g17893 ( .a(n21681), .o(n21682) );
no02f01 g17894 ( .a(n21682), .b(n21680), .o(n21683) );
no02f01 g17895 ( .a(n14296), .b(n11179), .o(n21684) );
ao12f01 g17896 ( .a(n14316), .b(n13571), .c(n11158), .o(n21685) );
in01f01 g17897 ( .a(n21685), .o(n21686) );
no03f01 g17898 ( .a(n21686), .b(n21684), .c(n13833), .o(n21687) );
oa12f01 g17899 ( .a(n21687), .b(n21683), .c(n11179), .o(n21688) );
in01f01 g17900 ( .a(n21688), .o(n21689) );
no02f01 g17901 ( .a(n14296), .b(n11158), .o(n21690) );
ao12f01 g17902 ( .a(n14317), .b(n13571), .c(n11179), .o(n21691) );
in01f01 g17903 ( .a(n21691), .o(n21692) );
no02f01 g17904 ( .a(n21692), .b(n21690), .o(n21693) );
oa12f01 g17905 ( .a(n21693), .b(n21683), .c(n11158), .o(n21694) );
no02f01 g17906 ( .a(n21694), .b(n21689), .o(n21695) );
no02f01 g17907 ( .a(n21657), .b(n21640), .o(n21696) );
in01f01 g17908 ( .a(n21696), .o(n21697) );
no02f01 g17909 ( .a(n21697), .b(n21654), .o(n21698) );
na02f01 g17910 ( .a(n21697), .b(n21654), .o(n21699) );
in01f01 g17911 ( .a(n21699), .o(n21700) );
no02f01 g17912 ( .a(n21700), .b(n21698), .o(n21701) );
in01f01 g17913 ( .a(n21701), .o(n21702) );
ao12f01 g17914 ( .a(n21695), .b(n21702), .c(n11158), .o(n21703) );
in01f01 g17915 ( .a(n21703), .o(n21704) );
no02f01 g17916 ( .a(n21662), .b(n11179), .o(n21705) );
no03f01 g17917 ( .a(n21705), .b(n21704), .c(n21677), .o(n21706) );
no02f01 g17918 ( .a(n21701), .b(n11158), .o(n21707) );
no02f01 g17919 ( .a(n21676), .b(n11158), .o(n21708) );
no02f01 g17920 ( .a(n21708), .b(n21707), .o(n21709) );
oa12f01 g17921 ( .a(n11179), .b(n21664), .c(n21661), .o(n21710) );
na02f01 g17922 ( .a(n21710), .b(n21709), .o(n21711) );
ao12f01 g17923 ( .a(n21711), .b(n21706), .c(n21667), .o(n21712) );
no02f01 g17924 ( .a(n21712), .b(n21662), .o(n21713) );
na02f01 g17925 ( .a(n21712), .b(n21662), .o(n21714) );
in01f01 g17926 ( .a(n21714), .o(n21715) );
no02f01 g17927 ( .a(n21715), .b(n21713), .o(n21716) );
in01f01 g17928 ( .a(delay_add_ln22_unr2_stage2_stallmux_q_31_), .o(n21717) );
no02f01 g17929 ( .a(n13530), .b(n21717), .o(n21718) );
no02f01 g17930 ( .a(n13531), .b(delay_add_ln22_unr2_stage2_stallmux_q_31_), .o(n21719) );
no02f01 g17931 ( .a(n21719), .b(n21718), .o(n21720) );
in01f01 g17932 ( .a(n21720), .o(n21721) );
no03f01 g17933 ( .a(n14265), .b(n14263), .c(n14259), .o(n21722) );
no03f01 g17934 ( .a(n21722), .b(n21721), .c(n14261), .o(n21723) );
oa12f01 g17935 ( .a(n21721), .b(n21722), .c(n14261), .o(n21724) );
in01f01 g17936 ( .a(n21724), .o(n21725) );
no02f01 g17937 ( .a(n21725), .b(n21723), .o(n21726) );
no02f01 g17938 ( .a(n21726), .b(n21716), .o(n21727) );
in01f01 g17939 ( .a(n21716), .o(n21728) );
in01f01 g17940 ( .a(n21723), .o(n21729) );
na02f01 g17941 ( .a(n21724), .b(n21729), .o(n21730) );
no02f01 g17942 ( .a(n21730), .b(n21728), .o(n21731) );
no02f01 g17943 ( .a(n21731), .b(n21727), .o(n21732) );
in01f01 g17944 ( .a(n21732), .o(n21733) );
in01f01 g17945 ( .a(n21709), .o(n21734) );
no02f01 g17946 ( .a(n21704), .b(n21677), .o(n21735) );
no02f01 g17947 ( .a(n21735), .b(n21734), .o(n21736) );
no02f01 g17948 ( .a(n21662), .b(n11158), .o(n21737) );
oa12f01 g17949 ( .a(n21736), .b(n21665), .c(n11158), .o(n21738) );
ao12f01 g17950 ( .a(n21661), .b(n21738), .c(n21667), .o(n21739) );
oa12f01 g17951 ( .a(n13377), .b(n21739), .c(n21737), .o(n21740) );
in01f01 g17952 ( .a(n21740), .o(n21741) );
no02f01 g17953 ( .a(n21736), .b(n21665), .o(n21742) );
na02f01 g17954 ( .a(n21736), .b(n21665), .o(n21743) );
in01f01 g17955 ( .a(n21743), .o(n21744) );
oa12f01 g17956 ( .a(n13298), .b(n21744), .c(n21742), .o(n21745) );
no04f01 g17957 ( .a(n21708), .b(n21707), .c(n21703), .d(n21677), .o(n21746) );
in01f01 g17958 ( .a(n21746), .o(n21747) );
oa22f01 g17959 ( .a(n21708), .b(n21677), .c(n21707), .d(n21703), .o(n21748) );
ao12f01 g17960 ( .a(n13243), .b(n21748), .c(n21747), .o(n21749) );
no02f01 g17961 ( .a(n21701), .b(n21695), .o(n21750) );
in01f01 g17962 ( .a(n21750), .o(n21751) );
na02f01 g17963 ( .a(n21701), .b(n21695), .o(n21752) );
ao12f01 g17964 ( .a(n12419), .b(n21752), .c(n21751), .o(n21753) );
in01f01 g17965 ( .a(n21753), .o(n21754) );
in01f01 g17966 ( .a(n12250), .o(n21755) );
in01f01 g17967 ( .a(n21683), .o(n21756) );
na02f01 g17968 ( .a(n21685), .b(n13831), .o(n21757) );
in01f01 g17969 ( .a(n13832), .o(n21758) );
na02f01 g17970 ( .a(n21691), .b(n21758), .o(n21759) );
no02f01 g17971 ( .a(n21759), .b(n21690), .o(n21760) );
oa12f01 g17972 ( .a(n21760), .b(n21757), .c(n21684), .o(n21761) );
na02f01 g17973 ( .a(n21761), .b(n21756), .o(n21762) );
in01f01 g17974 ( .a(n21762), .o(n21763) );
no02f01 g17975 ( .a(n21761), .b(n21756), .o(n21764) );
no02f01 g17976 ( .a(n21764), .b(n21763), .o(n21765) );
no02f01 g17977 ( .a(n21765), .b(n21755), .o(n21766) );
no02f01 g17978 ( .a(n12247), .b(n12245), .o(n21767) );
ao12f01 g17979 ( .a(n21759), .b(n21685), .c(n13831), .o(n21768) );
no02f01 g17980 ( .a(n21768), .b(n14296), .o(n21769) );
in01f01 g17981 ( .a(n21769), .o(n21770) );
na02f01 g17982 ( .a(n21768), .b(n14296), .o(n21771) );
ao12f01 g17983 ( .a(n21767), .b(n21771), .c(n21770), .o(n21772) );
in01f01 g17984 ( .a(n21772), .o(n21773) );
no02f01 g17985 ( .a(n14326), .b(n13838), .o(n21774) );
no02f01 g17986 ( .a(n21774), .b(n14325), .o(n21775) );
ao12f01 g17987 ( .a(n21775), .b(n14324), .c(n14314), .o(n21776) );
na03f01 g17988 ( .a(n21771), .b(n21770), .c(n21767), .o(n21777) );
in01f01 g17989 ( .a(n21777), .o(n21778) );
oa12f01 g17990 ( .a(n21773), .b(n21778), .c(n21776), .o(n21779) );
na02f01 g17991 ( .a(n21765), .b(n21755), .o(n21780) );
ao12f01 g17992 ( .a(n21766), .b(n21780), .c(n21779), .o(n21781) );
na03f01 g17993 ( .a(n21752), .b(n21751), .c(n12419), .o(n21782) );
in01f01 g17994 ( .a(n21782), .o(n21783) );
oa12f01 g17995 ( .a(n21754), .b(n21783), .c(n21781), .o(n21784) );
na03f01 g17996 ( .a(n21748), .b(n21747), .c(n13243), .o(n21785) );
ao12f01 g17997 ( .a(n21749), .b(n21785), .c(n21784), .o(n21786) );
no03f01 g17998 ( .a(n21744), .b(n21742), .c(n13298), .o(n21787) );
oa12f01 g17999 ( .a(n21745), .b(n21787), .c(n21786), .o(n21788) );
no03f01 g18000 ( .a(n21739), .b(n21737), .c(n13377), .o(n21789) );
in01f01 g18001 ( .a(n21789), .o(n21790) );
ao12f01 g18002 ( .a(n21741), .b(n21790), .c(n21788), .o(n21791) );
no02f01 g18003 ( .a(n21728), .b(n13539), .o(n21792) );
no02f01 g18004 ( .a(n21728), .b(n13461), .o(n21793) );
no02f01 g18005 ( .a(n21793), .b(n21792), .o(n21794) );
in01f01 g18006 ( .a(n21794), .o(n21795) );
no03f01 g18007 ( .a(n21795), .b(n21791), .c(n14269), .o(n21796) );
in01f01 g18008 ( .a(n21742), .o(n21797) );
ao12f01 g18009 ( .a(n13307), .b(n21743), .c(n21797), .o(n21798) );
in01f01 g18010 ( .a(n21749), .o(n21799) );
in01f01 g18011 ( .a(n21766), .o(n21800) );
oa12f01 g18012 ( .a(n13839), .b(n13828), .c(n13648), .o(n21801) );
ao12f01 g18013 ( .a(n14325), .b(n21774), .c(n21801), .o(n21802) );
ao12f01 g18014 ( .a(n21772), .b(n21777), .c(n21802), .o(n21803) );
in01f01 g18015 ( .a(n21780), .o(n21804) );
oa12f01 g18016 ( .a(n21800), .b(n21804), .c(n21803), .o(n21805) );
ao12f01 g18017 ( .a(n21753), .b(n21782), .c(n21805), .o(n21806) );
in01f01 g18018 ( .a(n21785), .o(n21807) );
oa12f01 g18019 ( .a(n21799), .b(n21807), .c(n21806), .o(n21808) );
na03f01 g18020 ( .a(n21743), .b(n21797), .c(n13307), .o(n21809) );
ao12f01 g18021 ( .a(n21798), .b(n21809), .c(n21808), .o(n21810) );
oa12f01 g18022 ( .a(n21740), .b(n21789), .c(n21810), .o(n21811) );
in01f01 g18023 ( .a(n13461), .o(n21812) );
ao12f01 g18024 ( .a(n21716), .b(n13546), .c(n21812), .o(n21813) );
ao12f01 g18025 ( .a(n21813), .b(n21794), .c(n21811), .o(n21814) );
ao12f01 g18026 ( .a(n21716), .b(n21814), .c(n14269), .o(n21815) );
no03f01 g18027 ( .a(n21815), .b(n21796), .c(n21733), .o(n21816) );
in01f01 g18028 ( .a(n21796), .o(n21817) );
in01f01 g18029 ( .a(n14268), .o(n21818) );
na02f01 g18030 ( .a(n21818), .b(n14266), .o(n21819) );
in01f01 g18031 ( .a(n21813), .o(n21820) );
oa12f01 g18032 ( .a(n21820), .b(n21795), .c(n21791), .o(n21821) );
oa12f01 g18033 ( .a(n21728), .b(n21821), .c(n21819), .o(n21822) );
ao12f01 g18034 ( .a(n21732), .b(n21822), .c(n21817), .o(n21823) );
oa12f01 g18035 ( .a(n11514), .b(n21823), .c(n21816), .o(n21824) );
in01f01 g18036 ( .a(n21793), .o(n21825) );
no02f01 g18037 ( .a(n21716), .b(n21812), .o(n21826) );
in01f01 g18038 ( .a(n21826), .o(n21827) );
na02f01 g18039 ( .a(n21827), .b(n21791), .o(n21828) );
no02f01 g18040 ( .a(n21716), .b(n13546), .o(n21829) );
no02f01 g18041 ( .a(n21829), .b(n21792), .o(n21830) );
in01f01 g18042 ( .a(n21830), .o(n21831) );
ao12f01 g18043 ( .a(n21831), .b(n21828), .c(n21825), .o(n21832) );
no02f01 g18044 ( .a(n21826), .b(n21811), .o(n21833) );
no03f01 g18045 ( .a(n21830), .b(n21833), .c(n21793), .o(n21834) );
no02f01 g18046 ( .a(n21834), .b(n21832), .o(n21835) );
no02f01 g18047 ( .a(n21835), .b(n11515), .o(n21836) );
no02f01 g18048 ( .a(n21826), .b(n21793), .o(n21837) );
na02f01 g18049 ( .a(n21837), .b(n21791), .o(n21838) );
in01f01 g18050 ( .a(n21837), .o(n21839) );
na02f01 g18051 ( .a(n21839), .b(n21811), .o(n21840) );
na02f01 g18052 ( .a(n21840), .b(n21838), .o(n21841) );
no02f01 g18053 ( .a(n21783), .b(n21753), .o(n21842) );
in01f01 g18054 ( .a(n21842), .o(n21843) );
no02f01 g18055 ( .a(n21843), .b(n21805), .o(n21844) );
no02f01 g18056 ( .a(n21842), .b(n21781), .o(n21845) );
no02f01 g18057 ( .a(n21845), .b(n21844), .o(n21846) );
no02f01 g18058 ( .a(n21846), .b(n11515), .o(n21847) );
in01f01 g18059 ( .a(n21847), .o(n21848) );
oa12f01 g18060 ( .a(n11514), .b(n14173), .c(n14087), .o(n21849) );
na02f01 g18061 ( .a(n14188), .b(n11514), .o(n21850) );
na02f01 g18062 ( .a(n21850), .b(n21849), .o(n21851) );
no02f01 g18063 ( .a(n14070), .b(n11515), .o(n21852) );
no02f01 g18064 ( .a(n14070), .b(n11514), .o(n21853) );
no02f01 g18065 ( .a(n14187), .b(n11514), .o(n21854) );
no02f01 g18066 ( .a(n21854), .b(n21853), .o(n21855) );
oa12f01 g18067 ( .a(n21855), .b(n21852), .c(n21851), .o(n21856) );
no02f01 g18068 ( .a(n14058), .b(n11515), .o(n21857) );
in01f01 g18069 ( .a(n21857), .o(n21858) );
no02f01 g18070 ( .a(n14047), .b(n11515), .o(n21859) );
in01f01 g18071 ( .a(n21859), .o(n21860) );
no02f01 g18072 ( .a(n14033), .b(n11515), .o(n21861) );
in01f01 g18073 ( .a(n21861), .o(n21862) );
na04f01 g18074 ( .a(n21862), .b(n21860), .c(n21858), .d(n21856), .o(n21863) );
no02f01 g18075 ( .a(n14019), .b(n11515), .o(n21864) );
no02f01 g18076 ( .a(n14033), .b(n11514), .o(n21865) );
no02f01 g18077 ( .a(n14047), .b(n11514), .o(n21866) );
no02f01 g18078 ( .a(n14058), .b(n11514), .o(n21867) );
no02f01 g18079 ( .a(n21867), .b(n21866), .o(n21868) );
in01f01 g18080 ( .a(n21868), .o(n21869) );
no02f01 g18081 ( .a(n21869), .b(n21865), .o(n21870) );
in01f01 g18082 ( .a(n21870), .o(n21871) );
no02f01 g18083 ( .a(n14019), .b(n11514), .o(n21872) );
no02f01 g18084 ( .a(n21872), .b(n21871), .o(n21873) );
oa12f01 g18085 ( .a(n21873), .b(n21864), .c(n21863), .o(n21874) );
no02f01 g18086 ( .a(n14004), .b(n11515), .o(n21875) );
in01f01 g18087 ( .a(n21875), .o(n21876) );
no02f01 g18088 ( .a(n14224), .b(n11515), .o(n21877) );
in01f01 g18089 ( .a(n21877), .o(n21878) );
no02f01 g18090 ( .a(n13984), .b(n11515), .o(n21879) );
in01f01 g18091 ( .a(n21879), .o(n21880) );
na04f01 g18092 ( .a(n21880), .b(n21878), .c(n21876), .d(n21874), .o(n21881) );
no02f01 g18093 ( .a(n13959), .b(n11515), .o(n21882) );
no02f01 g18094 ( .a(n13984), .b(n11514), .o(n21883) );
no02f01 g18095 ( .a(n14224), .b(n11514), .o(n21884) );
no02f01 g18096 ( .a(n14004), .b(n11514), .o(n21885) );
no02f01 g18097 ( .a(n21885), .b(n21884), .o(n21886) );
in01f01 g18098 ( .a(n21886), .o(n21887) );
no02f01 g18099 ( .a(n21887), .b(n21883), .o(n21888) );
in01f01 g18100 ( .a(n21888), .o(n21889) );
no02f01 g18101 ( .a(n13959), .b(n11514), .o(n21890) );
no02f01 g18102 ( .a(n21890), .b(n21889), .o(n21891) );
oa12f01 g18103 ( .a(n21891), .b(n21882), .c(n21881), .o(n21892) );
no02f01 g18104 ( .a(n13941), .b(n11515), .o(n21893) );
in01f01 g18105 ( .a(n21893), .o(n21894) );
no02f01 g18106 ( .a(n13925), .b(n11515), .o(n21895) );
in01f01 g18107 ( .a(n21895), .o(n21896) );
na03f01 g18108 ( .a(n21896), .b(n21894), .c(n21892), .o(n21897) );
no02f01 g18109 ( .a(n14246), .b(n11515), .o(n21898) );
no02f01 g18110 ( .a(n13906), .b(n11515), .o(n21899) );
no03f01 g18111 ( .a(n21899), .b(n21898), .c(n21897), .o(n21900) );
na02f01 g18112 ( .a(n13889), .b(n11515), .o(n21901) );
no02f01 g18113 ( .a(n13906), .b(n11514), .o(n21902) );
in01f01 g18114 ( .a(n21902), .o(n21903) );
no02f01 g18115 ( .a(n13925), .b(n11514), .o(n21904) );
no02f01 g18116 ( .a(n13941), .b(n11514), .o(n21905) );
no02f01 g18117 ( .a(n21905), .b(n21904), .o(n21906) );
na03f01 g18118 ( .a(n21906), .b(n21903), .c(n21901), .o(n21907) );
no02f01 g18119 ( .a(n21907), .b(n21900), .o(n21908) );
no02f01 g18120 ( .a(n14331), .b(n11515), .o(n21909) );
no02f01 g18121 ( .a(n21778), .b(n21772), .o(n21910) );
in01f01 g18122 ( .a(n21910), .o(n21911) );
no02f01 g18123 ( .a(n21911), .b(n21802), .o(n21912) );
no02f01 g18124 ( .a(n21910), .b(n21776), .o(n21913) );
no02f01 g18125 ( .a(n21913), .b(n21912), .o(n21914) );
no02f01 g18126 ( .a(n21914), .b(n11515), .o(n21915) );
no03f01 g18127 ( .a(n21915), .b(n21909), .c(n21908), .o(n21916) );
oa12f01 g18128 ( .a(n21777), .b(n21802), .c(n21772), .o(n21917) );
no02f01 g18129 ( .a(n21804), .b(n21766), .o(n21918) );
no02f01 g18130 ( .a(n21918), .b(n21917), .o(n21919) );
na02f01 g18131 ( .a(n21918), .b(n21917), .o(n21920) );
in01f01 g18132 ( .a(n21920), .o(n21921) );
no02f01 g18133 ( .a(n21921), .b(n21919), .o(n21922) );
oa12f01 g18134 ( .a(n21916), .b(n21922), .c(n11515), .o(n21923) );
no02f01 g18135 ( .a(n21922), .b(n11514), .o(n21924) );
no02f01 g18136 ( .a(n21914), .b(n11514), .o(n21925) );
no02f01 g18137 ( .a(n14331), .b(n11514), .o(n21926) );
no02f01 g18138 ( .a(n21926), .b(n21925), .o(n21927) );
in01f01 g18139 ( .a(n21927), .o(n21928) );
no02f01 g18140 ( .a(n21928), .b(n21924), .o(n21929) );
na02f01 g18141 ( .a(n21842), .b(n21781), .o(n21930) );
na02f01 g18142 ( .a(n21843), .b(n21805), .o(n21931) );
na02f01 g18143 ( .a(n21931), .b(n21930), .o(n21932) );
na02f01 g18144 ( .a(n21932), .b(n11515), .o(n21933) );
na03f01 g18145 ( .a(n21933), .b(n21929), .c(n21923), .o(n21934) );
no02f01 g18146 ( .a(n21807), .b(n21749), .o(n21935) );
na02f01 g18147 ( .a(n21935), .b(n21806), .o(n21936) );
na02f01 g18148 ( .a(n21785), .b(n21799), .o(n21937) );
na02f01 g18149 ( .a(n21937), .b(n21784), .o(n21938) );
na02f01 g18150 ( .a(n21938), .b(n21936), .o(n21939) );
na02f01 g18151 ( .a(n21939), .b(n11514), .o(n21940) );
na03f01 g18152 ( .a(n21940), .b(n21934), .c(n21848), .o(n21941) );
no02f01 g18153 ( .a(n21787), .b(n21798), .o(n21942) );
na02f01 g18154 ( .a(n21942), .b(n21786), .o(n21943) );
na02f01 g18155 ( .a(n21809), .b(n21745), .o(n21944) );
na02f01 g18156 ( .a(n21944), .b(n21808), .o(n21945) );
ao12f01 g18157 ( .a(n11515), .b(n21945), .c(n21943), .o(n21946) );
no02f01 g18158 ( .a(n21946), .b(n21941), .o(n21947) );
na02f01 g18159 ( .a(n21786), .b(n21745), .o(n21948) );
na02f01 g18160 ( .a(n21790), .b(n21740), .o(n21949) );
ao12f01 g18161 ( .a(n21949), .b(n21948), .c(n21809), .o(n21950) );
no02f01 g18162 ( .a(n21808), .b(n21798), .o(n21951) );
no02f01 g18163 ( .a(n21789), .b(n21741), .o(n21952) );
no03f01 g18164 ( .a(n21952), .b(n21951), .c(n21787), .o(n21953) );
no02f01 g18165 ( .a(n21953), .b(n21950), .o(n21954) );
oa12f01 g18166 ( .a(n21947), .b(n21954), .c(n11515), .o(n21955) );
ao12f01 g18167 ( .a(n21955), .b(n21841), .c(n11514), .o(n21956) );
no02f01 g18168 ( .a(n21839), .b(n21811), .o(n21957) );
no02f01 g18169 ( .a(n21837), .b(n21791), .o(n21958) );
no02f01 g18170 ( .a(n21958), .b(n21957), .o(n21959) );
oa12f01 g18171 ( .a(n21952), .b(n21951), .c(n21787), .o(n21960) );
na03f01 g18172 ( .a(n21949), .b(n21948), .c(n21809), .o(n21961) );
na02f01 g18173 ( .a(n21961), .b(n21960), .o(n21962) );
no02f01 g18174 ( .a(n21944), .b(n21808), .o(n21963) );
in01f01 g18175 ( .a(n21945), .o(n21964) );
no02f01 g18176 ( .a(n21964), .b(n21963), .o(n21965) );
no02f01 g18177 ( .a(n21937), .b(n21784), .o(n21966) );
no02f01 g18178 ( .a(n21935), .b(n21806), .o(n21967) );
no02f01 g18179 ( .a(n21967), .b(n21966), .o(n21968) );
no02f01 g18180 ( .a(n21968), .b(n11514), .o(n21969) );
in01f01 g18181 ( .a(n21969), .o(n21970) );
oa12f01 g18182 ( .a(n21970), .b(n21965), .c(n11514), .o(n21971) );
ao12f01 g18183 ( .a(n21971), .b(n21962), .c(n11515), .o(n21972) );
oa12f01 g18184 ( .a(n21972), .b(n21959), .c(n11514), .o(n21973) );
no02f01 g18185 ( .a(n21973), .b(n21956), .o(n21974) );
no02f01 g18186 ( .a(n21728), .b(n21819), .o(n21975) );
no02f01 g18187 ( .a(n21716), .b(n14269), .o(n21976) );
no02f01 g18188 ( .a(n21976), .b(n21975), .o(n21977) );
in01f01 g18189 ( .a(n21977), .o(n21978) );
na02f01 g18190 ( .a(n21978), .b(n21821), .o(n21979) );
na02f01 g18191 ( .a(n21977), .b(n21814), .o(n21980) );
ao12f01 g18192 ( .a(n11515), .b(n21980), .c(n21979), .o(n21981) );
no03f01 g18193 ( .a(n21981), .b(n21974), .c(n21836), .o(n21982) );
ao12f01 g18194 ( .a(n11514), .b(n21980), .c(n21979), .o(n21983) );
oa12f01 g18195 ( .a(n21830), .b(n21833), .c(n21793), .o(n21984) );
na03f01 g18196 ( .a(n21831), .b(n21828), .c(n21825), .o(n21985) );
ao12f01 g18197 ( .a(n11514), .b(n21985), .c(n21984), .o(n21986) );
no02f01 g18198 ( .a(n21986), .b(n21983), .o(n21987) );
in01f01 g18199 ( .a(n21987), .o(n21988) );
no02f01 g18200 ( .a(n21988), .b(n21982), .o(n21989) );
na03f01 g18201 ( .a(n21822), .b(n21817), .c(n21732), .o(n21990) );
oa12f01 g18202 ( .a(n21733), .b(n21815), .c(n21796), .o(n21991) );
ao12f01 g18203 ( .a(n11514), .b(n21991), .c(n21990), .o(n21992) );
oa12f01 g18204 ( .a(n21824), .b(n21992), .c(n21989), .o(n21993) );
in01f01 g18205 ( .a(n14270), .o(n21994) );
na02f01 g18206 ( .a(n21730), .b(n11179), .o(n21995) );
oa12f01 g18207 ( .a(n11158), .b(n21725), .c(n21723), .o(n21996) );
na02f01 g18208 ( .a(n21996), .b(n21995), .o(n21997) );
no03f01 g18209 ( .a(n14271), .b(n13547), .c(n13463), .o(n21998) );
oa12f01 g18210 ( .a(n21998), .b(n14275), .c(n13471), .o(n21999) );
ao12f01 g18211 ( .a(n21997), .b(n21999), .c(n21994), .o(n22000) );
no02f01 g18212 ( .a(n21726), .b(n11158), .o(n22001) );
ao12f01 g18213 ( .a(n11179), .b(n21724), .c(n21729), .o(n22002) );
no02f01 g18214 ( .a(n22002), .b(n22001), .o(n22003) );
na02f01 g18215 ( .a(n21819), .b(n11179), .o(n22004) );
na03f01 g18216 ( .a(n22004), .b(n13540), .c(n13462), .o(n22005) );
ao12f01 g18217 ( .a(n22005), .b(n14257), .c(n13439), .o(n22006) );
no03f01 g18218 ( .a(n22006), .b(n22003), .c(n14270), .o(n22007) );
oa12f01 g18219 ( .a(n21683), .b(n22007), .c(n22000), .o(n22008) );
ao12f01 g18220 ( .a(n14305), .b(n14255), .c(n13572), .o(n22009) );
oa12f01 g18221 ( .a(n22003), .b(n22006), .c(n14270), .o(n22010) );
na03f01 g18222 ( .a(n21999), .b(n21997), .c(n21994), .o(n22011) );
na03f01 g18223 ( .a(n22011), .b(n22010), .c(n21756), .o(n22012) );
na02f01 g18224 ( .a(n22012), .b(n14298), .o(n22013) );
oa12f01 g18225 ( .a(n22008), .b(n22013), .c(n22009), .o(n22014) );
in01f01 g18226 ( .a(n21676), .o(n22015) );
no02f01 g18227 ( .a(n13469), .b(n13468), .o(n22016) );
in01f01 g18228 ( .a(n22016), .o(n22017) );
na04f01 g18229 ( .a(n21996), .b(n21994), .c(n14257), .d(n22017), .o(n22018) );
no02f01 g18230 ( .a(n22005), .b(n22001), .o(n22019) );
ao12f01 g18231 ( .a(n22002), .b(n22019), .c(n22018), .o(n22020) );
no04f01 g18232 ( .a(n22002), .b(n14270), .c(n14275), .d(n13438), .o(n22021) );
no03f01 g18233 ( .a(n22021), .b(n22020), .c(n21997), .o(n22022) );
no04f01 g18234 ( .a(n22002), .b(n14270), .c(n14275), .d(n22016), .o(n22023) );
na02f01 g18235 ( .a(n21998), .b(n21995), .o(n22024) );
oa12f01 g18236 ( .a(n21996), .b(n22024), .c(n22023), .o(n22025) );
in01f01 g18237 ( .a(n22021), .o(n22026) );
ao12f01 g18238 ( .a(n22003), .b(n22026), .c(n22025), .o(n22027) );
no02f01 g18239 ( .a(n22027), .b(n22022), .o(n22028) );
ao12f01 g18240 ( .a(n22028), .b(n21702), .c(n22015), .o(n22029) );
oa12f01 g18241 ( .a(n22028), .b(n21702), .c(n22015), .o(n22030) );
oa12f01 g18242 ( .a(n22030), .b(n22029), .c(n22014), .o(n22031) );
na03f01 g18243 ( .a(n22026), .b(n22025), .c(n22003), .o(n22032) );
oa12f01 g18244 ( .a(n21997), .b(n22021), .c(n22020), .o(n22033) );
na02f01 g18245 ( .a(n22033), .b(n22032), .o(n22034) );
no02f01 g18246 ( .a(n22034), .b(n21665), .o(n22035) );
no02f01 g18247 ( .a(n22028), .b(n21666), .o(n22036) );
no02f01 g18248 ( .a(n22036), .b(n22035), .o(n22037) );
in01f01 g18249 ( .a(n22037), .o(n22038) );
na02f01 g18250 ( .a(n22038), .b(n22031), .o(n22039) );
ao12f01 g18251 ( .a(n13581), .b(n13577), .c(n13506), .o(n22040) );
no02f01 g18252 ( .a(n22040), .b(n13580), .o(n22041) );
no03f01 g18253 ( .a(n22007), .b(n22000), .c(n21683), .o(n22042) );
no02f01 g18254 ( .a(n22042), .b(n14304), .o(n22043) );
oa12f01 g18255 ( .a(n22043), .b(n14305), .c(n22041), .o(n22044) );
oa12f01 g18256 ( .a(n22034), .b(n21701), .c(n21676), .o(n22045) );
na03f01 g18257 ( .a(n22045), .b(n22044), .c(n22008), .o(n22046) );
na03f01 g18258 ( .a(n22037), .b(n22030), .c(n22046), .o(n22047) );
na02f01 g18259 ( .a(n22047), .b(n22039), .o(n22048) );
no02f01 g18260 ( .a(n22048), .b(n21993), .o(n22049) );
in01f01 g18261 ( .a(n21993), .o(n22050) );
ao12f01 g18262 ( .a(n22037), .b(n22030), .c(n22046), .o(n22051) );
no02f01 g18263 ( .a(n22038), .b(n22031), .o(n22052) );
no02f01 g18264 ( .a(n22052), .b(n22051), .o(n22053) );
no02f01 g18265 ( .a(n22053), .b(n22050), .o(n22054) );
no02f01 g18266 ( .a(n22054), .b(n22049), .o(n22055) );
in01f01 g18267 ( .a(n22055), .o(n22056) );
na02f01 g18268 ( .a(n21841), .b(n11514), .o(n22057) );
na02f01 g18269 ( .a(n21841), .b(n11515), .o(n22058) );
na02f01 g18270 ( .a(n22058), .b(n22057), .o(n22059) );
na02f01 g18271 ( .a(n21962), .b(n11514), .o(n22060) );
in01f01 g18272 ( .a(n22060), .o(n22061) );
na02f01 g18273 ( .a(n21962), .b(n11515), .o(n22062) );
no02f01 g18274 ( .a(n21971), .b(n21947), .o(n22063) );
ao12f01 g18275 ( .a(n22061), .b(n22063), .c(n22062), .o(n22064) );
no02f01 g18276 ( .a(n22064), .b(n22059), .o(n22065) );
in01f01 g18277 ( .a(n22064), .o(n22066) );
ao12f01 g18278 ( .a(n22066), .b(n22058), .c(n22057), .o(n22067) );
no02f01 g18279 ( .a(n22067), .b(n22065), .o(n22068) );
no02f01 g18280 ( .a(n22068), .b(n13517), .o(n22069) );
na02f01 g18281 ( .a(n22068), .b(n13517), .o(n22070) );
in01f01 g18282 ( .a(n22063), .o(n22071) );
na02f01 g18283 ( .a(n22062), .b(n22060), .o(n22072) );
na02f01 g18284 ( .a(n22072), .b(n22071), .o(n22073) );
in01f01 g18285 ( .a(n22072), .o(n22074) );
na02f01 g18286 ( .a(n22074), .b(n22063), .o(n22075) );
na02f01 g18287 ( .a(n22075), .b(n22073), .o(n22076) );
no02f01 g18288 ( .a(n22076), .b(n13354), .o(n22077) );
na02f01 g18289 ( .a(n13889), .b(n11514), .o(n22078) );
in01f01 g18290 ( .a(n21899), .o(n22079) );
na02f01 g18291 ( .a(n22079), .b(n22078), .o(n22080) );
no02f01 g18292 ( .a(n14246), .b(n11514), .o(n22081) );
in01f01 g18293 ( .a(n21906), .o(n22082) );
no03f01 g18294 ( .a(n22082), .b(n21902), .c(n22081), .o(n22083) );
oa12f01 g18295 ( .a(n22083), .b(n22080), .c(n21897), .o(n22084) );
na02f01 g18296 ( .a(n14335), .b(n11514), .o(n22085) );
in01f01 g18297 ( .a(n21915), .o(n22086) );
na03f01 g18298 ( .a(n22086), .b(n22085), .c(n22084), .o(n22087) );
no02f01 g18299 ( .a(n21922), .b(n11515), .o(n22088) );
no02f01 g18300 ( .a(n22088), .b(n22087), .o(n22089) );
oa12f01 g18301 ( .a(n21927), .b(n21922), .c(n11514), .o(n22090) );
no02f01 g18302 ( .a(n21846), .b(n11514), .o(n22091) );
no03f01 g18303 ( .a(n22091), .b(n22090), .c(n22089), .o(n22092) );
no02f01 g18304 ( .a(n21968), .b(n11515), .o(n22093) );
no03f01 g18305 ( .a(n22093), .b(n22092), .c(n21847), .o(n22094) );
no02f01 g18306 ( .a(n21969), .b(n22094), .o(n22095) );
in01f01 g18307 ( .a(n22095), .o(n22096) );
in01f01 g18308 ( .a(n21946), .o(n22097) );
na02f01 g18309 ( .a(n21945), .b(n21943), .o(n22098) );
na02f01 g18310 ( .a(n22098), .b(n11515), .o(n22099) );
na02f01 g18311 ( .a(n22099), .b(n22097), .o(n22100) );
no02f01 g18312 ( .a(n22100), .b(n22096), .o(n22101) );
ao12f01 g18313 ( .a(n22095), .b(n22099), .c(n22097), .o(n22102) );
no02f01 g18314 ( .a(n22102), .b(n22101), .o(n22103) );
na02f01 g18315 ( .a(n22103), .b(n13523), .o(n22104) );
na02f01 g18316 ( .a(n13037), .b(n13022), .o(n22105) );
na02f01 g18317 ( .a(n13018), .b(n12726), .o(n22106) );
na02f01 g18318 ( .a(n22106), .b(n22105), .o(n22107) );
no02f01 g18319 ( .a(n22092), .b(n21847), .o(n22108) );
no02f01 g18320 ( .a(n21969), .b(n22093), .o(n22109) );
in01f01 g18321 ( .a(n22109), .o(n22110) );
no02f01 g18322 ( .a(n22110), .b(n22108), .o(n22111) );
na02f01 g18323 ( .a(n22110), .b(n22108), .o(n22112) );
in01f01 g18324 ( .a(n22112), .o(n22113) );
no02f01 g18325 ( .a(n22113), .b(n22111), .o(n22114) );
na02f01 g18326 ( .a(n22114), .b(n22107), .o(n22115) );
no02f01 g18327 ( .a(n22103), .b(n13523), .o(n22116) );
ao12f01 g18328 ( .a(n22116), .b(n22115), .c(n22104), .o(n22117) );
na02f01 g18329 ( .a(n22076), .b(n13354), .o(n22118) );
ao12f01 g18330 ( .a(n22077), .b(n22118), .c(n22117), .o(n22119) );
ao12f01 g18331 ( .a(n22069), .b(n22119), .c(n22070), .o(n22120) );
na03f01 g18332 ( .a(n22095), .b(n22099), .c(n22097), .o(n22121) );
in01f01 g18333 ( .a(n22102), .o(n22122) );
na02f01 g18334 ( .a(n22122), .b(n22121), .o(n22123) );
na02f01 g18335 ( .a(n22123), .b(n13276), .o(n22124) );
in01f01 g18336 ( .a(n13105), .o(n22125) );
in01f01 g18337 ( .a(n21881), .o(n22126) );
no02f01 g18338 ( .a(n21889), .b(n22126), .o(n22127) );
no02f01 g18339 ( .a(n21890), .b(n21882), .o(n22128) );
no02f01 g18340 ( .a(n22128), .b(n22127), .o(n22129) );
na02f01 g18341 ( .a(n22128), .b(n22127), .o(n22130) );
in01f01 g18342 ( .a(n22130), .o(n22131) );
no02f01 g18343 ( .a(n22131), .b(n22129), .o(n22132) );
no02f01 g18344 ( .a(n22132), .b(n22125), .o(n22133) );
na02f01 g18345 ( .a(n21876), .b(n21874), .o(n22134) );
in01f01 g18346 ( .a(n22134), .o(n22135) );
ao12f01 g18347 ( .a(n21887), .b(n21878), .c(n22135), .o(n22136) );
in01f01 g18348 ( .a(n22136), .o(n22137) );
no02f01 g18349 ( .a(n21883), .b(n21879), .o(n22138) );
in01f01 g18350 ( .a(n22138), .o(n22139) );
no02f01 g18351 ( .a(n22139), .b(n22137), .o(n22140) );
no02f01 g18352 ( .a(n22138), .b(n22136), .o(n22141) );
no03f01 g18353 ( .a(n22141), .b(n22140), .c(n13092), .o(n22142) );
in01f01 g18354 ( .a(n21874), .o(n22143) );
no02f01 g18355 ( .a(n21885), .b(n21875), .o(n22144) );
no02f01 g18356 ( .a(n22144), .b(n22143), .o(n22145) );
na02f01 g18357 ( .a(n22144), .b(n22143), .o(n22146) );
in01f01 g18358 ( .a(n22146), .o(n22147) );
no03f01 g18359 ( .a(n22147), .b(n22145), .c(n13073), .o(n22148) );
no02f01 g18360 ( .a(n21872), .b(n21864), .o(n22149) );
ao12f01 g18361 ( .a(n22149), .b(n21870), .c(n21863), .o(n22150) );
in01f01 g18362 ( .a(n21863), .o(n22151) );
in01f01 g18363 ( .a(n22149), .o(n22152) );
no03f01 g18364 ( .a(n22152), .b(n21871), .c(n22151), .o(n22153) );
no02f01 g18365 ( .a(n22153), .b(n22150), .o(n22154) );
no02f01 g18366 ( .a(n22154), .b(n13065), .o(n22155) );
in01f01 g18367 ( .a(n21856), .o(n22156) );
no02f01 g18368 ( .a(n21857), .b(n22156), .o(n22157) );
no02f01 g18369 ( .a(n21867), .b(n22157), .o(n22158) );
no02f01 g18370 ( .a(n21866), .b(n21859), .o(n22159) );
no02f01 g18371 ( .a(n22159), .b(n22158), .o(n22160) );
na02f01 g18372 ( .a(n22159), .b(n22158), .o(n22161) );
in01f01 g18373 ( .a(n22161), .o(n22162) );
no02f01 g18374 ( .a(n22162), .b(n22160), .o(n22163) );
no02f01 g18375 ( .a(n22163), .b(n13047), .o(n22164) );
no02f01 g18376 ( .a(n21867), .b(n21857), .o(n22165) );
in01f01 g18377 ( .a(n22165), .o(n22166) );
no02f01 g18378 ( .a(n22166), .b(n21856), .o(n22167) );
na02f01 g18379 ( .a(n22166), .b(n21856), .o(n22168) );
in01f01 g18380 ( .a(n22168), .o(n22169) );
no02f01 g18381 ( .a(n22169), .b(n22167), .o(n22170) );
in01f01 g18382 ( .a(n22170), .o(n22171) );
no02f01 g18383 ( .a(n12928), .b(n12878), .o(n22172) );
no02f01 g18384 ( .a(n22172), .b(n12925), .o(n22173) );
na02f01 g18385 ( .a(n22172), .b(n12925), .o(n22174) );
in01f01 g18386 ( .a(n22174), .o(n22175) );
no02f01 g18387 ( .a(n22175), .b(n22173), .o(n22176) );
no02f01 g18388 ( .a(n22176), .b(n22171), .o(n22177) );
na02f01 g18389 ( .a(n22176), .b(n22171), .o(n22178) );
in01f01 g18390 ( .a(n21854), .o(n22179) );
na02f01 g18391 ( .a(n22179), .b(n21851), .o(n22180) );
in01f01 g18392 ( .a(n22180), .o(n22181) );
no02f01 g18393 ( .a(n21853), .b(n21852), .o(n22182) );
no02f01 g18394 ( .a(n22182), .b(n22181), .o(n22183) );
na02f01 g18395 ( .a(n22182), .b(n22181), .o(n22184) );
in01f01 g18396 ( .a(n22184), .o(n22185) );
no02f01 g18397 ( .a(n22185), .b(n22183), .o(n22186) );
in01f01 g18398 ( .a(n12924), .o(n22187) );
in01f01 g18399 ( .a(n12891), .o(n22188) );
no02f01 g18400 ( .a(n22188), .b(n12890), .o(n22189) );
no02f01 g18401 ( .a(n22189), .b(n22187), .o(n22190) );
na02f01 g18402 ( .a(n22189), .b(n22187), .o(n22191) );
in01f01 g18403 ( .a(n22191), .o(n22192) );
no02f01 g18404 ( .a(n22192), .b(n22190), .o(n22193) );
in01f01 g18405 ( .a(n22193), .o(n22194) );
no02f01 g18406 ( .a(n22194), .b(n22186), .o(n22195) );
na02f01 g18407 ( .a(n22179), .b(n21850), .o(n22196) );
na02f01 g18408 ( .a(n22196), .b(n21849), .o(n22197) );
in01f01 g18409 ( .a(n21849), .o(n22198) );
na03f01 g18410 ( .a(n22179), .b(n21850), .c(n22198), .o(n22199) );
na02f01 g18411 ( .a(n22199), .b(n22197), .o(n22200) );
no02f01 g18412 ( .a(n12908), .b(n12907), .o(n22201) );
no02f01 g18413 ( .a(n12921), .b(n12916), .o(n22202) );
no02f01 g18414 ( .a(n12922), .b(n12915), .o(n22203) );
no02f01 g18415 ( .a(n22203), .b(n22202), .o(n22204) );
no02f01 g18416 ( .a(n22204), .b(n22201), .o(n22205) );
na02f01 g18417 ( .a(n22204), .b(n22201), .o(n22206) );
in01f01 g18418 ( .a(n22206), .o(n22207) );
no02f01 g18419 ( .a(n22207), .b(n22205), .o(n22208) );
no02f01 g18420 ( .a(n22208), .b(n22200), .o(n22209) );
ao12f01 g18421 ( .a(n14172), .b(n14087), .c(n11514), .o(n22210) );
no03f01 g18422 ( .a(n14173), .b(n14086), .c(n11515), .o(n22211) );
no02f01 g18423 ( .a(n22211), .b(n22210), .o(n22212) );
no02f01 g18424 ( .a(n12906), .b(n12895), .o(n22213) );
in01f01 g18425 ( .a(n12906), .o(n22214) );
ao12f01 g18426 ( .a(n22214), .b(n12894), .c(n12893), .o(n22215) );
no02f01 g18427 ( .a(n22215), .b(n22213), .o(n22216) );
no02f01 g18428 ( .a(n22216), .b(n12900), .o(n22217) );
na02f01 g18429 ( .a(n22216), .b(n12900), .o(n22218) );
in01f01 g18430 ( .a(n22218), .o(n22219) );
no02f01 g18431 ( .a(n22219), .b(n22217), .o(n22220) );
in01f01 g18432 ( .a(n22220), .o(n22221) );
no02f01 g18433 ( .a(n22221), .b(n22212), .o(n22222) );
na02f01 g18434 ( .a(n14086), .b(n11515), .o(n22223) );
na02f01 g18435 ( .a(n14086), .b(n11514), .o(n22224) );
na02f01 g18436 ( .a(n22224), .b(n22223), .o(n22225) );
in01f01 g18437 ( .a(n12899), .o(n22226) );
no02f01 g18438 ( .a(n22226), .b(n12295), .o(n22227) );
no02f01 g18439 ( .a(n12899), .b(n12296), .o(n22228) );
no02f01 g18440 ( .a(n22228), .b(n22227), .o(n22229) );
no02f01 g18441 ( .a(n22229), .b(n22225), .o(n22230) );
na02f01 g18442 ( .a(n22221), .b(n22212), .o(n22231) );
oa12f01 g18443 ( .a(n22231), .b(n22230), .c(n22222), .o(n22232) );
na02f01 g18444 ( .a(n22208), .b(n22200), .o(n22233) );
ao12f01 g18445 ( .a(n22209), .b(n22233), .c(n22232), .o(n22234) );
na02f01 g18446 ( .a(n22194), .b(n22186), .o(n22235) );
ao12f01 g18447 ( .a(n22195), .b(n22235), .c(n22234), .o(n22236) );
ao12f01 g18448 ( .a(n22177), .b(n22236), .c(n22178), .o(n22237) );
na02f01 g18449 ( .a(n22163), .b(n13047), .o(n22238) );
ao12f01 g18450 ( .a(n22164), .b(n22238), .c(n22237), .o(n22239) );
ao12f01 g18451 ( .a(n21869), .b(n21860), .c(n22157), .o(n22240) );
no02f01 g18452 ( .a(n21865), .b(n21861), .o(n22241) );
no02f01 g18453 ( .a(n22241), .b(n22240), .o(n22242) );
na02f01 g18454 ( .a(n22241), .b(n22240), .o(n22243) );
in01f01 g18455 ( .a(n22243), .o(n22244) );
no02f01 g18456 ( .a(n22244), .b(n22242), .o(n22245) );
no02f01 g18457 ( .a(n22245), .b(n13054), .o(n22246) );
in01f01 g18458 ( .a(n22246), .o(n22247) );
na02f01 g18459 ( .a(n22154), .b(n13065), .o(n22248) );
na02f01 g18460 ( .a(n22245), .b(n13054), .o(n22249) );
na02f01 g18461 ( .a(n22249), .b(n22248), .o(n22250) );
ao12f01 g18462 ( .a(n22250), .b(n22247), .c(n22239), .o(n22251) );
in01f01 g18463 ( .a(n22145), .o(n22252) );
ao12f01 g18464 ( .a(n13074), .b(n22146), .c(n22252), .o(n22253) );
no03f01 g18465 ( .a(n22253), .b(n22251), .c(n22155), .o(n22254) );
in01f01 g18466 ( .a(n13085), .o(n22255) );
in01f01 g18467 ( .a(n21885), .o(n22256) );
na02f01 g18468 ( .a(n22256), .b(n22134), .o(n22257) );
no02f01 g18469 ( .a(n21884), .b(n21877), .o(n22258) );
in01f01 g18470 ( .a(n22258), .o(n22259) );
na02f01 g18471 ( .a(n22259), .b(n22257), .o(n22260) );
in01f01 g18472 ( .a(n22260), .o(n22261) );
no02f01 g18473 ( .a(n22259), .b(n22257), .o(n22262) );
no02f01 g18474 ( .a(n22262), .b(n22261), .o(n22263) );
na02f01 g18475 ( .a(n22263), .b(n22255), .o(n22264) );
in01f01 g18476 ( .a(n22264), .o(n22265) );
no03f01 g18477 ( .a(n22265), .b(n22254), .c(n22148), .o(n22266) );
no02f01 g18478 ( .a(n22263), .b(n22255), .o(n22267) );
in01f01 g18479 ( .a(n13092), .o(n22268) );
no02f01 g18480 ( .a(n22141), .b(n22140), .o(n22269) );
no02f01 g18481 ( .a(n22269), .b(n22268), .o(n22270) );
no03f01 g18482 ( .a(n22270), .b(n22267), .c(n22266), .o(n22271) );
na02f01 g18483 ( .a(n22132), .b(n22125), .o(n22272) );
in01f01 g18484 ( .a(n22272), .o(n22273) );
no03f01 g18485 ( .a(n22273), .b(n22271), .c(n22142), .o(n22274) );
in01f01 g18486 ( .a(n21892), .o(n22275) );
no02f01 g18487 ( .a(n21905), .b(n21893), .o(n22276) );
no02f01 g18488 ( .a(n22276), .b(n22275), .o(n22277) );
na02f01 g18489 ( .a(n22276), .b(n22275), .o(n22278) );
in01f01 g18490 ( .a(n22278), .o(n22279) );
no02f01 g18491 ( .a(n22279), .b(n22277), .o(n22280) );
no02f01 g18492 ( .a(n22280), .b(n13118), .o(n22281) );
no03f01 g18493 ( .a(n22281), .b(n22274), .c(n22133), .o(n22282) );
no02f01 g18494 ( .a(n21904), .b(n21895), .o(n22283) );
ao12f01 g18495 ( .a(n21905), .b(n21894), .c(n21892), .o(n22284) );
no02f01 g18496 ( .a(n22284), .b(n22283), .o(n22285) );
na02f01 g18497 ( .a(n22284), .b(n22283), .o(n22286) );
in01f01 g18498 ( .a(n22286), .o(n22287) );
no02f01 g18499 ( .a(n22287), .b(n22285), .o(n22288) );
in01f01 g18500 ( .a(n22288), .o(n22289) );
no02f01 g18501 ( .a(n22289), .b(n13130), .o(n22290) );
na02f01 g18502 ( .a(n22280), .b(n13118), .o(n22291) );
in01f01 g18503 ( .a(n22291), .o(n22292) );
no02f01 g18504 ( .a(n22292), .b(n22290), .o(n22293) );
in01f01 g18505 ( .a(n22293), .o(n22294) );
na02f01 g18506 ( .a(n22289), .b(n13130), .o(n22295) );
oa12f01 g18507 ( .a(n22295), .b(n22294), .c(n22282), .o(n22296) );
no03f01 g18508 ( .a(n21895), .b(n21893), .c(n22275), .o(n22297) );
no04f01 g18509 ( .a(n22082), .b(n21902), .c(n21899), .d(n22297), .o(n22298) );
no02f01 g18510 ( .a(n22082), .b(n22297), .o(n22299) );
ao12f01 g18511 ( .a(n22299), .b(n21903), .c(n22079), .o(n22300) );
no02f01 g18512 ( .a(n22300), .b(n22298), .o(n22301) );
no02f01 g18513 ( .a(n22301), .b(n13140), .o(n22302) );
in01f01 g18514 ( .a(n13150), .o(n22303) );
ao12f01 g18515 ( .a(n21899), .b(n22299), .c(n21903), .o(n22304) );
in01f01 g18516 ( .a(n22304), .o(n22305) );
no02f01 g18517 ( .a(n22081), .b(n21898), .o(n22306) );
no02f01 g18518 ( .a(n22306), .b(n22305), .o(n22307) );
na02f01 g18519 ( .a(n22306), .b(n22305), .o(n22308) );
in01f01 g18520 ( .a(n22308), .o(n22309) );
no02f01 g18521 ( .a(n22309), .b(n22307), .o(n22310) );
na02f01 g18522 ( .a(n22310), .b(n22303), .o(n22311) );
in01f01 g18523 ( .a(n22311), .o(n22312) );
na02f01 g18524 ( .a(n22301), .b(n13140), .o(n22313) );
in01f01 g18525 ( .a(n22313), .o(n22314) );
no02f01 g18526 ( .a(n22314), .b(n22312), .o(n22315) );
oa12f01 g18527 ( .a(n22315), .b(n22302), .c(n22296), .o(n22316) );
no02f01 g18528 ( .a(n22310), .b(n22303), .o(n22317) );
in01f01 g18529 ( .a(n22317), .o(n22318) );
no02f01 g18530 ( .a(n21925), .b(n21915), .o(n22319) );
in01f01 g18531 ( .a(n22319), .o(n22320) );
ao12f01 g18532 ( .a(n21926), .b(n22085), .c(n22084), .o(n22321) );
in01f01 g18533 ( .a(n22321), .o(n22322) );
no02f01 g18534 ( .a(n22322), .b(n22320), .o(n22323) );
no02f01 g18535 ( .a(n22321), .b(n22319), .o(n22324) );
no02f01 g18536 ( .a(n22324), .b(n22323), .o(n22325) );
no02f01 g18537 ( .a(n22325), .b(n13174), .o(n22326) );
in01f01 g18538 ( .a(n13158), .o(n22327) );
no02f01 g18539 ( .a(n21926), .b(n21909), .o(n22328) );
no02f01 g18540 ( .a(n22328), .b(n21908), .o(n22329) );
in01f01 g18541 ( .a(n22329), .o(n22330) );
na02f01 g18542 ( .a(n22328), .b(n21908), .o(n22331) );
ao12f01 g18543 ( .a(n22327), .b(n22331), .c(n22330), .o(n22332) );
no02f01 g18544 ( .a(n22332), .b(n22326), .o(n22333) );
na03f01 g18545 ( .a(n22333), .b(n22318), .c(n22316), .o(n22334) );
no02f01 g18546 ( .a(n22090), .b(n22089), .o(n22335) );
no02f01 g18547 ( .a(n22091), .b(n21847), .o(n22336) );
na02f01 g18548 ( .a(n22336), .b(n22335), .o(n22337) );
oa22f01 g18549 ( .a(n22091), .b(n21847), .c(n22090), .d(n22089), .o(n22338) );
na02f01 g18550 ( .a(n22338), .b(n22337), .o(n22339) );
na02f01 g18551 ( .a(n22339), .b(n13198), .o(n22340) );
no02f01 g18552 ( .a(n21928), .b(n21916), .o(n22341) );
no02f01 g18553 ( .a(n21924), .b(n22088), .o(n22342) );
no02f01 g18554 ( .a(n22342), .b(n22341), .o(n22343) );
na02f01 g18555 ( .a(n22342), .b(n22341), .o(n22344) );
in01f01 g18556 ( .a(n22344), .o(n22345) );
no02f01 g18557 ( .a(n22345), .b(n22343), .o(n22346) );
no02f01 g18558 ( .a(n22346), .b(n13201), .o(n22347) );
in01f01 g18559 ( .a(n22347), .o(n22348) );
na02f01 g18560 ( .a(n22348), .b(n22340), .o(n22349) );
na03f01 g18561 ( .a(n22338), .b(n22337), .c(n13192), .o(n22350) );
na02f01 g18562 ( .a(n22325), .b(n13174), .o(n22351) );
in01f01 g18563 ( .a(n22331), .o(n22352) );
no03f01 g18564 ( .a(n22352), .b(n22329), .c(n13158), .o(n22353) );
in01f01 g18565 ( .a(n22353), .o(n22354) );
ao12f01 g18566 ( .a(n22326), .b(n22354), .c(n22351), .o(n22355) );
no03f01 g18567 ( .a(n22345), .b(n22343), .c(n13183), .o(n22356) );
ao12f01 g18568 ( .a(n22356), .b(n22355), .c(n22348), .o(n22357) );
na02f01 g18569 ( .a(n22357), .b(n22350), .o(n22358) );
na02f01 g18570 ( .a(n22358), .b(n22340), .o(n22359) );
oa12f01 g18571 ( .a(n22359), .b(n22349), .c(n22334), .o(n22360) );
no02f01 g18572 ( .a(n22114), .b(n22107), .o(n22361) );
in01f01 g18573 ( .a(n22361), .o(n22362) );
na03f01 g18574 ( .a(n22362), .b(n22360), .c(n22124), .o(n22363) );
oa12f01 g18575 ( .a(n22118), .b(n22068), .c(n13517), .o(n22364) );
no02f01 g18576 ( .a(n22364), .b(n22363), .o(n22365) );
no02f01 g18577 ( .a(n22365), .b(n22120), .o(n22366) );
no02f01 g18578 ( .a(n21986), .b(n21836), .o(n22367) );
na02f01 g18579 ( .a(n22367), .b(n21974), .o(n22368) );
na02f01 g18580 ( .a(n22097), .b(n22094), .o(n22369) );
ao12f01 g18581 ( .a(n22369), .b(n21962), .c(n11514), .o(n22370) );
oa12f01 g18582 ( .a(n22370), .b(n21959), .c(n11515), .o(n22371) );
oa12f01 g18583 ( .a(n11515), .b(n22098), .c(n21939), .o(n22372) );
oa12f01 g18584 ( .a(n22372), .b(n21954), .c(n11514), .o(n22373) );
ao12f01 g18585 ( .a(n22373), .b(n21841), .c(n11515), .o(n22374) );
na02f01 g18586 ( .a(n22374), .b(n22371), .o(n22375) );
na02f01 g18587 ( .a(n21985), .b(n21984), .o(n22376) );
na02f01 g18588 ( .a(n22376), .b(n11514), .o(n22377) );
oa12f01 g18589 ( .a(n11515), .b(n21834), .c(n21832), .o(n22378) );
na02f01 g18590 ( .a(n22378), .b(n22377), .o(n22379) );
na02f01 g18591 ( .a(n22379), .b(n22375), .o(n22380) );
ao12f01 g18592 ( .a(n13510), .b(n22380), .c(n22368), .o(n22381) );
na03f01 g18593 ( .a(n22378), .b(n22374), .c(n22371), .o(n22382) );
no02f01 g18594 ( .a(n21977), .b(n21814), .o(n22383) );
no02f01 g18595 ( .a(n21978), .b(n21821), .o(n22384) );
oa12f01 g18596 ( .a(n11514), .b(n22384), .c(n22383), .o(n22385) );
oa12f01 g18597 ( .a(n11515), .b(n22384), .c(n22383), .o(n22386) );
na02f01 g18598 ( .a(n22386), .b(n22385), .o(n22387) );
na03f01 g18599 ( .a(n22387), .b(n22382), .c(n22377), .o(n22388) );
no03f01 g18600 ( .a(n21986), .b(n21973), .c(n21956), .o(n22389) );
no02f01 g18601 ( .a(n21983), .b(n21981), .o(n22390) );
oa12f01 g18602 ( .a(n22390), .b(n22389), .c(n21836), .o(n22391) );
ao12f01 g18603 ( .a(n14251), .b(n22391), .c(n22388), .o(n22392) );
no03f01 g18604 ( .a(n22392), .b(n22381), .c(n22366), .o(n22393) );
no03f01 g18605 ( .a(n14304), .b(n22040), .c(n13580), .o(n22394) );
ao12f01 g18606 ( .a(n21756), .b(n22011), .c(n22010), .o(n22395) );
no02f01 g18607 ( .a(n22042), .b(n22395), .o(n22396) );
oa12f01 g18608 ( .a(n22396), .b(n22394), .c(n14305), .o(n22397) );
na03f01 g18609 ( .a(n14298), .b(n14255), .c(n13572), .o(n22398) );
na02f01 g18610 ( .a(n22012), .b(n22008), .o(n22399) );
na03f01 g18611 ( .a(n22399), .b(n22398), .c(n14301), .o(n22400) );
na02f01 g18612 ( .a(n22400), .b(n22397), .o(n22401) );
no02f01 g18613 ( .a(n22401), .b(n21993), .o(n22402) );
in01f01 g18614 ( .a(n22402), .o(n22403) );
na03f01 g18615 ( .a(n14306), .b(n14255), .c(n13572), .o(n22404) );
na02f01 g18616 ( .a(n14302), .b(n14256), .o(n22405) );
na02f01 g18617 ( .a(n22405), .b(n22404), .o(n22406) );
ao12f01 g18618 ( .a(n11515), .b(n21991), .c(n21990), .o(n22407) );
oa22f01 g18619 ( .a(n21992), .b(n22407), .c(n21988), .d(n21982), .o(n22408) );
na03f01 g18620 ( .a(n22385), .b(n22375), .c(n22377), .o(n22409) );
oa12f01 g18621 ( .a(n11515), .b(n21823), .c(n21816), .o(n22410) );
na04f01 g18622 ( .a(n22410), .b(n21987), .c(n22409), .d(n21824), .o(n22411) );
ao12f01 g18623 ( .a(n22406), .b(n22411), .c(n22408), .o(n22412) );
no02f01 g18624 ( .a(n22412), .b(n22402), .o(n22413) );
na02f01 g18625 ( .a(n22401), .b(n21993), .o(n22414) );
in01f01 g18626 ( .a(n22392), .o(n22415) );
ao22f01 g18627 ( .a(n22410), .b(n21824), .c(n21987), .d(n22409), .o(n22416) );
no04f01 g18628 ( .a(n21992), .b(n21988), .c(n21982), .d(n22407), .o(n22417) );
oa12f01 g18629 ( .a(n14308), .b(n22417), .c(n22416), .o(n22418) );
na03f01 g18630 ( .a(n22391), .b(n22388), .c(n14251), .o(n22419) );
na03f01 g18631 ( .a(n22380), .b(n22368), .c(n13510), .o(n22420) );
na02f01 g18632 ( .a(n22420), .b(n22419), .o(n22421) );
na03f01 g18633 ( .a(n22421), .b(n22418), .c(n22415), .o(n22422) );
no03f01 g18634 ( .a(n22417), .b(n22416), .c(n14308), .o(n22423) );
in01f01 g18635 ( .a(n22423), .o(n22424) );
na03f01 g18636 ( .a(n22424), .b(n22422), .c(n22414), .o(n22425) );
ao22f01 g18637 ( .a(n22425), .b(n22403), .c(n22413), .d(n22393), .o(n22426) );
na03f01 g18638 ( .a(n22033), .b(n22032), .c(n21702), .o(n22427) );
oa12f01 g18639 ( .a(n21701), .b(n22027), .c(n22022), .o(n22428) );
na02f01 g18640 ( .a(n22428), .b(n22427), .o(n22429) );
na03f01 g18641 ( .a(n22429), .b(n22044), .c(n22008), .o(n22430) );
no03f01 g18642 ( .a(n22027), .b(n22022), .c(n21701), .o(n22431) );
ao12f01 g18643 ( .a(n21702), .b(n22033), .c(n22032), .o(n22432) );
no02f01 g18644 ( .a(n22432), .b(n22431), .o(n22433) );
na02f01 g18645 ( .a(n22433), .b(n22014), .o(n22434) );
na02f01 g18646 ( .a(n22434), .b(n22430), .o(n22435) );
in01f01 g18647 ( .a(n22435), .o(n22436) );
no02f01 g18648 ( .a(n22013), .b(n22009), .o(n22437) );
no03f01 g18649 ( .a(n22432), .b(n22437), .c(n22395), .o(n22438) );
no02f01 g18650 ( .a(n22034), .b(n21676), .o(n22439) );
no02f01 g18651 ( .a(n22028), .b(n22015), .o(n22440) );
no02f01 g18652 ( .a(n22440), .b(n22439), .o(n22441) );
in01f01 g18653 ( .a(n22441), .o(n22442) );
no03f01 g18654 ( .a(n22442), .b(n22438), .c(n22431), .o(n22443) );
na03f01 g18655 ( .a(n22428), .b(n22044), .c(n22008), .o(n22444) );
ao12f01 g18656 ( .a(n22441), .b(n22444), .c(n22427), .o(n22445) );
no02f01 g18657 ( .a(n22445), .b(n22443), .o(n22446) );
ao12f01 g18658 ( .a(n22050), .b(n22446), .c(n22436), .o(n22447) );
in01f01 g18659 ( .a(n22447), .o(n22448) );
na02f01 g18660 ( .a(n22448), .b(n22426), .o(n22449) );
na03f01 g18661 ( .a(n22441), .b(n22444), .c(n22427), .o(n22450) );
oa12f01 g18662 ( .a(n22442), .b(n22438), .c(n22431), .o(n22451) );
na02f01 g18663 ( .a(n22451), .b(n22450), .o(n22452) );
ao12f01 g18664 ( .a(n21993), .b(n22452), .c(n22435), .o(n22453) );
in01f01 g18665 ( .a(n22453), .o(n22454) );
ao12f01 g18666 ( .a(n22056), .b(n22454), .c(n22449), .o(n22455) );
in01f01 g18667 ( .a(n22065), .o(n22456) );
na02f01 g18668 ( .a(n22064), .b(n22059), .o(n22457) );
na02f01 g18669 ( .a(n22457), .b(n22456), .o(n22458) );
no02f01 g18670 ( .a(n22458), .b(n13424), .o(n22459) );
no02f01 g18671 ( .a(n22074), .b(n22063), .o(n22460) );
no02f01 g18672 ( .a(n22072), .b(n22071), .o(n22461) );
no02f01 g18673 ( .a(n22461), .b(n22460), .o(n22462) );
na02f01 g18674 ( .a(n22462), .b(n13520), .o(n22463) );
no02f01 g18675 ( .a(n22123), .b(n13276), .o(n22464) );
in01f01 g18676 ( .a(n22115), .o(n22465) );
oa12f01 g18677 ( .a(n22124), .b(n22465), .c(n22464), .o(n22466) );
no02f01 g18678 ( .a(n22462), .b(n13520), .o(n22467) );
oa12f01 g18679 ( .a(n22463), .b(n22467), .c(n22466), .o(n22468) );
no02f01 g18680 ( .a(n22468), .b(n22459), .o(n22469) );
oa22f01 g18681 ( .a(n22364), .b(n22363), .c(n22469), .d(n22069), .o(n22470) );
in01f01 g18682 ( .a(n22381), .o(n22471) );
na03f01 g18683 ( .a(n22415), .b(n22471), .c(n22470), .o(n22472) );
in01f01 g18684 ( .a(n22413), .o(n22473) );
in01f01 g18685 ( .a(n22414), .o(n22474) );
no03f01 g18686 ( .a(n22390), .b(n22389), .c(n21836), .o(n22475) );
ao12f01 g18687 ( .a(n22387), .b(n22382), .c(n22377), .o(n22476) );
no03f01 g18688 ( .a(n22476), .b(n22475), .c(n13586), .o(n22477) );
no02f01 g18689 ( .a(n22379), .b(n22375), .o(n22478) );
no02f01 g18690 ( .a(n22367), .b(n21974), .o(n22479) );
no03f01 g18691 ( .a(n22479), .b(n22478), .c(n13514), .o(n22480) );
no02f01 g18692 ( .a(n22480), .b(n22477), .o(n22481) );
no03f01 g18693 ( .a(n22481), .b(n22412), .c(n22392), .o(n22482) );
no03f01 g18694 ( .a(n22423), .b(n22482), .c(n22474), .o(n22483) );
oa22f01 g18695 ( .a(n22483), .b(n22402), .c(n22473), .d(n22472), .o(n22484) );
no02f01 g18696 ( .a(n22447), .b(n22484), .o(n22485) );
no03f01 g18697 ( .a(n22453), .b(n22485), .c(n22055), .o(n22486) );
oa12f01 g18698 ( .a(n4116), .b(n22486), .c(n22455), .o(n22487) );
oa12f01 g18699 ( .a(n22055), .b(n22453), .c(n22485), .o(n22488) );
na03f01 g18700 ( .a(n22454), .b(n22449), .c(n22056), .o(n22489) );
na03f01 g18701 ( .a(n22489), .b(n22488), .c(n2589), .o(n22490) );
na02f01 g18702 ( .a(n22490), .b(n22487), .o(n288) );
in01f01 g18703 ( .a(n18265), .o(n22492) );
no02f01 g18704 ( .a(n18317), .b(n22492), .o(n22493) );
no02f01 g18705 ( .a(n18283), .b(n18103), .o(n22494) );
no02f01 g18706 ( .a(n22494), .b(n18285), .o(n22495) );
no02f01 g18707 ( .a(n22495), .b(n22493), .o(n22496) );
na02f01 g18708 ( .a(n22495), .b(n22493), .o(n22497) );
in01f01 g18709 ( .a(n22497), .o(n22498) );
no02f01 g18710 ( .a(n22498), .b(n22496), .o(n22499) );
in01f01 g18711 ( .a(n22499), .o(n22500) );
no02f01 g18712 ( .a(n22500), .b(n18460), .o(n22501) );
in01f01 g18713 ( .a(n18221), .o(n22502) );
no02f01 g18714 ( .a(n22502), .b(n18156), .o(n22503) );
in01f01 g18715 ( .a(n22503), .o(n22504) );
in01f01 g18716 ( .a(n18242), .o(n22505) );
no02f01 g18717 ( .a(n22505), .b(n22504), .o(n22506) );
in01f01 g18718 ( .a(n22506), .o(n22507) );
no02f01 g18719 ( .a(n18261), .b(n18103), .o(n22508) );
no02f01 g18720 ( .a(n22508), .b(n18314), .o(n22509) );
oa12f01 g18721 ( .a(n22509), .b(n18263), .c(n22507), .o(n22510) );
in01f01 g18722 ( .a(n22510), .o(n22511) );
no02f01 g18723 ( .a(n18252), .b(n18103), .o(n22512) );
no02f01 g18724 ( .a(n22512), .b(n18254), .o(n22513) );
no02f01 g18725 ( .a(n22513), .b(n22511), .o(n22514) );
na02f01 g18726 ( .a(n22513), .b(n22511), .o(n22515) );
in01f01 g18727 ( .a(n22515), .o(n22516) );
no02f01 g18728 ( .a(n22516), .b(n22514), .o(n22517) );
no02f01 g18729 ( .a(n22517), .b(n18459), .o(n22518) );
no02f01 g18730 ( .a(n18230), .b(n18103), .o(n22519) );
no02f01 g18731 ( .a(n22519), .b(n18232), .o(n22520) );
no02f01 g18732 ( .a(n22520), .b(n22504), .o(n22521) );
na02f01 g18733 ( .a(n22520), .b(n22504), .o(n22522) );
in01f01 g18734 ( .a(n22522), .o(n22523) );
no02f01 g18735 ( .a(n22523), .b(n22521), .o(n22524) );
in01f01 g18736 ( .a(n22524), .o(n22525) );
no02f01 g18737 ( .a(n22525), .b(n18460), .o(n22526) );
no02f01 g18738 ( .a(n18216), .b(n18103), .o(n22527) );
in01f01 g18739 ( .a(n22527), .o(n22528) );
ao12f01 g18740 ( .a(n18218), .b(n22528), .c(n18210), .o(n22529) );
in01f01 g18741 ( .a(n22529), .o(n22530) );
no02f01 g18742 ( .a(n18154), .b(n18145), .o(n22531) );
no02f01 g18743 ( .a(n22531), .b(n18156), .o(n22532) );
no02f01 g18744 ( .a(n22532), .b(n22530), .o(n22533) );
na02f01 g18745 ( .a(n22532), .b(n22530), .o(n22534) );
in01f01 g18746 ( .a(n22534), .o(n22535) );
no02f01 g18747 ( .a(n22535), .b(n22533), .o(n22536) );
no02f01 g18748 ( .a(n22536), .b(n18459), .o(n22537) );
in01f01 g18749 ( .a(n22537), .o(n22538) );
no02f01 g18750 ( .a(n18206), .b(n18204), .o(n22539) );
no02f01 g18751 ( .a(n22539), .b(n18194), .o(n22540) );
na02f01 g18752 ( .a(n22539), .b(n18194), .o(n22541) );
in01f01 g18753 ( .a(n22541), .o(n22542) );
no02f01 g18754 ( .a(n22542), .b(n22540), .o(n22543) );
no02f01 g18755 ( .a(n22543), .b(n18460), .o(n22544) );
in01f01 g18756 ( .a(n22544), .o(n22545) );
no02f01 g18757 ( .a(n18192), .b(n18173), .o(n22546) );
no02f01 g18758 ( .a(n22546), .b(n18190), .o(n22547) );
na02f01 g18759 ( .a(n22546), .b(n18190), .o(n22548) );
in01f01 g18760 ( .a(n22548), .o(n22549) );
no02f01 g18761 ( .a(n22549), .b(n22547), .o(n22550) );
no02f01 g18762 ( .a(n22550), .b(n18459), .o(n22551) );
no02f01 g18763 ( .a(n18188), .b(n18178), .o(n22552) );
in01f01 g18764 ( .a(n22552), .o(n22553) );
no02f01 g18765 ( .a(n22553), .b(n18186), .o(n22554) );
na02f01 g18766 ( .a(n22553), .b(n18186), .o(n22555) );
in01f01 g18767 ( .a(n22555), .o(n22556) );
no02f01 g18768 ( .a(n22556), .b(n22554), .o(n22557) );
in01f01 g18769 ( .a(n22557), .o(n22558) );
no02f01 g18770 ( .a(n22558), .b(n18459), .o(n22559) );
in01f01 g18771 ( .a(n18185), .o(n22560) );
no03f01 g18772 ( .a(n22560), .b(n18184), .c(delay_sub_ln23_0_unr5_stage3_stallmux_q_0_), .o(n22561) );
no02f01 g18773 ( .a(n22560), .b(n18184), .o(n22562) );
no02f01 g18774 ( .a(n22562), .b(n4498), .o(n22563) );
no02f01 g18775 ( .a(n22563), .b(n22561), .o(n4448) );
na02f01 g18776 ( .a(n22558), .b(n18459), .o(n22565) );
oa12f01 g18777 ( .a(n22565), .b(n4448), .c(n22559), .o(n22566) );
na02f01 g18778 ( .a(n22550), .b(n18459), .o(n22567) );
ao12f01 g18779 ( .a(n22551), .b(n22567), .c(n22566), .o(n22568) );
na02f01 g18780 ( .a(n22543), .b(n18460), .o(n22569) );
in01f01 g18781 ( .a(n22569), .o(n22570) );
oa12f01 g18782 ( .a(n22545), .b(n22570), .c(n22568), .o(n22571) );
in01f01 g18783 ( .a(n18210), .o(n22572) );
no02f01 g18784 ( .a(n22527), .b(n18218), .o(n22573) );
in01f01 g18785 ( .a(n22573), .o(n22574) );
no02f01 g18786 ( .a(n22574), .b(n22572), .o(n22575) );
no02f01 g18787 ( .a(n22573), .b(n18210), .o(n22576) );
no02f01 g18788 ( .a(n22576), .b(n22575), .o(n22577) );
in01f01 g18789 ( .a(n22577), .o(n22578) );
no02f01 g18790 ( .a(n22578), .b(n18460), .o(n22579) );
no02f01 g18791 ( .a(n18206), .b(n18205), .o(n22580) );
no02f01 g18792 ( .a(n18207), .b(n18165), .o(n22581) );
no02f01 g18793 ( .a(n22581), .b(n22580), .o(n22582) );
na02f01 g18794 ( .a(n22581), .b(n22580), .o(n22583) );
in01f01 g18795 ( .a(n22583), .o(n22584) );
no02f01 g18796 ( .a(n22584), .b(n22582), .o(n22585) );
in01f01 g18797 ( .a(n22585), .o(n22586) );
no02f01 g18798 ( .a(n22586), .b(n18460), .o(n22587) );
no02f01 g18799 ( .a(n22587), .b(n22579), .o(n22588) );
na02f01 g18800 ( .a(n22588), .b(n22571), .o(n22589) );
no02f01 g18801 ( .a(n22577), .b(n18459), .o(n22590) );
no02f01 g18802 ( .a(n22585), .b(n18459), .o(n22591) );
no02f01 g18803 ( .a(n22591), .b(n22590), .o(n22592) );
na02f01 g18804 ( .a(n22592), .b(n22589), .o(n22593) );
na02f01 g18805 ( .a(n22536), .b(n18459), .o(n22594) );
na02f01 g18806 ( .a(n22594), .b(n22593), .o(n22595) );
na02f01 g18807 ( .a(n22595), .b(n22538), .o(n22596) );
in01f01 g18808 ( .a(n22596), .o(n22597) );
no02f01 g18809 ( .a(n22524), .b(n18459), .o(n22598) );
in01f01 g18810 ( .a(n22598), .o(n22599) );
ao12f01 g18811 ( .a(n22526), .b(n22599), .c(n22597), .o(n22600) );
no02f01 g18812 ( .a(n18314), .b(n22506), .o(n22601) );
no02f01 g18813 ( .a(n22508), .b(n18263), .o(n22602) );
no02f01 g18814 ( .a(n22602), .b(n22601), .o(n22603) );
na02f01 g18815 ( .a(n22602), .b(n22601), .o(n22604) );
in01f01 g18816 ( .a(n22604), .o(n22605) );
no02f01 g18817 ( .a(n22605), .b(n22603), .o(n22606) );
in01f01 g18818 ( .a(n22606), .o(n22607) );
no02f01 g18819 ( .a(n22607), .b(n18460), .o(n22608) );
in01f01 g18820 ( .a(n18232), .o(n22609) );
ao12f01 g18821 ( .a(n22519), .b(n22609), .c(n22503), .o(n22610) );
in01f01 g18822 ( .a(n22610), .o(n22611) );
no02f01 g18823 ( .a(n18239), .b(n18103), .o(n22612) );
no02f01 g18824 ( .a(n22612), .b(n18241), .o(n22613) );
in01f01 g18825 ( .a(n22613), .o(n22614) );
no02f01 g18826 ( .a(n22614), .b(n22611), .o(n22615) );
no02f01 g18827 ( .a(n22613), .b(n22610), .o(n22616) );
no02f01 g18828 ( .a(n22616), .b(n22615), .o(n22617) );
in01f01 g18829 ( .a(n22617), .o(n22618) );
no02f01 g18830 ( .a(n22618), .b(n18460), .o(n22619) );
no02f01 g18831 ( .a(n22619), .b(n22608), .o(n22620) );
na02f01 g18832 ( .a(n22620), .b(n22600), .o(n22621) );
no02f01 g18833 ( .a(n22606), .b(n18459), .o(n22622) );
no02f01 g18834 ( .a(n22617), .b(n18459), .o(n22623) );
no02f01 g18835 ( .a(n22623), .b(n22622), .o(n22624) );
na02f01 g18836 ( .a(n22624), .b(n22621), .o(n22625) );
na02f01 g18837 ( .a(n22517), .b(n18459), .o(n22626) );
na02f01 g18838 ( .a(n22626), .b(n22625), .o(n22627) );
in01f01 g18839 ( .a(n22627), .o(n22628) );
no02f01 g18840 ( .a(n22628), .b(n22518), .o(n22629) );
in01f01 g18841 ( .a(n22629), .o(n22630) );
no02f01 g18842 ( .a(n22499), .b(n18459), .o(n22631) );
no02f01 g18843 ( .a(n22631), .b(n22630), .o(n22632) );
no02f01 g18844 ( .a(n22494), .b(n18317), .o(n22633) );
oa12f01 g18845 ( .a(n22633), .b(n18285), .c(n18265), .o(n22634) );
no02f01 g18846 ( .a(n18273), .b(n18103), .o(n22635) );
no02f01 g18847 ( .a(n22635), .b(n18275), .o(n22636) );
in01f01 g18848 ( .a(n22636), .o(n22637) );
no02f01 g18849 ( .a(n22637), .b(n22634), .o(n22638) );
na02f01 g18850 ( .a(n22637), .b(n22634), .o(n22639) );
in01f01 g18851 ( .a(n22639), .o(n22640) );
no02f01 g18852 ( .a(n22640), .b(n22638), .o(n22641) );
in01f01 g18853 ( .a(n22641), .o(n22642) );
no02f01 g18854 ( .a(n22642), .b(n18460), .o(n22643) );
ao12f01 g18855 ( .a(n18320), .b(n18286), .c(n22492), .o(n22644) );
no02f01 g18856 ( .a(n18297), .b(n18103), .o(n22645) );
no02f01 g18857 ( .a(n22645), .b(n18299), .o(n22646) );
no02f01 g18858 ( .a(n22646), .b(n22644), .o(n22647) );
na02f01 g18859 ( .a(n22646), .b(n22644), .o(n22648) );
in01f01 g18860 ( .a(n22648), .o(n22649) );
no02f01 g18861 ( .a(n22649), .b(n22647), .o(n22650) );
in01f01 g18862 ( .a(n22650), .o(n22651) );
no02f01 g18863 ( .a(n22651), .b(n18460), .o(n22652) );
no04f01 g18864 ( .a(n22652), .b(n22643), .c(n22632), .d(n22501), .o(n22653) );
no02f01 g18865 ( .a(n22641), .b(n18459), .o(n22654) );
no02f01 g18866 ( .a(n22650), .b(n18459), .o(n22655) );
no02f01 g18867 ( .a(n22655), .b(n22654), .o(n22656) );
in01f01 g18868 ( .a(n22656), .o(n22657) );
no03f01 g18869 ( .a(n18299), .b(n18287), .c(n18265), .o(n22658) );
no02f01 g18870 ( .a(n22645), .b(n18320), .o(n22659) );
in01f01 g18871 ( .a(n22659), .o(n22660) );
no02f01 g18872 ( .a(n18308), .b(n18103), .o(n22661) );
no02f01 g18873 ( .a(n22661), .b(n18310), .o(n22662) );
in01f01 g18874 ( .a(n22662), .o(n22663) );
no03f01 g18875 ( .a(n22663), .b(n22660), .c(n22658), .o(n22664) );
no02f01 g18876 ( .a(n22660), .b(n22658), .o(n22665) );
no02f01 g18877 ( .a(n22662), .b(n22665), .o(n22666) );
no02f01 g18878 ( .a(n22666), .b(n22664), .o(n22667) );
in01f01 g18879 ( .a(n22667), .o(n22668) );
no02f01 g18880 ( .a(n22668), .b(n18460), .o(n22669) );
no02f01 g18881 ( .a(n18323), .b(n18313), .o(n22670) );
no02f01 g18882 ( .a(n18340), .b(n18103), .o(n22671) );
no02f01 g18883 ( .a(n22671), .b(n18342), .o(n22672) );
no02f01 g18884 ( .a(n22672), .b(n22670), .o(n22673) );
na02f01 g18885 ( .a(n22672), .b(n22670), .o(n22674) );
in01f01 g18886 ( .a(n22674), .o(n22675) );
no02f01 g18887 ( .a(n22675), .b(n22673), .o(n22676) );
in01f01 g18888 ( .a(n22676), .o(n22677) );
no02f01 g18889 ( .a(n22677), .b(n18460), .o(n22678) );
no02f01 g18890 ( .a(n22678), .b(n22669), .o(n22679) );
oa12f01 g18891 ( .a(n22679), .b(n22657), .c(n22653), .o(n22680) );
no02f01 g18892 ( .a(n22667), .b(n18459), .o(n22681) );
no02f01 g18893 ( .a(n22676), .b(n18459), .o(n22682) );
no02f01 g18894 ( .a(n22682), .b(n22681), .o(n22683) );
no02f01 g18895 ( .a(n18342), .b(n22670), .o(n22684) );
no02f01 g18896 ( .a(n22684), .b(n22671), .o(n22685) );
no02f01 g18897 ( .a(n18329), .b(n18103), .o(n22686) );
no02f01 g18898 ( .a(n22686), .b(n18331), .o(n22687) );
no02f01 g18899 ( .a(n22687), .b(n22685), .o(n22688) );
na02f01 g18900 ( .a(n22687), .b(n22685), .o(n22689) );
in01f01 g18901 ( .a(n22689), .o(n22690) );
no02f01 g18902 ( .a(n22690), .b(n22688), .o(n22691) );
in01f01 g18903 ( .a(n22691), .o(n22692) );
no02f01 g18904 ( .a(n22692), .b(n18460), .o(n22693) );
no02f01 g18905 ( .a(n18344), .b(n22670), .o(n22694) );
no02f01 g18906 ( .a(n22694), .b(n18365), .o(n22695) );
no02f01 g18907 ( .a(n18352), .b(n18103), .o(n22696) );
no02f01 g18908 ( .a(n22696), .b(n18354), .o(n22697) );
no02f01 g18909 ( .a(n22697), .b(n22695), .o(n22698) );
na02f01 g18910 ( .a(n22697), .b(n22695), .o(n22699) );
in01f01 g18911 ( .a(n22699), .o(n22700) );
no02f01 g18912 ( .a(n22700), .b(n22698), .o(n22701) );
in01f01 g18913 ( .a(n22701), .o(n22702) );
no02f01 g18914 ( .a(n22702), .b(n18460), .o(n22703) );
no02f01 g18915 ( .a(n22703), .b(n22693), .o(n22704) );
in01f01 g18916 ( .a(n22704), .o(n22705) );
ao12f01 g18917 ( .a(n22705), .b(n22683), .c(n22680), .o(n22706) );
no03f01 g18918 ( .a(n18354), .b(n18344), .c(n22670), .o(n22707) );
no02f01 g18919 ( .a(n22696), .b(n18365), .o(n22708) );
in01f01 g18920 ( .a(n22708), .o(n22709) );
no02f01 g18921 ( .a(n18360), .b(n18103), .o(n22710) );
no02f01 g18922 ( .a(n22710), .b(n18362), .o(n22711) );
in01f01 g18923 ( .a(n22711), .o(n22712) );
no03f01 g18924 ( .a(n22712), .b(n22709), .c(n22707), .o(n22713) );
no02f01 g18925 ( .a(n22709), .b(n22707), .o(n22714) );
no02f01 g18926 ( .a(n22711), .b(n22714), .o(n22715) );
no02f01 g18927 ( .a(n22715), .b(n22713), .o(n22716) );
in01f01 g18928 ( .a(n22716), .o(n22717) );
no02f01 g18929 ( .a(n22717), .b(n18460), .o(n22718) );
in01f01 g18930 ( .a(n18364), .o(n22719) );
in01f01 g18931 ( .a(n18367), .o(n22720) );
no02f01 g18932 ( .a(n22720), .b(n22719), .o(n22721) );
no02f01 g18933 ( .a(n18126), .b(n18103), .o(n22722) );
no02f01 g18934 ( .a(n18371), .b(n22722), .o(n22723) );
no02f01 g18935 ( .a(n22723), .b(n22721), .o(n22724) );
na02f01 g18936 ( .a(n22723), .b(n22721), .o(n22725) );
in01f01 g18937 ( .a(n22725), .o(n22726) );
no02f01 g18938 ( .a(n22726), .b(n22724), .o(n22727) );
in01f01 g18939 ( .a(n22727), .o(n22728) );
no02f01 g18940 ( .a(n22728), .b(n18460), .o(n22729) );
no02f01 g18941 ( .a(n22729), .b(n22718), .o(n22730) );
no02f01 g18942 ( .a(n22691), .b(n18459), .o(n22731) );
no02f01 g18943 ( .a(n22701), .b(n18459), .o(n22732) );
no02f01 g18944 ( .a(n22732), .b(n22731), .o(n22733) );
in01f01 g18945 ( .a(n22733), .o(n22734) );
no02f01 g18946 ( .a(n22716), .b(n18459), .o(n22735) );
no02f01 g18947 ( .a(n22727), .b(n18459), .o(n22736) );
no03f01 g18948 ( .a(n22736), .b(n22735), .c(n22734), .o(n22737) );
in01f01 g18949 ( .a(n22737), .o(n22738) );
ao12f01 g18950 ( .a(n22738), .b(n22730), .c(n22706), .o(n22739) );
no02f01 g18951 ( .a(n22720), .b(n22722), .o(n22740) );
oa12f01 g18952 ( .a(n22740), .b(n18371), .c(n18364), .o(n22741) );
in01f01 g18953 ( .a(n22741), .o(n22742) );
no02f01 g18954 ( .a(n18133), .b(n18103), .o(n22743) );
no02f01 g18955 ( .a(n22743), .b(n18369), .o(n22744) );
no02f01 g18956 ( .a(n22744), .b(n22742), .o(n22745) );
na02f01 g18957 ( .a(n22744), .b(n22742), .o(n22746) );
in01f01 g18958 ( .a(n22746), .o(n22747) );
no02f01 g18959 ( .a(n22747), .b(n22745), .o(n22748) );
no02f01 g18960 ( .a(n22748), .b(n18459), .o(n22749) );
na02f01 g18961 ( .a(n22748), .b(n18459), .o(n22750) );
in01f01 g18962 ( .a(n22750), .o(n22751) );
no02f01 g18963 ( .a(n22751), .b(n22749), .o(n22752) );
na02f01 g18964 ( .a(n22752), .b(n22739), .o(n22753) );
in01f01 g18965 ( .a(n22739), .o(n22754) );
in01f01 g18966 ( .a(n22752), .o(n22755) );
na02f01 g18967 ( .a(n22755), .b(n22754), .o(n22756) );
na02f01 g18968 ( .a(n22756), .b(n22753), .o(n293) );
in01f01 g18969 ( .a(n22316), .o(n22758) );
no02f01 g18970 ( .a(n22317), .b(n22758), .o(n22759) );
in01f01 g18971 ( .a(n22759), .o(n22760) );
no02f01 g18972 ( .a(n22353), .b(n22332), .o(n22761) );
no02f01 g18973 ( .a(n22761), .b(n22760), .o(n22762) );
na02f01 g18974 ( .a(n22761), .b(n22760), .o(n22763) );
in01f01 g18975 ( .a(n22763), .o(n22764) );
no02f01 g18976 ( .a(n22764), .b(n22762), .o(n22765) );
in01f01 g18977 ( .a(n22765), .o(n298) );
in01f01 g18978 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_23_), .o(n22767) );
in01f01 g18979 ( .a(delay_xor_ln21_unr9_stage4_stallmux_q_22_), .o(n22768) );
no02f01 g18980 ( .a(n_45224), .b(n22768), .o(n22769) );
no02f01 g18981 ( .a(n4997_1), .b(delay_xor_ln21_unr9_stage4_stallmux_q_15_), .o(n22770) );
no02f01 g18982 ( .a(n4997_1), .b(delay_xor_ln21_unr9_stage4_stallmux_q_12_), .o(n22771) );
no02f01 g18983 ( .a(n4997_1), .b(delay_xor_ln21_unr9_stage4_stallmux_q_8_), .o(n22772) );
in01f01 g18984 ( .a(delay_xor_ln21_unr9_stage4_stallmux_q_0_), .o(n22773) );
na02f01 g18985 ( .a(n_45224), .b(n22773), .o(n22774) );
in01f01 g18986 ( .a(delay_xor_ln21_unr9_stage4_stallmux_q_1_), .o(n22775) );
na02f01 g18987 ( .a(n_45224), .b(n22775), .o(n22776) );
na02f01 g18988 ( .a(n22776), .b(n22774), .o(n22777) );
no02f01 g18989 ( .a(n4997_1), .b(delay_xor_ln21_unr9_stage4_stallmux_q_4_), .o(n22778) );
no02f01 g18990 ( .a(n4997_1), .b(delay_xor_ln21_unr9_stage4_stallmux_q_3_), .o(n22779) );
no02f01 g18991 ( .a(n4997_1), .b(delay_xor_ln21_unr9_stage4_stallmux_q_2_), .o(n22780) );
no04f01 g18992 ( .a(n22780), .b(n22779), .c(n22778), .d(n22777), .o(n22781) );
in01f01 g18993 ( .a(n22781), .o(n22782) );
no02f01 g18994 ( .a(n4997_1), .b(delay_xor_ln21_unr9_stage4_stallmux_q_5_), .o(n22783) );
no02f01 g18995 ( .a(n22783), .b(n22782), .o(n22784) );
no02f01 g18996 ( .a(n4997_1), .b(delay_xor_ln21_unr9_stage4_stallmux_q_6_), .o(n22785) );
no02f01 g18997 ( .a(n4997_1), .b(delay_xor_ln21_unr9_stage4_stallmux_q_7_), .o(n22786) );
no02f01 g18998 ( .a(n22786), .b(n22785), .o(n22787) );
na02f01 g18999 ( .a(n22787), .b(n22784), .o(n22788) );
no02f01 g19000 ( .a(n22788), .b(n22772), .o(n22789) );
in01f01 g19001 ( .a(n22789), .o(n22790) );
no02f01 g19002 ( .a(n4997_1), .b(delay_xor_ln21_unr9_stage4_stallmux_q_9_), .o(n22791) );
no02f01 g19003 ( .a(n22791), .b(n22790), .o(n22792) );
in01f01 g19004 ( .a(n22792), .o(n22793) );
no02f01 g19005 ( .a(n4997_1), .b(delay_xor_ln21_unr9_stage4_stallmux_q_10_), .o(n22794) );
no02f01 g19006 ( .a(n22794), .b(n22793), .o(n22795) );
in01f01 g19007 ( .a(n22795), .o(n22796) );
no02f01 g19008 ( .a(n4997_1), .b(delay_xor_ln21_unr9_stage4_stallmux_q_11_), .o(n22797) );
no02f01 g19009 ( .a(n22797), .b(n22796), .o(n22798) );
in01f01 g19010 ( .a(n22798), .o(n22799) );
no02f01 g19011 ( .a(n22799), .b(n22771), .o(n22800) );
in01f01 g19012 ( .a(n22800), .o(n22801) );
no02f01 g19013 ( .a(n4997_1), .b(delay_xor_ln21_unr9_stage4_stallmux_q_13_), .o(n22802) );
no02f01 g19014 ( .a(n22802), .b(n22801), .o(n22803) );
in01f01 g19015 ( .a(n22803), .o(n22804) );
no02f01 g19016 ( .a(delay_xor_ln21_unr9_stage4_stallmux_q_14_), .b(n4997_1), .o(n22805) );
no02f01 g19017 ( .a(n22805), .b(n22804), .o(n22806) );
in01f01 g19018 ( .a(n22806), .o(n22807) );
no02f01 g19019 ( .a(n22807), .b(n22770), .o(n22808) );
in01f01 g19020 ( .a(n22808), .o(n22809) );
no02f01 g19021 ( .a(n4997_1), .b(delay_xor_ln21_unr9_stage4_stallmux_q_16_), .o(n22810) );
no02f01 g19022 ( .a(n22810), .b(n22809), .o(n22811) );
in01f01 g19023 ( .a(n22811), .o(n22812) );
no02f01 g19024 ( .a(n4997_1), .b(delay_xor_ln21_unr9_stage4_stallmux_q_17_), .o(n22813) );
no02f01 g19025 ( .a(n4997_1), .b(delay_xor_ln21_unr9_stage4_stallmux_q_18_), .o(n22814) );
no03f01 g19026 ( .a(n22814), .b(n22813), .c(n22812), .o(n22815) );
in01f01 g19027 ( .a(n22815), .o(n22816) );
no02f01 g19028 ( .a(n4997_1), .b(delay_xor_ln21_unr9_stage4_stallmux_q_19_), .o(n22817) );
no02f01 g19029 ( .a(n22817), .b(n22816), .o(n22818) );
in01f01 g19030 ( .a(n22818), .o(n22819) );
no02f01 g19031 ( .a(n4997_1), .b(delay_xor_ln21_unr9_stage4_stallmux_q_20_), .o(n22820) );
no02f01 g19032 ( .a(n4997_1), .b(delay_xor_ln21_unr9_stage4_stallmux_q_21_), .o(n22821) );
no03f01 g19033 ( .a(n22821), .b(n22820), .c(n22819), .o(n22822) );
no02f01 g19034 ( .a(n4997_1), .b(delay_xor_ln21_unr9_stage4_stallmux_q_22_), .o(n22823) );
no02f01 g19035 ( .a(n22823), .b(n22769), .o(n22824) );
in01f01 g19036 ( .a(n22824), .o(n22825) );
no02f01 g19037 ( .a(n22825), .b(n22822), .o(n22826) );
no02f01 g19038 ( .a(n22826), .b(n22769), .o(n22827) );
in01f01 g19039 ( .a(n22827), .o(n22828) );
in01f01 g19040 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_22_), .o(n22829) );
na02f01 g19041 ( .a(n22825), .b(n22822), .o(n22830) );
in01f01 g19042 ( .a(n22830), .o(n22831) );
no02f01 g19043 ( .a(n22831), .b(n22826), .o(n22832) );
in01f01 g19044 ( .a(n22832), .o(n22833) );
no02f01 g19045 ( .a(n22833), .b(n22829), .o(n22834) );
in01f01 g19046 ( .a(n22834), .o(n22835) );
ao12f01 g19047 ( .a(n22828), .b(n22835), .c(n22767), .o(n22836) );
in01f01 g19048 ( .a(n22836), .o(n22837) );
in01f01 g19049 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_21_), .o(n22838) );
no02f01 g19050 ( .a(n22820), .b(n22819), .o(n22839) );
na02f01 g19051 ( .a(n4997_1), .b(delay_xor_ln21_unr9_stage4_stallmux_q_21_), .o(n22840) );
in01f01 g19052 ( .a(n22840), .o(n22841) );
no02f01 g19053 ( .a(n22841), .b(n22821), .o(n22842) );
in01f01 g19054 ( .a(n22842), .o(n22843) );
na02f01 g19055 ( .a(n22843), .b(n22839), .o(n22844) );
in01f01 g19056 ( .a(n22844), .o(n22845) );
no02f01 g19057 ( .a(n22843), .b(n22839), .o(n22846) );
no02f01 g19058 ( .a(n22846), .b(n22845), .o(n22847) );
in01f01 g19059 ( .a(n22847), .o(n22848) );
no02f01 g19060 ( .a(n22848), .b(n22838), .o(n22849) );
in01f01 g19061 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_18_), .o(n22850) );
no02f01 g19062 ( .a(n22813), .b(n22812), .o(n22851) );
na02f01 g19063 ( .a(n4997_1), .b(delay_xor_ln21_unr9_stage4_stallmux_q_18_), .o(n22852) );
in01f01 g19064 ( .a(n22852), .o(n22853) );
no02f01 g19065 ( .a(n22853), .b(n22814), .o(n22854) );
in01f01 g19066 ( .a(n22854), .o(n22855) );
na02f01 g19067 ( .a(n22855), .b(n22851), .o(n22856) );
in01f01 g19068 ( .a(n22856), .o(n22857) );
no02f01 g19069 ( .a(n22855), .b(n22851), .o(n22858) );
no02f01 g19070 ( .a(n22858), .b(n22857), .o(n22859) );
in01f01 g19071 ( .a(n22859), .o(n22860) );
no02f01 g19072 ( .a(n22860), .b(n22850), .o(n22861) );
in01f01 g19073 ( .a(n22861), .o(n22862) );
in01f01 g19074 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_17_), .o(n22863) );
na02f01 g19075 ( .a(n4997_1), .b(delay_xor_ln21_unr9_stage4_stallmux_q_17_), .o(n22864) );
in01f01 g19076 ( .a(n22864), .o(n22865) );
no02f01 g19077 ( .a(n22865), .b(n22813), .o(n22866) );
in01f01 g19078 ( .a(n22866), .o(n22867) );
na02f01 g19079 ( .a(n22867), .b(n22811), .o(n22868) );
in01f01 g19080 ( .a(n22868), .o(n22869) );
no02f01 g19081 ( .a(n22867), .b(n22811), .o(n22870) );
no02f01 g19082 ( .a(n22870), .b(n22869), .o(n22871) );
in01f01 g19083 ( .a(n22871), .o(n22872) );
no02f01 g19084 ( .a(n22872), .b(n22863), .o(n22873) );
in01f01 g19085 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_16_), .o(n22874) );
na02f01 g19086 ( .a(n4997_1), .b(delay_xor_ln21_unr9_stage4_stallmux_q_16_), .o(n22875) );
in01f01 g19087 ( .a(n22875), .o(n22876) );
no02f01 g19088 ( .a(n22876), .b(n22810), .o(n22877) );
in01f01 g19089 ( .a(n22877), .o(n22878) );
no02f01 g19090 ( .a(n22878), .b(n22808), .o(n22879) );
na02f01 g19091 ( .a(n22878), .b(n22808), .o(n22880) );
in01f01 g19092 ( .a(n22880), .o(n22881) );
no02f01 g19093 ( .a(n22881), .b(n22879), .o(n22882) );
in01f01 g19094 ( .a(n22882), .o(n22883) );
no02f01 g19095 ( .a(n22883), .b(n22874), .o(n22884) );
na02f01 g19096 ( .a(n4997_1), .b(delay_xor_ln21_unr9_stage4_stallmux_q_15_), .o(n22885) );
in01f01 g19097 ( .a(n22885), .o(n22886) );
no02f01 g19098 ( .a(n22886), .b(n22770), .o(n22887) );
in01f01 g19099 ( .a(n22887), .o(n22888) );
no02f01 g19100 ( .a(n22888), .b(n22806), .o(n22889) );
na02f01 g19101 ( .a(n22888), .b(n22806), .o(n22890) );
in01f01 g19102 ( .a(n22890), .o(n22891) );
no02f01 g19103 ( .a(n22891), .b(n22889), .o(n22892) );
no02f01 g19104 ( .a(n22892), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_15_), .o(n22893) );
na02f01 g19105 ( .a(n4997_1), .b(delay_xor_ln21_unr9_stage4_stallmux_q_13_), .o(n22894) );
in01f01 g19106 ( .a(n22894), .o(n22895) );
no02f01 g19107 ( .a(n22895), .b(n22802), .o(n22896) );
in01f01 g19108 ( .a(n22896), .o(n22897) );
no02f01 g19109 ( .a(n22897), .b(n22800), .o(n22898) );
no02f01 g19110 ( .a(n22896), .b(n22801), .o(n22899) );
no02f01 g19111 ( .a(n22899), .b(n22898), .o(n22900) );
na02f01 g19112 ( .a(n22900), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_13_), .o(n22901) );
in01f01 g19113 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_12_), .o(n22902) );
na02f01 g19114 ( .a(n4997_1), .b(delay_xor_ln21_unr9_stage4_stallmux_q_12_), .o(n22903) );
in01f01 g19115 ( .a(n22903), .o(n22904) );
no02f01 g19116 ( .a(n22904), .b(n22771), .o(n22905) );
in01f01 g19117 ( .a(n22905), .o(n22906) );
no02f01 g19118 ( .a(n22906), .b(n22798), .o(n22907) );
no02f01 g19119 ( .a(n22905), .b(n22799), .o(n22908) );
no03f01 g19120 ( .a(n22908), .b(n22907), .c(n22902), .o(n22909) );
na02f01 g19121 ( .a(n4997_1), .b(delay_xor_ln21_unr9_stage4_stallmux_q_11_), .o(n22910) );
in01f01 g19122 ( .a(n22910), .o(n22911) );
no02f01 g19123 ( .a(n22911), .b(n22797), .o(n22912) );
no02f01 g19124 ( .a(n22912), .b(n22796), .o(n22913) );
na02f01 g19125 ( .a(n22912), .b(n22796), .o(n22914) );
in01f01 g19126 ( .a(n22914), .o(n22915) );
no02f01 g19127 ( .a(n22915), .b(n22913), .o(n22916) );
na02f01 g19128 ( .a(n22916), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_11_), .o(n22917) );
in01f01 g19129 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_10_), .o(n22918) );
na02f01 g19130 ( .a(n4997_1), .b(delay_xor_ln21_unr9_stage4_stallmux_q_10_), .o(n22919) );
in01f01 g19131 ( .a(n22919), .o(n22920) );
no02f01 g19132 ( .a(n22920), .b(n22794), .o(n22921) );
in01f01 g19133 ( .a(n22921), .o(n22922) );
no02f01 g19134 ( .a(n22922), .b(n22792), .o(n22923) );
no02f01 g19135 ( .a(n22921), .b(n22793), .o(n22924) );
no03f01 g19136 ( .a(n22924), .b(n22923), .c(n22918), .o(n22925) );
in01f01 g19137 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_9_), .o(n22926) );
na02f01 g19138 ( .a(n4997_1), .b(delay_xor_ln21_unr9_stage4_stallmux_q_9_), .o(n22927) );
in01f01 g19139 ( .a(n22927), .o(n22928) );
no02f01 g19140 ( .a(n22928), .b(n22791), .o(n22929) );
in01f01 g19141 ( .a(n22929), .o(n22930) );
no02f01 g19142 ( .a(n22930), .b(n22789), .o(n22931) );
no02f01 g19143 ( .a(n22929), .b(n22790), .o(n22932) );
no02f01 g19144 ( .a(n22932), .b(n22931), .o(n22933) );
in01f01 g19145 ( .a(n22933), .o(n22934) );
no02f01 g19146 ( .a(n22934), .b(n22926), .o(n22935) );
in01f01 g19147 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_8_), .o(n22936) );
na02f01 g19148 ( .a(n4997_1), .b(delay_xor_ln21_unr9_stage4_stallmux_q_8_), .o(n22937) );
in01f01 g19149 ( .a(n22937), .o(n22938) );
no02f01 g19150 ( .a(n22938), .b(n22772), .o(n22939) );
in01f01 g19151 ( .a(n22939), .o(n22940) );
ao12f01 g19152 ( .a(n22940), .b(n22787), .c(n22784), .o(n22941) );
no02f01 g19153 ( .a(n22939), .b(n22788), .o(n22942) );
no02f01 g19154 ( .a(n22942), .b(n22941), .o(n22943) );
in01f01 g19155 ( .a(n22943), .o(n22944) );
no02f01 g19156 ( .a(n22944), .b(n22936), .o(n22945) );
in01f01 g19157 ( .a(n22784), .o(n22946) );
no02f01 g19158 ( .a(n22785), .b(n22946), .o(n22947) );
na02f01 g19159 ( .a(n4997_1), .b(delay_xor_ln21_unr9_stage4_stallmux_q_7_), .o(n22948) );
in01f01 g19160 ( .a(n22948), .o(n22949) );
no02f01 g19161 ( .a(n22949), .b(n22786), .o(n22950) );
in01f01 g19162 ( .a(n22950), .o(n22951) );
na02f01 g19163 ( .a(n22951), .b(n22947), .o(n22952) );
in01f01 g19164 ( .a(n22952), .o(n22953) );
no02f01 g19165 ( .a(n22951), .b(n22947), .o(n22954) );
no02f01 g19166 ( .a(n22954), .b(n22953), .o(n22955) );
no02f01 g19167 ( .a(n22955), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_7_), .o(n22956) );
in01f01 g19168 ( .a(n22956), .o(n22957) );
na02f01 g19169 ( .a(n4997_1), .b(delay_xor_ln21_unr9_stage4_stallmux_q_6_), .o(n22958) );
in01f01 g19170 ( .a(n22958), .o(n22959) );
no02f01 g19171 ( .a(n22959), .b(n22785), .o(n22960) );
in01f01 g19172 ( .a(n22960), .o(n22961) );
no02f01 g19173 ( .a(n22961), .b(n22784), .o(n22962) );
no02f01 g19174 ( .a(n22960), .b(n22946), .o(n22963) );
no02f01 g19175 ( .a(n22963), .b(n22962), .o(n22964) );
no02f01 g19176 ( .a(n22964), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_6_), .o(n22965) );
in01f01 g19177 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_5_), .o(n22966) );
na02f01 g19178 ( .a(n4997_1), .b(delay_xor_ln21_unr9_stage4_stallmux_q_5_), .o(n22967) );
in01f01 g19179 ( .a(n22967), .o(n22968) );
no02f01 g19180 ( .a(n22968), .b(n22783), .o(n22969) );
in01f01 g19181 ( .a(n22969), .o(n22970) );
no02f01 g19182 ( .a(n22970), .b(n22781), .o(n22971) );
no02f01 g19183 ( .a(n22969), .b(n22782), .o(n22972) );
no02f01 g19184 ( .a(n22972), .b(n22971), .o(n22973) );
in01f01 g19185 ( .a(n22973), .o(n22974) );
no02f01 g19186 ( .a(n22974), .b(n22966), .o(n22975) );
in01f01 g19187 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_4_), .o(n22976) );
na02f01 g19188 ( .a(n4997_1), .b(delay_xor_ln21_unr9_stage4_stallmux_q_4_), .o(n22977) );
in01f01 g19189 ( .a(n22977), .o(n22978) );
no02f01 g19190 ( .a(n22978), .b(n22778), .o(n22979) );
in01f01 g19191 ( .a(n22979), .o(n22980) );
no02f01 g19192 ( .a(n4997_1), .b(delay_xor_ln21_unr9_stage4_stallmux_q_0_), .o(n22981) );
no02f01 g19193 ( .a(n4997_1), .b(delay_xor_ln21_unr9_stage4_stallmux_q_1_), .o(n22982) );
no02f01 g19194 ( .a(n22982), .b(n22981), .o(n22983) );
in01f01 g19195 ( .a(delay_xor_ln21_unr9_stage4_stallmux_q_2_), .o(n22984) );
na02f01 g19196 ( .a(n_45224), .b(n22984), .o(n22985) );
na02f01 g19197 ( .a(n22985), .b(n22983), .o(n22986) );
no02f01 g19198 ( .a(n22986), .b(n22779), .o(n22987) );
na02f01 g19199 ( .a(n22987), .b(n22980), .o(n22988) );
no02f01 g19200 ( .a(n22987), .b(n22980), .o(n22989) );
in01f01 g19201 ( .a(n22989), .o(n22990) );
na02f01 g19202 ( .a(n22990), .b(n22988), .o(n22991) );
no02f01 g19203 ( .a(n22991), .b(n22976), .o(n22992) );
in01f01 g19204 ( .a(n22992), .o(n22993) );
na02f01 g19205 ( .a(n4997_1), .b(delay_xor_ln21_unr9_stage4_stallmux_q_3_), .o(n22994) );
in01f01 g19206 ( .a(n22994), .o(n22995) );
no02f01 g19207 ( .a(n22995), .b(n22779), .o(n22996) );
no02f01 g19208 ( .a(n22996), .b(n22986), .o(n22997) );
no02f01 g19209 ( .a(n22780), .b(n22777), .o(n22998) );
no03f01 g19210 ( .a(n22995), .b(n22998), .c(n22779), .o(n22999) );
no02f01 g19211 ( .a(n22999), .b(n22997), .o(n23000) );
no02f01 g19212 ( .a(n23000), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_3_), .o(n23001) );
in01f01 g19213 ( .a(n23001), .o(n23002) );
no02f01 g19214 ( .a(n_45224), .b(n22984), .o(n23003) );
no02f01 g19215 ( .a(n23003), .b(n22780), .o(n23004) );
no02f01 g19216 ( .a(n23004), .b(n22777), .o(n23005) );
no03f01 g19217 ( .a(n23003), .b(n22780), .c(n22983), .o(n23006) );
no02f01 g19218 ( .a(n23006), .b(n23005), .o(n23007) );
na02f01 g19219 ( .a(n23007), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_2_), .o(n23008) );
in01f01 g19220 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_1_), .o(n23009) );
no02f01 g19221 ( .a(n_45224), .b(delay_xor_ln21_unr9_stage4_stallmux_q_0_), .o(n23010) );
in01f01 g19222 ( .a(n23010), .o(n23011) );
na02f01 g19223 ( .a(n_45224), .b(delay_xor_ln21_unr9_stage4_stallmux_q_0_), .o(n23012) );
na02f01 g19224 ( .a(n23012), .b(n23011), .o(n23013) );
no02f01 g19225 ( .a(n23013), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_0_), .o(n23014) );
no02f01 g19226 ( .a(n23014), .b(n23009), .o(n23015) );
na02f01 g19227 ( .a(n23014), .b(n23009), .o(n23016) );
na02f01 g19228 ( .a(n4997_1), .b(delay_xor_ln21_unr9_stage4_stallmux_q_1_), .o(n23017) );
na02f01 g19229 ( .a(n23017), .b(n22776), .o(n23018) );
no02f01 g19230 ( .a(n23018), .b(n22774), .o(n23019) );
ao12f01 g19231 ( .a(n22981), .b(n23017), .c(n22776), .o(n23020) );
no02f01 g19232 ( .a(n23020), .b(n23019), .o(n23021) );
ao12f01 g19233 ( .a(n23015), .b(n23021), .c(n23016), .o(n23022) );
no02f01 g19234 ( .a(n23007), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_2_), .o(n23023) );
oa12f01 g19235 ( .a(n23008), .b(n23023), .c(n23022), .o(n23024) );
in01f01 g19236 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_3_), .o(n23025) );
no03f01 g19237 ( .a(n22999), .b(n22997), .c(n23025), .o(n23026) );
oa12f01 g19238 ( .a(n23002), .b(n23026), .c(n23024), .o(n23027) );
ao12f01 g19239 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_4_), .b(n22990), .c(n22988), .o(n23028) );
oa12f01 g19240 ( .a(n22993), .b(n23028), .c(n23027), .o(n23029) );
no02f01 g19241 ( .a(n22973), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_5_), .o(n23030) );
in01f01 g19242 ( .a(n23030), .o(n23031) );
ao12f01 g19243 ( .a(n22975), .b(n23031), .c(n23029), .o(n23032) );
in01f01 g19244 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_7_), .o(n23033) );
no03f01 g19245 ( .a(n22954), .b(n22953), .c(n23033), .o(n23034) );
na02f01 g19246 ( .a(n22964), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_6_), .o(n23035) );
in01f01 g19247 ( .a(n23035), .o(n23036) );
no02f01 g19248 ( .a(n23036), .b(n23034), .o(n23037) );
oa12f01 g19249 ( .a(n23037), .b(n23032), .c(n22965), .o(n23038) );
na02f01 g19250 ( .a(n23038), .b(n22957), .o(n23039) );
no02f01 g19251 ( .a(n22943), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_8_), .o(n23040) );
no02f01 g19252 ( .a(n23040), .b(n23039), .o(n23041) );
no02f01 g19253 ( .a(n23041), .b(n22945), .o(n23042) );
no02f01 g19254 ( .a(n22933), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_9_), .o(n23043) );
no02f01 g19255 ( .a(n23043), .b(n23042), .o(n23044) );
no02f01 g19256 ( .a(n23044), .b(n22935), .o(n23045) );
no02f01 g19257 ( .a(n22924), .b(n22923), .o(n23046) );
no02f01 g19258 ( .a(n23046), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_10_), .o(n23047) );
no02f01 g19259 ( .a(n23047), .b(n23045), .o(n23048) );
no02f01 g19260 ( .a(n22916), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_11_), .o(n23049) );
in01f01 g19261 ( .a(n23049), .o(n23050) );
oa12f01 g19262 ( .a(n23050), .b(n23048), .c(n22925), .o(n23051) );
no02f01 g19263 ( .a(n22908), .b(n22907), .o(n23052) );
no02f01 g19264 ( .a(n23052), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_12_), .o(n23053) );
ao12f01 g19265 ( .a(n23053), .b(n23051), .c(n22917), .o(n23054) );
no02f01 g19266 ( .a(n22900), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_13_), .o(n23055) );
in01f01 g19267 ( .a(n23055), .o(n23056) );
oa12f01 g19268 ( .a(n23056), .b(n23054), .c(n22909), .o(n23057) );
na02f01 g19269 ( .a(n23057), .b(n22901), .o(n23058) );
na02f01 g19270 ( .a(delay_xor_ln21_unr9_stage4_stallmux_q_14_), .b(n4997_1), .o(n23059) );
in01f01 g19271 ( .a(n23059), .o(n23060) );
no02f01 g19272 ( .a(n23060), .b(n22805), .o(n23061) );
no02f01 g19273 ( .a(n23061), .b(n22804), .o(n23062) );
na02f01 g19274 ( .a(n23061), .b(n22804), .o(n23063) );
in01f01 g19275 ( .a(n23063), .o(n23064) );
no02f01 g19276 ( .a(n23064), .b(n23062), .o(n23065) );
no02f01 g19277 ( .a(n23065), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_14_), .o(n23066) );
in01f01 g19278 ( .a(n23066), .o(n23067) );
in01f01 g19279 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_15_), .o(n23068) );
no03f01 g19280 ( .a(n22891), .b(n22889), .c(n23068), .o(n23069) );
na02f01 g19281 ( .a(n23065), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_14_), .o(n23070) );
in01f01 g19282 ( .a(n23070), .o(n23071) );
no02f01 g19283 ( .a(n23071), .b(n23069), .o(n23072) );
in01f01 g19284 ( .a(n23072), .o(n23073) );
ao12f01 g19285 ( .a(n23073), .b(n23067), .c(n23058), .o(n23074) );
no02f01 g19286 ( .a(n22882), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_16_), .o(n23075) );
no03f01 g19287 ( .a(n23075), .b(n23074), .c(n22893), .o(n23076) );
no02f01 g19288 ( .a(n23076), .b(n22884), .o(n23077) );
no02f01 g19289 ( .a(n22871), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_17_), .o(n23078) );
no02f01 g19290 ( .a(n23078), .b(n23077), .o(n23079) );
no02f01 g19291 ( .a(n22859), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_18_), .o(n23080) );
in01f01 g19292 ( .a(n23080), .o(n23081) );
oa12f01 g19293 ( .a(n23081), .b(n23079), .c(n22873), .o(n23082) );
na02f01 g19294 ( .a(n4997_1), .b(delay_xor_ln21_unr9_stage4_stallmux_q_19_), .o(n23083) );
in01f01 g19295 ( .a(n23083), .o(n23084) );
no02f01 g19296 ( .a(n23084), .b(n22817), .o(n23085) );
no02f01 g19297 ( .a(n23085), .b(n22816), .o(n23086) );
na02f01 g19298 ( .a(n23085), .b(n22816), .o(n23087) );
in01f01 g19299 ( .a(n23087), .o(n23088) );
no02f01 g19300 ( .a(n23088), .b(n23086), .o(n23089) );
no02f01 g19301 ( .a(n23089), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_19_), .o(n23090) );
ao12f01 g19302 ( .a(n23090), .b(n23082), .c(n22862), .o(n23091) );
na02f01 g19303 ( .a(n23089), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_19_), .o(n23092) );
in01f01 g19304 ( .a(n23092), .o(n23093) );
na02f01 g19305 ( .a(n4997_1), .b(delay_xor_ln21_unr9_stage4_stallmux_q_20_), .o(n23094) );
in01f01 g19306 ( .a(n23094), .o(n23095) );
no02f01 g19307 ( .a(n23095), .b(n22820), .o(n23096) );
in01f01 g19308 ( .a(n23096), .o(n23097) );
na02f01 g19309 ( .a(n23097), .b(n22818), .o(n23098) );
in01f01 g19310 ( .a(n23098), .o(n23099) );
no02f01 g19311 ( .a(n23097), .b(n22818), .o(n23100) );
no02f01 g19312 ( .a(n23100), .b(n23099), .o(n23101) );
no02f01 g19313 ( .a(n23101), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_20_), .o(n23102) );
in01f01 g19314 ( .a(n23102), .o(n23103) );
oa12f01 g19315 ( .a(n23103), .b(n23093), .c(n23091), .o(n23104) );
na02f01 g19316 ( .a(n23101), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_20_), .o(n23105) );
no02f01 g19317 ( .a(n22847), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_21_), .o(n23106) );
ao12f01 g19318 ( .a(n23106), .b(n23105), .c(n23104), .o(n23107) );
no02f01 g19319 ( .a(n23107), .b(n22849), .o(n23108) );
no02f01 g19320 ( .a(n22827), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_23_), .o(n23109) );
no02f01 g19321 ( .a(n22832), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_22_), .o(n23110) );
no02f01 g19322 ( .a(n23110), .b(n23109), .o(n23111) );
in01f01 g19323 ( .a(n23111), .o(n23112) );
oa12f01 g19324 ( .a(n22837), .b(n23112), .c(n23108), .o(n23113) );
no02f01 g19325 ( .a(n22827), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_24_), .o(n23114) );
no02f01 g19326 ( .a(n22827), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_25_), .o(n23115) );
no02f01 g19327 ( .a(n23115), .b(n23114), .o(n23116) );
na02f01 g19328 ( .a(n23116), .b(n23113), .o(n23117) );
no02f01 g19329 ( .a(n22827), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_26_), .o(n23118) );
no02f01 g19330 ( .a(n23118), .b(n23117), .o(n23119) );
no02f01 g19331 ( .a(n22827), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_27_), .o(n23120) );
in01f01 g19332 ( .a(n23120), .o(n23121) );
na02f01 g19333 ( .a(n23121), .b(n23119), .o(n23122) );
no02f01 g19334 ( .a(n22827), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_29_), .o(n23123) );
no02f01 g19335 ( .a(n22827), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_28_), .o(n23124) );
no02f01 g19336 ( .a(n23124), .b(n23123), .o(n23125) );
in01f01 g19337 ( .a(n23125), .o(n23126) );
no02f01 g19338 ( .a(n22827), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_30_), .o(n23127) );
no03f01 g19339 ( .a(n23127), .b(n23126), .c(n23122), .o(n23128) );
in01f01 g19340 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_27_), .o(n23129) );
in01f01 g19341 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_26_), .o(n23130) );
ao12f01 g19342 ( .a(n22828), .b(n23130), .c(n23129), .o(n23131) );
in01f01 g19343 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_24_), .o(n23132) );
in01f01 g19344 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_25_), .o(n23133) );
ao12f01 g19345 ( .a(n22828), .b(n23133), .c(n23132), .o(n23134) );
no02f01 g19346 ( .a(n23134), .b(n23131), .o(n23135) );
in01f01 g19347 ( .a(n23135), .o(n23136) );
in01f01 g19348 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_29_), .o(n23137) );
in01f01 g19349 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_28_), .o(n23138) );
ao12f01 g19350 ( .a(n22828), .b(n23138), .c(n23137), .o(n23139) );
na02f01 g19351 ( .a(n22827), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_30_), .o(n23140) );
in01f01 g19352 ( .a(n23140), .o(n23141) );
no04f01 g19353 ( .a(n23141), .b(n23139), .c(n23136), .d(n23128), .o(n23142) );
no02f01 g19354 ( .a(n22827), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_31_), .o(n23143) );
na02f01 g19355 ( .a(n22827), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_31_), .o(n23144) );
in01f01 g19356 ( .a(n23144), .o(n23145) );
no02f01 g19357 ( .a(n23145), .b(n23143), .o(n23146) );
no02f01 g19358 ( .a(n23146), .b(n23142), .o(n23147) );
na02f01 g19359 ( .a(n23146), .b(n23142), .o(n23148) );
in01f01 g19360 ( .a(n23148), .o(n23149) );
no02f01 g19361 ( .a(n23149), .b(n23147), .o(n23150) );
in01f01 g19362 ( .a(n23150), .o(n23151) );
na02f01 g19363 ( .a(n23135), .b(n23122), .o(n23152) );
oa12f01 g19364 ( .a(n23125), .b(n23152), .c(n23139), .o(n23153) );
in01f01 g19365 ( .a(n23153), .o(n23154) );
no02f01 g19366 ( .a(n23141), .b(n23127), .o(n23155) );
in01f01 g19367 ( .a(n23155), .o(n23156) );
no02f01 g19368 ( .a(n23156), .b(n23154), .o(n23157) );
no02f01 g19369 ( .a(n23155), .b(n23153), .o(n23158) );
no02f01 g19370 ( .a(n23158), .b(n23157), .o(n23159) );
no02f01 g19371 ( .a(n23159), .b(n5119), .o(n23160) );
in01f01 g19372 ( .a(n23160), .o(n23161) );
in01f01 g19373 ( .a(n23134), .o(n23162) );
na02f01 g19374 ( .a(n23162), .b(n23117), .o(n23163) );
no02f01 g19375 ( .a(n22828), .b(n23130), .o(n23164) );
no02f01 g19376 ( .a(n23164), .b(n23118), .o(n23165) );
in01f01 g19377 ( .a(n23165), .o(n23166) );
na02f01 g19378 ( .a(n23166), .b(n23163), .o(n23167) );
in01f01 g19379 ( .a(n23167), .o(n23168) );
no02f01 g19380 ( .a(n23166), .b(n23163), .o(n23169) );
no02f01 g19381 ( .a(n23169), .b(n23168), .o(n23170) );
no02f01 g19382 ( .a(n22828), .b(n23133), .o(n23171) );
no02f01 g19383 ( .a(n23171), .b(n23115), .o(n23172) );
in01f01 g19384 ( .a(n23114), .o(n23173) );
no02f01 g19385 ( .a(n22828), .b(n23132), .o(n23174) );
ao12f01 g19386 ( .a(n23174), .b(n23173), .c(n23113), .o(n23175) );
na02f01 g19387 ( .a(n23175), .b(n23172), .o(n23176) );
in01f01 g19388 ( .a(n23172), .o(n23177) );
in01f01 g19389 ( .a(n22849), .o(n23178) );
na02f01 g19390 ( .a(n23105), .b(n23104), .o(n23179) );
in01f01 g19391 ( .a(n23106), .o(n23180) );
na02f01 g19392 ( .a(n23180), .b(n23179), .o(n23181) );
na02f01 g19393 ( .a(n23181), .b(n23178), .o(n23182) );
ao12f01 g19394 ( .a(n22836), .b(n23111), .c(n23182), .o(n23183) );
no02f01 g19395 ( .a(n23114), .b(n23183), .o(n23184) );
oa12f01 g19396 ( .a(n23177), .b(n23174), .c(n23184), .o(n23185) );
na02f01 g19397 ( .a(n23185), .b(n23176), .o(n23186) );
no02f01 g19398 ( .a(n23110), .b(n22834), .o(n23187) );
na02f01 g19399 ( .a(n23187), .b(n23108), .o(n23188) );
in01f01 g19400 ( .a(n23188), .o(n23189) );
no02f01 g19401 ( .a(n23187), .b(n23108), .o(n23190) );
no02f01 g19402 ( .a(n23190), .b(n23189), .o(n23191) );
no02f01 g19403 ( .a(n23191), .b(n5142), .o(n23192) );
na02f01 g19404 ( .a(n22827), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_23_), .o(n23193) );
in01f01 g19405 ( .a(n23193), .o(n23194) );
no02f01 g19406 ( .a(n23194), .b(n23109), .o(n23195) );
no03f01 g19407 ( .a(n23107), .b(n22849), .c(n22834), .o(n23196) );
oa12f01 g19408 ( .a(n23195), .b(n23196), .c(n23110), .o(n23197) );
no03f01 g19409 ( .a(n23196), .b(n23195), .c(n23110), .o(n23198) );
in01f01 g19410 ( .a(n23198), .o(n23199) );
ao12f01 g19411 ( .a(n5142), .b(n23199), .c(n23197), .o(n23200) );
no02f01 g19412 ( .a(n23200), .b(n23192), .o(n23201) );
no02f01 g19413 ( .a(n23174), .b(n23114), .o(n23202) );
in01f01 g19414 ( .a(n23202), .o(n23203) );
na02f01 g19415 ( .a(n23203), .b(n23113), .o(n23204) );
no02f01 g19416 ( .a(n23203), .b(n23113), .o(n23205) );
in01f01 g19417 ( .a(n23205), .o(n23206) );
na02f01 g19418 ( .a(n23206), .b(n23204), .o(n23207) );
na02f01 g19419 ( .a(n23207), .b(n5119), .o(n23208) );
no02f01 g19420 ( .a(n23069), .b(n22893), .o(n23209) );
in01f01 g19421 ( .a(n23209), .o(n23210) );
na03f01 g19422 ( .a(n23070), .b(n23057), .c(n22901), .o(n23211) );
ao12f01 g19423 ( .a(n23210), .b(n23211), .c(n23067), .o(n23212) );
in01f01 g19424 ( .a(n23212), .o(n23213) );
na03f01 g19425 ( .a(n23211), .b(n23210), .c(n23067), .o(n23214) );
na02f01 g19426 ( .a(n23214), .b(n23213), .o(n23215) );
na02f01 g19427 ( .a(n23215), .b(n5119), .o(n23216) );
na02f01 g19428 ( .a(n23056), .b(n22901), .o(n23217) );
no03f01 g19429 ( .a(n23217), .b(n23054), .c(n22909), .o(n23218) );
oa12f01 g19430 ( .a(n23217), .b(n23054), .c(n22909), .o(n23219) );
in01f01 g19431 ( .a(n23219), .o(n23220) );
no02f01 g19432 ( .a(n23220), .b(n23218), .o(n23221) );
no02f01 g19433 ( .a(n23053), .b(n22909), .o(n23222) );
na03f01 g19434 ( .a(n23222), .b(n23051), .c(n22917), .o(n23223) );
ao12f01 g19435 ( .a(n23222), .b(n23051), .c(n22917), .o(n23224) );
in01f01 g19436 ( .a(n23224), .o(n23225) );
na02f01 g19437 ( .a(n23225), .b(n23223), .o(n23226) );
no02f01 g19438 ( .a(n23047), .b(n22925), .o(n23227) );
no02f01 g19439 ( .a(n23227), .b(n23045), .o(n23228) );
in01f01 g19440 ( .a(n23228), .o(n23229) );
na02f01 g19441 ( .a(n23227), .b(n23045), .o(n23230) );
na02f01 g19442 ( .a(n23230), .b(n23229), .o(n23231) );
na02f01 g19443 ( .a(n23231), .b(n5119), .o(n23232) );
na02f01 g19444 ( .a(n23050), .b(n22917), .o(n23233) );
no03f01 g19445 ( .a(n23233), .b(n23048), .c(n22925), .o(n23234) );
oa12f01 g19446 ( .a(n23233), .b(n23048), .c(n22925), .o(n23235) );
in01f01 g19447 ( .a(n23235), .o(n23236) );
no02f01 g19448 ( .a(n23236), .b(n23234), .o(n23237) );
oa12f01 g19449 ( .a(n23232), .b(n23237), .c(n5142), .o(n23238) );
ao12f01 g19450 ( .a(n23238), .b(n23226), .c(n5119), .o(n23239) );
oa12f01 g19451 ( .a(n23239), .b(n23221), .c(n5142), .o(n23240) );
no02f01 g19452 ( .a(n23071), .b(n23066), .o(n23241) );
ao12f01 g19453 ( .a(n23241), .b(n23057), .c(n22901), .o(n23242) );
in01f01 g19454 ( .a(n23242), .o(n23243) );
na03f01 g19455 ( .a(n23241), .b(n23057), .c(n22901), .o(n23244) );
na02f01 g19456 ( .a(n23244), .b(n23243), .o(n23245) );
ao12f01 g19457 ( .a(n23240), .b(n23245), .c(n5119), .o(n23246) );
na02f01 g19458 ( .a(n23246), .b(n23216), .o(n23247) );
no02f01 g19459 ( .a(n23075), .b(n22884), .o(n23248) );
no03f01 g19460 ( .a(n23248), .b(n23074), .c(n22893), .o(n23249) );
in01f01 g19461 ( .a(n23249), .o(n23250) );
oa12f01 g19462 ( .a(n23248), .b(n23074), .c(n22893), .o(n23251) );
na02f01 g19463 ( .a(n23251), .b(n23250), .o(n23252) );
ao12f01 g19464 ( .a(n23247), .b(n23252), .c(n5119), .o(n23253) );
no02f01 g19465 ( .a(n23078), .b(n22873), .o(n23254) );
na02f01 g19466 ( .a(n23254), .b(n23077), .o(n23255) );
in01f01 g19467 ( .a(n23255), .o(n23256) );
no02f01 g19468 ( .a(n23254), .b(n23077), .o(n23257) );
no02f01 g19469 ( .a(n23257), .b(n23256), .o(n23258) );
ao12f01 g19470 ( .a(n5142), .b(n23258), .c(n23253), .o(n23259) );
no02f01 g19471 ( .a(n23080), .b(n22861), .o(n23260) );
in01f01 g19472 ( .a(n23260), .o(n23261) );
no03f01 g19473 ( .a(n23261), .b(n23079), .c(n22873), .o(n23262) );
in01f01 g19474 ( .a(n23262), .o(n23263) );
oa12f01 g19475 ( .a(n23261), .b(n23079), .c(n22873), .o(n23264) );
na02f01 g19476 ( .a(n23264), .b(n23263), .o(n23265) );
ao12f01 g19477 ( .a(n23259), .b(n23265), .c(n5119), .o(n23266) );
na02f01 g19478 ( .a(n23082), .b(n22862), .o(n23267) );
no02f01 g19479 ( .a(n23093), .b(n23090), .o(n23268) );
in01f01 g19480 ( .a(n23268), .o(n23269) );
na02f01 g19481 ( .a(n23269), .b(n23267), .o(n23270) );
in01f01 g19482 ( .a(n23270), .o(n23271) );
no02f01 g19483 ( .a(n23269), .b(n23267), .o(n23272) );
no02f01 g19484 ( .a(n23272), .b(n23271), .o(n23273) );
oa12f01 g19485 ( .a(n23266), .b(n23273), .c(n5142), .o(n23274) );
no02f01 g19486 ( .a(n23093), .b(n23091), .o(n23275) );
na02f01 g19487 ( .a(n23105), .b(n23103), .o(n23276) );
in01f01 g19488 ( .a(n23276), .o(n23277) );
na02f01 g19489 ( .a(n23277), .b(n23275), .o(n23278) );
no02f01 g19490 ( .a(n23277), .b(n23275), .o(n23279) );
in01f01 g19491 ( .a(n23279), .o(n23280) );
na02f01 g19492 ( .a(n23280), .b(n23278), .o(n23281) );
ao12f01 g19493 ( .a(n23274), .b(n23281), .c(n5119), .o(n23282) );
no02f01 g19494 ( .a(n23106), .b(n22849), .o(n23283) );
in01f01 g19495 ( .a(n23283), .o(n23284) );
no02f01 g19496 ( .a(n23284), .b(n23179), .o(n23285) );
na02f01 g19497 ( .a(n23284), .b(n23179), .o(n23286) );
in01f01 g19498 ( .a(n23286), .o(n23287) );
no02f01 g19499 ( .a(n23287), .b(n23285), .o(n23288) );
oa12f01 g19500 ( .a(n23282), .b(n23288), .c(n5142), .o(n23289) );
in01f01 g19501 ( .a(n23285), .o(n23290) );
na02f01 g19502 ( .a(n23286), .b(n23290), .o(n23291) );
in01f01 g19503 ( .a(n23278), .o(n23292) );
no02f01 g19504 ( .a(n23279), .b(n23292), .o(n23293) );
in01f01 g19505 ( .a(n23272), .o(n23294) );
na02f01 g19506 ( .a(n23294), .b(n23270), .o(n23295) );
in01f01 g19507 ( .a(n23264), .o(n23296) );
no02f01 g19508 ( .a(n23296), .b(n23262), .o(n23297) );
no02f01 g19509 ( .a(n23297), .b(n5119), .o(n23298) );
ao12f01 g19510 ( .a(n23298), .b(n23295), .c(n5142), .o(n23299) );
oa12f01 g19511 ( .a(n23299), .b(n23293), .c(n5119), .o(n23300) );
ao12f01 g19512 ( .a(n23300), .b(n23291), .c(n5142), .o(n23301) );
na02f01 g19513 ( .a(n23301), .b(n23289), .o(n23302) );
na03f01 g19514 ( .a(n23302), .b(n23208), .c(n23201), .o(n23303) );
ao12f01 g19515 ( .a(n23303), .b(n23186), .c(n5119), .o(n23304) );
in01f01 g19516 ( .a(n23186), .o(n23305) );
in01f01 g19517 ( .a(n23197), .o(n23306) );
no02f01 g19518 ( .a(n23198), .b(n23306), .o(n23307) );
ao12f01 g19519 ( .a(n5119), .b(n23307), .c(n23191), .o(n23308) );
in01f01 g19520 ( .a(n23204), .o(n23309) );
no02f01 g19521 ( .a(n23205), .b(n23309), .o(n23310) );
no02f01 g19522 ( .a(n23310), .b(n5119), .o(n23311) );
no02f01 g19523 ( .a(n23311), .b(n23308), .o(n23312) );
oa12f01 g19524 ( .a(n23312), .b(n23305), .c(n5119), .o(n23313) );
oa22f01 g19525 ( .a(n23313), .b(n23304), .c(n23170), .d(n5142), .o(n23314) );
no03f01 g19526 ( .a(n23134), .b(n23164), .c(n23119), .o(n23315) );
no02f01 g19527 ( .a(n22828), .b(n23129), .o(n23316) );
no02f01 g19528 ( .a(n23316), .b(n23120), .o(n23317) );
no02f01 g19529 ( .a(n23317), .b(n23315), .o(n23318) );
na02f01 g19530 ( .a(n23317), .b(n23315), .o(n23319) );
in01f01 g19531 ( .a(n23319), .o(n23320) );
no02f01 g19532 ( .a(n23320), .b(n23318), .o(n23321) );
no02f01 g19533 ( .a(n23321), .b(n5142), .o(n23322) );
no02f01 g19534 ( .a(n22828), .b(n23138), .o(n23323) );
no02f01 g19535 ( .a(n23323), .b(n23124), .o(n23324) );
in01f01 g19536 ( .a(n23324), .o(n23325) );
na02f01 g19537 ( .a(n23325), .b(n23152), .o(n23326) );
in01f01 g19538 ( .a(n23326), .o(n23327) );
no02f01 g19539 ( .a(n23325), .b(n23152), .o(n23328) );
no02f01 g19540 ( .a(n23328), .b(n23327), .o(n23329) );
no02f01 g19541 ( .a(n23329), .b(n5142), .o(n23330) );
no03f01 g19542 ( .a(n23330), .b(n23322), .c(n23314), .o(n23331) );
no02f01 g19543 ( .a(n23321), .b(n5119), .o(n23332) );
no02f01 g19544 ( .a(n23170), .b(n5119), .o(n23333) );
no02f01 g19545 ( .a(n23333), .b(n23332), .o(n23334) );
oa12f01 g19546 ( .a(n23334), .b(n23329), .c(n5119), .o(n23335) );
no02f01 g19547 ( .a(n23335), .b(n23331), .o(n23336) );
no02f01 g19548 ( .a(n22828), .b(n23137), .o(n23337) );
no02f01 g19549 ( .a(n23337), .b(n23123), .o(n23338) );
no02f01 g19550 ( .a(n23323), .b(n23136), .o(n23339) );
oa12f01 g19551 ( .a(n23339), .b(n23124), .c(n23122), .o(n23340) );
in01f01 g19552 ( .a(n23340), .o(n23341) );
no02f01 g19553 ( .a(n23341), .b(n23338), .o(n23342) );
na02f01 g19554 ( .a(n23341), .b(n23338), .o(n23343) );
in01f01 g19555 ( .a(n23343), .o(n23344) );
no02f01 g19556 ( .a(n23344), .b(n23342), .o(n23345) );
no02f01 g19557 ( .a(n23345), .b(n5119), .o(n23346) );
in01f01 g19558 ( .a(n23346), .o(n23347) );
na02f01 g19559 ( .a(n23347), .b(n23336), .o(n23348) );
no02f01 g19560 ( .a(n23345), .b(n5142), .o(n23349) );
in01f01 g19561 ( .a(n23349), .o(n23350) );
no02f01 g19562 ( .a(n23159), .b(n5142), .o(n23351) );
in01f01 g19563 ( .a(n23351), .o(n23352) );
na03f01 g19564 ( .a(n23352), .b(n23350), .c(n23348), .o(n23353) );
ao22f01 g19565 ( .a(n23353), .b(n23161), .c(n23151), .d(n5119), .o(n23354) );
no02f01 g19566 ( .a(n23150), .b(n5119), .o(n23355) );
no03f01 g19567 ( .a(n23355), .b(n23354), .c(n23151), .o(n23356) );
na02f01 g19568 ( .a(n23353), .b(n23161), .o(n23357) );
no02f01 g19569 ( .a(n23150), .b(n5119), .o(n23359) );
no02f01 g19570 ( .a(n23359), .b(n23356), .o(n23360) );
in01f01 g19571 ( .a(delay_xor_ln22_unr9_stage4_stallmux_q_22_), .o(n23361) );
no02f01 g19572 ( .a(n_45224), .b(n23361), .o(n23362) );
in01f01 g19573 ( .a(delay_xor_ln22_unr9_stage4_stallmux_q_2_), .o(n23363) );
na02f01 g19574 ( .a(n_45224), .b(n23363), .o(n23364) );
in01f01 g19575 ( .a(n_45622), .o(n23365) );
in01f01 g19576 ( .a(n_45209), .o(n23366) );
oa12f01 g19577 ( .a(n_45224), .b(n23366), .c(n23365), .o(n23367) );
na02f01 g19578 ( .a(n23367), .b(n23364), .o(n23368) );
in01f01 g19579 ( .a(delay_xor_ln22_unr9_stage4_stallmux_q_3_), .o(n23369) );
na02f01 g19580 ( .a(n_45224), .b(n23369), .o(n23370) );
no02f01 g19581 ( .a(n4997_1), .b(delay_xor_ln22_unr9_stage4_stallmux_q_4_), .o(n23371) );
in01f01 g19582 ( .a(n23371), .o(n23372) );
na02f01 g19583 ( .a(n23372), .b(n23370), .o(n23373) );
no02f01 g19584 ( .a(n23373), .b(n23368), .o(n23374) );
no02f01 g19585 ( .a(n4997_1), .b(delay_xor_ln22_unr9_stage4_stallmux_q_7_), .o(n23375) );
no02f01 g19586 ( .a(n4997_1), .b(delay_xor_ln22_unr9_stage4_stallmux_q_5_), .o(n23376) );
no02f01 g19587 ( .a(delay_xor_ln22_unr9_stage4_stallmux_q_6_), .b(n4997_1), .o(n23377) );
no03f01 g19588 ( .a(n23377), .b(n23376), .c(n23375), .o(n23378) );
na02f01 g19589 ( .a(n23378), .b(n23374), .o(n23379) );
no02f01 g19590 ( .a(delay_xor_ln22_unr9_stage4_stallmux_q_8_), .b(n4997_1), .o(n23380) );
no02f01 g19591 ( .a(n23380), .b(n23379), .o(n23381) );
in01f01 g19592 ( .a(n23381), .o(n23382) );
no02f01 g19593 ( .a(n4997_1), .b(delay_xor_ln22_unr9_stage4_stallmux_q_9_), .o(n23383) );
no02f01 g19594 ( .a(n23383), .b(n23382), .o(n23384) );
no02f01 g19595 ( .a(n4997_1), .b(delay_xor_ln22_unr9_stage4_stallmux_q_11_), .o(n23385) );
no02f01 g19596 ( .a(n4997_1), .b(delay_xor_ln22_unr9_stage4_stallmux_q_12_), .o(n23386) );
no02f01 g19597 ( .a(n4997_1), .b(delay_xor_ln22_unr9_stage4_stallmux_q_10_), .o(n23387) );
no03f01 g19598 ( .a(n23387), .b(n23386), .c(n23385), .o(n23388) );
na02f01 g19599 ( .a(n23388), .b(n23384), .o(n23389) );
in01f01 g19600 ( .a(n23389), .o(n23390) );
no02f01 g19601 ( .a(n4997_1), .b(delay_xor_ln22_unr9_stage4_stallmux_q_13_), .o(n23391) );
no02f01 g19602 ( .a(n4997_1), .b(delay_xor_ln22_unr9_stage4_stallmux_q_14_), .o(n23392) );
no02f01 g19603 ( .a(n23392), .b(n23391), .o(n23393) );
na02f01 g19604 ( .a(n23393), .b(n23390), .o(n23394) );
no02f01 g19605 ( .a(n4997_1), .b(delay_xor_ln22_unr9_stage4_stallmux_q_15_), .o(n23395) );
no02f01 g19606 ( .a(n23395), .b(n23394), .o(n23396) );
in01f01 g19607 ( .a(n23396), .o(n23397) );
no02f01 g19608 ( .a(n4997_1), .b(delay_xor_ln22_unr9_stage4_stallmux_q_16_), .o(n23398) );
no02f01 g19609 ( .a(n23398), .b(n23397), .o(n23399) );
in01f01 g19610 ( .a(n23399), .o(n23400) );
no02f01 g19611 ( .a(n4997_1), .b(delay_xor_ln22_unr9_stage4_stallmux_q_17_), .o(n23401) );
no02f01 g19612 ( .a(n23401), .b(n23400), .o(n23402) );
in01f01 g19613 ( .a(n23402), .o(n23403) );
no02f01 g19614 ( .a(n4997_1), .b(delay_xor_ln22_unr9_stage4_stallmux_q_18_), .o(n23404) );
no02f01 g19615 ( .a(n23404), .b(n23403), .o(n23405) );
in01f01 g19616 ( .a(n23405), .o(n23406) );
no02f01 g19617 ( .a(n4997_1), .b(delay_xor_ln22_unr9_stage4_stallmux_q_19_), .o(n23407) );
no02f01 g19618 ( .a(n23407), .b(n23406), .o(n23408) );
in01f01 g19619 ( .a(n23408), .o(n23409) );
no02f01 g19620 ( .a(n4997_1), .b(delay_xor_ln22_unr9_stage4_stallmux_q_20_), .o(n23410) );
no02f01 g19621 ( .a(n23410), .b(n23409), .o(n23411) );
in01f01 g19622 ( .a(n23411), .o(n23412) );
no02f01 g19623 ( .a(n4997_1), .b(delay_xor_ln22_unr9_stage4_stallmux_q_21_), .o(n23413) );
no02f01 g19624 ( .a(n23413), .b(n23412), .o(n23414) );
no02f01 g19625 ( .a(n4997_1), .b(delay_xor_ln22_unr9_stage4_stallmux_q_22_), .o(n23415) );
no02f01 g19626 ( .a(n23415), .b(n23362), .o(n23416) );
in01f01 g19627 ( .a(n23416), .o(n23417) );
no02f01 g19628 ( .a(n23417), .b(n23414), .o(n23418) );
no02f01 g19629 ( .a(n23418), .b(n23362), .o(n23419) );
in01f01 g19630 ( .a(n23419), .o(n23420) );
no02f01 g19631 ( .a(n23420), .b(delay_add_ln22_unr8_stage4_stallmux_q_31_), .o(n23421) );
na02f01 g19632 ( .a(n23420), .b(delay_add_ln22_unr8_stage4_stallmux_q_31_), .o(n23422) );
in01f01 g19633 ( .a(n23422), .o(n23423) );
no02f01 g19634 ( .a(n23423), .b(n23421), .o(n23424) );
in01f01 g19635 ( .a(n23424), .o(n23425) );
in01f01 g19636 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_21_), .o(n23426) );
na02f01 g19637 ( .a(n4997_1), .b(delay_xor_ln22_unr9_stage4_stallmux_q_21_), .o(n23427) );
in01f01 g19638 ( .a(n23427), .o(n23428) );
no02f01 g19639 ( .a(n23428), .b(n23413), .o(n23429) );
no02f01 g19640 ( .a(n23429), .b(n23412), .o(n23430) );
na02f01 g19641 ( .a(n23429), .b(n23412), .o(n23431) );
in01f01 g19642 ( .a(n23431), .o(n23432) );
no02f01 g19643 ( .a(n23432), .b(n23430), .o(n23433) );
no02f01 g19644 ( .a(n23433), .b(n23426), .o(n23434) );
in01f01 g19645 ( .a(n23434), .o(n23435) );
in01f01 g19646 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_20_), .o(n23436) );
na02f01 g19647 ( .a(n4997_1), .b(delay_xor_ln22_unr9_stage4_stallmux_q_20_), .o(n23437) );
in01f01 g19648 ( .a(n23437), .o(n23438) );
no02f01 g19649 ( .a(n23438), .b(n23410), .o(n23439) );
no02f01 g19650 ( .a(n23439), .b(n23409), .o(n23440) );
na02f01 g19651 ( .a(n23439), .b(n23409), .o(n23441) );
in01f01 g19652 ( .a(n23441), .o(n23442) );
no02f01 g19653 ( .a(n23442), .b(n23440), .o(n23443) );
no02f01 g19654 ( .a(n23443), .b(n23436), .o(n23444) );
in01f01 g19655 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_19_), .o(n23445) );
na02f01 g19656 ( .a(n4997_1), .b(delay_xor_ln22_unr9_stage4_stallmux_q_19_), .o(n23446) );
in01f01 g19657 ( .a(n23446), .o(n23447) );
no02f01 g19658 ( .a(n23447), .b(n23407), .o(n23448) );
no02f01 g19659 ( .a(n23448), .b(n23406), .o(n23449) );
na02f01 g19660 ( .a(n23448), .b(n23406), .o(n23450) );
in01f01 g19661 ( .a(n23450), .o(n23451) );
no02f01 g19662 ( .a(n23451), .b(n23449), .o(n23452) );
no02f01 g19663 ( .a(n23452), .b(n23445), .o(n23453) );
in01f01 g19664 ( .a(n23453), .o(n23454) );
in01f01 g19665 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_17_), .o(n23455) );
na02f01 g19666 ( .a(n4997_1), .b(delay_xor_ln22_unr9_stage4_stallmux_q_17_), .o(n23456) );
in01f01 g19667 ( .a(n23456), .o(n23457) );
no02f01 g19668 ( .a(n23457), .b(n23401), .o(n23458) );
in01f01 g19669 ( .a(n23458), .o(n23459) );
no02f01 g19670 ( .a(n23459), .b(n23399), .o(n23460) );
no02f01 g19671 ( .a(n23458), .b(n23400), .o(n23461) );
no02f01 g19672 ( .a(n23461), .b(n23460), .o(n23462) );
no02f01 g19673 ( .a(n23462), .b(n23455), .o(n23463) );
in01f01 g19674 ( .a(n23463), .o(n23464) );
na02f01 g19675 ( .a(n23462), .b(n23455), .o(n23465) );
in01f01 g19676 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_16_), .o(n23466) );
na02f01 g19677 ( .a(n4997_1), .b(delay_xor_ln22_unr9_stage4_stallmux_q_16_), .o(n23467) );
in01f01 g19678 ( .a(n23467), .o(n23468) );
no02f01 g19679 ( .a(n23468), .b(n23398), .o(n23469) );
no02f01 g19680 ( .a(n23469), .b(n23397), .o(n23470) );
na02f01 g19681 ( .a(n23469), .b(n23397), .o(n23471) );
in01f01 g19682 ( .a(n23471), .o(n23472) );
no02f01 g19683 ( .a(n23472), .b(n23470), .o(n23473) );
no02f01 g19684 ( .a(n23473), .b(n23466), .o(n23474) );
in01f01 g19685 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_15_), .o(n23475) );
na02f01 g19686 ( .a(n4997_1), .b(delay_xor_ln22_unr9_stage4_stallmux_q_15_), .o(n23476) );
in01f01 g19687 ( .a(n23476), .o(n23477) );
no02f01 g19688 ( .a(n23477), .b(n23395), .o(n23478) );
in01f01 g19689 ( .a(n23478), .o(n23479) );
ao12f01 g19690 ( .a(n23479), .b(n23393), .c(n23390), .o(n23480) );
no02f01 g19691 ( .a(n23478), .b(n23394), .o(n23481) );
no02f01 g19692 ( .a(n23481), .b(n23480), .o(n23482) );
no02f01 g19693 ( .a(n23482), .b(n23475), .o(n23483) );
in01f01 g19694 ( .a(n23483), .o(n23484) );
in01f01 g19695 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_14_), .o(n23485) );
na02f01 g19696 ( .a(n4997_1), .b(delay_xor_ln22_unr9_stage4_stallmux_q_14_), .o(n23486) );
in01f01 g19697 ( .a(n23486), .o(n23487) );
no02f01 g19698 ( .a(n23487), .b(n23392), .o(n23488) );
no02f01 g19699 ( .a(n23488), .b(n23391), .o(n23489) );
no02f01 g19700 ( .a(n23391), .b(n23389), .o(n23490) );
in01f01 g19701 ( .a(n23490), .o(n23491) );
ao22f01 g19702 ( .a(n23491), .b(n23488), .c(n23489), .d(n23390), .o(n23492) );
no02f01 g19703 ( .a(n23492), .b(n23485), .o(n23493) );
in01f01 g19704 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_13_), .o(n23494) );
na02f01 g19705 ( .a(n4997_1), .b(delay_xor_ln22_unr9_stage4_stallmux_q_13_), .o(n23495) );
in01f01 g19706 ( .a(n23495), .o(n23496) );
no02f01 g19707 ( .a(n23496), .b(n23391), .o(n23497) );
in01f01 g19708 ( .a(n23497), .o(n23498) );
no02f01 g19709 ( .a(n23498), .b(n23390), .o(n23499) );
no02f01 g19710 ( .a(n23497), .b(n23389), .o(n23500) );
no02f01 g19711 ( .a(n23500), .b(n23499), .o(n23501) );
no02f01 g19712 ( .a(n23501), .b(n23494), .o(n23502) );
in01f01 g19713 ( .a(n23502), .o(n23503) );
in01f01 g19714 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_12_), .o(n23504) );
in01f01 g19715 ( .a(n23384), .o(n23505) );
no02f01 g19716 ( .a(n23387), .b(n23505), .o(n23506) );
in01f01 g19717 ( .a(n23506), .o(n23507) );
no02f01 g19718 ( .a(n23507), .b(n23385), .o(n23508) );
in01f01 g19719 ( .a(n23508), .o(n23509) );
na02f01 g19720 ( .a(n4997_1), .b(delay_xor_ln22_unr9_stage4_stallmux_q_12_), .o(n23510) );
in01f01 g19721 ( .a(n23510), .o(n23511) );
no02f01 g19722 ( .a(n23511), .b(n23386), .o(n23512) );
no02f01 g19723 ( .a(n23512), .b(n23509), .o(n23513) );
na02f01 g19724 ( .a(n23512), .b(n23509), .o(n23514) );
in01f01 g19725 ( .a(n23514), .o(n23515) );
no02f01 g19726 ( .a(n23515), .b(n23513), .o(n23516) );
no02f01 g19727 ( .a(n23516), .b(n23504), .o(n23517) );
in01f01 g19728 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_11_), .o(n23518) );
na02f01 g19729 ( .a(n4997_1), .b(delay_xor_ln22_unr9_stage4_stallmux_q_11_), .o(n23519) );
in01f01 g19730 ( .a(n23519), .o(n23520) );
no02f01 g19731 ( .a(n23520), .b(n23385), .o(n23521) );
no02f01 g19732 ( .a(n23521), .b(n23507), .o(n23522) );
na02f01 g19733 ( .a(n23521), .b(n23507), .o(n23523) );
in01f01 g19734 ( .a(n23523), .o(n23524) );
no02f01 g19735 ( .a(n23524), .b(n23522), .o(n23525) );
no02f01 g19736 ( .a(n23525), .b(n23518), .o(n23526) );
in01f01 g19737 ( .a(n23526), .o(n23527) );
in01f01 g19738 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_10_), .o(n23528) );
na02f01 g19739 ( .a(n4997_1), .b(delay_xor_ln22_unr9_stage4_stallmux_q_10_), .o(n23529) );
in01f01 g19740 ( .a(n23529), .o(n23530) );
no02f01 g19741 ( .a(n23530), .b(n23387), .o(n23531) );
in01f01 g19742 ( .a(n23531), .o(n23532) );
no02f01 g19743 ( .a(n23532), .b(n23384), .o(n23533) );
no02f01 g19744 ( .a(n23531), .b(n23505), .o(n23534) );
no02f01 g19745 ( .a(n23534), .b(n23533), .o(n23535) );
no02f01 g19746 ( .a(n23535), .b(n23528), .o(n23536) );
in01f01 g19747 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_9_), .o(n23537) );
na02f01 g19748 ( .a(n4997_1), .b(delay_xor_ln22_unr9_stage4_stallmux_q_9_), .o(n23538) );
in01f01 g19749 ( .a(n23538), .o(n23539) );
no02f01 g19750 ( .a(n23539), .b(n23383), .o(n23540) );
no02f01 g19751 ( .a(n23540), .b(n23382), .o(n23541) );
na02f01 g19752 ( .a(n23540), .b(n23382), .o(n23542) );
in01f01 g19753 ( .a(n23542), .o(n23543) );
no02f01 g19754 ( .a(n23543), .b(n23541), .o(n23544) );
no02f01 g19755 ( .a(n23544), .b(n23537), .o(n23545) );
in01f01 g19756 ( .a(n23545), .o(n23546) );
in01f01 g19757 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_8_), .o(n23547) );
na02f01 g19758 ( .a(delay_xor_ln22_unr9_stage4_stallmux_q_8_), .b(n4997_1), .o(n23548) );
in01f01 g19759 ( .a(n23548), .o(n23549) );
no02f01 g19760 ( .a(n23549), .b(n23380), .o(n23550) );
in01f01 g19761 ( .a(n23550), .o(n23551) );
ao12f01 g19762 ( .a(n23551), .b(n23378), .c(n23374), .o(n23552) );
no02f01 g19763 ( .a(n23550), .b(n23379), .o(n23553) );
no02f01 g19764 ( .a(n23553), .b(n23552), .o(n23554) );
no02f01 g19765 ( .a(n23554), .b(n23547), .o(n23555) );
in01f01 g19766 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_7_), .o(n23556) );
na02f01 g19767 ( .a(n4997_1), .b(delay_xor_ln22_unr9_stage4_stallmux_q_7_), .o(n23557) );
in01f01 g19768 ( .a(n23557), .o(n23558) );
no02f01 g19769 ( .a(n23558), .b(n23375), .o(n23559) );
in01f01 g19770 ( .a(n23559), .o(n23560) );
no03f01 g19771 ( .a(n23376), .b(n23373), .c(n23368), .o(n23561) );
in01f01 g19772 ( .a(n23561), .o(n23562) );
no02f01 g19773 ( .a(n23562), .b(n23377), .o(n23563) );
na02f01 g19774 ( .a(n23563), .b(n23560), .o(n23564) );
in01f01 g19775 ( .a(n23564), .o(n23565) );
no02f01 g19776 ( .a(n23563), .b(n23560), .o(n23566) );
no02f01 g19777 ( .a(n23566), .b(n23565), .o(n23567) );
no02f01 g19778 ( .a(n23567), .b(n23556), .o(n23568) );
in01f01 g19779 ( .a(n23568), .o(n23569) );
in01f01 g19780 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_6_), .o(n23570) );
na02f01 g19781 ( .a(delay_xor_ln22_unr9_stage4_stallmux_q_6_), .b(n4997_1), .o(n23571) );
in01f01 g19782 ( .a(n23571), .o(n23572) );
no02f01 g19783 ( .a(n23572), .b(n23377), .o(n23573) );
in01f01 g19784 ( .a(n23573), .o(n23574) );
no02f01 g19785 ( .a(n23574), .b(n23561), .o(n23575) );
na02f01 g19786 ( .a(n23574), .b(n23561), .o(n23576) );
in01f01 g19787 ( .a(n23576), .o(n23577) );
no02f01 g19788 ( .a(n23577), .b(n23575), .o(n23578) );
no02f01 g19789 ( .a(n23578), .b(n23570), .o(n23579) );
in01f01 g19790 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_5_), .o(n23580) );
na02f01 g19791 ( .a(n4997_1), .b(delay_xor_ln22_unr9_stage4_stallmux_q_5_), .o(n23581) );
in01f01 g19792 ( .a(n23581), .o(n23582) );
no02f01 g19793 ( .a(n23582), .b(n23376), .o(n23583) );
in01f01 g19794 ( .a(n23583), .o(n23584) );
no02f01 g19795 ( .a(n23584), .b(n23374), .o(n23585) );
no03f01 g19796 ( .a(n23583), .b(n23373), .c(n23368), .o(n23586) );
no02f01 g19797 ( .a(n23586), .b(n23585), .o(n23587) );
no02f01 g19798 ( .a(n23587), .b(n23580), .o(n23588) );
in01f01 g19799 ( .a(n23588), .o(n23589) );
in01f01 g19800 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_4_), .o(n23590) );
na02f01 g19801 ( .a(n4997_1), .b(delay_xor_ln22_unr9_stage4_stallmux_q_4_), .o(n23591) );
na02f01 g19802 ( .a(n23591), .b(n23372), .o(n23592) );
in01f01 g19803 ( .a(n23592), .o(n23593) );
no02f01 g19804 ( .a(n4997_1), .b(delay_xor_ln22_unr9_stage4_stallmux_q_2_), .o(n23594) );
ao12f01 g19805 ( .a(n4997_1), .b(n_45209), .c(n_45622), .o(n23595) );
no02f01 g19806 ( .a(n23595), .b(n23594), .o(n23596) );
na02f01 g19807 ( .a(n23370), .b(n23596), .o(n23597) );
no02f01 g19808 ( .a(n23597), .b(n23593), .o(n23598) );
in01f01 g19809 ( .a(n23597), .o(n23599) );
no02f01 g19810 ( .a(n23599), .b(n23592), .o(n23600) );
no02f01 g19811 ( .a(n23600), .b(n23598), .o(n23601) );
no02f01 g19812 ( .a(n23601), .b(n23590), .o(n23602) );
in01f01 g19813 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_3_), .o(n23603) );
na02f01 g19814 ( .a(n4997_1), .b(delay_xor_ln22_unr9_stage4_stallmux_q_3_), .o(n23604) );
na02f01 g19815 ( .a(n23604), .b(n23370), .o(n23605) );
no02f01 g19816 ( .a(n23605), .b(n23596), .o(n23606) );
no02f01 g19817 ( .a(n4997_1), .b(delay_xor_ln22_unr9_stage4_stallmux_q_3_), .o(n23607) );
no02f01 g19818 ( .a(n_45224), .b(n23369), .o(n23608) );
no02f01 g19819 ( .a(n23608), .b(n23607), .o(n23609) );
no02f01 g19820 ( .a(n23609), .b(n23368), .o(n23610) );
no02f01 g19821 ( .a(n23610), .b(n23606), .o(n23611) );
no02f01 g19822 ( .a(n23611), .b(n23603), .o(n23612) );
in01f01 g19823 ( .a(n23612), .o(n23613) );
in01f01 g19824 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_2_), .o(n23614) );
no02f01 g19825 ( .a(n_45224), .b(n23363), .o(n23615) );
oa12f01 g19826 ( .a(n23367), .b(n23615), .c(n23594), .o(n23616) );
na02f01 g19827 ( .a(n4997_1), .b(delay_xor_ln22_unr9_stage4_stallmux_q_2_), .o(n23617) );
na03f01 g19828 ( .a(n23617), .b(n23595), .c(n23364), .o(n23618) );
ao12f01 g19829 ( .a(n23614), .b(n23618), .c(n23616), .o(n23619) );
in01f01 g19830 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_0_), .o(n23620) );
no02f01 g19831 ( .a(n_45209), .b(n_45224), .o(n23621) );
na02f01 g19832 ( .a(n_45209), .b(n_45224), .o(n23622) );
in01f01 g19833 ( .a(n23622), .o(n23623) );
no03f01 g19834 ( .a(n23623), .b(n23621), .c(n23620), .o(n23624) );
na02f01 g19835 ( .a(n23624), .b(delay_add_ln22_unr8_stage4_stallmux_q_1_), .o(n23625) );
no03f01 g19836 ( .a(n_45209), .b(n4997_1), .c(n23365), .o(n23626) );
na02f01 g19837 ( .a(n_45224), .b(n23365), .o(n23627) );
na02f01 g19838 ( .a(n4997_1), .b(n_45622), .o(n23628) );
ao22f01 g19839 ( .a(n23628), .b(n23627), .c(n23366), .d(n_45224), .o(n23629) );
oa22f01 g19840 ( .a(n23629), .b(n23626), .c(n23624), .d(delay_add_ln22_unr8_stage4_stallmux_q_1_), .o(n23630) );
ao12f01 g19841 ( .a(n23595), .b(n23617), .c(n23364), .o(n23631) );
no03f01 g19842 ( .a(n23615), .b(n23367), .c(n23594), .o(n23632) );
no03f01 g19843 ( .a(n23632), .b(n23631), .c(delay_add_ln22_unr8_stage4_stallmux_q_2_), .o(n23633) );
ao12f01 g19844 ( .a(n23633), .b(n23630), .c(n23625), .o(n23634) );
no03f01 g19845 ( .a(n23610), .b(n23606), .c(delay_add_ln22_unr8_stage4_stallmux_q_3_), .o(n23635) );
in01f01 g19846 ( .a(n23635), .o(n23636) );
oa12f01 g19847 ( .a(n23636), .b(n23634), .c(n23619), .o(n23637) );
no03f01 g19848 ( .a(n23600), .b(n23598), .c(delay_add_ln22_unr8_stage4_stallmux_q_4_), .o(n23638) );
ao12f01 g19849 ( .a(n23638), .b(n23637), .c(n23613), .o(n23639) );
na02f01 g19850 ( .a(n23587), .b(n23580), .o(n23640) );
oa12f01 g19851 ( .a(n23640), .b(n23639), .c(n23602), .o(n23641) );
no03f01 g19852 ( .a(n23577), .b(n23575), .c(delay_add_ln22_unr8_stage4_stallmux_q_6_), .o(n23642) );
ao12f01 g19853 ( .a(n23642), .b(n23641), .c(n23589), .o(n23643) );
no03f01 g19854 ( .a(n23566), .b(n23565), .c(delay_add_ln22_unr8_stage4_stallmux_q_7_), .o(n23644) );
in01f01 g19855 ( .a(n23644), .o(n23645) );
oa12f01 g19856 ( .a(n23645), .b(n23643), .c(n23579), .o(n23646) );
na02f01 g19857 ( .a(n23554), .b(n23547), .o(n23647) );
in01f01 g19858 ( .a(n23647), .o(n23648) );
ao12f01 g19859 ( .a(n23648), .b(n23646), .c(n23569), .o(n23649) );
na02f01 g19860 ( .a(n23544), .b(n23537), .o(n23650) );
oa12f01 g19861 ( .a(n23650), .b(n23649), .c(n23555), .o(n23651) );
na02f01 g19862 ( .a(n23535), .b(n23528), .o(n23652) );
in01f01 g19863 ( .a(n23652), .o(n23653) );
ao12f01 g19864 ( .a(n23653), .b(n23651), .c(n23546), .o(n23654) );
na02f01 g19865 ( .a(n23525), .b(n23518), .o(n23655) );
oa12f01 g19866 ( .a(n23655), .b(n23654), .c(n23536), .o(n23656) );
na02f01 g19867 ( .a(n23516), .b(n23504), .o(n23657) );
in01f01 g19868 ( .a(n23657), .o(n23658) );
ao12f01 g19869 ( .a(n23658), .b(n23656), .c(n23527), .o(n23659) );
na02f01 g19870 ( .a(n23501), .b(n23494), .o(n23660) );
oa12f01 g19871 ( .a(n23660), .b(n23659), .c(n23517), .o(n23661) );
na02f01 g19872 ( .a(n23492), .b(n23485), .o(n23662) );
in01f01 g19873 ( .a(n23662), .o(n23663) );
ao12f01 g19874 ( .a(n23663), .b(n23661), .c(n23503), .o(n23664) );
na02f01 g19875 ( .a(n23482), .b(n23475), .o(n23665) );
oa12f01 g19876 ( .a(n23665), .b(n23664), .c(n23493), .o(n23666) );
na02f01 g19877 ( .a(n23473), .b(n23466), .o(n23667) );
in01f01 g19878 ( .a(n23667), .o(n23668) );
ao12f01 g19879 ( .a(n23668), .b(n23666), .c(n23484), .o(n23669) );
oa12f01 g19880 ( .a(n23465), .b(n23669), .c(n23474), .o(n23670) );
na02f01 g19881 ( .a(n4997_1), .b(delay_xor_ln22_unr9_stage4_stallmux_q_18_), .o(n23671) );
in01f01 g19882 ( .a(n23671), .o(n23672) );
no02f01 g19883 ( .a(n23672), .b(n23404), .o(n23673) );
no02f01 g19884 ( .a(n23673), .b(n23403), .o(n23674) );
na02f01 g19885 ( .a(n23673), .b(n23403), .o(n23675) );
in01f01 g19886 ( .a(n23675), .o(n23676) );
no02f01 g19887 ( .a(n23676), .b(n23674), .o(n23677) );
in01f01 g19888 ( .a(n23677), .o(n23678) );
no02f01 g19889 ( .a(n23678), .b(delay_add_ln22_unr8_stage4_stallmux_q_18_), .o(n23679) );
ao12f01 g19890 ( .a(n23679), .b(n23670), .c(n23464), .o(n23680) );
na02f01 g19891 ( .a(n23678), .b(delay_add_ln22_unr8_stage4_stallmux_q_18_), .o(n23681) );
in01f01 g19892 ( .a(n23681), .o(n23682) );
na02f01 g19893 ( .a(n23452), .b(n23445), .o(n23683) );
oa12f01 g19894 ( .a(n23683), .b(n23682), .c(n23680), .o(n23684) );
na02f01 g19895 ( .a(n23443), .b(n23436), .o(n23685) );
in01f01 g19896 ( .a(n23685), .o(n23686) );
ao12f01 g19897 ( .a(n23686), .b(n23684), .c(n23454), .o(n23687) );
na02f01 g19898 ( .a(n23433), .b(n23426), .o(n23688) );
oa12f01 g19899 ( .a(n23688), .b(n23687), .c(n23444), .o(n23689) );
in01f01 g19900 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_22_), .o(n23690) );
na02f01 g19901 ( .a(n23417), .b(n23414), .o(n23691) );
in01f01 g19902 ( .a(n23691), .o(n23692) );
no02f01 g19903 ( .a(n23692), .b(n23418), .o(n23693) );
no02f01 g19904 ( .a(n23693), .b(n23690), .o(n23694) );
in01f01 g19905 ( .a(n23694), .o(n23695) );
in01f01 g19906 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_23_), .o(n23696) );
no02f01 g19907 ( .a(n23419), .b(n23696), .o(n23697) );
in01f01 g19908 ( .a(n23697), .o(n23698) );
na04f01 g19909 ( .a(n23698), .b(n23695), .c(n23689), .d(n23435), .o(n23699) );
no02f01 g19910 ( .a(n23420), .b(delay_add_ln22_unr8_stage4_stallmux_q_23_), .o(n23700) );
na02f01 g19911 ( .a(n23693), .b(n23690), .o(n23701) );
in01f01 g19912 ( .a(n23701), .o(n23702) );
no02f01 g19913 ( .a(n23702), .b(n23700), .o(n23703) );
na02f01 g19914 ( .a(n23703), .b(n23699), .o(n23704) );
no02f01 g19915 ( .a(n23420), .b(delay_add_ln22_unr8_stage4_stallmux_q_26_), .o(n23705) );
ao12f01 g19916 ( .a(n23420), .b(delay_add_ln22_unr8_stage4_stallmux_q_24_), .c(delay_add_ln22_unr8_stage4_stallmux_q_25_), .o(n23706) );
no02f01 g19917 ( .a(n23706), .b(n23705), .o(n23707) );
in01f01 g19918 ( .a(n23707), .o(n23708) );
no02f01 g19919 ( .a(n23708), .b(n23704), .o(n23709) );
no02f01 g19920 ( .a(n23420), .b(delay_add_ln22_unr8_stage4_stallmux_q_27_), .o(n23710) );
in01f01 g19921 ( .a(n23710), .o(n23711) );
na02f01 g19922 ( .a(n23711), .b(n23709), .o(n23712) );
no02f01 g19923 ( .a(n23420), .b(delay_add_ln22_unr8_stage4_stallmux_q_28_), .o(n23713) );
no02f01 g19924 ( .a(n23713), .b(n23712), .o(n23714) );
no02f01 g19925 ( .a(n23420), .b(delay_add_ln22_unr8_stage4_stallmux_q_29_), .o(n23715) );
in01f01 g19926 ( .a(n23715), .o(n23716) );
na02f01 g19927 ( .a(n23716), .b(n23714), .o(n23717) );
no02f01 g19928 ( .a(n23420), .b(delay_add_ln22_unr8_stage4_stallmux_q_30_), .o(n23718) );
in01f01 g19929 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_26_), .o(n23719) );
in01f01 g19930 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_27_), .o(n23720) );
ao12f01 g19931 ( .a(n23419), .b(n23720), .c(n23719), .o(n23721) );
in01f01 g19932 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_25_), .o(n23722) );
in01f01 g19933 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_24_), .o(n23723) );
ao12f01 g19934 ( .a(n23419), .b(n23723), .c(n23722), .o(n23724) );
no02f01 g19935 ( .a(n23724), .b(n23721), .o(n23725) );
in01f01 g19936 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_28_), .o(n23726) );
no02f01 g19937 ( .a(n23419), .b(n23726), .o(n23727) );
in01f01 g19938 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_29_), .o(n23728) );
no02f01 g19939 ( .a(n23419), .b(n23728), .o(n23729) );
no02f01 g19940 ( .a(n23729), .b(n23727), .o(n23730) );
na02f01 g19941 ( .a(n23730), .b(n23725), .o(n23731) );
na02f01 g19942 ( .a(n23420), .b(delay_add_ln22_unr8_stage4_stallmux_q_30_), .o(n23732) );
in01f01 g19943 ( .a(n23732), .o(n23733) );
no02f01 g19944 ( .a(n23733), .b(n23731), .o(n23734) );
oa12f01 g19945 ( .a(n23734), .b(n23718), .c(n23717), .o(n23735) );
no02f01 g19946 ( .a(n23735), .b(n23425), .o(n23736) );
na02f01 g19947 ( .a(n23735), .b(n23425), .o(n23737) );
in01f01 g19948 ( .a(n23737), .o(n23738) );
no02f01 g19949 ( .a(n23738), .b(n23736), .o(n23739) );
no02f01 g19950 ( .a(n23739), .b(n23360), .o(n23740) );
in01f01 g19951 ( .a(n23360), .o(n23741) );
in01f01 g19952 ( .a(n23739), .o(n23742) );
no02f01 g19953 ( .a(n23742), .b(n23741), .o(n23743) );
no02f01 g19954 ( .a(n23743), .b(n23740), .o(n23744) );
na03f01 g19955 ( .a(n23695), .b(n23689), .c(n23435), .o(n23745) );
no02f01 g19956 ( .a(n23700), .b(n23697), .o(n23746) );
in01f01 g19957 ( .a(n23746), .o(n23747) );
na03f01 g19958 ( .a(n23747), .b(n23701), .c(n23745), .o(n23748) );
in01f01 g19959 ( .a(n23444), .o(n23749) );
in01f01 g19960 ( .a(n23465), .o(n23750) );
in01f01 g19961 ( .a(n23474), .o(n23751) );
in01f01 g19962 ( .a(n23493), .o(n23752) );
in01f01 g19963 ( .a(n23517), .o(n23753) );
in01f01 g19964 ( .a(n23536), .o(n23754) );
in01f01 g19965 ( .a(n23555), .o(n23755) );
in01f01 g19966 ( .a(n23579), .o(n23756) );
in01f01 g19967 ( .a(n23602), .o(n23757) );
in01f01 g19968 ( .a(n23619), .o(n23758) );
in01f01 g19969 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_1_), .o(n23759) );
in01f01 g19970 ( .a(n23621), .o(n23760) );
na03f01 g19971 ( .a(n23622), .b(n23760), .c(delay_add_ln22_unr8_stage4_stallmux_q_0_), .o(n23761) );
no02f01 g19972 ( .a(n23761), .b(n23759), .o(n23762) );
in01f01 g19973 ( .a(n23626), .o(n23763) );
no02f01 g19974 ( .a(n4997_1), .b(n_45622), .o(n23764) );
no02f01 g19975 ( .a(n_45224), .b(n23365), .o(n23765) );
oa22f01 g19976 ( .a(n23765), .b(n23764), .c(n_45209), .d(n4997_1), .o(n23766) );
ao22f01 g19977 ( .a(n23766), .b(n23763), .c(n23761), .d(n23759), .o(n23767) );
na03f01 g19978 ( .a(n23618), .b(n23616), .c(n23614), .o(n23768) );
oa12f01 g19979 ( .a(n23768), .b(n23767), .c(n23762), .o(n23769) );
ao12f01 g19980 ( .a(n23635), .b(n23769), .c(n23758), .o(n23770) );
in01f01 g19981 ( .a(n23638), .o(n23771) );
oa12f01 g19982 ( .a(n23771), .b(n23770), .c(n23612), .o(n23772) );
in01f01 g19983 ( .a(n23640), .o(n23773) );
ao12f01 g19984 ( .a(n23773), .b(n23772), .c(n23757), .o(n23774) );
in01f01 g19985 ( .a(n23642), .o(n23775) );
oa12f01 g19986 ( .a(n23775), .b(n23774), .c(n23588), .o(n23776) );
ao12f01 g19987 ( .a(n23644), .b(n23776), .c(n23756), .o(n23777) );
oa12f01 g19988 ( .a(n23647), .b(n23777), .c(n23568), .o(n23778) );
in01f01 g19989 ( .a(n23650), .o(n23779) );
ao12f01 g19990 ( .a(n23779), .b(n23778), .c(n23755), .o(n23780) );
oa12f01 g19991 ( .a(n23652), .b(n23780), .c(n23545), .o(n23781) );
in01f01 g19992 ( .a(n23655), .o(n23782) );
ao12f01 g19993 ( .a(n23782), .b(n23781), .c(n23754), .o(n23783) );
oa12f01 g19994 ( .a(n23657), .b(n23783), .c(n23526), .o(n23784) );
in01f01 g19995 ( .a(n23660), .o(n23785) );
ao12f01 g19996 ( .a(n23785), .b(n23784), .c(n23753), .o(n23786) );
oa12f01 g19997 ( .a(n23662), .b(n23786), .c(n23502), .o(n23787) );
in01f01 g19998 ( .a(n23665), .o(n23788) );
ao12f01 g19999 ( .a(n23788), .b(n23787), .c(n23752), .o(n23789) );
oa12f01 g20000 ( .a(n23667), .b(n23789), .c(n23483), .o(n23790) );
ao12f01 g20001 ( .a(n23750), .b(n23790), .c(n23751), .o(n23791) );
in01f01 g20002 ( .a(n23679), .o(n23792) );
oa12f01 g20003 ( .a(n23792), .b(n23791), .c(n23463), .o(n23793) );
in01f01 g20004 ( .a(n23683), .o(n23794) );
ao12f01 g20005 ( .a(n23794), .b(n23681), .c(n23793), .o(n23795) );
oa12f01 g20006 ( .a(n23685), .b(n23795), .c(n23453), .o(n23796) );
in01f01 g20007 ( .a(n23688), .o(n23797) );
ao12f01 g20008 ( .a(n23797), .b(n23796), .c(n23749), .o(n23798) );
no03f01 g20009 ( .a(n23694), .b(n23798), .c(n23434), .o(n23799) );
oa12f01 g20010 ( .a(n23746), .b(n23702), .c(n23799), .o(n23800) );
na02f01 g20011 ( .a(n23800), .b(n23748), .o(n23801) );
no02f01 g20012 ( .a(n23797), .b(n23434), .o(n23802) );
na03f01 g20013 ( .a(n23802), .b(n23796), .c(n23749), .o(n23803) );
in01f01 g20014 ( .a(n23802), .o(n23804) );
oa12f01 g20015 ( .a(n23804), .b(n23687), .c(n23444), .o(n23805) );
na02f01 g20016 ( .a(n23805), .b(n23803), .o(n23806) );
na02f01 g20017 ( .a(n23357), .b(n23151), .o(n23807) );
in01f01 g20018 ( .a(n23807), .o(n23808) );
no02f01 g20019 ( .a(n23357), .b(n23151), .o(n23809) );
oa12f01 g20020 ( .a(n23806), .b(n23809), .c(n23808), .o(n23810) );
no03f01 g20021 ( .a(n23804), .b(n23687), .c(n23444), .o(n23811) );
ao12f01 g20022 ( .a(n23802), .b(n23796), .c(n23749), .o(n23812) );
no02f01 g20023 ( .a(n23812), .b(n23811), .o(n23813) );
in01f01 g20024 ( .a(n23809), .o(n23814) );
na03f01 g20025 ( .a(n23814), .b(n23807), .c(n23813), .o(n23815) );
no02f01 g20026 ( .a(n23686), .b(n23444), .o(n23816) );
in01f01 g20027 ( .a(n23816), .o(n23817) );
no03f01 g20028 ( .a(n23817), .b(n23795), .c(n23453), .o(n23818) );
ao12f01 g20029 ( .a(n23816), .b(n23684), .c(n23454), .o(n23819) );
no02f01 g20030 ( .a(n23819), .b(n23818), .o(n23820) );
na02f01 g20031 ( .a(n23350), .b(n23348), .o(n23821) );
no02f01 g20032 ( .a(n23351), .b(n23160), .o(n23822) );
no02f01 g20033 ( .a(n23822), .b(n23821), .o(n23823) );
in01f01 g20034 ( .a(n23823), .o(n23824) );
na02f01 g20035 ( .a(n23822), .b(n23821), .o(n23825) );
ao12f01 g20036 ( .a(n23820), .b(n23825), .c(n23824), .o(n23826) );
no02f01 g20037 ( .a(n23794), .b(n23453), .o(n23827) );
in01f01 g20038 ( .a(n23827), .o(n23828) );
na03f01 g20039 ( .a(n23681), .b(n23670), .c(n23464), .o(n23829) );
na03f01 g20040 ( .a(n23829), .b(n23828), .c(n23792), .o(n23830) );
no03f01 g20041 ( .a(n23682), .b(n23791), .c(n23463), .o(n23831) );
oa12f01 g20042 ( .a(n23827), .b(n23831), .c(n23679), .o(n23832) );
na02f01 g20043 ( .a(n23832), .b(n23830), .o(n23833) );
no02f01 g20044 ( .a(n23349), .b(n23346), .o(n23834) );
na02f01 g20045 ( .a(n23834), .b(n23336), .o(n23835) );
in01f01 g20046 ( .a(n23835), .o(n23836) );
no02f01 g20047 ( .a(n23834), .b(n23336), .o(n23837) );
oa12f01 g20048 ( .a(n23833), .b(n23837), .c(n23836), .o(n23838) );
no02f01 g20049 ( .a(n23322), .b(n23314), .o(n23839) );
in01f01 g20050 ( .a(n23334), .o(n23840) );
no02f01 g20051 ( .a(n23840), .b(n23839), .o(n23841) );
no02f01 g20052 ( .a(n23841), .b(n23329), .o(n23842) );
in01f01 g20053 ( .a(n23329), .o(n23843) );
no03f01 g20054 ( .a(n23840), .b(n23843), .c(n23839), .o(n23844) );
no02f01 g20055 ( .a(n23682), .b(n23679), .o(n23845) );
na03f01 g20056 ( .a(n23845), .b(n23670), .c(n23464), .o(n23846) );
in01f01 g20057 ( .a(n23845), .o(n23847) );
oa12f01 g20058 ( .a(n23847), .b(n23791), .c(n23463), .o(n23848) );
na02f01 g20059 ( .a(n23848), .b(n23846), .o(n23849) );
oa12f01 g20060 ( .a(n23849), .b(n23844), .c(n23842), .o(n23850) );
in01f01 g20061 ( .a(n23850), .o(n23851) );
in01f01 g20062 ( .a(n23170), .o(n23852) );
na02f01 g20063 ( .a(n23186), .b(n5119), .o(n23853) );
na04f01 g20064 ( .a(n23302), .b(n23208), .c(n23201), .d(n23853), .o(n23854) );
in01f01 g20065 ( .a(n23312), .o(n23855) );
ao12f01 g20066 ( .a(n23855), .b(n23186), .c(n5142), .o(n23856) );
ao22f01 g20067 ( .a(n23856), .b(n23854), .c(n23852), .d(n5119), .o(n23857) );
in01f01 g20068 ( .a(n23318), .o(n23858) );
na02f01 g20069 ( .a(n23319), .b(n23858), .o(n23859) );
na02f01 g20070 ( .a(n23859), .b(n5119), .o(n23860) );
na02f01 g20071 ( .a(n23859), .b(n5142), .o(n23861) );
na02f01 g20072 ( .a(n23861), .b(n23860), .o(n23862) );
no03f01 g20073 ( .a(n23862), .b(n23333), .c(n23857), .o(n23863) );
in01f01 g20074 ( .a(n23333), .o(n23864) );
no02f01 g20075 ( .a(n23332), .b(n23322), .o(n23865) );
ao12f01 g20076 ( .a(n23865), .b(n23864), .c(n23314), .o(n23866) );
no02f01 g20077 ( .a(n23750), .b(n23463), .o(n23867) );
na03f01 g20078 ( .a(n23867), .b(n23790), .c(n23751), .o(n23868) );
in01f01 g20079 ( .a(n23867), .o(n23869) );
oa12f01 g20080 ( .a(n23869), .b(n23669), .c(n23474), .o(n23870) );
na02f01 g20081 ( .a(n23870), .b(n23868), .o(n23871) );
oa12f01 g20082 ( .a(n23871), .b(n23866), .c(n23863), .o(n23872) );
no03f01 g20083 ( .a(n23313), .b(n23304), .c(n23852), .o(n23873) );
in01f01 g20084 ( .a(n23873), .o(n23874) );
oa12f01 g20085 ( .a(n23852), .b(n23313), .c(n23304), .o(n23875) );
no02f01 g20086 ( .a(n23668), .b(n23474), .o(n23876) );
in01f01 g20087 ( .a(n23876), .o(n23877) );
no03f01 g20088 ( .a(n23877), .b(n23789), .c(n23483), .o(n23878) );
ao12f01 g20089 ( .a(n23876), .b(n23666), .c(n23484), .o(n23879) );
no02f01 g20090 ( .a(n23879), .b(n23878), .o(n23880) );
ao12f01 g20091 ( .a(n23880), .b(n23875), .c(n23874), .o(n23881) );
in01f01 g20092 ( .a(n23208), .o(n23882) );
in01f01 g20093 ( .a(n23298), .o(n23883) );
oa12f01 g20094 ( .a(n23883), .b(n23273), .c(n5119), .o(n23884) );
ao12f01 g20095 ( .a(n23884), .b(n23281), .c(n5142), .o(n23885) );
oa12f01 g20096 ( .a(n23885), .b(n23288), .c(n5119), .o(n23886) );
no03f01 g20097 ( .a(n23289), .b(n23200), .c(n23192), .o(n23887) );
no04f01 g20098 ( .a(n23887), .b(n23311), .c(n23308), .d(n23886), .o(n23888) );
no03f01 g20099 ( .a(n23888), .b(n23882), .c(n23305), .o(n23889) );
in01f01 g20100 ( .a(n23190), .o(n23890) );
na02f01 g20101 ( .a(n23890), .b(n23188), .o(n23891) );
na02f01 g20102 ( .a(n23199), .b(n23197), .o(n23892) );
oa12f01 g20103 ( .a(n5142), .b(n23892), .c(n23891), .o(n23893) );
na02f01 g20104 ( .a(n23207), .b(n5142), .o(n23894) );
na02f01 g20105 ( .a(n23891), .b(n5119), .o(n23895) );
oa12f01 g20106 ( .a(n5119), .b(n23198), .c(n23306), .o(n23896) );
in01f01 g20107 ( .a(n23214), .o(n23897) );
no02f01 g20108 ( .a(n23897), .b(n23212), .o(n23898) );
no02f01 g20109 ( .a(n23898), .b(n5142), .o(n23899) );
in01f01 g20110 ( .a(n23218), .o(n23900) );
na02f01 g20111 ( .a(n23219), .b(n23900), .o(n23901) );
in01f01 g20112 ( .a(n23223), .o(n23902) );
no02f01 g20113 ( .a(n23224), .b(n23902), .o(n23903) );
in01f01 g20114 ( .a(n23230), .o(n23904) );
no02f01 g20115 ( .a(n23904), .b(n23228), .o(n23905) );
no02f01 g20116 ( .a(n23905), .b(n5142), .o(n23906) );
in01f01 g20117 ( .a(n23234), .o(n23907) );
na02f01 g20118 ( .a(n23235), .b(n23907), .o(n23908) );
ao12f01 g20119 ( .a(n23906), .b(n23908), .c(n5119), .o(n23909) );
oa12f01 g20120 ( .a(n23909), .b(n23903), .c(n5142), .o(n23910) );
ao12f01 g20121 ( .a(n23910), .b(n23901), .c(n5119), .o(n23911) );
in01f01 g20122 ( .a(n23244), .o(n23912) );
no02f01 g20123 ( .a(n23912), .b(n23242), .o(n23913) );
oa12f01 g20124 ( .a(n23911), .b(n23913), .c(n5142), .o(n23914) );
no02f01 g20125 ( .a(n23914), .b(n23899), .o(n23915) );
in01f01 g20126 ( .a(n23251), .o(n23916) );
no02f01 g20127 ( .a(n23916), .b(n23249), .o(n23917) );
oa12f01 g20128 ( .a(n23915), .b(n23917), .c(n5142), .o(n23918) );
in01f01 g20129 ( .a(n23257), .o(n23919) );
na02f01 g20130 ( .a(n23919), .b(n23255), .o(n23920) );
oa12f01 g20131 ( .a(n5119), .b(n23920), .c(n23918), .o(n23921) );
oa12f01 g20132 ( .a(n23921), .b(n23297), .c(n5142), .o(n23922) );
ao12f01 g20133 ( .a(n23922), .b(n23295), .c(n5119), .o(n23923) );
oa12f01 g20134 ( .a(n23923), .b(n23293), .c(n5142), .o(n23924) );
ao12f01 g20135 ( .a(n23924), .b(n23291), .c(n5119), .o(n23925) );
na03f01 g20136 ( .a(n23925), .b(n23896), .c(n23895), .o(n23926) );
na04f01 g20137 ( .a(n23926), .b(n23894), .c(n23893), .d(n23301), .o(n23927) );
ao12f01 g20138 ( .a(n23186), .b(n23927), .c(n23208), .o(n23928) );
no02f01 g20139 ( .a(n23788), .b(n23483), .o(n23929) );
in01f01 g20140 ( .a(n23929), .o(n23930) );
oa12f01 g20141 ( .a(n23930), .b(n23664), .c(n23493), .o(n23931) );
na03f01 g20142 ( .a(n23929), .b(n23787), .c(n23752), .o(n23932) );
na02f01 g20143 ( .a(n23932), .b(n23931), .o(n23933) );
no03f01 g20144 ( .a(n23933), .b(n23928), .c(n23889), .o(n23934) );
na03f01 g20145 ( .a(n23927), .b(n23208), .c(n23186), .o(n23935) );
oa12f01 g20146 ( .a(n23305), .b(n23888), .c(n23882), .o(n23936) );
ao12f01 g20147 ( .a(n23929), .b(n23787), .c(n23752), .o(n23937) );
no03f01 g20148 ( .a(n23930), .b(n23664), .c(n23493), .o(n23938) );
no02f01 g20149 ( .a(n23938), .b(n23937), .o(n23939) );
ao12f01 g20150 ( .a(n23939), .b(n23936), .c(n23935), .o(n23940) );
no02f01 g20151 ( .a(n23663), .b(n23493), .o(n23941) );
ao12f01 g20152 ( .a(n23941), .b(n23661), .c(n23503), .o(n23942) );
in01f01 g20153 ( .a(n23941), .o(n23943) );
no03f01 g20154 ( .a(n23943), .b(n23786), .c(n23502), .o(n23944) );
no02f01 g20155 ( .a(n23944), .b(n23942), .o(n23945) );
no02f01 g20156 ( .a(n23308), .b(n23886), .o(n23946) );
na03f01 g20157 ( .a(n23946), .b(n23926), .c(n23310), .o(n23947) );
na02f01 g20158 ( .a(n23893), .b(n23301), .o(n23948) );
oa12f01 g20159 ( .a(n23207), .b(n23948), .c(n23887), .o(n23949) );
ao12f01 g20160 ( .a(n23945), .b(n23949), .c(n23947), .o(n23950) );
oa12f01 g20161 ( .a(n23943), .b(n23786), .c(n23502), .o(n23951) );
na03f01 g20162 ( .a(n23941), .b(n23661), .c(n23503), .o(n23952) );
na02f01 g20163 ( .a(n23952), .b(n23951), .o(n23953) );
no03f01 g20164 ( .a(n23948), .b(n23887), .c(n23207), .o(n23954) );
ao12f01 g20165 ( .a(n23310), .b(n23946), .c(n23926), .o(n23955) );
no03f01 g20166 ( .a(n23955), .b(n23954), .c(n23953), .o(n23956) );
no02f01 g20167 ( .a(n23785), .b(n23502), .o(n23957) );
na03f01 g20168 ( .a(n23957), .b(n23784), .c(n23753), .o(n23958) );
in01f01 g20169 ( .a(n23957), .o(n23959) );
oa12f01 g20170 ( .a(n23959), .b(n23659), .c(n23517), .o(n23960) );
na02f01 g20171 ( .a(n23960), .b(n23958), .o(n23961) );
no02f01 g20172 ( .a(n23191), .b(n5119), .o(n23962) );
ao22f01 g20173 ( .a(n23301), .b(n23289), .c(n23891), .d(n5119), .o(n23963) );
no03f01 g20174 ( .a(n23963), .b(n23962), .c(n23892), .o(n23964) );
na02f01 g20175 ( .a(n23891), .b(n5142), .o(n23965) );
oa22f01 g20176 ( .a(n23886), .b(n23925), .c(n23191), .d(n5142), .o(n23966) );
ao12f01 g20177 ( .a(n23307), .b(n23966), .c(n23965), .o(n23967) );
oa12f01 g20178 ( .a(n23961), .b(n23967), .c(n23964), .o(n23968) );
oa12f01 g20179 ( .a(n23891), .b(n23886), .c(n23925), .o(n23969) );
na03f01 g20180 ( .a(n23301), .b(n23289), .c(n23191), .o(n23970) );
no02f01 g20181 ( .a(n23658), .b(n23517), .o(n23971) );
ao12f01 g20182 ( .a(n23971), .b(n23656), .c(n23527), .o(n23972) );
in01f01 g20183 ( .a(n23971), .o(n23973) );
no03f01 g20184 ( .a(n23973), .b(n23783), .c(n23526), .o(n23974) );
no02f01 g20185 ( .a(n23974), .b(n23972), .o(n23975) );
ao12f01 g20186 ( .a(n23975), .b(n23970), .c(n23969), .o(n23976) );
na02f01 g20187 ( .a(n23885), .b(n23924), .o(n23977) );
na02f01 g20188 ( .a(n23977), .b(n23291), .o(n23978) );
no02f01 g20189 ( .a(n23300), .b(n23282), .o(n23979) );
na02f01 g20190 ( .a(n23979), .b(n23288), .o(n23980) );
na02f01 g20191 ( .a(n23980), .b(n23978), .o(n23981) );
no03f01 g20192 ( .a(n23884), .b(n23281), .c(n23923), .o(n23982) );
ao12f01 g20193 ( .a(n23293), .b(n23299), .c(n23274), .o(n23983) );
na02f01 g20194 ( .a(n23651), .b(n23546), .o(n23984) );
no02f01 g20195 ( .a(n23653), .b(n23536), .o(n23985) );
in01f01 g20196 ( .a(n23985), .o(n23986) );
na02f01 g20197 ( .a(n23986), .b(n23984), .o(n23987) );
no02f01 g20198 ( .a(n23780), .b(n23545), .o(n23988) );
na02f01 g20199 ( .a(n23985), .b(n23988), .o(n23989) );
na02f01 g20200 ( .a(n23989), .b(n23987), .o(n23990) );
no03f01 g20201 ( .a(n23990), .b(n23983), .c(n23982), .o(n23991) );
na02f01 g20202 ( .a(n23883), .b(n23922), .o(n23992) );
na02f01 g20203 ( .a(n23992), .b(n23295), .o(n23993) );
no02f01 g20204 ( .a(n23298), .b(n23266), .o(n23994) );
na02f01 g20205 ( .a(n23994), .b(n23273), .o(n23995) );
na02f01 g20206 ( .a(n23995), .b(n23993), .o(n23996) );
na02f01 g20207 ( .a(n23297), .b(n23259), .o(n23997) );
na02f01 g20208 ( .a(n23265), .b(n23921), .o(n23998) );
na02f01 g20209 ( .a(n23998), .b(n23997), .o(n23999) );
na02f01 g20210 ( .a(n23646), .b(n23569), .o(n24000) );
no02f01 g20211 ( .a(n23648), .b(n23555), .o(n24001) );
in01f01 g20212 ( .a(n24001), .o(n24002) );
no02f01 g20213 ( .a(n24002), .b(n24000), .o(n24003) );
na02f01 g20214 ( .a(n24002), .b(n24000), .o(n24004) );
in01f01 g20215 ( .a(n24004), .o(n24005) );
no02f01 g20216 ( .a(n24005), .b(n24003), .o(n24006) );
in01f01 g20217 ( .a(n24006), .o(n24007) );
no02f01 g20218 ( .a(n23258), .b(n23918), .o(n24008) );
no02f01 g20219 ( .a(n23920), .b(n23253), .o(n24009) );
no02f01 g20220 ( .a(n24009), .b(n24008), .o(n24010) );
no02f01 g20221 ( .a(n23246), .b(n23215), .o(n24011) );
no02f01 g20222 ( .a(n23914), .b(n23898), .o(n24012) );
na02f01 g20223 ( .a(n23772), .b(n23757), .o(n24013) );
no02f01 g20224 ( .a(n23773), .b(n23588), .o(n24014) );
in01f01 g20225 ( .a(n24014), .o(n24015) );
no02f01 g20226 ( .a(n24015), .b(n24013), .o(n24016) );
na02f01 g20227 ( .a(n24015), .b(n24013), .o(n24017) );
in01f01 g20228 ( .a(n24017), .o(n24018) );
no02f01 g20229 ( .a(n24018), .b(n24016), .o(n24019) );
in01f01 g20230 ( .a(n24019), .o(n24020) );
no03f01 g20231 ( .a(n24020), .b(n24012), .c(n24011), .o(n24021) );
na02f01 g20232 ( .a(n23245), .b(n23911), .o(n24022) );
na02f01 g20233 ( .a(n23913), .b(n23240), .o(n24023) );
na02f01 g20234 ( .a(n23637), .b(n23613), .o(n24024) );
no02f01 g20235 ( .a(n23638), .b(n23602), .o(n24025) );
in01f01 g20236 ( .a(n24025), .o(n24026) );
no02f01 g20237 ( .a(n24026), .b(n24024), .o(n24027) );
na02f01 g20238 ( .a(n24026), .b(n24024), .o(n24028) );
in01f01 g20239 ( .a(n24028), .o(n24029) );
no02f01 g20240 ( .a(n24029), .b(n24027), .o(n24030) );
ao12f01 g20241 ( .a(n24030), .b(n24023), .c(n24022), .o(n24031) );
no02f01 g20242 ( .a(n23239), .b(n23901), .o(n24032) );
no02f01 g20243 ( .a(n23910), .b(n23221), .o(n24033) );
na02f01 g20244 ( .a(n23769), .b(n23758), .o(n24034) );
no02f01 g20245 ( .a(n23635), .b(n23612), .o(n24035) );
in01f01 g20246 ( .a(n24035), .o(n24036) );
no02f01 g20247 ( .a(n24036), .b(n24034), .o(n24037) );
na02f01 g20248 ( .a(n24036), .b(n24034), .o(n24038) );
in01f01 g20249 ( .a(n24038), .o(n24039) );
no02f01 g20250 ( .a(n24039), .b(n24037), .o(n24040) );
in01f01 g20251 ( .a(n24040), .o(n24041) );
oa12f01 g20252 ( .a(n24041), .b(n24033), .c(n24032), .o(n24042) );
na02f01 g20253 ( .a(n23909), .b(n23226), .o(n24043) );
na02f01 g20254 ( .a(n23238), .b(n23903), .o(n24044) );
na02f01 g20255 ( .a(n23630), .b(n23625), .o(n24045) );
no02f01 g20256 ( .a(n23633), .b(n23619), .o(n24046) );
in01f01 g20257 ( .a(n24046), .o(n24047) );
no02f01 g20258 ( .a(n24047), .b(n24045), .o(n24048) );
na02f01 g20259 ( .a(n24047), .b(n24045), .o(n24049) );
in01f01 g20260 ( .a(n24049), .o(n24050) );
no02f01 g20261 ( .a(n24050), .b(n24048), .o(n24051) );
na03f01 g20262 ( .a(n24051), .b(n24044), .c(n24043), .o(n24052) );
na02f01 g20263 ( .a(n23237), .b(n23906), .o(n24053) );
na02f01 g20264 ( .a(n23908), .b(n23232), .o(n24054) );
na02f01 g20265 ( .a(n24054), .b(n24053), .o(n24055) );
no03f01 g20266 ( .a(n23623), .b(n23621), .c(delay_add_ln22_unr8_stage4_stallmux_q_0_), .o(n24056) );
ao12f01 g20267 ( .a(n23620), .b(n23622), .c(n23760), .o(n24057) );
no02f01 g20268 ( .a(n24057), .b(n24056), .o(n24058) );
no02f01 g20269 ( .a(n24058), .b(n23905), .o(n24059) );
in01f01 g20270 ( .a(n24059), .o(n24060) );
no03f01 g20271 ( .a(n23629), .b(n23626), .c(delay_add_ln22_unr8_stage4_stallmux_q_1_), .o(n24061) );
ao12f01 g20272 ( .a(n23759), .b(n23766), .c(n23763), .o(n24062) );
no03f01 g20273 ( .a(n24062), .b(n24061), .c(n23624), .o(n24063) );
no02f01 g20274 ( .a(n24062), .b(n24061), .o(n24064) );
no02f01 g20275 ( .a(n24064), .b(n23761), .o(n24065) );
no02f01 g20276 ( .a(n24065), .b(n24063), .o(n24066) );
na02f01 g20277 ( .a(n24066), .b(n24060), .o(n24067) );
na02f01 g20278 ( .a(n24067), .b(n24055), .o(n24068) );
no02f01 g20279 ( .a(n24066), .b(n24060), .o(n24069) );
in01f01 g20280 ( .a(n24069), .o(n24070) );
na02f01 g20281 ( .a(n24070), .b(n24068), .o(n24071) );
ao12f01 g20282 ( .a(n24051), .b(n24044), .c(n24043), .o(n24072) );
ao12f01 g20283 ( .a(n24072), .b(n24071), .c(n24052), .o(n24073) );
no03f01 g20284 ( .a(n24041), .b(n24033), .c(n24032), .o(n24074) );
oa12f01 g20285 ( .a(n24042), .b(n24074), .c(n24073), .o(n24075) );
na03f01 g20286 ( .a(n24030), .b(n24023), .c(n24022), .o(n24076) );
ao12f01 g20287 ( .a(n24031), .b(n24076), .c(n24075), .o(n24077) );
oa12f01 g20288 ( .a(n24020), .b(n24012), .c(n24011), .o(n24078) );
oa12f01 g20289 ( .a(n24078), .b(n24077), .c(n24021), .o(n24079) );
na03f01 g20290 ( .a(n23252), .b(n23246), .c(n23216), .o(n24080) );
oa12f01 g20291 ( .a(n23917), .b(n23914), .c(n23899), .o(n24081) );
no02f01 g20292 ( .a(n23774), .b(n23588), .o(n24082) );
no02f01 g20293 ( .a(n23642), .b(n23579), .o(n24083) );
no02f01 g20294 ( .a(n24083), .b(n24082), .o(n24084) );
na02f01 g20295 ( .a(n24083), .b(n24082), .o(n24085) );
in01f01 g20296 ( .a(n24085), .o(n24086) );
no02f01 g20297 ( .a(n24086), .b(n24084), .o(n24087) );
na03f01 g20298 ( .a(n24087), .b(n24081), .c(n24080), .o(n24088) );
na02f01 g20299 ( .a(n24088), .b(n24079), .o(n24089) );
ao12f01 g20300 ( .a(n24087), .b(n24081), .c(n24080), .o(n24090) );
na02f01 g20301 ( .a(n23776), .b(n23756), .o(n24091) );
no02f01 g20302 ( .a(n23644), .b(n23568), .o(n24092) );
in01f01 g20303 ( .a(n24092), .o(n24093) );
no02f01 g20304 ( .a(n24093), .b(n24091), .o(n24094) );
na02f01 g20305 ( .a(n24093), .b(n24091), .o(n24095) );
in01f01 g20306 ( .a(n24095), .o(n24096) );
no02f01 g20307 ( .a(n24096), .b(n24094), .o(n24097) );
in01f01 g20308 ( .a(n24097), .o(n24098) );
no02f01 g20309 ( .a(n24098), .b(n24090), .o(n24099) );
ao12f01 g20310 ( .a(n24010), .b(n24099), .c(n24089), .o(n24100) );
no03f01 g20311 ( .a(n23917), .b(n23914), .c(n23899), .o(n24101) );
ao12f01 g20312 ( .a(n23252), .b(n23246), .c(n23216), .o(n24102) );
in01f01 g20313 ( .a(n24087), .o(n24103) );
oa12f01 g20314 ( .a(n24103), .b(n24102), .c(n24101), .o(n24104) );
ao12f01 g20315 ( .a(n24097), .b(n24104), .c(n24089), .o(n24105) );
oa22f01 g20316 ( .a(n24105), .b(n24100), .c(n24007), .d(n23999), .o(n24106) );
ao12f01 g20317 ( .a(n24006), .b(n23998), .c(n23997), .o(n24107) );
in01f01 g20318 ( .a(n24107), .o(n24108) );
no02f01 g20319 ( .a(n23649), .b(n23555), .o(n24109) );
no02f01 g20320 ( .a(n23779), .b(n23545), .o(n24110) );
no02f01 g20321 ( .a(n24110), .b(n24109), .o(n24111) );
na02f01 g20322 ( .a(n24110), .b(n24109), .o(n24112) );
in01f01 g20323 ( .a(n24112), .o(n24113) );
no02f01 g20324 ( .a(n24113), .b(n24111), .o(n24114) );
na03f01 g20325 ( .a(n24114), .b(n24108), .c(n24106), .o(n24115) );
ao12f01 g20326 ( .a(n24114), .b(n24108), .c(n24106), .o(n24116) );
ao12f01 g20327 ( .a(n24116), .b(n24115), .c(n23996), .o(n24117) );
oa12f01 g20328 ( .a(n23990), .b(n23983), .c(n23982), .o(n24118) );
oa12f01 g20329 ( .a(n24118), .b(n24117), .c(n23991), .o(n24119) );
no02f01 g20330 ( .a(n23782), .b(n23526), .o(n24120) );
na03f01 g20331 ( .a(n24120), .b(n23781), .c(n23754), .o(n24121) );
in01f01 g20332 ( .a(n24120), .o(n24122) );
oa12f01 g20333 ( .a(n24122), .b(n23654), .c(n23536), .o(n24123) );
na02f01 g20334 ( .a(n24123), .b(n24121), .o(n24124) );
ao12f01 g20335 ( .a(n23981), .b(n24124), .c(n24119), .o(n24125) );
no02f01 g20336 ( .a(n24124), .b(n24119), .o(n24126) );
ao12f01 g20337 ( .a(n23191), .b(n23301), .c(n23289), .o(n24127) );
no03f01 g20338 ( .a(n23886), .b(n23925), .c(n23891), .o(n24128) );
oa12f01 g20339 ( .a(n23973), .b(n23783), .c(n23526), .o(n24129) );
na03f01 g20340 ( .a(n23971), .b(n23656), .c(n23527), .o(n24130) );
na02f01 g20341 ( .a(n24130), .b(n24129), .o(n24131) );
no03f01 g20342 ( .a(n24131), .b(n24128), .c(n24127), .o(n24132) );
no03f01 g20343 ( .a(n24132), .b(n24126), .c(n24125), .o(n24133) );
no03f01 g20344 ( .a(n23959), .b(n23659), .c(n23517), .o(n24134) );
ao12f01 g20345 ( .a(n23957), .b(n23784), .c(n23753), .o(n24135) );
no02f01 g20346 ( .a(n24135), .b(n24134), .o(n24136) );
na03f01 g20347 ( .a(n23966), .b(n23965), .c(n23307), .o(n24137) );
oa12f01 g20348 ( .a(n23892), .b(n23963), .c(n23962), .o(n24138) );
na03f01 g20349 ( .a(n24138), .b(n24137), .c(n24136), .o(n24139) );
oa12f01 g20350 ( .a(n24139), .b(n24133), .c(n23976), .o(n24140) );
ao12f01 g20351 ( .a(n23956), .b(n24140), .c(n23968), .o(n24141) );
no03f01 g20352 ( .a(n24141), .b(n23950), .c(n23940), .o(n24142) );
in01f01 g20353 ( .a(n23875), .o(n24143) );
na03f01 g20354 ( .a(n23876), .b(n23666), .c(n23484), .o(n24144) );
oa12f01 g20355 ( .a(n23877), .b(n23789), .c(n23483), .o(n24145) );
na02f01 g20356 ( .a(n24145), .b(n24144), .o(n24146) );
no03f01 g20357 ( .a(n24146), .b(n24143), .c(n23873), .o(n24147) );
no03f01 g20358 ( .a(n24147), .b(n24142), .c(n23934), .o(n24148) );
na03f01 g20359 ( .a(n23865), .b(n23864), .c(n23314), .o(n24149) );
oa12f01 g20360 ( .a(n23862), .b(n23333), .c(n23857), .o(n24150) );
no03f01 g20361 ( .a(n23869), .b(n23669), .c(n23474), .o(n24151) );
ao12f01 g20362 ( .a(n23867), .b(n23790), .c(n23751), .o(n24152) );
no02f01 g20363 ( .a(n24152), .b(n24151), .o(n24153) );
na03f01 g20364 ( .a(n24153), .b(n24150), .c(n24149), .o(n24154) );
oa12f01 g20365 ( .a(n24154), .b(n24148), .c(n23881), .o(n24155) );
no03f01 g20366 ( .a(n23849), .b(n23844), .c(n23842), .o(n24156) );
ao12f01 g20367 ( .a(n24156), .b(n24155), .c(n23872), .o(n24157) );
no03f01 g20368 ( .a(n23837), .b(n23836), .c(n23833), .o(n24158) );
in01f01 g20369 ( .a(n24158), .o(n24159) );
oa12f01 g20370 ( .a(n24159), .b(n24157), .c(n23851), .o(n24160) );
na03f01 g20371 ( .a(n23816), .b(n23684), .c(n23454), .o(n24161) );
oa12f01 g20372 ( .a(n23817), .b(n23795), .c(n23453), .o(n24162) );
na02f01 g20373 ( .a(n24162), .b(n24161), .o(n24163) );
in01f01 g20374 ( .a(n23825), .o(n24164) );
no03f01 g20375 ( .a(n24164), .b(n23823), .c(n24163), .o(n24165) );
ao12f01 g20376 ( .a(n24165), .b(n24160), .c(n23838), .o(n24166) );
oa12f01 g20377 ( .a(n23815), .b(n24166), .c(n23826), .o(n24167) );
na02f01 g20378 ( .a(n24167), .b(n23810), .o(n24168) );
no02f01 g20379 ( .a(n23702), .b(n23694), .o(n24169) );
in01f01 g20380 ( .a(n24169), .o(n24170) );
no03f01 g20381 ( .a(n24170), .b(n23798), .c(n23434), .o(n24171) );
ao12f01 g20382 ( .a(n24169), .b(n23689), .c(n23435), .o(n24172) );
no02f01 g20383 ( .a(n24172), .b(n24171), .o(n24173) );
no02f01 g20384 ( .a(n24173), .b(n23360), .o(n24174) );
no03f01 g20385 ( .a(n24174), .b(n24168), .c(n23801), .o(n24175) );
na02f01 g20386 ( .a(n24173), .b(n23360), .o(n24176) );
no03f01 g20387 ( .a(n23746), .b(n23702), .c(n23799), .o(n24177) );
ao12f01 g20388 ( .a(n23747), .b(n23701), .c(n23745), .o(n24178) );
no02f01 g20389 ( .a(n24178), .b(n24177), .o(n24179) );
ao12f01 g20390 ( .a(n24179), .b(n24167), .c(n23810), .o(n24180) );
oa12f01 g20391 ( .a(n24176), .b(n24180), .c(n23741), .o(n24181) );
no04f01 g20392 ( .a(n23697), .b(n23694), .c(n23798), .d(n23434), .o(n24182) );
in01f01 g20393 ( .a(n23703), .o(n24183) );
no02f01 g20394 ( .a(n24183), .b(n24182), .o(n24184) );
no02f01 g20395 ( .a(n23420), .b(delay_add_ln22_unr8_stage4_stallmux_q_24_), .o(n24185) );
in01f01 g20396 ( .a(n24185), .o(n24186) );
na02f01 g20397 ( .a(n24186), .b(n24184), .o(n24187) );
no02f01 g20398 ( .a(n23419), .b(n23723), .o(n24188) );
in01f01 g20399 ( .a(n24188), .o(n24189) );
no02f01 g20400 ( .a(n23420), .b(delay_add_ln22_unr8_stage4_stallmux_q_25_), .o(n24190) );
no02f01 g20401 ( .a(n23419), .b(n23722), .o(n24191) );
no02f01 g20402 ( .a(n24191), .b(n24190), .o(n24192) );
na03f01 g20403 ( .a(n24192), .b(n24189), .c(n24187), .o(n24193) );
no02f01 g20404 ( .a(n24185), .b(n23704), .o(n24194) );
in01f01 g20405 ( .a(n24192), .o(n24195) );
oa12f01 g20406 ( .a(n24195), .b(n24188), .c(n24194), .o(n24196) );
na02f01 g20407 ( .a(n24196), .b(n24193), .o(n24197) );
no02f01 g20408 ( .a(n24188), .b(n24185), .o(n24198) );
in01f01 g20409 ( .a(n24198), .o(n24199) );
ao12f01 g20410 ( .a(n24199), .b(n23703), .c(n23699), .o(n24200) );
no03f01 g20411 ( .a(n24198), .b(n24183), .c(n24182), .o(n24201) );
no02f01 g20412 ( .a(n24201), .b(n24200), .o(n24202) );
in01f01 g20413 ( .a(n24202), .o(n24203) );
ao12f01 g20414 ( .a(n23741), .b(n24203), .c(n24197), .o(n24204) );
in01f01 g20415 ( .a(n23724), .o(n24205) );
ao12f01 g20416 ( .a(n23706), .b(n24205), .c(n23704), .o(n24206) );
in01f01 g20417 ( .a(n24206), .o(n24207) );
no02f01 g20418 ( .a(n23419), .b(n23719), .o(n24208) );
no02f01 g20419 ( .a(n24208), .b(n23705), .o(n24209) );
no02f01 g20420 ( .a(n24209), .b(n24207), .o(n24210) );
in01f01 g20421 ( .a(n24210), .o(n24211) );
na02f01 g20422 ( .a(n24209), .b(n24207), .o(n24212) );
na02f01 g20423 ( .a(n24212), .b(n24211), .o(n24213) );
no02f01 g20424 ( .a(n24213), .b(n23741), .o(n24214) );
no03f01 g20425 ( .a(n23724), .b(n24208), .c(n23709), .o(n24215) );
no02f01 g20426 ( .a(n23419), .b(n23720), .o(n24216) );
no02f01 g20427 ( .a(n24216), .b(n23710), .o(n24217) );
no02f01 g20428 ( .a(n24217), .b(n24215), .o(n24218) );
na02f01 g20429 ( .a(n24217), .b(n24215), .o(n24219) );
in01f01 g20430 ( .a(n24219), .o(n24220) );
no02f01 g20431 ( .a(n24220), .b(n24218), .o(n24221) );
in01f01 g20432 ( .a(n24221), .o(n24222) );
no02f01 g20433 ( .a(n24222), .b(n23741), .o(n24223) );
no02f01 g20434 ( .a(n24223), .b(n24214), .o(n24224) );
in01f01 g20435 ( .a(n24224), .o(n24225) );
no04f01 g20436 ( .a(n24225), .b(n24204), .c(n24181), .d(n24175), .o(n24226) );
in01f01 g20437 ( .a(n23725), .o(n24227) );
no02f01 g20438 ( .a(n23727), .b(n24227), .o(n24228) );
oa12f01 g20439 ( .a(n24228), .b(n23713), .c(n23712), .o(n24229) );
in01f01 g20440 ( .a(n24229), .o(n24230) );
no02f01 g20441 ( .a(n23729), .b(n23715), .o(n24231) );
no02f01 g20442 ( .a(n24231), .b(n24230), .o(n24232) );
in01f01 g20443 ( .a(n24232), .o(n24233) );
na02f01 g20444 ( .a(n24231), .b(n24230), .o(n24234) );
na02f01 g20445 ( .a(n24234), .b(n24233), .o(n24235) );
no02f01 g20446 ( .a(n24235), .b(n23741), .o(n24236) );
na02f01 g20447 ( .a(n23725), .b(n23712), .o(n24237) );
in01f01 g20448 ( .a(n24237), .o(n24238) );
no02f01 g20449 ( .a(n23727), .b(n23713), .o(n24239) );
no02f01 g20450 ( .a(n24239), .b(n24238), .o(n24240) );
na02f01 g20451 ( .a(n24239), .b(n24238), .o(n24241) );
in01f01 g20452 ( .a(n24241), .o(n24242) );
no02f01 g20453 ( .a(n24242), .b(n24240), .o(n24243) );
in01f01 g20454 ( .a(n24243), .o(n24244) );
no02f01 g20455 ( .a(n24244), .b(n23741), .o(n24245) );
no02f01 g20456 ( .a(n24245), .b(n24236), .o(n24246) );
in01f01 g20457 ( .a(n24246), .o(n24247) );
no02f01 g20458 ( .a(n23733), .b(n23718), .o(n24248) );
ao12f01 g20459 ( .a(n23731), .b(n23716), .c(n23714), .o(n24249) );
no02f01 g20460 ( .a(n24249), .b(n24248), .o(n24250) );
na02f01 g20461 ( .a(n24249), .b(n24248), .o(n24251) );
in01f01 g20462 ( .a(n24251), .o(n24252) );
no02f01 g20463 ( .a(n24252), .b(n24250), .o(n24253) );
in01f01 g20464 ( .a(n24253), .o(n24254) );
no02f01 g20465 ( .a(n24254), .b(n23741), .o(n24255) );
no02f01 g20466 ( .a(n24255), .b(n24247), .o(n24256) );
in01f01 g20467 ( .a(n24234), .o(n24257) );
no02f01 g20468 ( .a(n24257), .b(n24232), .o(n24258) );
ao12f01 g20469 ( .a(n23360), .b(n24243), .c(n24258), .o(n24259) );
oa12f01 g20470 ( .a(n23741), .b(n24259), .c(n24254), .o(n24260) );
in01f01 g20471 ( .a(n24212), .o(n24261) );
no02f01 g20472 ( .a(n24261), .b(n24210), .o(n24262) );
no02f01 g20473 ( .a(n24203), .b(n24197), .o(n24263) );
in01f01 g20474 ( .a(n24263), .o(n24264) );
no02f01 g20475 ( .a(n24264), .b(n24222), .o(n24265) );
ao12f01 g20476 ( .a(n23360), .b(n24265), .c(n24262), .o(n24266) );
in01f01 g20477 ( .a(n24266), .o(n24267) );
na02f01 g20478 ( .a(n24267), .b(n24260), .o(n24268) );
ao12f01 g20479 ( .a(n24268), .b(n24256), .c(n24226), .o(n24269) );
na02f01 g20480 ( .a(n24269), .b(n23744), .o(n24270) );
in01f01 g20481 ( .a(n24270), .o(n24271) );
no02f01 g20482 ( .a(n24269), .b(n23744), .o(n24272) );
no02f01 g20483 ( .a(n24272), .b(n24271), .o(n24273) );
no02f01 g20484 ( .a(n24273), .b(n5529), .o(n24274) );
no02f01 g20485 ( .a(n24253), .b(n23360), .o(n24275) );
no02f01 g20486 ( .a(n24275), .b(n24255), .o(n24276) );
ao12f01 g20487 ( .a(n23813), .b(n23814), .c(n23807), .o(n24277) );
no03f01 g20488 ( .a(n23809), .b(n23808), .c(n23806), .o(n24278) );
oa12f01 g20489 ( .a(n24163), .b(n24164), .c(n23823), .o(n24279) );
no03f01 g20490 ( .a(n23831), .b(n23827), .c(n23679), .o(n24280) );
ao12f01 g20491 ( .a(n23828), .b(n23829), .c(n23792), .o(n24281) );
no02f01 g20492 ( .a(n24281), .b(n24280), .o(n24282) );
in01f01 g20493 ( .a(n23837), .o(n24283) );
ao12f01 g20494 ( .a(n24282), .b(n24283), .c(n23835), .o(n24284) );
ao12f01 g20495 ( .a(n24153), .b(n24150), .c(n24149), .o(n24285) );
oa12f01 g20496 ( .a(n24146), .b(n24143), .c(n23873), .o(n24286) );
na03f01 g20497 ( .a(n23939), .b(n23936), .c(n23935), .o(n24287) );
oa12f01 g20498 ( .a(n23933), .b(n23928), .c(n23889), .o(n24288) );
oa12f01 g20499 ( .a(n23953), .b(n23955), .c(n23954), .o(n24289) );
na03f01 g20500 ( .a(n23949), .b(n23947), .c(n23945), .o(n24290) );
ao12f01 g20501 ( .a(n24136), .b(n24138), .c(n24137), .o(n24291) );
oa12f01 g20502 ( .a(n24131), .b(n24128), .c(n24127), .o(n24292) );
no02f01 g20503 ( .a(n23979), .b(n23288), .o(n24293) );
no02f01 g20504 ( .a(n23977), .b(n23291), .o(n24294) );
no02f01 g20505 ( .a(n24294), .b(n24293), .o(n24295) );
na03f01 g20506 ( .a(n23299), .b(n23293), .c(n23274), .o(n24296) );
oa12f01 g20507 ( .a(n23281), .b(n23884), .c(n23923), .o(n24297) );
no02f01 g20508 ( .a(n23985), .b(n23988), .o(n24298) );
no02f01 g20509 ( .a(n23986), .b(n23984), .o(n24299) );
no02f01 g20510 ( .a(n24299), .b(n24298), .o(n24300) );
na03f01 g20511 ( .a(n24300), .b(n24297), .c(n24296), .o(n24301) );
no02f01 g20512 ( .a(n23994), .b(n23273), .o(n24302) );
no02f01 g20513 ( .a(n23992), .b(n23295), .o(n24303) );
no02f01 g20514 ( .a(n24303), .b(n24302), .o(n24304) );
no02f01 g20515 ( .a(n23265), .b(n23921), .o(n24305) );
no02f01 g20516 ( .a(n23297), .b(n23259), .o(n24306) );
no03f01 g20517 ( .a(n24007), .b(n24306), .c(n24305), .o(n24307) );
na02f01 g20518 ( .a(n23920), .b(n23253), .o(n24308) );
na02f01 g20519 ( .a(n23258), .b(n23918), .o(n24309) );
na02f01 g20520 ( .a(n24309), .b(n24308), .o(n24310) );
na02f01 g20521 ( .a(n23914), .b(n23898), .o(n24311) );
na02f01 g20522 ( .a(n23246), .b(n23215), .o(n24312) );
na03f01 g20523 ( .a(n24019), .b(n24312), .c(n24311), .o(n24313) );
no02f01 g20524 ( .a(n23913), .b(n23240), .o(n24314) );
no02f01 g20525 ( .a(n23245), .b(n23911), .o(n24315) );
in01f01 g20526 ( .a(n24030), .o(n24316) );
oa12f01 g20527 ( .a(n24316), .b(n24315), .c(n24314), .o(n24317) );
na02f01 g20528 ( .a(n23910), .b(n23221), .o(n24318) );
na02f01 g20529 ( .a(n23239), .b(n23901), .o(n24319) );
ao12f01 g20530 ( .a(n24040), .b(n24319), .c(n24318), .o(n24320) );
no02f01 g20531 ( .a(n23238), .b(n23903), .o(n24321) );
no02f01 g20532 ( .a(n23909), .b(n23226), .o(n24322) );
in01f01 g20533 ( .a(n24051), .o(n24323) );
no03f01 g20534 ( .a(n24323), .b(n24322), .c(n24321), .o(n24324) );
ao12f01 g20535 ( .a(n24069), .b(n24067), .c(n24055), .o(n24325) );
oa12f01 g20536 ( .a(n24323), .b(n24322), .c(n24321), .o(n24326) );
oa12f01 g20537 ( .a(n24326), .b(n24325), .c(n24324), .o(n24327) );
na03f01 g20538 ( .a(n24040), .b(n24319), .c(n24318), .o(n24328) );
ao12f01 g20539 ( .a(n24320), .b(n24328), .c(n24327), .o(n24329) );
no03f01 g20540 ( .a(n24316), .b(n24315), .c(n24314), .o(n24330) );
oa12f01 g20541 ( .a(n24317), .b(n24330), .c(n24329), .o(n24331) );
ao12f01 g20542 ( .a(n24019), .b(n24312), .c(n24311), .o(n24332) );
ao12f01 g20543 ( .a(n24332), .b(n24331), .c(n24313), .o(n24333) );
no03f01 g20544 ( .a(n24103), .b(n24102), .c(n24101), .o(n24334) );
no02f01 g20545 ( .a(n24334), .b(n24333), .o(n24335) );
na02f01 g20546 ( .a(n24097), .b(n24104), .o(n24336) );
oa12f01 g20547 ( .a(n24310), .b(n24336), .c(n24335), .o(n24337) );
oa12f01 g20548 ( .a(n24098), .b(n24090), .c(n24335), .o(n24338) );
ao12f01 g20549 ( .a(n24307), .b(n24338), .c(n24337), .o(n24339) );
in01f01 g20550 ( .a(n24114), .o(n24340) );
no03f01 g20551 ( .a(n24340), .b(n24107), .c(n24339), .o(n24341) );
oa12f01 g20552 ( .a(n24340), .b(n24107), .c(n24339), .o(n24342) );
oa12f01 g20553 ( .a(n24342), .b(n24341), .c(n24304), .o(n24343) );
ao12f01 g20554 ( .a(n24300), .b(n24297), .c(n24296), .o(n24344) );
ao12f01 g20555 ( .a(n24344), .b(n24343), .c(n24301), .o(n24345) );
no03f01 g20556 ( .a(n24122), .b(n23654), .c(n23536), .o(n24346) );
ao12f01 g20557 ( .a(n24120), .b(n23781), .c(n23754), .o(n24347) );
no02f01 g20558 ( .a(n24347), .b(n24346), .o(n24348) );
oa12f01 g20559 ( .a(n24295), .b(n24348), .c(n24345), .o(n24349) );
na02f01 g20560 ( .a(n24348), .b(n24345), .o(n24350) );
na03f01 g20561 ( .a(n23975), .b(n23970), .c(n23969), .o(n24351) );
na03f01 g20562 ( .a(n24351), .b(n24350), .c(n24349), .o(n24352) );
no03f01 g20563 ( .a(n23967), .b(n23964), .c(n23961), .o(n24353) );
ao12f01 g20564 ( .a(n24353), .b(n24352), .c(n24292), .o(n24354) );
oa12f01 g20565 ( .a(n24290), .b(n24354), .c(n24291), .o(n24355) );
na03f01 g20566 ( .a(n24355), .b(n24289), .c(n24288), .o(n24356) );
na03f01 g20567 ( .a(n23880), .b(n23875), .c(n23874), .o(n24357) );
na03f01 g20568 ( .a(n24357), .b(n24356), .c(n24287), .o(n24358) );
no03f01 g20569 ( .a(n23871), .b(n23866), .c(n23863), .o(n24359) );
ao12f01 g20570 ( .a(n24359), .b(n24358), .c(n24286), .o(n24360) );
in01f01 g20571 ( .a(n24156), .o(n24361) );
oa12f01 g20572 ( .a(n24361), .b(n24360), .c(n24285), .o(n24362) );
ao12f01 g20573 ( .a(n24158), .b(n24362), .c(n23850), .o(n24363) );
na03f01 g20574 ( .a(n23825), .b(n23824), .c(n23820), .o(n24364) );
oa12f01 g20575 ( .a(n24364), .b(n24363), .c(n24284), .o(n24365) );
ao12f01 g20576 ( .a(n24278), .b(n24365), .c(n24279), .o(n24366) );
no02f01 g20577 ( .a(n24366), .b(n24277), .o(n24367) );
in01f01 g20578 ( .a(n24174), .o(n24368) );
na03f01 g20579 ( .a(n24368), .b(n24367), .c(n24179), .o(n24369) );
in01f01 g20580 ( .a(n24176), .o(n24370) );
oa12f01 g20581 ( .a(n23801), .b(n24366), .c(n24277), .o(n24371) );
ao12f01 g20582 ( .a(n24370), .b(n24371), .c(n23360), .o(n24372) );
in01f01 g20583 ( .a(n24204), .o(n24373) );
na04f01 g20584 ( .a(n24224), .b(n24373), .c(n24372), .d(n24369), .o(n24374) );
na02f01 g20585 ( .a(n24267), .b(n24374), .o(n24375) );
ao12f01 g20586 ( .a(n24259), .b(n24375), .c(n24246), .o(n24376) );
na02f01 g20587 ( .a(n24376), .b(n24276), .o(n24377) );
in01f01 g20588 ( .a(n24276), .o(n24378) );
in01f01 g20589 ( .a(n24259), .o(n24379) );
no02f01 g20590 ( .a(n24266), .b(n24226), .o(n24380) );
oa12f01 g20591 ( .a(n24379), .b(n24380), .c(n24247), .o(n24381) );
na02f01 g20592 ( .a(n24381), .b(n24378), .o(n24382) );
na02f01 g20593 ( .a(n24382), .b(n24377), .o(n24383) );
na02f01 g20594 ( .a(n24383), .b(n5529), .o(n24384) );
no03f01 g20595 ( .a(n24195), .b(n24188), .c(n24194), .o(n24385) );
ao12f01 g20596 ( .a(n24192), .b(n24189), .c(n24187), .o(n24386) );
no02f01 g20597 ( .a(n24386), .b(n24385), .o(n24387) );
no02f01 g20598 ( .a(n24387), .b(n23360), .o(n24388) );
no02f01 g20599 ( .a(n24197), .b(n23741), .o(n24389) );
no02f01 g20600 ( .a(n24389), .b(n24388), .o(n24390) );
in01f01 g20601 ( .a(n24390), .o(n24391) );
no02f01 g20602 ( .a(n24202), .b(n23360), .o(n24392) );
no02f01 g20603 ( .a(n24203), .b(n23741), .o(n24393) );
no03f01 g20604 ( .a(n24393), .b(n24181), .c(n24175), .o(n24394) );
no03f01 g20605 ( .a(n24394), .b(n24392), .c(n24391), .o(n24395) );
in01f01 g20606 ( .a(n24392), .o(n24396) );
in01f01 g20607 ( .a(n24393), .o(n24397) );
na03f01 g20608 ( .a(n24397), .b(n24372), .c(n24369), .o(n24398) );
ao12f01 g20609 ( .a(n24390), .b(n24398), .c(n24396), .o(n24399) );
oa12f01 g20610 ( .a(n5527), .b(n24399), .c(n24395), .o(n24400) );
na02f01 g20611 ( .a(n24176), .b(n24368), .o(n24401) );
no02f01 g20612 ( .a(n24401), .b(n24168), .o(n24402) );
no02f01 g20613 ( .a(n24370), .b(n24174), .o(n24403) );
no02f01 g20614 ( .a(n24403), .b(n24367), .o(n24404) );
no02f01 g20615 ( .a(n24404), .b(n24402), .o(n24405) );
no02f01 g20616 ( .a(n24166), .b(n23826), .o(n24406) );
no02f01 g20617 ( .a(n24278), .b(n24277), .o(n24407) );
na02f01 g20618 ( .a(n24407), .b(n24406), .o(n24408) );
na02f01 g20619 ( .a(n24365), .b(n24279), .o(n24409) );
na02f01 g20620 ( .a(n23815), .b(n23810), .o(n24410) );
na02f01 g20621 ( .a(n24410), .b(n24409), .o(n24411) );
ao12f01 g20622 ( .a(n5527), .b(n24411), .c(n24408), .o(n24412) );
no02f01 g20623 ( .a(n24363), .b(n24284), .o(n24413) );
no02f01 g20624 ( .a(n24165), .b(n23826), .o(n24414) );
na02f01 g20625 ( .a(n24414), .b(n24413), .o(n24415) );
na02f01 g20626 ( .a(n24160), .b(n23838), .o(n24416) );
na02f01 g20627 ( .a(n24364), .b(n24279), .o(n24417) );
na02f01 g20628 ( .a(n24417), .b(n24416), .o(n24418) );
na02f01 g20629 ( .a(n24418), .b(n24415), .o(n24419) );
na02f01 g20630 ( .a(n24419), .b(n5529), .o(n24420) );
no02f01 g20631 ( .a(n24360), .b(n24285), .o(n24421) );
in01f01 g20632 ( .a(n24421), .o(n24422) );
na02f01 g20633 ( .a(n24361), .b(n23850), .o(n24423) );
no02f01 g20634 ( .a(n24423), .b(n24422), .o(n24424) );
no02f01 g20635 ( .a(n24156), .b(n23851), .o(n24425) );
no02f01 g20636 ( .a(n24425), .b(n24421), .o(n24426) );
no02f01 g20637 ( .a(n24426), .b(n24424), .o(n24427) );
no02f01 g20638 ( .a(n24427), .b(n5527), .o(n24428) );
no04f01 g20639 ( .a(n24359), .b(n24148), .c(n23881), .d(n24285), .o(n24429) );
ao22f01 g20640 ( .a(n24154), .b(n23872), .c(n24358), .d(n24286), .o(n24430) );
no02f01 g20641 ( .a(n24430), .b(n24429), .o(n24431) );
no02f01 g20642 ( .a(n24431), .b(n5529), .o(n24432) );
in01f01 g20643 ( .a(n24432), .o(n24433) );
no02f01 g20644 ( .a(n23940), .b(n23934), .o(n24434) );
na02f01 g20645 ( .a(n24140), .b(n23968), .o(n24435) );
oa12f01 g20646 ( .a(n24290), .b(n24435), .c(n23950), .o(n24436) );
no02f01 g20647 ( .a(n24436), .b(n24434), .o(n24437) );
na02f01 g20648 ( .a(n24288), .b(n24287), .o(n24438) );
no02f01 g20649 ( .a(n24354), .b(n24291), .o(n24439) );
ao12f01 g20650 ( .a(n23956), .b(n24439), .c(n24289), .o(n24440) );
no02f01 g20651 ( .a(n24440), .b(n24438), .o(n24441) );
no02f01 g20652 ( .a(n24441), .b(n24437), .o(n24442) );
no02f01 g20653 ( .a(n24442), .b(n5527), .o(n24443) );
na02f01 g20654 ( .a(n24290), .b(n24289), .o(n24444) );
na02f01 g20655 ( .a(n24444), .b(n24435), .o(n24445) );
no02f01 g20656 ( .a(n23956), .b(n23950), .o(n24446) );
na02f01 g20657 ( .a(n24446), .b(n24439), .o(n24447) );
na02f01 g20658 ( .a(n24447), .b(n24445), .o(n24448) );
na02f01 g20659 ( .a(n24448), .b(n5529), .o(n24449) );
no02f01 g20660 ( .a(n24126), .b(n24125), .o(n24450) );
na02f01 g20661 ( .a(n24351), .b(n24292), .o(n24451) );
na02f01 g20662 ( .a(n24451), .b(n24450), .o(n24452) );
na02f01 g20663 ( .a(n24350), .b(n24349), .o(n24453) );
no02f01 g20664 ( .a(n24132), .b(n23976), .o(n24454) );
na02f01 g20665 ( .a(n24454), .b(n24453), .o(n24455) );
na02f01 g20666 ( .a(n24455), .b(n24452), .o(n24456) );
na02f01 g20667 ( .a(n24348), .b(n24295), .o(n24457) );
na02f01 g20668 ( .a(n24124), .b(n23981), .o(n24458) );
na02f01 g20669 ( .a(n24458), .b(n24457), .o(n24459) );
na02f01 g20670 ( .a(n24459), .b(n24119), .o(n24460) );
no02f01 g20671 ( .a(n24124), .b(n23981), .o(n24461) );
no02f01 g20672 ( .a(n24348), .b(n24295), .o(n24462) );
no02f01 g20673 ( .a(n24462), .b(n24461), .o(n24463) );
na02f01 g20674 ( .a(n24463), .b(n24345), .o(n24464) );
na02f01 g20675 ( .a(n24464), .b(n24460), .o(n24465) );
oa12f01 g20676 ( .a(n5529), .b(n24465), .c(n24456), .o(n24466) );
in01f01 g20677 ( .a(n24466), .o(n24467) );
no02f01 g20678 ( .a(n24133), .b(n23976), .o(n24468) );
no02f01 g20679 ( .a(n24353), .b(n24291), .o(n24469) );
no02f01 g20680 ( .a(n24469), .b(n24468), .o(n24470) );
na02f01 g20681 ( .a(n24352), .b(n24292), .o(n24471) );
na02f01 g20682 ( .a(n24139), .b(n23968), .o(n24472) );
no02f01 g20683 ( .a(n24472), .b(n24471), .o(n24473) );
no02f01 g20684 ( .a(n24473), .b(n24470), .o(n24474) );
no02f01 g20685 ( .a(n24474), .b(n5527), .o(n24475) );
no02f01 g20686 ( .a(n24475), .b(n24467), .o(n24476) );
na02f01 g20687 ( .a(n24476), .b(n24449), .o(n24477) );
no02f01 g20688 ( .a(n24477), .b(n24443), .o(n24478) );
na02f01 g20689 ( .a(n24356), .b(n24287), .o(n24479) );
no02f01 g20690 ( .a(n24147), .b(n23881), .o(n24480) );
na02f01 g20691 ( .a(n24480), .b(n24479), .o(n24481) );
no02f01 g20692 ( .a(n24142), .b(n23934), .o(n24482) );
na02f01 g20693 ( .a(n24357), .b(n24286), .o(n24483) );
na02f01 g20694 ( .a(n24483), .b(n24482), .o(n24484) );
na02f01 g20695 ( .a(n24484), .b(n24481), .o(n24485) );
na02f01 g20696 ( .a(n24485), .b(n5529), .o(n24486) );
na02f01 g20697 ( .a(n24485), .b(n5527), .o(n24487) );
na02f01 g20698 ( .a(n24440), .b(n24438), .o(n24488) );
na02f01 g20699 ( .a(n24436), .b(n24434), .o(n24489) );
na02f01 g20700 ( .a(n24489), .b(n24488), .o(n24490) );
na02f01 g20701 ( .a(n24490), .b(n5527), .o(n24491) );
na02f01 g20702 ( .a(n24491), .b(n24487), .o(n24492) );
ao12f01 g20703 ( .a(n24492), .b(n24486), .c(n24478), .o(n24493) );
no02f01 g20704 ( .a(n24431), .b(n5527), .o(n24494) );
oa12f01 g20705 ( .a(n24433), .b(n24494), .c(n24493), .o(n24495) );
no02f01 g20706 ( .a(n24427), .b(n5529), .o(n24496) );
no02f01 g20707 ( .a(n24496), .b(n24495), .o(n24497) );
na02f01 g20708 ( .a(n24362), .b(n23850), .o(n24498) );
na02f01 g20709 ( .a(n24159), .b(n23838), .o(n24499) );
no02f01 g20710 ( .a(n24499), .b(n24498), .o(n24500) );
no02f01 g20711 ( .a(n24157), .b(n23851), .o(n24501) );
no02f01 g20712 ( .a(n24158), .b(n24284), .o(n24502) );
no02f01 g20713 ( .a(n24502), .b(n24501), .o(n24503) );
no02f01 g20714 ( .a(n24503), .b(n24500), .o(n24504) );
no02f01 g20715 ( .a(n24504), .b(n5527), .o(n24505) );
no03f01 g20716 ( .a(n24505), .b(n24497), .c(n24428), .o(n24506) );
na02f01 g20717 ( .a(n24506), .b(n24420), .o(n24507) );
no02f01 g20718 ( .a(n24507), .b(n24412), .o(n24508) );
oa12f01 g20719 ( .a(n24508), .b(n24405), .c(n5527), .o(n24509) );
na02f01 g20720 ( .a(n24403), .b(n24367), .o(n24510) );
na02f01 g20721 ( .a(n24401), .b(n24168), .o(n24511) );
na02f01 g20722 ( .a(n24511), .b(n24510), .o(n24512) );
no02f01 g20723 ( .a(n24410), .b(n24409), .o(n24513) );
no02f01 g20724 ( .a(n24407), .b(n24406), .o(n24514) );
oa12f01 g20725 ( .a(n5527), .b(n24514), .c(n24513), .o(n24515) );
no02f01 g20726 ( .a(n24417), .b(n24416), .o(n24516) );
no02f01 g20727 ( .a(n24414), .b(n24413), .o(n24517) );
no02f01 g20728 ( .a(n24517), .b(n24516), .o(n24518) );
no02f01 g20729 ( .a(n24518), .b(n5529), .o(n24519) );
no02f01 g20730 ( .a(n24504), .b(n5529), .o(n24520) );
no02f01 g20731 ( .a(n24520), .b(n24519), .o(n24521) );
na02f01 g20732 ( .a(n24521), .b(n24515), .o(n24522) );
ao12f01 g20733 ( .a(n24522), .b(n24512), .c(n5527), .o(n24523) );
no02f01 g20734 ( .a(n24174), .b(n24168), .o(n24524) );
no02f01 g20735 ( .a(n23801), .b(n23741), .o(n24525) );
no02f01 g20736 ( .a(n24179), .b(n23360), .o(n24526) );
no02f01 g20737 ( .a(n24526), .b(n24525), .o(n24527) );
oa12f01 g20738 ( .a(n24527), .b(n24370), .c(n24524), .o(n24528) );
na02f01 g20739 ( .a(n24368), .b(n24367), .o(n24529) );
in01f01 g20740 ( .a(n24527), .o(n24530) );
na03f01 g20741 ( .a(n24530), .b(n24176), .c(n24529), .o(n24531) );
na02f01 g20742 ( .a(n24531), .b(n24528), .o(n24532) );
ao22f01 g20743 ( .a(n24532), .b(n5529), .c(n24523), .d(n24509), .o(n24533) );
no02f01 g20744 ( .a(n24393), .b(n24392), .o(n24534) );
oa12f01 g20745 ( .a(n24534), .b(n24181), .c(n24175), .o(n24535) );
in01f01 g20746 ( .a(n24534), .o(n24536) );
na03f01 g20747 ( .a(n24536), .b(n24372), .c(n24369), .o(n24537) );
na02f01 g20748 ( .a(n24537), .b(n24535), .o(n24538) );
na02f01 g20749 ( .a(n24538), .b(n5529), .o(n24539) );
na02f01 g20750 ( .a(n24539), .b(n24533), .o(n24540) );
ao12f01 g20751 ( .a(n24536), .b(n24372), .c(n24369), .o(n24541) );
no03f01 g20752 ( .a(n24534), .b(n24181), .c(n24175), .o(n24542) );
no02f01 g20753 ( .a(n24542), .b(n24541), .o(n24543) );
no02f01 g20754 ( .a(n24543), .b(n5529), .o(n24544) );
ao12f01 g20755 ( .a(n24530), .b(n24176), .c(n24529), .o(n24545) );
no03f01 g20756 ( .a(n24527), .b(n24370), .c(n24524), .o(n24546) );
no02f01 g20757 ( .a(n24546), .b(n24545), .o(n24547) );
no02f01 g20758 ( .a(n24547), .b(n5529), .o(n24548) );
no02f01 g20759 ( .a(n24548), .b(n24544), .o(n24549) );
no03f01 g20760 ( .a(n24204), .b(n24181), .c(n24175), .o(n24550) );
no02f01 g20761 ( .a(n24263), .b(n23360), .o(n24551) );
no02f01 g20762 ( .a(n24262), .b(n23360), .o(n24552) );
no02f01 g20763 ( .a(n24552), .b(n24214), .o(n24553) );
in01f01 g20764 ( .a(n24553), .o(n24554) );
no03f01 g20765 ( .a(n24554), .b(n24551), .c(n24550), .o(n24555) );
na03f01 g20766 ( .a(n24373), .b(n24372), .c(n24369), .o(n24556) );
in01f01 g20767 ( .a(n24551), .o(n24557) );
ao12f01 g20768 ( .a(n24553), .b(n24557), .c(n24556), .o(n24558) );
oa12f01 g20769 ( .a(n5527), .b(n24558), .c(n24555), .o(n24559) );
na04f01 g20770 ( .a(n24559), .b(n24549), .c(n24540), .d(n24400), .o(n24560) );
no02f01 g20771 ( .a(n24558), .b(n24555), .o(n24561) );
no02f01 g20772 ( .a(n24561), .b(n5527), .o(n24562) );
no02f01 g20773 ( .a(n24399), .b(n24395), .o(n24563) );
no02f01 g20774 ( .a(n24563), .b(n5527), .o(n24564) );
no02f01 g20775 ( .a(n24564), .b(n24562), .o(n24565) );
na02f01 g20776 ( .a(n24565), .b(n24560), .o(n24566) );
no02f01 g20777 ( .a(n24258), .b(n23360), .o(n24567) );
no02f01 g20778 ( .a(n24567), .b(n24236), .o(n24568) );
no02f01 g20779 ( .a(n24243), .b(n23360), .o(n24569) );
no03f01 g20780 ( .a(n24266), .b(n24569), .c(n24226), .o(n24570) );
no03f01 g20781 ( .a(n24570), .b(n24568), .c(n24245), .o(n24571) );
in01f01 g20782 ( .a(n24245), .o(n24572) );
in01f01 g20783 ( .a(n24568), .o(n24573) );
in01f01 g20784 ( .a(n24569), .o(n24574) );
na03f01 g20785 ( .a(n24267), .b(n24574), .c(n24374), .o(n24575) );
ao12f01 g20786 ( .a(n24573), .b(n24575), .c(n24572), .o(n24576) );
oa12f01 g20787 ( .a(n5529), .b(n24576), .c(n24571), .o(n24577) );
in01f01 g20788 ( .a(n24214), .o(n24578) );
no02f01 g20789 ( .a(n24221), .b(n23360), .o(n24579) );
no02f01 g20790 ( .a(n24579), .b(n24223), .o(n24580) );
in01f01 g20791 ( .a(n24580), .o(n24581) );
in01f01 g20792 ( .a(n24552), .o(n24582) );
na03f01 g20793 ( .a(n24557), .b(n24582), .c(n24556), .o(n24583) );
ao12f01 g20794 ( .a(n24581), .b(n24583), .c(n24578), .o(n24584) );
no03f01 g20795 ( .a(n24551), .b(n24552), .c(n24550), .o(n24585) );
no03f01 g20796 ( .a(n24585), .b(n24580), .c(n24214), .o(n24586) );
oa12f01 g20797 ( .a(n5529), .b(n24586), .c(n24584), .o(n24587) );
no02f01 g20798 ( .a(n24569), .b(n24245), .o(n24588) );
in01f01 g20799 ( .a(n24588), .o(n24589) );
na02f01 g20800 ( .a(n24589), .b(n24375), .o(n24590) );
na02f01 g20801 ( .a(n24588), .b(n24380), .o(n24591) );
na02f01 g20802 ( .a(n24591), .b(n24590), .o(n24592) );
na02f01 g20803 ( .a(n24592), .b(n5529), .o(n24593) );
na03f01 g20804 ( .a(n24593), .b(n24587), .c(n24577), .o(n24594) );
na03f01 g20805 ( .a(n24575), .b(n24573), .c(n24572), .o(n24595) );
oa12f01 g20806 ( .a(n24568), .b(n24570), .c(n24245), .o(n24596) );
ao12f01 g20807 ( .a(n5529), .b(n24596), .c(n24595), .o(n24597) );
no02f01 g20808 ( .a(n24586), .b(n24584), .o(n24598) );
no02f01 g20809 ( .a(n24598), .b(n5529), .o(n24599) );
no02f01 g20810 ( .a(n24588), .b(n24380), .o(n24600) );
no02f01 g20811 ( .a(n24589), .b(n24375), .o(n24601) );
no02f01 g20812 ( .a(n24601), .b(n24600), .o(n24602) );
no02f01 g20813 ( .a(n24602), .b(n5529), .o(n24603) );
no03f01 g20814 ( .a(n24603), .b(n24599), .c(n24597), .o(n24604) );
oa12f01 g20815 ( .a(n24604), .b(n24594), .c(n24566), .o(n24605) );
no02f01 g20816 ( .a(n24381), .b(n24378), .o(n24606) );
no02f01 g20817 ( .a(n24376), .b(n24276), .o(n24607) );
no02f01 g20818 ( .a(n24607), .b(n24606), .o(n24608) );
no02f01 g20819 ( .a(n24608), .b(n5529), .o(n24609) );
oa12f01 g20820 ( .a(n24384), .b(n24609), .c(n24605), .o(n24610) );
no02f01 g20821 ( .a(n24273), .b(n5527), .o(n24611) );
in01f01 g20822 ( .a(n24611), .o(n24612) );
ao12f01 g20823 ( .a(n24274), .b(n24612), .c(n24610), .o(n24613) );
no02f01 g20824 ( .a(n23739), .b(n5119), .o(n24614) );
no02f01 g20825 ( .a(n24221), .b(n5142), .o(n24615) );
no02f01 g20826 ( .a(n24202), .b(n5142), .o(n24616) );
na02f01 g20827 ( .a(n23990), .b(n5119), .o(n24617) );
oa12f01 g20828 ( .a(n24617), .b(n24348), .c(n5142), .o(n24618) );
ao12f01 g20829 ( .a(n24618), .b(n24131), .c(n5119), .o(n24619) );
oa12f01 g20830 ( .a(n24619), .b(n24136), .c(n5142), .o(n24620) );
ao12f01 g20831 ( .a(n24620), .b(n23953), .c(n5119), .o(n24621) );
oa12f01 g20832 ( .a(n24621), .b(n23939), .c(n5142), .o(n24622) );
ao12f01 g20833 ( .a(n24622), .b(n24146), .c(n5119), .o(n24623) );
na02f01 g20834 ( .a(n24623), .b(n24153), .o(n24624) );
oa12f01 g20835 ( .a(n5119), .b(n24624), .c(n23849), .o(n24625) );
oa12f01 g20836 ( .a(n24625), .b(n24282), .c(n5142), .o(n24626) );
ao12f01 g20837 ( .a(n5142), .b(n24162), .c(n24161), .o(n24627) );
no04f01 g20838 ( .a(n24627), .b(n24626), .c(n23812), .d(n23811), .o(n24628) );
ao12f01 g20839 ( .a(n5119), .b(n23805), .c(n23803), .o(n24629) );
oa12f01 g20840 ( .a(n5142), .b(n23849), .c(n23833), .o(n24630) );
oa12f01 g20841 ( .a(n24630), .b(n23820), .c(n5119), .o(n24631) );
no03f01 g20842 ( .a(n24631), .b(n24629), .c(n24628), .o(n24632) );
na03f01 g20843 ( .a(n24169), .b(n23689), .c(n23435), .o(n24633) );
oa12f01 g20844 ( .a(n24170), .b(n23798), .c(n23434), .o(n24634) );
ao12f01 g20845 ( .a(n5142), .b(n24634), .c(n24633), .o(n24635) );
no04f01 g20846 ( .a(n24635), .b(n24632), .c(n24178), .d(n24177), .o(n24636) );
na02f01 g20847 ( .a(n24634), .b(n24633), .o(n24637) );
na02f01 g20848 ( .a(n24637), .b(n5142), .o(n24638) );
oa12f01 g20849 ( .a(n24638), .b(n24179), .c(n5119), .o(n24639) );
no02f01 g20850 ( .a(n24639), .b(n24636), .o(n24640) );
no03f01 g20851 ( .a(n24640), .b(n24616), .c(n24197), .o(n24641) );
ao12f01 g20852 ( .a(n5119), .b(n24202), .c(n24387), .o(n24642) );
oa22f01 g20853 ( .a(n24642), .b(n24641), .c(n24262), .d(n5142), .o(n24643) );
no02f01 g20854 ( .a(n24643), .b(n24615), .o(n24644) );
oa12f01 g20855 ( .a(n24644), .b(n24243), .c(n5142), .o(n24645) );
no02f01 g20856 ( .a(n24258), .b(n5142), .o(n24646) );
no02f01 g20857 ( .a(n24646), .b(n24645), .o(n24647) );
ao12f01 g20858 ( .a(n5119), .b(n24221), .c(n24262), .o(n24648) );
ao12f01 g20859 ( .a(n24648), .b(n24244), .c(n5142), .o(n24649) );
na02f01 g20860 ( .a(n24235), .b(n5142), .o(n24650) );
na02f01 g20861 ( .a(n24650), .b(n24649), .o(n24651) );
oa22f01 g20862 ( .a(n24651), .b(n24647), .c(n24253), .d(n5142), .o(n24652) );
no02f01 g20863 ( .a(n24253), .b(n5119), .o(n24653) );
in01f01 g20864 ( .a(n24653), .o(n24654) );
ao22f01 g20865 ( .a(n24654), .b(n24652), .c(n23742), .d(n5119), .o(n24655) );
no03f01 g20866 ( .a(n24655), .b(n24614), .c(n23742), .o(n24656) );
na02f01 g20867 ( .a(n24654), .b(n24652), .o(n24657) );
no02f01 g20868 ( .a(n23739), .b(n5119), .o(n24659) );
no02f01 g20869 ( .a(n24659), .b(n24656), .o(n24660) );
in01f01 g20870 ( .a(n24660), .o(n24661) );
ao12f01 g20871 ( .a(n24661), .b(n23321), .c(n23170), .o(n24662) );
ao12f01 g20872 ( .a(n24661), .b(n23310), .c(n23305), .o(n24663) );
no02f01 g20873 ( .a(n24663), .b(n24662), .o(n24664) );
na03f01 g20874 ( .a(n24654), .b(n24652), .c(n23739), .o(n24665) );
na02f01 g20875 ( .a(n24657), .b(n23742), .o(n24666) );
na03f01 g20876 ( .a(n24666), .b(n24665), .c(n23291), .o(n24667) );
in01f01 g20877 ( .a(n24616), .o(n24668) );
no03f01 g20878 ( .a(n23847), .b(n23791), .c(n23463), .o(n24669) );
ao12f01 g20879 ( .a(n23845), .b(n23670), .c(n23464), .o(n24670) );
no02f01 g20880 ( .a(n24670), .b(n24669), .o(n24671) );
oa12f01 g20881 ( .a(n5119), .b(n24124), .c(n23990), .o(n24672) );
oa12f01 g20882 ( .a(n24672), .b(n23975), .c(n5142), .o(n24673) );
ao12f01 g20883 ( .a(n24673), .b(n23961), .c(n5119), .o(n24674) );
oa12f01 g20884 ( .a(n24674), .b(n23945), .c(n5142), .o(n24675) );
ao12f01 g20885 ( .a(n24675), .b(n23933), .c(n5119), .o(n24676) );
oa12f01 g20886 ( .a(n24676), .b(n23880), .c(n5142), .o(n24677) );
oa12f01 g20887 ( .a(n5119), .b(n24677), .c(n23871), .o(n24678) );
oa12f01 g20888 ( .a(n24678), .b(n24671), .c(n5142), .o(n24679) );
ao12f01 g20889 ( .a(n24679), .b(n23833), .c(n5119), .o(n24680) );
oa12f01 g20890 ( .a(n5119), .b(n23819), .c(n23818), .o(n24681) );
na04f01 g20891 ( .a(n24681), .b(n24680), .c(n23805), .d(n23803), .o(n24682) );
oa12f01 g20892 ( .a(n5142), .b(n23812), .c(n23811), .o(n24683) );
ao12f01 g20893 ( .a(n5119), .b(n24671), .c(n24282), .o(n24684) );
ao12f01 g20894 ( .a(n24684), .b(n24163), .c(n5142), .o(n24685) );
na03f01 g20895 ( .a(n24685), .b(n24683), .c(n24682), .o(n24686) );
oa12f01 g20896 ( .a(n5119), .b(n24172), .c(n24171), .o(n24687) );
na04f01 g20897 ( .a(n24687), .b(n24686), .c(n23800), .d(n23748), .o(n24688) );
no02f01 g20898 ( .a(n24173), .b(n5119), .o(n24689) );
ao12f01 g20899 ( .a(n24689), .b(n23801), .c(n5142), .o(n24690) );
na02f01 g20900 ( .a(n24690), .b(n24688), .o(n24691) );
na03f01 g20901 ( .a(n24691), .b(n24668), .c(n24387), .o(n24692) );
oa12f01 g20902 ( .a(n5142), .b(n24203), .c(n24197), .o(n24693) );
ao22f01 g20903 ( .a(n24693), .b(n24692), .c(n24213), .d(n5119), .o(n24694) );
oa12f01 g20904 ( .a(n24694), .b(n24221), .c(n5142), .o(n24695) );
ao12f01 g20905 ( .a(n24695), .b(n24244), .c(n5119), .o(n24696) );
na02f01 g20906 ( .a(n24235), .b(n5119), .o(n24697) );
na02f01 g20907 ( .a(n24697), .b(n24696), .o(n24698) );
in01f01 g20908 ( .a(n24648), .o(n24699) );
oa12f01 g20909 ( .a(n24699), .b(n24243), .c(n5119), .o(n24700) );
no02f01 g20910 ( .a(n24258), .b(n5119), .o(n24701) );
no02f01 g20911 ( .a(n24701), .b(n24700), .o(n24702) );
na02f01 g20912 ( .a(n24702), .b(n24698), .o(n24703) );
no02f01 g20913 ( .a(n24703), .b(n24254), .o(n24704) );
no02f01 g20914 ( .a(n24651), .b(n24647), .o(n24705) );
no02f01 g20915 ( .a(n24705), .b(n24253), .o(n24706) );
no03f01 g20916 ( .a(n24706), .b(n24704), .c(n23293), .o(n24707) );
na02f01 g20917 ( .a(n24650), .b(n24697), .o(n24708) );
oa12f01 g20918 ( .a(n24708), .b(n24700), .c(n24696), .o(n24709) );
no02f01 g20919 ( .a(n24701), .b(n24646), .o(n24710) );
na03f01 g20920 ( .a(n24710), .b(n24649), .c(n24645), .o(n24711) );
na03f01 g20921 ( .a(n24711), .b(n24709), .c(n23295), .o(n24712) );
ao12f01 g20922 ( .a(n24243), .b(n24699), .c(n24695), .o(n24713) );
no03f01 g20923 ( .a(n24648), .b(n24644), .c(n24244), .o(n24714) );
no03f01 g20924 ( .a(n24714), .b(n24713), .c(n23297), .o(n24715) );
na02f01 g20925 ( .a(n24213), .b(n5142), .o(n24716) );
in01f01 g20926 ( .a(n24716), .o(n24717) );
no03f01 g20927 ( .a(n24717), .b(n24694), .c(n24222), .o(n24718) );
ao12f01 g20928 ( .a(n24221), .b(n24716), .c(n24643), .o(n24719) );
no03f01 g20929 ( .a(n24719), .b(n24718), .c(n23258), .o(n24720) );
in01f01 g20930 ( .a(n24720), .o(n24721) );
no03f01 g20931 ( .a(n24642), .b(n24641), .c(n24213), .o(n24722) );
ao12f01 g20932 ( .a(n24262), .b(n24693), .c(n24692), .o(n24723) );
no03f01 g20933 ( .a(n24723), .b(n24722), .c(n23917), .o(n24724) );
na02f01 g20934 ( .a(n23801), .b(n5142), .o(n24725) );
oa12f01 g20935 ( .a(n5142), .b(n24201), .c(n24200), .o(n24726) );
na04f01 g20936 ( .a(n24726), .b(n24725), .c(n24638), .d(n24688), .o(n24727) );
na03f01 g20937 ( .a(n24727), .b(n24668), .c(n24197), .o(n24728) );
no02f01 g20938 ( .a(n24179), .b(n5119), .o(n24729) );
oa12f01 g20939 ( .a(n24198), .b(n24183), .c(n24182), .o(n24730) );
na03f01 g20940 ( .a(n24199), .b(n23703), .c(n23699), .o(n24731) );
ao12f01 g20941 ( .a(n5119), .b(n24731), .c(n24730), .o(n24732) );
no04f01 g20942 ( .a(n24732), .b(n24729), .c(n24689), .d(n24636), .o(n24733) );
oa12f01 g20943 ( .a(n24387), .b(n24733), .c(n24616), .o(n24734) );
ao12f01 g20944 ( .a(n23215), .b(n24734), .c(n24728), .o(n24735) );
no02f01 g20945 ( .a(n24635), .b(n24632), .o(n24736) );
no03f01 g20946 ( .a(n24689), .b(n24736), .c(n23801), .o(n24737) );
na02f01 g20947 ( .a(n24687), .b(n24686), .o(n24738) );
ao12f01 g20948 ( .a(n24179), .b(n24638), .c(n24738), .o(n24739) );
no02f01 g20949 ( .a(n24739), .b(n24737), .o(n24740) );
no02f01 g20950 ( .a(n23820), .b(n5119), .o(n24741) );
ao12f01 g20951 ( .a(n24627), .b(n24630), .c(n24626), .o(n24742) );
no03f01 g20952 ( .a(n24742), .b(n24741), .c(n23806), .o(n24743) );
na02f01 g20953 ( .a(n24163), .b(n5142), .o(n24744) );
oa22f01 g20954 ( .a(n24684), .b(n24680), .c(n23820), .d(n5142), .o(n24745) );
ao12f01 g20955 ( .a(n23813), .b(n24745), .c(n24744), .o(n24746) );
oa12f01 g20956 ( .a(n23237), .b(n24746), .c(n24743), .o(n24747) );
na03f01 g20957 ( .a(n24630), .b(n24626), .c(n23820), .o(n24748) );
oa12f01 g20958 ( .a(n24163), .b(n24684), .c(n24680), .o(n24749) );
na03f01 g20959 ( .a(n24749), .b(n24748), .c(n23231), .o(n24750) );
ao12f01 g20960 ( .a(n23231), .b(n24749), .c(n24748), .o(n24751) );
oa12f01 g20961 ( .a(n5119), .b(n24624), .c(n23849), .o(n24752) );
no02f01 g20962 ( .a(n24752), .b(n23833), .o(n24753) );
in01f01 g20963 ( .a(n24624), .o(n24754) );
ao12f01 g20964 ( .a(n5142), .b(n24754), .c(n24671), .o(n24755) );
no02f01 g20965 ( .a(n24755), .b(n24282), .o(n24756) );
no02f01 g20966 ( .a(n23043), .b(n22935), .o(n24757) );
no02f01 g20967 ( .a(n24757), .b(n23042), .o(n24758) );
na02f01 g20968 ( .a(n24757), .b(n23042), .o(n24759) );
in01f01 g20969 ( .a(n24759), .o(n24760) );
no02f01 g20970 ( .a(n24760), .b(n24758), .o(n24761) );
no03f01 g20971 ( .a(n24761), .b(n24756), .c(n24753), .o(n24762) );
oa12f01 g20972 ( .a(n24761), .b(n24756), .c(n24753), .o(n24763) );
no02f01 g20973 ( .a(n24678), .b(n23849), .o(n24764) );
ao12f01 g20974 ( .a(n24671), .b(n24624), .c(n5119), .o(n24765) );
no02f01 g20975 ( .a(n23040), .b(n22945), .o(n24766) );
no02f01 g20976 ( .a(n24766), .b(n23039), .o(n24767) );
na02f01 g20977 ( .a(n24766), .b(n23039), .o(n24768) );
in01f01 g20978 ( .a(n24768), .o(n24769) );
no02f01 g20979 ( .a(n24769), .b(n24767), .o(n24770) );
no03f01 g20980 ( .a(n24770), .b(n24765), .c(n24764), .o(n24771) );
in01f01 g20981 ( .a(n24771), .o(n24772) );
na03f01 g20982 ( .a(n24624), .b(n24671), .c(n5119), .o(n24773) );
na02f01 g20983 ( .a(n24678), .b(n23849), .o(n24774) );
in01f01 g20984 ( .a(n24770), .o(n24775) );
ao12f01 g20985 ( .a(n24775), .b(n24774), .c(n24773), .o(n24776) );
na02f01 g20986 ( .a(n24622), .b(n23880), .o(n24777) );
na02f01 g20987 ( .a(n24676), .b(n24146), .o(n24778) );
in01f01 g20988 ( .a(n23032), .o(n24779) );
no02f01 g20989 ( .a(n23036), .b(n22965), .o(n24780) );
in01f01 g20990 ( .a(n24780), .o(n24781) );
no02f01 g20991 ( .a(n24781), .b(n24779), .o(n24782) );
no02f01 g20992 ( .a(n24780), .b(n23032), .o(n24783) );
no02f01 g20993 ( .a(n24783), .b(n24782), .o(n24784) );
in01f01 g20994 ( .a(n24784), .o(n24785) );
ao12f01 g20995 ( .a(n24785), .b(n24778), .c(n24777), .o(n24786) );
no02f01 g20996 ( .a(n24621), .b(n23933), .o(n24787) );
no02f01 g20997 ( .a(n24675), .b(n23939), .o(n24788) );
in01f01 g20998 ( .a(n23029), .o(n24789) );
no02f01 g20999 ( .a(n23030), .b(n22975), .o(n24790) );
no02f01 g21000 ( .a(n24790), .b(n24789), .o(n24791) );
na02f01 g21001 ( .a(n24790), .b(n24789), .o(n24792) );
in01f01 g21002 ( .a(n24792), .o(n24793) );
no02f01 g21003 ( .a(n24793), .b(n24791), .o(n24794) );
no03f01 g21004 ( .a(n24794), .b(n24788), .c(n24787), .o(n24795) );
no02f01 g21005 ( .a(n24674), .b(n23953), .o(n24796) );
no02f01 g21006 ( .a(n24620), .b(n23945), .o(n24797) );
in01f01 g21007 ( .a(n23027), .o(n24798) );
no03f01 g21008 ( .a(n23028), .b(n24798), .c(n22992), .o(n24799) );
no02f01 g21009 ( .a(n23028), .b(n22992), .o(n24800) );
no02f01 g21010 ( .a(n24800), .b(n23027), .o(n24801) );
no02f01 g21011 ( .a(n24801), .b(n24799), .o(n24802) );
no03f01 g21012 ( .a(n24802), .b(n24797), .c(n24796), .o(n24803) );
in01f01 g21013 ( .a(n24803), .o(n24804) );
no02f01 g21014 ( .a(n24673), .b(n24136), .o(n24805) );
no02f01 g21015 ( .a(n24619), .b(n23961), .o(n24806) );
no03f01 g21016 ( .a(n23026), .b(n23024), .c(n23001), .o(n24807) );
in01f01 g21017 ( .a(n23024), .o(n24808) );
no02f01 g21018 ( .a(n23026), .b(n23001), .o(n24809) );
no02f01 g21019 ( .a(n24809), .b(n24808), .o(n24810) );
no02f01 g21020 ( .a(n24810), .b(n24807), .o(n24811) );
oa12f01 g21021 ( .a(n24811), .b(n24806), .c(n24805), .o(n24812) );
no02f01 g21022 ( .a(n24672), .b(n24131), .o(n24813) );
no02f01 g21023 ( .a(n24618), .b(n23975), .o(n24814) );
in01f01 g21024 ( .a(n23008), .o(n24815) );
in01f01 g21025 ( .a(n23022), .o(n24816) );
no03f01 g21026 ( .a(n23023), .b(n24816), .c(n24815), .o(n24817) );
in01f01 g21027 ( .a(n23023), .o(n24818) );
ao12f01 g21028 ( .a(n23022), .b(n24818), .c(n23008), .o(n24819) );
no02f01 g21029 ( .a(n24819), .b(n24817), .o(n24820) );
no03f01 g21030 ( .a(n24820), .b(n24814), .c(n24813), .o(n24821) );
in01f01 g21031 ( .a(n24821), .o(n24822) );
na02f01 g21032 ( .a(n24618), .b(n23975), .o(n24823) );
na02f01 g21033 ( .a(n24672), .b(n24131), .o(n24824) );
in01f01 g21034 ( .a(n24820), .o(n24825) );
ao12f01 g21035 ( .a(n24825), .b(n24824), .c(n24823), .o(n24826) );
in01f01 g21036 ( .a(n23014), .o(n24827) );
no02f01 g21037 ( .a(n23021), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_1_), .o(n24828) );
no03f01 g21038 ( .a(n23020), .b(n23019), .c(n23009), .o(n24829) );
no03f01 g21039 ( .a(n24829), .b(n24828), .c(n24827), .o(n24830) );
no02f01 g21040 ( .a(n24829), .b(n24828), .o(n24831) );
no02f01 g21041 ( .a(n24831), .b(n23014), .o(n24832) );
no02f01 g21042 ( .a(n24832), .b(n24830), .o(n24833) );
in01f01 g21043 ( .a(n24833), .o(n24834) );
in01f01 g21044 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_0_), .o(n24835) );
no02f01 g21045 ( .a(n23013), .b(n24835), .o(n24836) );
ao12f01 g21046 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_0_), .b(n23012), .c(n23011), .o(n24837) );
no02f01 g21047 ( .a(n24837), .b(n24836), .o(n24838) );
no02f01 g21048 ( .a(n24838), .b(n24300), .o(n24839) );
in01f01 g21049 ( .a(n24839), .o(n24840) );
no02f01 g21050 ( .a(n24840), .b(n24834), .o(n24841) );
in01f01 g21051 ( .a(n24841), .o(n24842) );
no02f01 g21052 ( .a(n24300), .b(n5142), .o(n24843) );
no02f01 g21053 ( .a(n24843), .b(n24348), .o(n24844) );
no02f01 g21054 ( .a(n24617), .b(n24124), .o(n24845) );
no02f01 g21055 ( .a(n24845), .b(n24844), .o(n24846) );
no02f01 g21056 ( .a(n24839), .b(n24833), .o(n24847) );
ao12f01 g21057 ( .a(n24847), .b(n24846), .c(n24842), .o(n24848) );
oa12f01 g21058 ( .a(n24822), .b(n24848), .c(n24826), .o(n24849) );
no03f01 g21059 ( .a(n24811), .b(n24806), .c(n24805), .o(n24850) );
ao12f01 g21060 ( .a(n24850), .b(n24849), .c(n24812), .o(n24851) );
na02f01 g21061 ( .a(n24620), .b(n23945), .o(n24852) );
na02f01 g21062 ( .a(n24674), .b(n23953), .o(n24853) );
in01f01 g21063 ( .a(n24802), .o(n24854) );
ao12f01 g21064 ( .a(n24854), .b(n24853), .c(n24852), .o(n24855) );
oa12f01 g21065 ( .a(n24804), .b(n24855), .c(n24851), .o(n24856) );
oa12f01 g21066 ( .a(n24794), .b(n24788), .c(n24787), .o(n24857) );
ao12f01 g21067 ( .a(n24795), .b(n24857), .c(n24856), .o(n24858) );
na03f01 g21068 ( .a(n24785), .b(n24778), .c(n24777), .o(n24859) );
ao12f01 g21069 ( .a(n24786), .b(n24859), .c(n24858), .o(n24860) );
no02f01 g21070 ( .a(n24623), .b(n23871), .o(n24861) );
no02f01 g21071 ( .a(n24677), .b(n24153), .o(n24862) );
ao12f01 g21072 ( .a(n22965), .b(n23035), .c(n23032), .o(n24863) );
in01f01 g21073 ( .a(n24863), .o(n24864) );
no02f01 g21074 ( .a(n23034), .b(n22956), .o(n24865) );
no02f01 g21075 ( .a(n24865), .b(n24864), .o(n24866) );
na02f01 g21076 ( .a(n24865), .b(n24864), .o(n24867) );
in01f01 g21077 ( .a(n24867), .o(n24868) );
no02f01 g21078 ( .a(n24868), .b(n24866), .o(n24869) );
oa12f01 g21079 ( .a(n24869), .b(n24862), .c(n24861), .o(n24870) );
no03f01 g21080 ( .a(n24869), .b(n24862), .c(n24861), .o(n24871) );
ao12f01 g21081 ( .a(n24871), .b(n24870), .c(n24860), .o(n24872) );
oa12f01 g21082 ( .a(n24772), .b(n24872), .c(n24776), .o(n24873) );
ao12f01 g21083 ( .a(n24762), .b(n24873), .c(n24763), .o(n24874) );
oa12f01 g21084 ( .a(n24750), .b(n24874), .c(n24751), .o(n24875) );
no03f01 g21085 ( .a(n24746), .b(n24743), .c(n23237), .o(n24876) );
oa12f01 g21086 ( .a(n24747), .b(n24876), .c(n24875), .o(n24877) );
no02f01 g21087 ( .a(n24631), .b(n24629), .o(n24878) );
na03f01 g21088 ( .a(n24878), .b(n24682), .c(n24173), .o(n24879) );
na02f01 g21089 ( .a(n24685), .b(n24683), .o(n24880) );
oa12f01 g21090 ( .a(n24637), .b(n24880), .c(n24628), .o(n24881) );
ao12f01 g21091 ( .a(n23226), .b(n24881), .c(n24879), .o(n24882) );
no02f01 g21092 ( .a(n24882), .b(n24877), .o(n24883) );
na03f01 g21093 ( .a(n24881), .b(n24879), .c(n23226), .o(n24884) );
na02f01 g21094 ( .a(n24884), .b(n23221), .o(n24885) );
oa12f01 g21095 ( .a(n24740), .b(n24885), .c(n24883), .o(n24886) );
no03f01 g21096 ( .a(n24880), .b(n24628), .c(n24637), .o(n24887) );
ao12f01 g21097 ( .a(n24173), .b(n24878), .c(n24682), .o(n24888) );
no03f01 g21098 ( .a(n24888), .b(n24887), .c(n23903), .o(n24889) );
oa12f01 g21099 ( .a(n23901), .b(n24889), .c(n24883), .o(n24890) );
na03f01 g21100 ( .a(n24690), .b(n24688), .c(n24202), .o(n24891) );
oa12f01 g21101 ( .a(n24203), .b(n24639), .c(n24636), .o(n24892) );
na02f01 g21102 ( .a(n24892), .b(n24891), .o(n24893) );
ao22f01 g21103 ( .a(n24893), .b(n23913), .c(n24890), .d(n24886), .o(n24894) );
no02f01 g21104 ( .a(n24893), .b(n23913), .o(n24895) );
no03f01 g21105 ( .a(n24733), .b(n24616), .c(n24387), .o(n24896) );
ao12f01 g21106 ( .a(n24197), .b(n24727), .c(n24668), .o(n24897) );
no03f01 g21107 ( .a(n24897), .b(n24896), .c(n23898), .o(n24898) );
no03f01 g21108 ( .a(n24898), .b(n24895), .c(n24894), .o(n24899) );
na03f01 g21109 ( .a(n24693), .b(n24692), .c(n24262), .o(n24900) );
oa12f01 g21110 ( .a(n24213), .b(n24642), .c(n24641), .o(n24901) );
ao12f01 g21111 ( .a(n23252), .b(n24901), .c(n24900), .o(n24902) );
no03f01 g21112 ( .a(n24902), .b(n24899), .c(n24735), .o(n24903) );
oa12f01 g21113 ( .a(n23258), .b(n24719), .c(n24718), .o(n24904) );
oa12f01 g21114 ( .a(n24904), .b(n24903), .c(n24724), .o(n24905) );
oa12f01 g21115 ( .a(n24244), .b(n24648), .c(n24644), .o(n24906) );
na03f01 g21116 ( .a(n24699), .b(n24695), .c(n24243), .o(n24907) );
ao12f01 g21117 ( .a(n23265), .b(n24907), .c(n24906), .o(n24908) );
ao12f01 g21118 ( .a(n24908), .b(n24905), .c(n24721), .o(n24909) );
ao12f01 g21119 ( .a(n24710), .b(n24649), .c(n24645), .o(n24910) );
no03f01 g21120 ( .a(n24708), .b(n24700), .c(n24696), .o(n24911) );
oa12f01 g21121 ( .a(n23273), .b(n24911), .c(n24910), .o(n24912) );
oa12f01 g21122 ( .a(n24912), .b(n24909), .c(n24715), .o(n24913) );
na02f01 g21123 ( .a(n24705), .b(n24253), .o(n24914) );
na02f01 g21124 ( .a(n24703), .b(n24254), .o(n24915) );
ao12f01 g21125 ( .a(n23281), .b(n24915), .c(n24914), .o(n24916) );
ao12f01 g21126 ( .a(n24916), .b(n24913), .c(n24712), .o(n24917) );
in01f01 g21127 ( .a(n24665), .o(n24918) );
ao12f01 g21128 ( .a(n23739), .b(n24654), .c(n24652), .o(n24919) );
oa12f01 g21129 ( .a(n23288), .b(n24919), .c(n24918), .o(n24920) );
oa12f01 g21130 ( .a(n24920), .b(n24917), .c(n24707), .o(n24921) );
na02f01 g21131 ( .a(n24921), .b(n24667), .o(n24922) );
ao12f01 g21132 ( .a(n24660), .b(n24922), .c(n23892), .o(n24923) );
in01f01 g21133 ( .a(n24614), .o(n24924) );
ao22f01 g21134 ( .a(n24702), .b(n24698), .c(n24254), .d(n5119), .o(n24925) );
oa22f01 g21135 ( .a(n24653), .b(n24925), .c(n23739), .d(n5142), .o(n24926) );
na03f01 g21136 ( .a(n24926), .b(n24924), .c(n23739), .o(n24927) );
in01f01 g21137 ( .a(n24659), .o(n24928) );
na03f01 g21138 ( .a(n24928), .b(n24927), .c(n23891), .o(n24929) );
na04f01 g21139 ( .a(n24929), .b(n24921), .c(n24667), .d(n23307), .o(n24930) );
oa12f01 g21140 ( .a(n23191), .b(n24659), .c(n24656), .o(n24931) );
na02f01 g21141 ( .a(n24931), .b(n24930), .o(n24932) );
no02f01 g21142 ( .a(n24932), .b(n24923), .o(n24933) );
in01f01 g21143 ( .a(n24933), .o(n24934) );
no02f01 g21144 ( .a(n24660), .b(n23852), .o(n24935) );
in01f01 g21145 ( .a(n24935), .o(n24936) );
ao12f01 g21146 ( .a(n24660), .b(n23207), .c(n23186), .o(n24937) );
no02f01 g21147 ( .a(n24660), .b(n23859), .o(n24938) );
no02f01 g21148 ( .a(n24938), .b(n24937), .o(n24939) );
na02f01 g21149 ( .a(n24939), .b(n24936), .o(n24940) );
oa12f01 g21150 ( .a(n24664), .b(n24940), .c(n24934), .o(n24941) );
in01f01 g21151 ( .a(n23345), .o(n24942) );
ao12f01 g21152 ( .a(n24660), .b(n24942), .c(n23843), .o(n24943) );
in01f01 g21153 ( .a(n24943), .o(n24944) );
no02f01 g21154 ( .a(n24942), .b(n23843), .o(n24945) );
no02f01 g21155 ( .a(n24945), .b(n24661), .o(n24946) );
ao12f01 g21156 ( .a(n24946), .b(n24944), .c(n24941), .o(n24947) );
in01f01 g21157 ( .a(n24947), .o(n24948) );
in01f01 g21158 ( .a(n23159), .o(n24949) );
no02f01 g21159 ( .a(n24660), .b(n24949), .o(n24950) );
no02f01 g21160 ( .a(n24661), .b(n23159), .o(n24951) );
no02f01 g21161 ( .a(n24951), .b(n24950), .o(n24952) );
in01f01 g21162 ( .a(n24952), .o(n24953) );
no02f01 g21163 ( .a(n24953), .b(n24948), .o(n24954) );
no02f01 g21164 ( .a(n24952), .b(n24947), .o(n24955) );
no02f01 g21165 ( .a(n24955), .b(n24954), .o(n24956) );
in01f01 g21166 ( .a(n24956), .o(n24957) );
no02f01 g21167 ( .a(n24957), .b(n24613), .o(n24958) );
in01f01 g21168 ( .a(n24274), .o(n24959) );
no02f01 g21169 ( .a(n24608), .b(n5527), .o(n24960) );
na03f01 g21170 ( .a(n24398), .b(n24396), .c(n24390), .o(n24961) );
oa12f01 g21171 ( .a(n24391), .b(n24394), .c(n24392), .o(n24962) );
ao12f01 g21172 ( .a(n5529), .b(n24962), .c(n24961), .o(n24963) );
oa12f01 g21173 ( .a(n5529), .b(n24514), .c(n24513), .o(n24964) );
no02f01 g21174 ( .a(n24518), .b(n5527), .o(n24965) );
na02f01 g21175 ( .a(n24486), .b(n24478), .o(n24966) );
no02f01 g21176 ( .a(n24483), .b(n24482), .o(n24967) );
no02f01 g21177 ( .a(n24480), .b(n24479), .o(n24968) );
no02f01 g21178 ( .a(n24968), .b(n24967), .o(n24969) );
no02f01 g21179 ( .a(n24969), .b(n5529), .o(n24970) );
no02f01 g21180 ( .a(n24442), .b(n5529), .o(n24971) );
no02f01 g21181 ( .a(n24971), .b(n24970), .o(n24972) );
na02f01 g21182 ( .a(n24972), .b(n24966), .o(n24973) );
in01f01 g21183 ( .a(n24494), .o(n24974) );
ao12f01 g21184 ( .a(n24432), .b(n24974), .c(n24973), .o(n24975) );
na02f01 g21185 ( .a(n24425), .b(n24421), .o(n24976) );
na02f01 g21186 ( .a(n24423), .b(n24422), .o(n24977) );
na02f01 g21187 ( .a(n24977), .b(n24976), .o(n24978) );
na02f01 g21188 ( .a(n24978), .b(n5527), .o(n24979) );
ao12f01 g21189 ( .a(n24428), .b(n24979), .c(n24975), .o(n24980) );
na02f01 g21190 ( .a(n24502), .b(n24501), .o(n24981) );
na02f01 g21191 ( .a(n24499), .b(n24498), .o(n24982) );
na02f01 g21192 ( .a(n24982), .b(n24981), .o(n24983) );
na02f01 g21193 ( .a(n24983), .b(n5529), .o(n24984) );
na02f01 g21194 ( .a(n24984), .b(n24980), .o(n24985) );
no02f01 g21195 ( .a(n24985), .b(n24965), .o(n24986) );
na02f01 g21196 ( .a(n24986), .b(n24964), .o(n24987) );
ao12f01 g21197 ( .a(n24987), .b(n24512), .c(n5529), .o(n24988) );
ao12f01 g21198 ( .a(n5529), .b(n24411), .c(n24408), .o(n24989) );
na02f01 g21199 ( .a(n24419), .b(n5527), .o(n24990) );
na02f01 g21200 ( .a(n24983), .b(n5527), .o(n24991) );
na02f01 g21201 ( .a(n24991), .b(n24990), .o(n24992) );
no02f01 g21202 ( .a(n24992), .b(n24989), .o(n24993) );
oa12f01 g21203 ( .a(n24993), .b(n24405), .c(n5529), .o(n24994) );
oa22f01 g21204 ( .a(n24547), .b(n5527), .c(n24994), .d(n24988), .o(n24995) );
ao12f01 g21205 ( .a(n24995), .b(n24538), .c(n5529), .o(n24996) );
na02f01 g21206 ( .a(n24532), .b(n5527), .o(n24997) );
oa12f01 g21207 ( .a(n24997), .b(n24543), .c(n5529), .o(n24998) );
na03f01 g21208 ( .a(n24553), .b(n24557), .c(n24556), .o(n24999) );
oa12f01 g21209 ( .a(n24554), .b(n24551), .c(n24550), .o(n25000) );
ao12f01 g21210 ( .a(n5529), .b(n25000), .c(n24999), .o(n25001) );
no04f01 g21211 ( .a(n25001), .b(n24998), .c(n24996), .d(n24963), .o(n25002) );
na02f01 g21212 ( .a(n25000), .b(n24999), .o(n25003) );
na02f01 g21213 ( .a(n25003), .b(n5529), .o(n25004) );
na02f01 g21214 ( .a(n24962), .b(n24961), .o(n25005) );
na02f01 g21215 ( .a(n25005), .b(n5529), .o(n25006) );
na02f01 g21216 ( .a(n25006), .b(n25004), .o(n25007) );
no02f01 g21217 ( .a(n25007), .b(n25002), .o(n25008) );
ao12f01 g21218 ( .a(n5527), .b(n24596), .c(n24595), .o(n25009) );
oa12f01 g21219 ( .a(n24580), .b(n24585), .c(n24214), .o(n25010) );
na03f01 g21220 ( .a(n24583), .b(n24581), .c(n24578), .o(n25011) );
ao12f01 g21221 ( .a(n5527), .b(n25011), .c(n25010), .o(n25012) );
no02f01 g21222 ( .a(n24602), .b(n5527), .o(n25013) );
no03f01 g21223 ( .a(n25013), .b(n25012), .c(n25009), .o(n25014) );
oa12f01 g21224 ( .a(n5527), .b(n24576), .c(n24571), .o(n25015) );
na02f01 g21225 ( .a(n25011), .b(n25010), .o(n25016) );
na02f01 g21226 ( .a(n25016), .b(n5527), .o(n25017) );
na02f01 g21227 ( .a(n24592), .b(n5527), .o(n25018) );
na03f01 g21228 ( .a(n25018), .b(n25017), .c(n25015), .o(n25019) );
ao12f01 g21229 ( .a(n25019), .b(n25014), .c(n25008), .o(n25020) );
na02f01 g21230 ( .a(n24383), .b(n5527), .o(n25021) );
ao12f01 g21231 ( .a(n24960), .b(n25021), .c(n25020), .o(n25022) );
oa12f01 g21232 ( .a(n24959), .b(n24611), .c(n25022), .o(n25023) );
no02f01 g21233 ( .a(n24956), .b(n25023), .o(n25024) );
no02f01 g21234 ( .a(n25024), .b(n24958), .o(n25025) );
in01f01 g21235 ( .a(n25025), .o(n25026) );
no02f01 g21236 ( .a(n24660), .b(n23843), .o(n25027) );
no02f01 g21237 ( .a(n24661), .b(n23329), .o(n25028) );
no02f01 g21238 ( .a(n25028), .b(n25027), .o(n25029) );
in01f01 g21239 ( .a(n25029), .o(n25030) );
na02f01 g21240 ( .a(n25030), .b(n24941), .o(n25031) );
in01f01 g21241 ( .a(n24941), .o(n25032) );
na02f01 g21242 ( .a(n25029), .b(n25032), .o(n25033) );
na02f01 g21243 ( .a(n25033), .b(n25031), .o(n25034) );
no02f01 g21244 ( .a(n25034), .b(n24613), .o(n25035) );
in01f01 g21245 ( .a(n25027), .o(n25036) );
ao12f01 g21246 ( .a(n25028), .b(n25036), .c(n24941), .o(n25037) );
no02f01 g21247 ( .a(n24661), .b(n23345), .o(n25038) );
no02f01 g21248 ( .a(n24660), .b(n24942), .o(n25039) );
no02f01 g21249 ( .a(n25039), .b(n25038), .o(n25040) );
na02f01 g21250 ( .a(n25040), .b(n25037), .o(n25041) );
in01f01 g21251 ( .a(n25041), .o(n25042) );
no02f01 g21252 ( .a(n25040), .b(n25037), .o(n25043) );
no02f01 g21253 ( .a(n25043), .b(n25042), .o(n25044) );
in01f01 g21254 ( .a(n25044), .o(n25045) );
no02f01 g21255 ( .a(n25045), .b(n24613), .o(n25046) );
no02f01 g21256 ( .a(n25046), .b(n25035), .o(n25047) );
no02f01 g21257 ( .a(n24661), .b(n23310), .o(n25048) );
no02f01 g21258 ( .a(n24660), .b(n23207), .o(n25049) );
no02f01 g21259 ( .a(n25049), .b(n25048), .o(n25050) );
no03f01 g21260 ( .a(n25050), .b(n24932), .c(n24923), .o(n25051) );
no03f01 g21261 ( .a(n24919), .b(n24918), .c(n23288), .o(n25052) );
na03f01 g21262 ( .a(n24915), .b(n24914), .c(n23281), .o(n25053) );
no03f01 g21263 ( .a(n24911), .b(n24910), .c(n23273), .o(n25054) );
na03f01 g21264 ( .a(n24907), .b(n24906), .c(n23265), .o(n25055) );
na03f01 g21265 ( .a(n24901), .b(n24900), .c(n23252), .o(n25056) );
oa12f01 g21266 ( .a(n23898), .b(n24897), .c(n24896), .o(n25057) );
na03f01 g21267 ( .a(n24638), .b(n24738), .c(n24179), .o(n25058) );
oa12f01 g21268 ( .a(n23801), .b(n24689), .c(n24736), .o(n25059) );
na02f01 g21269 ( .a(n25059), .b(n25058), .o(n25060) );
na03f01 g21270 ( .a(n24745), .b(n24744), .c(n23813), .o(n25061) );
oa12f01 g21271 ( .a(n23806), .b(n24742), .c(n24741), .o(n25062) );
ao12f01 g21272 ( .a(n23908), .b(n25062), .c(n25061), .o(n25063) );
no03f01 g21273 ( .a(n24684), .b(n24680), .c(n24163), .o(n25064) );
ao12f01 g21274 ( .a(n23820), .b(n24630), .c(n24626), .o(n25065) );
no03f01 g21275 ( .a(n25065), .b(n25064), .c(n23905), .o(n25066) );
oa12f01 g21276 ( .a(n23905), .b(n25065), .c(n25064), .o(n25067) );
na02f01 g21277 ( .a(n24755), .b(n24282), .o(n25068) );
na02f01 g21278 ( .a(n24752), .b(n23833), .o(n25069) );
in01f01 g21279 ( .a(n24761), .o(n25070) );
na03f01 g21280 ( .a(n25070), .b(n25069), .c(n25068), .o(n25071) );
ao12f01 g21281 ( .a(n25070), .b(n25069), .c(n25068), .o(n25072) );
oa12f01 g21282 ( .a(n24770), .b(n24765), .c(n24764), .o(n25073) );
in01f01 g21283 ( .a(n24786), .o(n25074) );
in01f01 g21284 ( .a(n24795), .o(n25075) );
na02f01 g21285 ( .a(n24619), .b(n23961), .o(n25076) );
na02f01 g21286 ( .a(n24673), .b(n24136), .o(n25077) );
in01f01 g21287 ( .a(n24811), .o(n25078) );
ao12f01 g21288 ( .a(n25078), .b(n25077), .c(n25076), .o(n25079) );
oa12f01 g21289 ( .a(n24820), .b(n24814), .c(n24813), .o(n25080) );
na02f01 g21290 ( .a(n24617), .b(n24124), .o(n25081) );
na02f01 g21291 ( .a(n24843), .b(n24348), .o(n25082) );
na02f01 g21292 ( .a(n25082), .b(n25081), .o(n25083) );
in01f01 g21293 ( .a(n24847), .o(n25084) );
oa12f01 g21294 ( .a(n25084), .b(n25083), .c(n24841), .o(n25085) );
ao12f01 g21295 ( .a(n24821), .b(n25085), .c(n25080), .o(n25086) );
in01f01 g21296 ( .a(n24850), .o(n25087) );
oa12f01 g21297 ( .a(n25087), .b(n25086), .c(n25079), .o(n25088) );
oa12f01 g21298 ( .a(n24802), .b(n24797), .c(n24796), .o(n25089) );
ao12f01 g21299 ( .a(n24803), .b(n25089), .c(n25088), .o(n25090) );
na02f01 g21300 ( .a(n24675), .b(n23939), .o(n25091) );
na02f01 g21301 ( .a(n24621), .b(n23933), .o(n25092) );
in01f01 g21302 ( .a(n24794), .o(n25093) );
ao12f01 g21303 ( .a(n25093), .b(n25092), .c(n25091), .o(n25094) );
oa12f01 g21304 ( .a(n25075), .b(n25094), .c(n25090), .o(n25095) );
no02f01 g21305 ( .a(n24676), .b(n24146), .o(n25096) );
no02f01 g21306 ( .a(n24622), .b(n23880), .o(n25097) );
no03f01 g21307 ( .a(n24784), .b(n25097), .c(n25096), .o(n25098) );
oa12f01 g21308 ( .a(n25074), .b(n25098), .c(n25095), .o(n25099) );
na02f01 g21309 ( .a(n24677), .b(n24153), .o(n25100) );
na02f01 g21310 ( .a(n24623), .b(n23871), .o(n25101) );
in01f01 g21311 ( .a(n24869), .o(n25102) );
ao12f01 g21312 ( .a(n25102), .b(n25101), .c(n25100), .o(n25103) );
in01f01 g21313 ( .a(n24871), .o(n25104) );
oa12f01 g21314 ( .a(n25104), .b(n25103), .c(n25099), .o(n25105) );
ao12f01 g21315 ( .a(n24771), .b(n25105), .c(n25073), .o(n25106) );
oa12f01 g21316 ( .a(n25071), .b(n25106), .c(n25072), .o(n25107) );
ao12f01 g21317 ( .a(n25066), .b(n25107), .c(n25067), .o(n25108) );
na03f01 g21318 ( .a(n25062), .b(n25061), .c(n23908), .o(n25109) );
ao12f01 g21319 ( .a(n25063), .b(n25109), .c(n25108), .o(n25110) );
oa12f01 g21320 ( .a(n23903), .b(n24888), .c(n24887), .o(n25111) );
na02f01 g21321 ( .a(n25111), .b(n25110), .o(n25112) );
no02f01 g21322 ( .a(n24889), .b(n23901), .o(n25113) );
ao12f01 g21323 ( .a(n25060), .b(n25113), .c(n25112), .o(n25114) );
ao12f01 g21324 ( .a(n23221), .b(n24884), .c(n25112), .o(n25115) );
no03f01 g21325 ( .a(n24639), .b(n24636), .c(n24203), .o(n25116) );
ao12f01 g21326 ( .a(n24202), .b(n24690), .c(n24688), .o(n25117) );
no02f01 g21327 ( .a(n25117), .b(n25116), .o(n25118) );
oa22f01 g21328 ( .a(n25118), .b(n23245), .c(n25115), .d(n25114), .o(n25119) );
na02f01 g21329 ( .a(n25118), .b(n23245), .o(n25120) );
na03f01 g21330 ( .a(n24734), .b(n24728), .c(n23215), .o(n25121) );
na03f01 g21331 ( .a(n25121), .b(n25120), .c(n25119), .o(n25122) );
oa12f01 g21332 ( .a(n23917), .b(n24723), .c(n24722), .o(n25123) );
na03f01 g21333 ( .a(n25123), .b(n25122), .c(n25057), .o(n25124) );
na03f01 g21334 ( .a(n24716), .b(n24643), .c(n24221), .o(n25125) );
oa12f01 g21335 ( .a(n24222), .b(n24717), .c(n24694), .o(n25126) );
ao12f01 g21336 ( .a(n23920), .b(n25126), .c(n25125), .o(n25127) );
ao12f01 g21337 ( .a(n25127), .b(n25124), .c(n25056), .o(n25128) );
oa12f01 g21338 ( .a(n23297), .b(n24714), .c(n24713), .o(n25129) );
oa12f01 g21339 ( .a(n25129), .b(n25128), .c(n24720), .o(n25130) );
ao12f01 g21340 ( .a(n23295), .b(n24711), .c(n24709), .o(n25131) );
ao12f01 g21341 ( .a(n25131), .b(n25130), .c(n25055), .o(n25132) );
oa12f01 g21342 ( .a(n23293), .b(n24706), .c(n24704), .o(n25133) );
oa12f01 g21343 ( .a(n25133), .b(n25132), .c(n25054), .o(n25134) );
ao12f01 g21344 ( .a(n23291), .b(n24666), .c(n24665), .o(n25135) );
ao12f01 g21345 ( .a(n25135), .b(n25134), .c(n25053), .o(n25136) );
no02f01 g21346 ( .a(n25136), .b(n25052), .o(n25137) );
oa12f01 g21347 ( .a(n24661), .b(n25137), .c(n23307), .o(n25138) );
no03f01 g21348 ( .a(n24659), .b(n24656), .c(n23191), .o(n25139) );
no04f01 g21349 ( .a(n25139), .b(n25136), .c(n25052), .d(n23892), .o(n25140) );
ao12f01 g21350 ( .a(n23891), .b(n24928), .c(n24927), .o(n25141) );
no02f01 g21351 ( .a(n25141), .b(n25140), .o(n25142) );
in01f01 g21352 ( .a(n25050), .o(n25143) );
ao12f01 g21353 ( .a(n25143), .b(n25142), .c(n25138), .o(n25144) );
no02f01 g21354 ( .a(n25144), .b(n25051), .o(n25145) );
na02f01 g21355 ( .a(n25145), .b(n25023), .o(n25146) );
no02f01 g21356 ( .a(n24660), .b(n23186), .o(n25147) );
no02f01 g21357 ( .a(n24661), .b(n23305), .o(n25148) );
no02f01 g21358 ( .a(n25148), .b(n25147), .o(n25149) );
in01f01 g21359 ( .a(n25149), .o(n25150) );
no03f01 g21360 ( .a(n25049), .b(n24932), .c(n24923), .o(n25151) );
no03f01 g21361 ( .a(n25151), .b(n25150), .c(n25048), .o(n25152) );
in01f01 g21362 ( .a(n25048), .o(n25153) );
in01f01 g21363 ( .a(n25049), .o(n25154) );
na03f01 g21364 ( .a(n25154), .b(n25142), .c(n25138), .o(n25155) );
ao12f01 g21365 ( .a(n25149), .b(n25155), .c(n25153), .o(n25156) );
no02f01 g21366 ( .a(n25156), .b(n25152), .o(n25157) );
na02f01 g21367 ( .a(n25157), .b(n25023), .o(n25158) );
na02f01 g21368 ( .a(n25158), .b(n25146), .o(n25159) );
no02f01 g21369 ( .a(n24661), .b(n23321), .o(n25160) );
no02f01 g21370 ( .a(n25160), .b(n24938), .o(n25161) );
in01f01 g21371 ( .a(n25161), .o(n25162) );
no02f01 g21372 ( .a(n24661), .b(n23170), .o(n25163) );
no03f01 g21373 ( .a(n24937), .b(n24932), .c(n24923), .o(n25164) );
no03f01 g21374 ( .a(n25164), .b(n24663), .c(n25163), .o(n25165) );
no02f01 g21375 ( .a(n25165), .b(n24935), .o(n25166) );
no02f01 g21376 ( .a(n25166), .b(n25162), .o(n25167) );
in01f01 g21377 ( .a(n25167), .o(n25168) );
na02f01 g21378 ( .a(n25166), .b(n25162), .o(n25169) );
na02f01 g21379 ( .a(n25169), .b(n25168), .o(n25170) );
no02f01 g21380 ( .a(n25170), .b(n24613), .o(n25171) );
in01f01 g21381 ( .a(n24663), .o(n25172) );
in01f01 g21382 ( .a(n24937), .o(n25173) );
na03f01 g21383 ( .a(n25173), .b(n25142), .c(n25138), .o(n25174) );
no02f01 g21384 ( .a(n24935), .b(n25163), .o(n25175) );
ao12f01 g21385 ( .a(n25175), .b(n25174), .c(n25172), .o(n25176) );
in01f01 g21386 ( .a(n25175), .o(n25177) );
no03f01 g21387 ( .a(n25177), .b(n25164), .c(n24663), .o(n25178) );
no02f01 g21388 ( .a(n25178), .b(n25176), .o(n25179) );
na02f01 g21389 ( .a(n25179), .b(n25023), .o(n25180) );
in01f01 g21390 ( .a(n25180), .o(n25181) );
no03f01 g21391 ( .a(n25181), .b(n25171), .c(n25159), .o(n25182) );
in01f01 g21392 ( .a(n25182), .o(n25183) );
na02f01 g21393 ( .a(n24920), .b(n24667), .o(n25184) );
no03f01 g21394 ( .a(n25184), .b(n24917), .c(n24707), .o(n25185) );
no02f01 g21395 ( .a(n25135), .b(n25052), .o(n25186) );
ao12f01 g21396 ( .a(n25186), .b(n25134), .c(n25053), .o(n25187) );
no02f01 g21397 ( .a(n25187), .b(n25185), .o(n25188) );
na02f01 g21398 ( .a(n25188), .b(n25023), .o(n25189) );
no02f01 g21399 ( .a(n24611), .b(n24274), .o(n25190) );
no02f01 g21400 ( .a(n25190), .b(n24610), .o(n25191) );
in01f01 g21401 ( .a(n25190), .o(n25192) );
no02f01 g21402 ( .a(n25192), .b(n25022), .o(n25193) );
na02f01 g21403 ( .a(n24913), .b(n24712), .o(n25194) );
na02f01 g21404 ( .a(n25133), .b(n25053), .o(n25195) );
no02f01 g21405 ( .a(n25195), .b(n25194), .o(n25196) );
no02f01 g21406 ( .a(n25132), .b(n25054), .o(n25197) );
no02f01 g21407 ( .a(n24916), .b(n24707), .o(n25198) );
no02f01 g21408 ( .a(n25198), .b(n25197), .o(n25199) );
no02f01 g21409 ( .a(n25199), .b(n25196), .o(n25200) );
oa12f01 g21410 ( .a(n25200), .b(n25193), .c(n25191), .o(n25201) );
na03f01 g21411 ( .a(n24929), .b(n24921), .c(n24667), .o(n25202) );
na02f01 g21412 ( .a(n24660), .b(n23892), .o(n25203) );
no02f01 g21413 ( .a(n24660), .b(n23892), .o(n25204) );
in01f01 g21414 ( .a(n25204), .o(n25205) );
na02f01 g21415 ( .a(n25205), .b(n25203), .o(n25206) );
ao12f01 g21416 ( .a(n25206), .b(n24931), .c(n25202), .o(n25207) );
no03f01 g21417 ( .a(n25139), .b(n25136), .c(n25052), .o(n25208) );
in01f01 g21418 ( .a(n25203), .o(n25209) );
no02f01 g21419 ( .a(n25204), .b(n25209), .o(n25210) );
no03f01 g21420 ( .a(n25210), .b(n25141), .c(n25208), .o(n25211) );
no02f01 g21421 ( .a(n25211), .b(n25207), .o(n25212) );
no02f01 g21422 ( .a(n25141), .b(n25139), .o(n25213) );
ao12f01 g21423 ( .a(n25213), .b(n24921), .c(n24667), .o(n25214) );
na02f01 g21424 ( .a(n24931), .b(n24929), .o(n25215) );
no03f01 g21425 ( .a(n25215), .b(n25136), .c(n25052), .o(n25216) );
no02f01 g21426 ( .a(n25216), .b(n25214), .o(n25217) );
oa12f01 g21427 ( .a(n25023), .b(n25217), .c(n25212), .o(n25218) );
na03f01 g21428 ( .a(n25218), .b(n25201), .c(n25189), .o(n25219) );
no02f01 g21429 ( .a(n24609), .b(n24960), .o(n25220) );
na02f01 g21430 ( .a(n25220), .b(n25020), .o(n25221) );
na02f01 g21431 ( .a(n25021), .b(n24384), .o(n25222) );
na02f01 g21432 ( .a(n25222), .b(n24605), .o(n25223) );
na02f01 g21433 ( .a(n24912), .b(n24712), .o(n25224) );
no03f01 g21434 ( .a(n25224), .b(n24909), .c(n24715), .o(n25225) );
no02f01 g21435 ( .a(n25131), .b(n25054), .o(n25226) );
ao12f01 g21436 ( .a(n25226), .b(n25130), .c(n25055), .o(n25227) );
no02f01 g21437 ( .a(n25227), .b(n25225), .o(n25228) );
in01f01 g21438 ( .a(n25228), .o(n25229) );
ao12f01 g21439 ( .a(n25229), .b(n25223), .c(n25221), .o(n25230) );
in01f01 g21440 ( .a(n25230), .o(n25231) );
no02f01 g21441 ( .a(n24603), .b(n24599), .o(n25232) );
no02f01 g21442 ( .a(n24597), .b(n25009), .o(n25233) );
no03f01 g21443 ( .a(n25012), .b(n25007), .c(n25002), .o(n25234) );
na02f01 g21444 ( .a(n25234), .b(n24593), .o(n25235) );
na03f01 g21445 ( .a(n25235), .b(n25233), .c(n25232), .o(n25236) );
in01f01 g21446 ( .a(n25232), .o(n25237) );
in01f01 g21447 ( .a(n25233), .o(n25238) );
na03f01 g21448 ( .a(n24587), .b(n24565), .c(n24560), .o(n25239) );
no02f01 g21449 ( .a(n25239), .b(n25013), .o(n25240) );
oa12f01 g21450 ( .a(n25238), .b(n25240), .c(n25237), .o(n25241) );
na02f01 g21451 ( .a(n24905), .b(n24721), .o(n25242) );
na02f01 g21452 ( .a(n25129), .b(n25055), .o(n25243) );
no02f01 g21453 ( .a(n25243), .b(n25242), .o(n25244) );
no02f01 g21454 ( .a(n25128), .b(n24720), .o(n25245) );
no02f01 g21455 ( .a(n24908), .b(n24715), .o(n25246) );
no02f01 g21456 ( .a(n25246), .b(n25245), .o(n25247) );
no02f01 g21457 ( .a(n25247), .b(n25244), .o(n25248) );
in01f01 g21458 ( .a(n25248), .o(n25249) );
ao12f01 g21459 ( .a(n25249), .b(n25241), .c(n25236), .o(n25250) );
na02f01 g21460 ( .a(n25124), .b(n25056), .o(n25251) );
no03f01 g21461 ( .a(n25127), .b(n25251), .c(n24720), .o(n25252) );
no02f01 g21462 ( .a(n24903), .b(n24724), .o(n25253) );
ao12f01 g21463 ( .a(n25253), .b(n24904), .c(n24721), .o(n25254) );
no02f01 g21464 ( .a(n25254), .b(n25252), .o(n25255) );
in01f01 g21465 ( .a(n25255), .o(n25256) );
no02f01 g21466 ( .a(n24603), .b(n25013), .o(n25257) );
na03f01 g21467 ( .a(n25257), .b(n25239), .c(n25017), .o(n25258) );
in01f01 g21468 ( .a(n25257), .o(n25259) );
oa12f01 g21469 ( .a(n25259), .b(n25234), .c(n24599), .o(n25260) );
ao12f01 g21470 ( .a(n25256), .b(n25260), .c(n25258), .o(n25261) );
no03f01 g21471 ( .a(n25259), .b(n25234), .c(n24599), .o(n25262) );
ao12f01 g21472 ( .a(n25257), .b(n25239), .c(n25017), .o(n25263) );
no03f01 g21473 ( .a(n25263), .b(n25262), .c(n25255), .o(n25264) );
na02f01 g21474 ( .a(n25017), .b(n24587), .o(n25265) );
na02f01 g21475 ( .a(n25265), .b(n25008), .o(n25266) );
no02f01 g21476 ( .a(n24599), .b(n25012), .o(n25267) );
na02f01 g21477 ( .a(n25267), .b(n24566), .o(n25268) );
na02f01 g21478 ( .a(n25268), .b(n25266), .o(n25269) );
no02f01 g21479 ( .a(n24899), .b(n24735), .o(n25270) );
na02f01 g21480 ( .a(n25123), .b(n25056), .o(n25271) );
no02f01 g21481 ( .a(n25271), .b(n25270), .o(n25272) );
na02f01 g21482 ( .a(n25122), .b(n25057), .o(n25273) );
no02f01 g21483 ( .a(n24902), .b(n24724), .o(n25274) );
no02f01 g21484 ( .a(n25274), .b(n25273), .o(n25275) );
no02f01 g21485 ( .a(n25275), .b(n25272), .o(n25276) );
no02f01 g21486 ( .a(n25276), .b(n25269), .o(n25277) );
no02f01 g21487 ( .a(n25277), .b(n25264), .o(n25278) );
no03f01 g21488 ( .a(n25278), .b(n25261), .c(n25250), .o(n25279) );
no03f01 g21489 ( .a(n25240), .b(n25238), .c(n25237), .o(n25280) );
ao12f01 g21490 ( .a(n25233), .b(n25235), .c(n25232), .o(n25281) );
no03f01 g21491 ( .a(n25248), .b(n25281), .c(n25280), .o(n25282) );
in01f01 g21492 ( .a(n25282), .o(n25283) );
na03f01 g21493 ( .a(n25229), .b(n25223), .c(n25221), .o(n25284) );
na02f01 g21494 ( .a(n25284), .b(n25283), .o(n25285) );
oa12f01 g21495 ( .a(n25231), .b(n25285), .c(n25279), .o(n25286) );
no02f01 g21496 ( .a(n25286), .b(n25219), .o(n25287) );
oa12f01 g21497 ( .a(n25210), .b(n25141), .c(n25208), .o(n25288) );
na03f01 g21498 ( .a(n25206), .b(n24931), .c(n25202), .o(n25289) );
na02f01 g21499 ( .a(n25289), .b(n25288), .o(n25290) );
oa12f01 g21500 ( .a(n25215), .b(n25136), .c(n25052), .o(n25291) );
na03f01 g21501 ( .a(n25213), .b(n24921), .c(n24667), .o(n25292) );
na02f01 g21502 ( .a(n25292), .b(n25291), .o(n25293) );
ao12f01 g21503 ( .a(n24613), .b(n25293), .c(n25290), .o(n25294) );
no02f01 g21504 ( .a(n25188), .b(n25023), .o(n25295) );
no03f01 g21505 ( .a(n25200), .b(n25193), .c(n25191), .o(n25296) );
oa12f01 g21506 ( .a(n25189), .b(n25296), .c(n25295), .o(n25297) );
ao12f01 g21507 ( .a(n25023), .b(n25217), .c(n25212), .o(n25298) );
in01f01 g21508 ( .a(n25298), .o(n25299) );
ao12f01 g21509 ( .a(n25294), .b(n25299), .c(n25297), .o(n25300) );
no02f01 g21510 ( .a(n25300), .b(n25287), .o(n25301) );
in01f01 g21511 ( .a(n25261), .o(n25302) );
no02f01 g21512 ( .a(n24998), .b(n24996), .o(n25303) );
ao12f01 g21513 ( .a(n24564), .b(n25303), .c(n24400), .o(n25304) );
no02f01 g21514 ( .a(n24562), .b(n25001), .o(n25305) );
in01f01 g21515 ( .a(n25305), .o(n25306) );
na02f01 g21516 ( .a(n25306), .b(n25304), .o(n25307) );
no02f01 g21517 ( .a(n25306), .b(n25304), .o(n25308) );
in01f01 g21518 ( .a(n25308), .o(n25309) );
na02f01 g21519 ( .a(n25121), .b(n25057), .o(n25310) );
no02f01 g21520 ( .a(n25115), .b(n25114), .o(n25311) );
no02f01 g21521 ( .a(n25118), .b(n23245), .o(n25312) );
ao12f01 g21522 ( .a(n25312), .b(n25120), .c(n25311), .o(n25313) );
no02f01 g21523 ( .a(n25313), .b(n25310), .o(n25314) );
no02f01 g21524 ( .a(n24898), .b(n24735), .o(n25315) );
na02f01 g21525 ( .a(n24890), .b(n24886), .o(n25316) );
na02f01 g21526 ( .a(n24893), .b(n23913), .o(n25317) );
oa12f01 g21527 ( .a(n25317), .b(n24895), .c(n25316), .o(n25318) );
no02f01 g21528 ( .a(n25318), .b(n25315), .o(n25319) );
no02f01 g21529 ( .a(n25319), .b(n25314), .o(n25320) );
in01f01 g21530 ( .a(n25320), .o(n25321) );
ao12f01 g21531 ( .a(n25321), .b(n25309), .c(n25307), .o(n25322) );
in01f01 g21532 ( .a(n24539), .o(n25323) );
no02f01 g21533 ( .a(n24544), .b(n25323), .o(n25324) );
no02f01 g21534 ( .a(n24548), .b(n24533), .o(n25325) );
no02f01 g21535 ( .a(n25325), .b(n25324), .o(n25326) );
no04f01 g21536 ( .a(n24548), .b(n24544), .c(n25323), .d(n24533), .o(n25327) );
no02f01 g21537 ( .a(n25327), .b(n25326), .o(n25328) );
na02f01 g21538 ( .a(n24512), .b(n5529), .o(n25329) );
na02f01 g21539 ( .a(n24512), .b(n5527), .o(n25330) );
na02f01 g21540 ( .a(n24521), .b(n24507), .o(n25331) );
na02f01 g21541 ( .a(n25331), .b(n24964), .o(n25332) );
ao22f01 g21542 ( .a(n25332), .b(n24515), .c(n25330), .d(n25329), .o(n25333) );
no02f01 g21543 ( .a(n24405), .b(n5527), .o(n25334) );
no02f01 g21544 ( .a(n24405), .b(n5529), .o(n25335) );
ao12f01 g21545 ( .a(n24412), .b(n24521), .c(n24507), .o(n25336) );
no04f01 g21546 ( .a(n25336), .b(n24989), .c(n25335), .d(n25334), .o(n25337) );
na02f01 g21547 ( .a(n25109), .b(n24747), .o(n25338) );
na02f01 g21548 ( .a(n25338), .b(n24875), .o(n25339) );
na03f01 g21549 ( .a(n25109), .b(n25108), .c(n24747), .o(n25340) );
na02f01 g21550 ( .a(n25340), .b(n25339), .o(n25341) );
in01f01 g21551 ( .a(n25341), .o(n25342) );
no03f01 g21552 ( .a(n25342), .b(n25337), .c(n25333), .o(n25343) );
in01f01 g21553 ( .a(n25343), .o(n25344) );
no02f01 g21554 ( .a(n24992), .b(n24986), .o(n25345) );
no02f01 g21555 ( .a(n24989), .b(n24412), .o(n25346) );
no02f01 g21556 ( .a(n25346), .b(n25345), .o(n25347) );
na02f01 g21557 ( .a(n24515), .b(n24964), .o(n25348) );
no02f01 g21558 ( .a(n25348), .b(n25331), .o(n25349) );
no02f01 g21559 ( .a(n24751), .b(n25066), .o(n25350) );
no02f01 g21560 ( .a(n25350), .b(n24874), .o(n25351) );
na02f01 g21561 ( .a(n25350), .b(n24874), .o(n25352) );
in01f01 g21562 ( .a(n25352), .o(n25353) );
no02f01 g21563 ( .a(n25353), .b(n25351), .o(n25354) );
no03f01 g21564 ( .a(n25354), .b(n25349), .c(n25347), .o(n25355) );
ao22f01 g21565 ( .a(n24991), .b(n24985), .c(n24990), .d(n24420), .o(n25356) );
no04f01 g21566 ( .a(n24520), .b(n24519), .c(n24506), .d(n24965), .o(n25357) );
no02f01 g21567 ( .a(n25072), .b(n24762), .o(n25358) );
no02f01 g21568 ( .a(n25358), .b(n25106), .o(n25359) );
na02f01 g21569 ( .a(n25358), .b(n25106), .o(n25360) );
in01f01 g21570 ( .a(n25360), .o(n25361) );
no02f01 g21571 ( .a(n25361), .b(n25359), .o(n25362) );
no03f01 g21572 ( .a(n25362), .b(n25357), .c(n25356), .o(n25363) );
in01f01 g21573 ( .a(n25363), .o(n25364) );
na02f01 g21574 ( .a(n24978), .b(n5529), .o(n25365) );
oa12f01 g21575 ( .a(n25365), .b(n24496), .c(n24495), .o(n25366) );
no02f01 g21576 ( .a(n24520), .b(n24505), .o(n25367) );
na02f01 g21577 ( .a(n25367), .b(n25366), .o(n25368) );
na02f01 g21578 ( .a(n24991), .b(n24984), .o(n25369) );
na02f01 g21579 ( .a(n25369), .b(n24980), .o(n25370) );
na02f01 g21580 ( .a(n25370), .b(n25368), .o(n25371) );
no02f01 g21581 ( .a(n24776), .b(n24771), .o(n25372) );
no02f01 g21582 ( .a(n25372), .b(n24872), .o(n25373) );
na02f01 g21583 ( .a(n25372), .b(n24872), .o(n25374) );
in01f01 g21584 ( .a(n25374), .o(n25375) );
no02f01 g21585 ( .a(n25375), .b(n25373), .o(n25376) );
no02f01 g21586 ( .a(n25376), .b(n25371), .o(n25377) );
ao12f01 g21587 ( .a(n24975), .b(n24979), .c(n25365), .o(n25378) );
no03f01 g21588 ( .a(n24496), .b(n24495), .c(n24428), .o(n25379) );
no02f01 g21589 ( .a(n25379), .b(n25378), .o(n25380) );
oa12f01 g21590 ( .a(n24491), .b(n24477), .c(n24443), .o(n25381) );
in01f01 g21591 ( .a(n25381), .o(n25382) );
ao12f01 g21592 ( .a(n25382), .b(n24487), .c(n24486), .o(n25383) );
no02f01 g21593 ( .a(n24969), .b(n5527), .o(n25384) );
no03f01 g21594 ( .a(n25381), .b(n24970), .c(n25384), .o(n25385) );
no02f01 g21595 ( .a(n25094), .b(n24795), .o(n25386) );
no02f01 g21596 ( .a(n25386), .b(n25090), .o(n25387) );
na02f01 g21597 ( .a(n25386), .b(n25090), .o(n25388) );
in01f01 g21598 ( .a(n25388), .o(n25389) );
no02f01 g21599 ( .a(n25389), .b(n25387), .o(n25390) );
no03f01 g21600 ( .a(n25390), .b(n25385), .c(n25383), .o(n25391) );
in01f01 g21601 ( .a(n24477), .o(n25392) );
oa12f01 g21602 ( .a(n25392), .b(n24971), .c(n24443), .o(n25393) );
na02f01 g21603 ( .a(n24490), .b(n5529), .o(n25394) );
na03f01 g21604 ( .a(n24491), .b(n24477), .c(n25394), .o(n25395) );
no02f01 g21605 ( .a(n24855), .b(n24803), .o(n25396) );
no02f01 g21606 ( .a(n25396), .b(n24851), .o(n25397) );
na02f01 g21607 ( .a(n25396), .b(n24851), .o(n25398) );
in01f01 g21608 ( .a(n25398), .o(n25399) );
no02f01 g21609 ( .a(n25399), .b(n25397), .o(n25400) );
in01f01 g21610 ( .a(n25400), .o(n25401) );
na03f01 g21611 ( .a(n25401), .b(n25395), .c(n25393), .o(n25402) );
in01f01 g21612 ( .a(n24476), .o(n25403) );
na02f01 g21613 ( .a(n24448), .b(n5527), .o(n25404) );
ao12f01 g21614 ( .a(n25403), .b(n25404), .c(n24449), .o(n25405) );
no02f01 g21615 ( .a(n24446), .b(n24439), .o(n25406) );
no02f01 g21616 ( .a(n24444), .b(n24435), .o(n25407) );
no02f01 g21617 ( .a(n25407), .b(n25406), .o(n25408) );
no02f01 g21618 ( .a(n25408), .b(n5527), .o(n25409) );
no02f01 g21619 ( .a(n25408), .b(n5529), .o(n25410) );
no03f01 g21620 ( .a(n25410), .b(n24476), .c(n25409), .o(n25411) );
no03f01 g21621 ( .a(n24850), .b(n24849), .c(n25079), .o(n25412) );
ao12f01 g21622 ( .a(n25086), .b(n25087), .c(n24812), .o(n25413) );
no02f01 g21623 ( .a(n25413), .b(n25412), .o(n25414) );
oa12f01 g21624 ( .a(n25414), .b(n25411), .c(n25405), .o(n25415) );
no02f01 g21625 ( .a(n24463), .b(n24345), .o(n25416) );
no02f01 g21626 ( .a(n24459), .b(n24119), .o(n25417) );
no02f01 g21627 ( .a(n25417), .b(n25416), .o(n25418) );
na02f01 g21628 ( .a(n25418), .b(n5529), .o(n25419) );
na02f01 g21629 ( .a(n25418), .b(n5527), .o(n25420) );
no02f01 g21630 ( .a(n24838), .b(n23990), .o(n25421) );
in01f01 g21631 ( .a(n24838), .o(n25422) );
no02f01 g21632 ( .a(n25422), .b(n24300), .o(n25423) );
no02f01 g21633 ( .a(n25423), .b(n25421), .o(n25424) );
in01f01 g21634 ( .a(n25424), .o(n25425) );
na03f01 g21635 ( .a(n25425), .b(n25420), .c(n25419), .o(n25426) );
no02f01 g21636 ( .a(n25083), .b(n24833), .o(n25427) );
no02f01 g21637 ( .a(n24846), .b(n24834), .o(n25428) );
no02f01 g21638 ( .a(n25428), .b(n25427), .o(n25429) );
no02f01 g21639 ( .a(n25429), .b(n24839), .o(n25430) );
na02f01 g21640 ( .a(n25429), .b(n24839), .o(n25431) );
in01f01 g21641 ( .a(n25431), .o(n25432) );
no02f01 g21642 ( .a(n25432), .b(n25430), .o(n25433) );
in01f01 g21643 ( .a(n25433), .o(n25434) );
na02f01 g21644 ( .a(n25434), .b(n25426), .o(n25435) );
in01f01 g21645 ( .a(n25435), .o(n25436) );
no02f01 g21646 ( .a(n24454), .b(n24453), .o(n25437) );
no02f01 g21647 ( .a(n24451), .b(n24450), .o(n25438) );
no02f01 g21648 ( .a(n25438), .b(n25437), .o(n25439) );
ao12f01 g21649 ( .a(n25439), .b(n24465), .c(n5529), .o(n25440) );
no03f01 g21650 ( .a(n25418), .b(n24456), .c(n5527), .o(n25441) );
no02f01 g21651 ( .a(n25441), .b(n25440), .o(n25442) );
oa12f01 g21652 ( .a(n25442), .b(n25434), .c(n25426), .o(n25443) );
in01f01 g21653 ( .a(n25443), .o(n25444) );
no02f01 g21654 ( .a(n25444), .b(n25436), .o(n25445) );
no03f01 g21655 ( .a(n25085), .b(n24826), .c(n24821), .o(n25446) );
ao12f01 g21656 ( .a(n24848), .b(n25080), .c(n24822), .o(n25447) );
no02f01 g21657 ( .a(n25447), .b(n25446), .o(n25448) );
na03f01 g21658 ( .a(n25448), .b(n25443), .c(n25435), .o(n25449) );
no02f01 g21659 ( .a(n24474), .b(n5529), .o(n25450) );
no03f01 g21660 ( .a(n25450), .b(n24475), .c(n24466), .o(n25451) );
na02f01 g21661 ( .a(n24472), .b(n24471), .o(n25452) );
na02f01 g21662 ( .a(n24469), .b(n24468), .o(n25453) );
na02f01 g21663 ( .a(n25453), .b(n25452), .o(n25454) );
na02f01 g21664 ( .a(n25454), .b(n5529), .o(n25455) );
na02f01 g21665 ( .a(n25454), .b(n5527), .o(n25456) );
ao12f01 g21666 ( .a(n24467), .b(n25456), .c(n25455), .o(n25457) );
no02f01 g21667 ( .a(n25457), .b(n25451), .o(n25458) );
na02f01 g21668 ( .a(n25458), .b(n25449), .o(n25459) );
oa12f01 g21669 ( .a(n25459), .b(n25448), .c(n25445), .o(n25460) );
no03f01 g21670 ( .a(n25414), .b(n25411), .c(n25405), .o(n25461) );
ao12f01 g21671 ( .a(n25461), .b(n25460), .c(n25415), .o(n25462) );
ao12f01 g21672 ( .a(n25401), .b(n25395), .c(n25393), .o(n25463) );
oa12f01 g21673 ( .a(n25402), .b(n25463), .c(n25462), .o(n25464) );
oa12f01 g21674 ( .a(n25390), .b(n25385), .c(n25383), .o(n25465) );
ao12f01 g21675 ( .a(n25391), .b(n25465), .c(n25464), .o(n25466) );
no02f01 g21676 ( .a(n24494), .b(n24432), .o(n25467) );
na02f01 g21677 ( .a(n25467), .b(n24493), .o(n25468) );
oa12f01 g21678 ( .a(n24973), .b(n24494), .c(n24432), .o(n25469) );
no03f01 g21679 ( .a(n25098), .b(n25095), .c(n24786), .o(n25470) );
ao12f01 g21680 ( .a(n24858), .b(n24859), .c(n25074), .o(n25471) );
no02f01 g21681 ( .a(n25471), .b(n25470), .o(n25472) );
in01f01 g21682 ( .a(n25472), .o(n25473) );
ao12f01 g21683 ( .a(n25473), .b(n25469), .c(n25468), .o(n25474) );
no02f01 g21684 ( .a(n25474), .b(n25466), .o(n25475) );
na03f01 g21685 ( .a(n25473), .b(n25469), .c(n25468), .o(n25476) );
no03f01 g21686 ( .a(n24871), .b(n25103), .c(n24860), .o(n25477) );
ao12f01 g21687 ( .a(n25099), .b(n25104), .c(n24870), .o(n25478) );
no02f01 g21688 ( .a(n25478), .b(n25477), .o(n25479) );
na02f01 g21689 ( .a(n25479), .b(n25476), .o(n25480) );
oa12f01 g21690 ( .a(n25380), .b(n25480), .c(n25475), .o(n25481) );
in01f01 g21691 ( .a(n25476), .o(n25482) );
in01f01 g21692 ( .a(n25479), .o(n25483) );
oa12f01 g21693 ( .a(n25483), .b(n25482), .c(n25475), .o(n25484) );
ao22f01 g21694 ( .a(n25484), .b(n25481), .c(n25376), .d(n25371), .o(n25485) );
oa12f01 g21695 ( .a(n25362), .b(n25357), .c(n25356), .o(n25486) );
oa12f01 g21696 ( .a(n25486), .b(n25485), .c(n25377), .o(n25487) );
na02f01 g21697 ( .a(n25348), .b(n25331), .o(n25488) );
na02f01 g21698 ( .a(n25346), .b(n25345), .o(n25489) );
in01f01 g21699 ( .a(n25354), .o(n25490) );
ao12f01 g21700 ( .a(n25490), .b(n25489), .c(n25488), .o(n25491) );
ao12f01 g21701 ( .a(n25491), .b(n25487), .c(n25364), .o(n25492) );
oa12f01 g21702 ( .a(n25342), .b(n25337), .c(n25333), .o(n25493) );
oa12f01 g21703 ( .a(n25493), .b(n25492), .c(n25355), .o(n25494) );
no02f01 g21704 ( .a(n24547), .b(n5527), .o(n25495) );
oa22f01 g21705 ( .a(n24548), .b(n25495), .c(n24994), .d(n24988), .o(n25496) );
na02f01 g21706 ( .a(n24532), .b(n5529), .o(n25497) );
na04f01 g21707 ( .a(n24997), .b(n25497), .c(n24523), .d(n24509), .o(n25498) );
na02f01 g21708 ( .a(n24884), .b(n25111), .o(n25499) );
na02f01 g21709 ( .a(n25499), .b(n25110), .o(n25500) );
no02f01 g21710 ( .a(n24889), .b(n24882), .o(n25501) );
na02f01 g21711 ( .a(n25501), .b(n24877), .o(n25502) );
na02f01 g21712 ( .a(n25502), .b(n25500), .o(n25503) );
ao12f01 g21713 ( .a(n25503), .b(n25498), .c(n25496), .o(n25504) );
ao12f01 g21714 ( .a(n25504), .b(n25494), .c(n25344), .o(n25505) );
na03f01 g21715 ( .a(n25503), .b(n25498), .c(n25496), .o(n25506) );
ao12f01 g21716 ( .a(n24882), .b(n24884), .c(n24877), .o(n25507) );
no02f01 g21717 ( .a(n24740), .b(n23901), .o(n25508) );
no02f01 g21718 ( .a(n25060), .b(n23221), .o(n25509) );
no03f01 g21719 ( .a(n25509), .b(n25508), .c(n25507), .o(n25510) );
in01f01 g21720 ( .a(n25507), .o(n25511) );
na02f01 g21721 ( .a(n25060), .b(n23221), .o(n25512) );
na02f01 g21722 ( .a(n24740), .b(n23901), .o(n25513) );
ao12f01 g21723 ( .a(n25511), .b(n25513), .c(n25512), .o(n25514) );
no02f01 g21724 ( .a(n25514), .b(n25510), .o(n25515) );
na02f01 g21725 ( .a(n25515), .b(n25506), .o(n25516) );
oa12f01 g21726 ( .a(n25328), .b(n25516), .c(n25505), .o(n25517) );
in01f01 g21727 ( .a(n25506), .o(n25518) );
in01f01 g21728 ( .a(n25515), .o(n25519) );
oa12f01 g21729 ( .a(n25519), .b(n25518), .c(n25505), .o(n25520) );
na03f01 g21730 ( .a(n25006), .b(n25303), .c(n24400), .o(n25521) );
oa22f01 g21731 ( .a(n24564), .b(n24963), .c(n24998), .d(n24996), .o(n25522) );
ao12f01 g21732 ( .a(n25311), .b(n25120), .c(n25317), .o(n25523) );
no03f01 g21733 ( .a(n24895), .b(n25312), .c(n25316), .o(n25524) );
no02f01 g21734 ( .a(n25524), .b(n25523), .o(n25525) );
in01f01 g21735 ( .a(n25525), .o(n25526) );
ao12f01 g21736 ( .a(n25526), .b(n25522), .c(n25521), .o(n25527) );
ao12f01 g21737 ( .a(n25527), .b(n25520), .c(n25517), .o(n25528) );
in01f01 g21738 ( .a(n25307), .o(n25529) );
no03f01 g21739 ( .a(n25320), .b(n25308), .c(n25529), .o(n25530) );
na03f01 g21740 ( .a(n25526), .b(n25522), .c(n25521), .o(n25531) );
in01f01 g21741 ( .a(n25531), .o(n25532) );
no03f01 g21742 ( .a(n25532), .b(n25530), .c(n25528), .o(n25533) );
no02f01 g21743 ( .a(n25533), .b(n25322), .o(n25534) );
na02f01 g21744 ( .a(n25276), .b(n25269), .o(n25535) );
no02f01 g21745 ( .a(n25250), .b(n25230), .o(n25536) );
na04f01 g21746 ( .a(n25536), .b(n25535), .c(n25534), .d(n25302), .o(n25537) );
no02f01 g21747 ( .a(n25537), .b(n25219), .o(n25538) );
in01f01 g21748 ( .a(n25145), .o(n25539) );
na03f01 g21749 ( .a(n25155), .b(n25149), .c(n25153), .o(n25540) );
oa12f01 g21750 ( .a(n25150), .b(n25151), .c(n25048), .o(n25541) );
na02f01 g21751 ( .a(n25541), .b(n25540), .o(n25542) );
no02f01 g21752 ( .a(n25542), .b(n25539), .o(n25543) );
ao12f01 g21753 ( .a(n25023), .b(n25543), .c(n25179), .o(n25544) );
oa12f01 g21754 ( .a(n24613), .b(n25544), .c(n25170), .o(n25545) );
in01f01 g21755 ( .a(n25034), .o(n25546) );
ao12f01 g21756 ( .a(n25023), .b(n25044), .c(n25546), .o(n25547) );
in01f01 g21757 ( .a(n25547), .o(n25548) );
na02f01 g21758 ( .a(n25548), .b(n25545), .o(n25549) );
ao12f01 g21759 ( .a(n25549), .b(n25538), .c(n25182), .o(n25550) );
oa12f01 g21760 ( .a(n25550), .b(n25301), .c(n25183), .o(n25551) );
na03f01 g21761 ( .a(n25551), .b(n25047), .c(n25026), .o(n25552) );
in01f01 g21762 ( .a(n25047), .o(n25553) );
na03f01 g21763 ( .a(n25186), .b(n25134), .c(n25053), .o(n25554) );
oa12f01 g21764 ( .a(n25184), .b(n24917), .c(n24707), .o(n25555) );
na02f01 g21765 ( .a(n25555), .b(n25554), .o(n25556) );
no02f01 g21766 ( .a(n25556), .b(n24613), .o(n25557) );
na02f01 g21767 ( .a(n25192), .b(n25022), .o(n25558) );
na02f01 g21768 ( .a(n25190), .b(n24610), .o(n25559) );
in01f01 g21769 ( .a(n25200), .o(n25560) );
ao12f01 g21770 ( .a(n25560), .b(n25559), .c(n25558), .o(n25561) );
no03f01 g21771 ( .a(n25294), .b(n25561), .c(n25557), .o(n25562) );
oa12f01 g21772 ( .a(n25248), .b(n25281), .c(n25280), .o(n25563) );
na02f01 g21773 ( .a(n25260), .b(n25258), .o(n25564) );
oa22f01 g21774 ( .a(n25276), .b(n25269), .c(n25564), .d(n25255), .o(n25565) );
na03f01 g21775 ( .a(n25565), .b(n25302), .c(n25563), .o(n25566) );
in01f01 g21776 ( .a(n25284), .o(n25567) );
no02f01 g21777 ( .a(n25567), .b(n25282), .o(n25568) );
ao12f01 g21778 ( .a(n25230), .b(n25568), .c(n25566), .o(n25569) );
na02f01 g21779 ( .a(n25569), .b(n25562), .o(n25570) );
na02f01 g21780 ( .a(n25556), .b(n24613), .o(n25571) );
na03f01 g21781 ( .a(n25560), .b(n25559), .c(n25558), .o(n25572) );
ao12f01 g21782 ( .a(n25557), .b(n25572), .c(n25571), .o(n25573) );
oa12f01 g21783 ( .a(n25218), .b(n25298), .c(n25573), .o(n25574) );
na02f01 g21784 ( .a(n25574), .b(n25570), .o(n25575) );
na02f01 g21785 ( .a(n25538), .b(n25182), .o(n25576) );
in01f01 g21786 ( .a(n25549), .o(n25577) );
na02f01 g21787 ( .a(n25577), .b(n25576), .o(n25578) );
ao12f01 g21788 ( .a(n25578), .b(n25575), .c(n25182), .o(n25579) );
oa12f01 g21789 ( .a(n25025), .b(n25579), .c(n25553), .o(n25580) );
na02f01 g21790 ( .a(n25580), .b(n25552), .o(n303) );
na02f01 g21791 ( .a(n22401), .b(n11514), .o(n25582) );
na02f01 g21792 ( .a(n22401), .b(n11515), .o(n25583) );
na02f01 g21793 ( .a(n25583), .b(n25582), .o(n25584) );
ao12f01 g21794 ( .a(n13588), .b(n22406), .c(n11515), .o(n25585) );
oa12f01 g21795 ( .a(n25585), .b(n14309), .c(n14253), .o(n25586) );
no02f01 g21796 ( .a(n25586), .b(n25584), .o(n25587) );
ao12f01 g21797 ( .a(n22399), .b(n22398), .c(n14301), .o(n25588) );
no03f01 g21798 ( .a(n22396), .b(n22394), .c(n14305), .o(n25589) );
no02f01 g21799 ( .a(n25589), .b(n25588), .o(n25590) );
no02f01 g21800 ( .a(n25590), .b(n11515), .o(n25591) );
no02f01 g21801 ( .a(n25590), .b(n11514), .o(n25592) );
no02f01 g21802 ( .a(n25592), .b(n25591), .o(n25593) );
ao12f01 g21803 ( .a(n14253), .b(n22406), .c(n11514), .o(n25594) );
oa12f01 g21804 ( .a(n14252), .b(n14308), .c(n11514), .o(n25595) );
no02f01 g21805 ( .a(n25595), .b(n25594), .o(n25596) );
no02f01 g21806 ( .a(n25596), .b(n25593), .o(n25597) );
no02f01 g21807 ( .a(n25597), .b(n25587), .o(n25598) );
na02f01 g21808 ( .a(n25598), .b(n21914), .o(n25599) );
no02f01 g21809 ( .a(n25598), .b(n21914), .o(n25600) );
in01f01 g21810 ( .a(n25600), .o(n25601) );
na02f01 g21811 ( .a(n13965), .b(n13909), .o(n25602) );
na03f01 g21812 ( .a(n14331), .b(n14313), .c(n14311), .o(n25603) );
na02f01 g21813 ( .a(n25603), .b(n14247), .o(n25604) );
ao12f01 g21814 ( .a(n25604), .b(n14239), .c(n25602), .o(n25605) );
oa12f01 g21815 ( .a(n14335), .b(n14312), .c(n14333), .o(n25606) );
ao12f01 g21816 ( .a(n14336), .b(n25606), .c(n13890), .o(n25607) );
no02f01 g21817 ( .a(n25607), .b(n25605), .o(n25608) );
na02f01 g21818 ( .a(n25608), .b(n25601), .o(n25609) );
na02f01 g21819 ( .a(n25609), .b(n25599), .o(n25610) );
ao12f01 g21820 ( .a(n11515), .b(n22434), .c(n22430), .o(n25611) );
ao12f01 g21821 ( .a(n11514), .b(n22434), .c(n22430), .o(n25612) );
no02f01 g21822 ( .a(n25612), .b(n25611), .o(n25613) );
oa12f01 g21823 ( .a(n25582), .b(n25586), .c(n25592), .o(n25614) );
na02f01 g21824 ( .a(n25614), .b(n25613), .o(n25615) );
ao12f01 g21825 ( .a(n25591), .b(n25596), .c(n25583), .o(n25616) );
oa12f01 g21826 ( .a(n25616), .b(n25612), .c(n25611), .o(n25617) );
ao12f01 g21827 ( .a(n21922), .b(n25617), .c(n25615), .o(n25618) );
na03f01 g21828 ( .a(n25617), .b(n25615), .c(n21922), .o(n25619) );
in01f01 g21829 ( .a(n25619), .o(n25620) );
no02f01 g21830 ( .a(n25620), .b(n25618), .o(n25621) );
na02f01 g21831 ( .a(n25621), .b(n25610), .o(n25622) );
no02f01 g21832 ( .a(n25621), .b(n25610), .o(n25623) );
in01f01 g21833 ( .a(n25623), .o(n25624) );
na02f01 g21834 ( .a(n25624), .b(n25622), .o(n6047) );
na02f01 g21835 ( .a(n6047), .b(n4116), .o(n25626) );
na03f01 g21836 ( .a(n25624), .b(n25622), .c(n2589), .o(n25627) );
na02f01 g21837 ( .a(n25627), .b(n25626), .o(n308) );
na02f01 g21838 ( .a(n10876), .b(n10809), .o(n25629) );
in01f01 g21839 ( .a(n25629), .o(n25630) );
ao12f01 g21840 ( .a(n10926), .b(n10899), .c(n25630), .o(n25631) );
no02f01 g21841 ( .a(n10910), .b(n3521), .o(n25632) );
no02f01 g21842 ( .a(n25632), .b(n10912), .o(n25633) );
na02f01 g21843 ( .a(n25633), .b(n25631), .o(n25634) );
in01f01 g21844 ( .a(n25631), .o(n25635) );
in01f01 g21845 ( .a(n25633), .o(n25636) );
na02f01 g21846 ( .a(n25636), .b(n25635), .o(n25637) );
na02f01 g21847 ( .a(n25637), .b(n25634), .o(n313) );
no02f01 g21848 ( .a(n22381), .b(n22366), .o(n25639) );
oa12f01 g21849 ( .a(n22415), .b(n22421), .c(n25639), .o(n25640) );
no02f01 g21850 ( .a(n22423), .b(n22412), .o(n25641) );
na02f01 g21851 ( .a(n25641), .b(n25640), .o(n25642) );
na02f01 g21852 ( .a(n22471), .b(n22470), .o(n25643) );
ao12f01 g21853 ( .a(n22392), .b(n22481), .c(n25643), .o(n25644) );
in01f01 g21854 ( .a(n25641), .o(n25645) );
na02f01 g21855 ( .a(n25645), .b(n25644), .o(n25646) );
na03f01 g21856 ( .a(n25646), .b(n25642), .c(n2589), .o(n25647) );
na02f01 g21857 ( .a(n25646), .b(n25642), .o(n804) );
na02f01 g21858 ( .a(n804), .b(n4116), .o(n25649) );
na02f01 g21859 ( .a(n25649), .b(n25647), .o(n318) );
in01f01 g21860 ( .a(n22749), .o(n25651) );
oa12f01 g21861 ( .a(n25651), .b(n22751), .c(n22739), .o(n25652) );
no02f01 g21862 ( .a(n22720), .b(n18134), .o(n25653) );
oa12f01 g21863 ( .a(n25653), .b(n18373), .c(n18364), .o(n25654) );
in01f01 g21864 ( .a(n25654), .o(n25655) );
no02f01 g21865 ( .a(n18375), .b(n18143), .o(n25656) );
no02f01 g21866 ( .a(n25656), .b(n25655), .o(n25657) );
na02f01 g21867 ( .a(n25656), .b(n25655), .o(n25658) );
in01f01 g21868 ( .a(n25658), .o(n25659) );
no02f01 g21869 ( .a(n25659), .b(n25657), .o(n25660) );
in01f01 g21870 ( .a(n25660), .o(n25661) );
no02f01 g21871 ( .a(n25661), .b(n18459), .o(n25662) );
no02f01 g21872 ( .a(n25660), .b(n18460), .o(n25663) );
no02f01 g21873 ( .a(n25663), .b(n25662), .o(n25664) );
in01f01 g21874 ( .a(n25664), .o(n25665) );
na02f01 g21875 ( .a(n25665), .b(n25652), .o(n25666) );
in01f01 g21876 ( .a(n25652), .o(n25667) );
na02f01 g21877 ( .a(n25664), .b(n25667), .o(n25668) );
na02f01 g21878 ( .a(n25668), .b(n25666), .o(n323) );
na02f01 g21879 ( .a(n25290), .b(n5527), .o(n25670) );
na02f01 g21880 ( .a(n25290), .b(n5529), .o(n25671) );
na02f01 g21881 ( .a(n25671), .b(n25670), .o(n25672) );
oa12f01 g21882 ( .a(n5529), .b(n25247), .c(n25244), .o(n25673) );
oa12f01 g21883 ( .a(n5527), .b(n25254), .c(n25252), .o(n25674) );
oa12f01 g21884 ( .a(n25316), .b(n24895), .c(n25312), .o(n25675) );
na03f01 g21885 ( .a(n25120), .b(n25317), .c(n25311), .o(n25676) );
ao12f01 g21886 ( .a(n5527), .b(n25676), .c(n25675), .o(n25677) );
na03f01 g21887 ( .a(n25513), .b(n25512), .c(n25511), .o(n25678) );
oa12f01 g21888 ( .a(n25507), .b(n25509), .c(n25508), .o(n25679) );
ao12f01 g21889 ( .a(n5527), .b(n25679), .c(n25678), .o(n25680) );
oa12f01 g21890 ( .a(n5529), .b(n25503), .c(n25341), .o(n25681) );
in01f01 g21891 ( .a(n25681), .o(n25682) );
no03f01 g21892 ( .a(n25682), .b(n25680), .c(n25677), .o(n25683) );
oa12f01 g21893 ( .a(n5527), .b(n25524), .c(n25523), .o(n25684) );
oa12f01 g21894 ( .a(n5527), .b(n25514), .c(n25510), .o(n25685) );
na02f01 g21895 ( .a(n25685), .b(n25684), .o(n25686) );
oa12f01 g21896 ( .a(n5529), .b(n25319), .c(n25314), .o(n25687) );
oa12f01 g21897 ( .a(n25687), .b(n25686), .c(n25683), .o(n25688) );
na02f01 g21898 ( .a(n25274), .b(n25273), .o(n25689) );
na02f01 g21899 ( .a(n25271), .b(n25270), .o(n25690) );
ao12f01 g21900 ( .a(n5527), .b(n25690), .c(n25689), .o(n25691) );
no02f01 g21901 ( .a(n25691), .b(n25688), .o(n25692) );
oa12f01 g21902 ( .a(n5527), .b(n25319), .c(n25314), .o(n25693) );
oa12f01 g21903 ( .a(n5527), .b(n25275), .c(n25272), .o(n25694) );
na02f01 g21904 ( .a(n25694), .b(n25693), .o(n25695) );
oa12f01 g21905 ( .a(n5529), .b(n25254), .c(n25252), .o(n25696) );
oa12f01 g21906 ( .a(n25696), .b(n25695), .c(n25692), .o(n25697) );
oa12f01 g21907 ( .a(n5527), .b(n25247), .c(n25244), .o(n25698) );
na03f01 g21908 ( .a(n25698), .b(n25697), .c(n25674), .o(n25699) );
oa12f01 g21909 ( .a(n5529), .b(n25227), .c(n25225), .o(n25700) );
na03f01 g21910 ( .a(n25700), .b(n25699), .c(n25673), .o(n25701) );
na02f01 g21911 ( .a(n25198), .b(n25197), .o(n25702) );
na02f01 g21912 ( .a(n25195), .b(n25194), .o(n25703) );
ao12f01 g21913 ( .a(n5527), .b(n25703), .c(n25702), .o(n25704) );
no02f01 g21914 ( .a(n25704), .b(n25701), .o(n25705) );
oa12f01 g21915 ( .a(n25705), .b(n25188), .c(n5527), .o(n25706) );
ao12f01 g21916 ( .a(n25706), .b(n25293), .c(n5529), .o(n25707) );
oa12f01 g21917 ( .a(n5527), .b(n25199), .c(n25196), .o(n25708) );
oa12f01 g21918 ( .a(n5527), .b(n25227), .c(n25225), .o(n25709) );
na02f01 g21919 ( .a(n25709), .b(n25708), .o(n25710) );
ao12f01 g21920 ( .a(n25710), .b(n25556), .c(n5527), .o(n25711) );
oa12f01 g21921 ( .a(n25711), .b(n25217), .c(n5529), .o(n25712) );
no02f01 g21922 ( .a(n25712), .b(n25707), .o(n25713) );
in01f01 g21923 ( .a(n25713), .o(n25714) );
na02f01 g21924 ( .a(n25714), .b(n25672), .o(n25715) );
no02f01 g21925 ( .a(n25212), .b(n5529), .o(n25716) );
no02f01 g21926 ( .a(n25212), .b(n5527), .o(n25717) );
no02f01 g21927 ( .a(n25717), .b(n25716), .o(n25718) );
na02f01 g21928 ( .a(n25713), .b(n25718), .o(n25719) );
ao12f01 g21929 ( .a(n25439), .b(n25719), .c(n25715), .o(n25720) );
no02f01 g21930 ( .a(n25713), .b(n25718), .o(n25721) );
no02f01 g21931 ( .a(n25714), .b(n25672), .o(n25722) );
no03f01 g21932 ( .a(n25722), .b(n25721), .c(n24456), .o(n25723) );
no02f01 g21933 ( .a(n25723), .b(n25720), .o(n25724) );
na02f01 g21934 ( .a(n25293), .b(n5529), .o(n25725) );
na02f01 g21935 ( .a(n25293), .b(n5527), .o(n25726) );
na02f01 g21936 ( .a(n25726), .b(n25725), .o(n25727) );
in01f01 g21937 ( .a(n25673), .o(n25728) );
na03f01 g21938 ( .a(n24904), .b(n25253), .c(n24721), .o(n25729) );
oa12f01 g21939 ( .a(n25251), .b(n25127), .c(n24720), .o(n25730) );
ao12f01 g21940 ( .a(n5529), .b(n25730), .c(n25729), .o(n25731) );
oa12f01 g21941 ( .a(n5529), .b(n25524), .c(n25523), .o(n25732) );
oa12f01 g21942 ( .a(n5529), .b(n25514), .c(n25510), .o(n25733) );
na03f01 g21943 ( .a(n25681), .b(n25733), .c(n25732), .o(n25734) );
ao12f01 g21944 ( .a(n5529), .b(n25676), .c(n25675), .o(n25735) );
ao12f01 g21945 ( .a(n5529), .b(n25679), .c(n25678), .o(n25736) );
no02f01 g21946 ( .a(n25736), .b(n25735), .o(n25737) );
na02f01 g21947 ( .a(n25318), .b(n25315), .o(n25738) );
na02f01 g21948 ( .a(n25313), .b(n25310), .o(n25739) );
ao12f01 g21949 ( .a(n5527), .b(n25739), .c(n25738), .o(n25740) );
ao12f01 g21950 ( .a(n25740), .b(n25737), .c(n25734), .o(n25741) );
oa12f01 g21951 ( .a(n5529), .b(n25275), .c(n25272), .o(n25742) );
na02f01 g21952 ( .a(n25742), .b(n25741), .o(n25743) );
ao12f01 g21953 ( .a(n5529), .b(n25739), .c(n25738), .o(n25744) );
ao12f01 g21954 ( .a(n5529), .b(n25690), .c(n25689), .o(n25745) );
no02f01 g21955 ( .a(n25745), .b(n25744), .o(n25746) );
ao12f01 g21956 ( .a(n5527), .b(n25730), .c(n25729), .o(n25747) );
ao12f01 g21957 ( .a(n25747), .b(n25746), .c(n25743), .o(n25748) );
na02f01 g21958 ( .a(n25246), .b(n25245), .o(n25749) );
na02f01 g21959 ( .a(n25243), .b(n25242), .o(n25750) );
ao12f01 g21960 ( .a(n5529), .b(n25750), .c(n25749), .o(n25751) );
no03f01 g21961 ( .a(n25751), .b(n25748), .c(n25731), .o(n25752) );
na03f01 g21962 ( .a(n25226), .b(n25130), .c(n25055), .o(n25753) );
oa12f01 g21963 ( .a(n25224), .b(n24909), .c(n24715), .o(n25754) );
ao12f01 g21964 ( .a(n5527), .b(n25754), .c(n25753), .o(n25755) );
no03f01 g21965 ( .a(n25755), .b(n25752), .c(n25728), .o(n25756) );
oa12f01 g21966 ( .a(n5529), .b(n25199), .c(n25196), .o(n25757) );
na02f01 g21967 ( .a(n25757), .b(n25756), .o(n25758) );
ao12f01 g21968 ( .a(n25758), .b(n25556), .c(n5529), .o(n25759) );
ao12f01 g21969 ( .a(n5529), .b(n25703), .c(n25702), .o(n25760) );
ao12f01 g21970 ( .a(n5529), .b(n25754), .c(n25753), .o(n25761) );
no02f01 g21971 ( .a(n25761), .b(n25760), .o(n25762) );
oa12f01 g21972 ( .a(n25762), .b(n25188), .c(n5529), .o(n25763) );
no02f01 g21973 ( .a(n25763), .b(n25759), .o(n25764) );
in01f01 g21974 ( .a(n25764), .o(n25765) );
no02f01 g21975 ( .a(n25765), .b(n25727), .o(n25766) );
no02f01 g21976 ( .a(n25217), .b(n5527), .o(n25767) );
no02f01 g21977 ( .a(n25217), .b(n5529), .o(n25768) );
no02f01 g21978 ( .a(n25768), .b(n25767), .o(n25769) );
no02f01 g21979 ( .a(n25764), .b(n25769), .o(n25770) );
no02f01 g21980 ( .a(n25770), .b(n25766), .o(n25771) );
no02f01 g21981 ( .a(n25771), .b(n25418), .o(n25772) );
no02f01 g21982 ( .a(n25710), .b(n25705), .o(n25773) );
no02f01 g21983 ( .a(n25188), .b(n5527), .o(n25774) );
no02f01 g21984 ( .a(n25188), .b(n5529), .o(n25775) );
no02f01 g21985 ( .a(n25775), .b(n25774), .o(n25776) );
no02f01 g21986 ( .a(n25776), .b(n25773), .o(n25777) );
na02f01 g21987 ( .a(n25776), .b(n25773), .o(n25778) );
in01f01 g21988 ( .a(n25778), .o(n25779) );
no02f01 g21989 ( .a(n25779), .b(n25777), .o(n25780) );
no02f01 g21990 ( .a(n25752), .b(n25728), .o(n25781) );
na02f01 g21991 ( .a(n25709), .b(n25700), .o(n25782) );
na02f01 g21992 ( .a(n25782), .b(n25781), .o(n25783) );
na02f01 g21993 ( .a(n25699), .b(n25673), .o(n25784) );
no02f01 g21994 ( .a(n25761), .b(n25755), .o(n25785) );
na02f01 g21995 ( .a(n25785), .b(n25784), .o(n25786) );
no02f01 g21996 ( .a(n24105), .b(n24100), .o(n25787) );
no02f01 g21997 ( .a(n24107), .b(n24307), .o(n25788) );
no02f01 g21998 ( .a(n25788), .b(n25787), .o(n25789) );
na02f01 g21999 ( .a(n25788), .b(n25787), .o(n25790) );
in01f01 g22000 ( .a(n25790), .o(n25791) );
no02f01 g22001 ( .a(n25791), .b(n25789), .o(n25792) );
ao12f01 g22002 ( .a(n25792), .b(n25786), .c(n25783), .o(n25793) );
in01f01 g22003 ( .a(n25793), .o(n25794) );
na02f01 g22004 ( .a(n25697), .b(n25674), .o(n25795) );
na02f01 g22005 ( .a(n25698), .b(n25673), .o(n25796) );
no02f01 g22006 ( .a(n25796), .b(n25795), .o(n25797) );
no02f01 g22007 ( .a(n25748), .b(n25731), .o(n25798) );
ao12f01 g22008 ( .a(n25798), .b(n25698), .c(n25673), .o(n25799) );
no02f01 g22009 ( .a(n25799), .b(n25797), .o(n25800) );
ao22f01 g22010 ( .a(n25694), .b(n25742), .c(n25693), .d(n25688), .o(n25801) );
no04f01 g22011 ( .a(n25745), .b(n25744), .c(n25691), .d(n25741), .o(n25802) );
no02f01 g22012 ( .a(n24332), .b(n24021), .o(n25803) );
no02f01 g22013 ( .a(n25803), .b(n24077), .o(n25804) );
na02f01 g22014 ( .a(n25803), .b(n24077), .o(n25805) );
in01f01 g22015 ( .a(n25805), .o(n25806) );
no02f01 g22016 ( .a(n25806), .b(n25804), .o(n25807) );
in01f01 g22017 ( .a(n25807), .o(n25808) );
oa12f01 g22018 ( .a(n25808), .b(n25802), .c(n25801), .o(n25809) );
no03f01 g22019 ( .a(n25808), .b(n25802), .c(n25801), .o(n25810) );
na04f01 g22020 ( .a(n25693), .b(n25687), .c(n25737), .d(n25734), .o(n25811) );
oa22f01 g22021 ( .a(n25744), .b(n25740), .c(n25686), .d(n25683), .o(n25812) );
no02f01 g22022 ( .a(n24330), .b(n24031), .o(n25813) );
no02f01 g22023 ( .a(n25813), .b(n24329), .o(n25814) );
na02f01 g22024 ( .a(n25813), .b(n24329), .o(n25815) );
in01f01 g22025 ( .a(n25815), .o(n25816) );
no02f01 g22026 ( .a(n25816), .b(n25814), .o(n25817) );
ao12f01 g22027 ( .a(n25817), .b(n25812), .c(n25811), .o(n25818) );
oa12f01 g22028 ( .a(n25681), .b(n25736), .c(n25680), .o(n25819) );
na03f01 g22029 ( .a(n25685), .b(n25682), .c(n25733), .o(n25820) );
no02f01 g22030 ( .a(n24072), .b(n24324), .o(n25821) );
no02f01 g22031 ( .a(n25821), .b(n24325), .o(n25822) );
na02f01 g22032 ( .a(n25821), .b(n24325), .o(n25823) );
in01f01 g22033 ( .a(n25823), .o(n25824) );
no02f01 g22034 ( .a(n25824), .b(n25822), .o(n25825) );
ao12f01 g22035 ( .a(n25825), .b(n25820), .c(n25819), .o(n25826) );
na03f01 g22036 ( .a(n25825), .b(n25820), .c(n25819), .o(n25827) );
no02f01 g22037 ( .a(n25341), .b(n5529), .o(n25828) );
no02f01 g22038 ( .a(n25341), .b(n5527), .o(n25829) );
no02f01 g22039 ( .a(n25829), .b(n25828), .o(n25830) );
in01f01 g22040 ( .a(n24058), .o(n25831) );
no02f01 g22041 ( .a(n25831), .b(n23905), .o(n25832) );
no02f01 g22042 ( .a(n24058), .b(n23231), .o(n25833) );
no02f01 g22043 ( .a(n25833), .b(n25832), .o(n25834) );
in01f01 g22044 ( .a(n25834), .o(n25835) );
na02f01 g22045 ( .a(n25835), .b(n25830), .o(n25836) );
in01f01 g22046 ( .a(n24066), .o(n25837) );
no02f01 g22047 ( .a(n25837), .b(n24055), .o(n25838) );
na02f01 g22048 ( .a(n25837), .b(n24055), .o(n25839) );
in01f01 g22049 ( .a(n25839), .o(n25840) );
no03f01 g22050 ( .a(n25840), .b(n25838), .c(n24059), .o(n25841) );
in01f01 g22051 ( .a(n25838), .o(n25842) );
ao12f01 g22052 ( .a(n24060), .b(n25839), .c(n25842), .o(n25843) );
no02f01 g22053 ( .a(n25843), .b(n25841), .o(n25844) );
no02f01 g22054 ( .a(n25844), .b(n25836), .o(n25845) );
na02f01 g22055 ( .a(n25844), .b(n25836), .o(n25846) );
oa12f01 g22056 ( .a(n25503), .b(n25342), .c(n5527), .o(n25847) );
na04f01 g22057 ( .a(n25502), .b(n25500), .c(n25341), .d(n5529), .o(n25848) );
na02f01 g22058 ( .a(n25848), .b(n25847), .o(n25849) );
ao12f01 g22059 ( .a(n25845), .b(n25849), .c(n25846), .o(n25850) );
in01f01 g22060 ( .a(n25850), .o(n25851) );
ao12f01 g22061 ( .a(n25826), .b(n25851), .c(n25827), .o(n25852) );
oa12f01 g22062 ( .a(n25685), .b(n25682), .c(n25680), .o(n25853) );
no03f01 g22063 ( .a(n25853), .b(n25735), .c(n25677), .o(n25854) );
ao12f01 g22064 ( .a(n25736), .b(n25681), .c(n25733), .o(n25855) );
ao12f01 g22065 ( .a(n25855), .b(n25684), .c(n25732), .o(n25856) );
no03f01 g22066 ( .a(n24074), .b(n24327), .c(n24320), .o(n25857) );
ao12f01 g22067 ( .a(n24073), .b(n24328), .c(n24042), .o(n25858) );
no02f01 g22068 ( .a(n25858), .b(n25857), .o(n25859) );
in01f01 g22069 ( .a(n25859), .o(n25860) );
no03f01 g22070 ( .a(n25860), .b(n25856), .c(n25854), .o(n25861) );
oa12f01 g22071 ( .a(n25860), .b(n25856), .c(n25854), .o(n25862) );
oa12f01 g22072 ( .a(n25862), .b(n25861), .c(n25852), .o(n25863) );
na03f01 g22073 ( .a(n25817), .b(n25812), .c(n25811), .o(n25864) );
ao12f01 g22074 ( .a(n25818), .b(n25864), .c(n25863), .o(n25865) );
oa12f01 g22075 ( .a(n25809), .b(n25865), .c(n25810), .o(n25866) );
oa22f01 g22076 ( .a(n25747), .b(n25731), .c(n25695), .d(n25692), .o(n25867) );
na04f01 g22077 ( .a(n25696), .b(n25746), .c(n25743), .d(n25674), .o(n25868) );
no03f01 g22078 ( .a(n24090), .b(n24334), .c(n24079), .o(n25869) );
ao12f01 g22079 ( .a(n24333), .b(n24104), .c(n24088), .o(n25870) );
no02f01 g22080 ( .a(n25870), .b(n25869), .o(n25871) );
na03f01 g22081 ( .a(n25871), .b(n25868), .c(n25867), .o(n25872) );
na02f01 g22082 ( .a(n25872), .b(n25866), .o(n25873) );
ao12f01 g22083 ( .a(n25871), .b(n25868), .c(n25867), .o(n25874) );
ao12f01 g22084 ( .a(n24334), .b(n24104), .c(n24333), .o(n25875) );
no02f01 g22085 ( .a(n24098), .b(n24310), .o(n25876) );
no02f01 g22086 ( .a(n24097), .b(n24010), .o(n25877) );
no02f01 g22087 ( .a(n25877), .b(n25876), .o(n25878) );
in01f01 g22088 ( .a(n25878), .o(n25879) );
no02f01 g22089 ( .a(n25879), .b(n25875), .o(n25880) );
na02f01 g22090 ( .a(n25879), .b(n25875), .o(n25881) );
in01f01 g22091 ( .a(n25881), .o(n25882) );
no02f01 g22092 ( .a(n25882), .b(n25880), .o(n25883) );
in01f01 g22093 ( .a(n25883), .o(n25884) );
no02f01 g22094 ( .a(n25884), .b(n25874), .o(n25885) );
ao12f01 g22095 ( .a(n25800), .b(n25885), .c(n25873), .o(n25886) );
ao22f01 g22096 ( .a(n25696), .b(n25674), .c(n25746), .d(n25743), .o(n25887) );
no04f01 g22097 ( .a(n25747), .b(n25695), .c(n25692), .d(n25731), .o(n25888) );
in01f01 g22098 ( .a(n25871), .o(n25889) );
oa12f01 g22099 ( .a(n25889), .b(n25888), .c(n25887), .o(n25890) );
ao12f01 g22100 ( .a(n25883), .b(n25890), .c(n25873), .o(n25891) );
na03f01 g22101 ( .a(n25792), .b(n25786), .c(n25783), .o(n25892) );
oa12f01 g22102 ( .a(n25892), .b(n25891), .c(n25886), .o(n25893) );
ao22f01 g22103 ( .a(n25709), .b(n25701), .c(n25708), .d(n25757), .o(n25894) );
na02f01 g22104 ( .a(n25709), .b(n25701), .o(n25895) );
na02f01 g22105 ( .a(n25708), .b(n25757), .o(n25896) );
no02f01 g22106 ( .a(n25896), .b(n25895), .o(n25897) );
no02f01 g22107 ( .a(n24107), .b(n24339), .o(n25898) );
no02f01 g22108 ( .a(n24114), .b(n24304), .o(n25899) );
no02f01 g22109 ( .a(n24340), .b(n23996), .o(n25900) );
no02f01 g22110 ( .a(n25900), .b(n25899), .o(n25901) );
no02f01 g22111 ( .a(n25901), .b(n25898), .o(n25902) );
na02f01 g22112 ( .a(n25901), .b(n25898), .o(n25903) );
in01f01 g22113 ( .a(n25903), .o(n25904) );
no02f01 g22114 ( .a(n25904), .b(n25902), .o(n25905) );
in01f01 g22115 ( .a(n25905), .o(n25906) );
no03f01 g22116 ( .a(n25906), .b(n25897), .c(n25894), .o(n25907) );
ao12f01 g22117 ( .a(n25907), .b(n25893), .c(n25794), .o(n25908) );
na02f01 g22118 ( .a(n25896), .b(n25895), .o(n25909) );
na04f01 g22119 ( .a(n25709), .b(n25708), .c(n25757), .d(n25701), .o(n25910) );
ao12f01 g22120 ( .a(n25905), .b(n25910), .c(n25909), .o(n25911) );
no02f01 g22121 ( .a(n24344), .b(n23991), .o(n25912) );
no02f01 g22122 ( .a(n25912), .b(n24117), .o(n25913) );
na02f01 g22123 ( .a(n25912), .b(n24117), .o(n25914) );
in01f01 g22124 ( .a(n25914), .o(n25915) );
no02f01 g22125 ( .a(n25915), .b(n25913), .o(n25916) );
in01f01 g22126 ( .a(n25916), .o(n25917) );
no03f01 g22127 ( .a(n25917), .b(n25911), .c(n25908), .o(n25918) );
oa12f01 g22128 ( .a(n25917), .b(n25911), .c(n25908), .o(n25919) );
oa12f01 g22129 ( .a(n25919), .b(n25918), .c(n25780), .o(n25920) );
na02f01 g22130 ( .a(n25771), .b(n25418), .o(n25921) );
ao12f01 g22131 ( .a(n25772), .b(n25921), .c(n25920), .o(n25922) );
no02f01 g22132 ( .a(n25922), .b(n25724), .o(n25923) );
na02f01 g22133 ( .a(n25922), .b(n25724), .o(n25924) );
in01f01 g22134 ( .a(n25924), .o(n25925) );
no02f01 g22135 ( .a(n25925), .b(n25923), .o(n25926) );
na02f01 g22136 ( .a(n25926), .b(n6037), .o(n25927) );
in01f01 g22137 ( .a(n25926), .o(n1285) );
na02f01 g22138 ( .a(n1285), .b(n5873), .o(n25929) );
na02f01 g22139 ( .a(n25929), .b(n25927), .o(n328) );
in01f01 g22140 ( .a(n14153), .o(n25931) );
in01f01 g22141 ( .a(n14154), .o(n25932) );
oa12f01 g22142 ( .a(n25931), .b(n25932), .c(n14115), .o(n25933) );
in01f01 g22143 ( .a(n14115), .o(n25934) );
na03f01 g22144 ( .a(n14154), .b(n14153), .c(n25934), .o(n25935) );
na02f01 g22145 ( .a(n25935), .b(n25933), .o(n333) );
oa12f01 g22146 ( .a(n14149), .b(n14144), .c(n14143), .o(n25937) );
na02f01 g22147 ( .a(n14148), .b(n14145), .o(n25938) );
na02f01 g22148 ( .a(n25938), .b(n25937), .o(n338) );
ao12f01 g22149 ( .a(n_17093), .b(n17433), .c(n17416), .o(n25940) );
in01f01 g22150 ( .a(n25940), .o(n25941) );
no02f01 g22151 ( .a(n16879), .b(delay_add_ln22_unr11_stage5_stallmux_q_31_), .o(n25942) );
na02f01 g22152 ( .a(n16879), .b(delay_add_ln22_unr11_stage5_stallmux_q_31_), .o(n25943) );
in01f01 g22153 ( .a(n25943), .o(n25944) );
no02f01 g22154 ( .a(n25944), .b(n25942), .o(n25945) );
in01f01 g22155 ( .a(n25945), .o(n25946) );
no03f01 g22156 ( .a(n17428), .b(n17420), .c(n17410), .o(n25947) );
ao12f01 g22157 ( .a(n16882), .b(n17426), .c(n17421), .o(n25948) );
no02f01 g22158 ( .a(n25948), .b(n17374), .o(n25949) );
in01f01 g22159 ( .a(n25949), .o(n25950) );
no03f01 g22160 ( .a(n25950), .b(n25947), .c(n25946), .o(n25951) );
no02f01 g22161 ( .a(n25950), .b(n25947), .o(n25952) );
no02f01 g22162 ( .a(n25952), .b(n25945), .o(n25953) );
no02f01 g22163 ( .a(n25953), .b(n25951), .o(n25954) );
ao12f01 g22164 ( .a(n_17093), .b(n25954), .c(n25941), .o(n25955) );
no02f01 g22165 ( .a(n17435), .b(n17474), .o(n25956) );
no02f01 g22166 ( .a(n25954), .b(n7550), .o(n25957) );
in01f01 g22167 ( .a(n25957), .o(n25958) );
ao12f01 g22168 ( .a(n25955), .b(n25958), .c(n25956), .o(n25959) );
no02f01 g22169 ( .a(n25954), .b(n_17093), .o(n25960) );
no02f01 g22170 ( .a(n25960), .b(n25957), .o(n25961) );
no02f01 g22171 ( .a(n25961), .b(n25959), .o(n25962) );
in01f01 g22172 ( .a(n25962), .o(n25963) );
na02f01 g22173 ( .a(n25961), .b(n25959), .o(n25964) );
na02f01 g22174 ( .a(n25964), .b(n25963), .o(n25965) );
na04f01 g22175 ( .a(n16777), .b(n16763), .c(n16588), .d(n16585), .o(n25966) );
no02f01 g22176 ( .a(n16549), .b(delay_xor_ln21_unr12_stage5_stallmux_q_18_), .o(n25967) );
no02f01 g22177 ( .a(n25967), .b(n25966), .o(n25968) );
no02f01 g22178 ( .a(n16549), .b(delay_xor_ln21_unr12_stage5_stallmux_q_19_), .o(n25969) );
na02f01 g22179 ( .a(n16549), .b(delay_xor_ln21_unr12_stage5_stallmux_q_19_), .o(n25970) );
in01f01 g22180 ( .a(n25970), .o(n25971) );
no02f01 g22181 ( .a(n25971), .b(n25969), .o(n25972) );
in01f01 g22182 ( .a(n25972), .o(n25973) );
no02f01 g22183 ( .a(n25973), .b(n25968), .o(n25974) );
no03f01 g22184 ( .a(n25972), .b(n25967), .c(n25966), .o(n25975) );
no02f01 g22185 ( .a(n25975), .b(n25974), .o(n25976) );
no02f01 g22186 ( .a(n25976), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_19_), .o(n25977) );
na02f01 g22187 ( .a(n16549), .b(delay_xor_ln21_unr12_stage5_stallmux_q_18_), .o(n25978) );
in01f01 g22188 ( .a(n25978), .o(n25979) );
no02f01 g22189 ( .a(n25979), .b(n25967), .o(n25980) );
no02f01 g22190 ( .a(n25980), .b(n25966), .o(n25981) );
na02f01 g22191 ( .a(n25980), .b(n25966), .o(n25982) );
in01f01 g22192 ( .a(n25982), .o(n25983) );
no02f01 g22193 ( .a(n25983), .b(n25981), .o(n25984) );
no02f01 g22194 ( .a(n25984), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_18_), .o(n25985) );
no02f01 g22195 ( .a(n25985), .b(n25977), .o(n25986) );
in01f01 g22196 ( .a(n25986), .o(n25987) );
no03f01 g22197 ( .a(n25987), .b(n16785), .c(n16831), .o(n25988) );
in01f01 g22198 ( .a(n25977), .o(n25989) );
ao12f01 g22199 ( .a(n16785), .b(n16786), .c(n16772), .o(n25990) );
in01f01 g22200 ( .a(n25990), .o(n25991) );
na02f01 g22201 ( .a(n25976), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_19_), .o(n25992) );
in01f01 g22202 ( .a(n25992), .o(n25993) );
na02f01 g22203 ( .a(n25984), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_18_), .o(n25994) );
in01f01 g22204 ( .a(n25994), .o(n25995) );
no02f01 g22205 ( .a(n25995), .b(n25993), .o(n25996) );
oa12f01 g22206 ( .a(n25996), .b(n25991), .c(n25985), .o(n25997) );
na02f01 g22207 ( .a(n25997), .b(n25989), .o(n25998) );
in01f01 g22208 ( .a(n25998), .o(n25999) );
no02f01 g22209 ( .a(n25999), .b(n25988), .o(n26000) );
in01f01 g22210 ( .a(n26000), .o(n26001) );
ao12f01 g22211 ( .a(n25969), .b(n25970), .c(n25968), .o(n26002) );
in01f01 g22212 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_21_), .o(n26003) );
in01f01 g22213 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_20_), .o(n26004) );
ao12f01 g22214 ( .a(n26002), .b(n26004), .c(n26003), .o(n26005) );
in01f01 g22215 ( .a(n26005), .o(n26006) );
no02f01 g22216 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_23_), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_22_), .o(n26007) );
oa12f01 g22217 ( .a(n26006), .b(n26007), .c(n26002), .o(n26008) );
in01f01 g22218 ( .a(n26002), .o(n26009) );
no02f01 g22219 ( .a(n26009), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_22_), .o(n26010) );
no02f01 g22220 ( .a(n26009), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_23_), .o(n26011) );
ao12f01 g22221 ( .a(n26009), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_20_), .c(delay_sub_ln21_0_unr11_stage5_stallmux_q_21_), .o(n26012) );
no03f01 g22222 ( .a(n26012), .b(n26011), .c(n26010), .o(n26013) );
oa12f01 g22223 ( .a(n26013), .b(n26008), .c(n26001), .o(n26014) );
no02f01 g22224 ( .a(n26009), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_26_), .o(n26015) );
ao12f01 g22225 ( .a(n26009), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_24_), .c(delay_sub_ln21_0_unr11_stage5_stallmux_q_25_), .o(n26016) );
no03f01 g22226 ( .a(n26016), .b(n26015), .c(n26014), .o(n26017) );
no02f01 g22227 ( .a(n26009), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_27_), .o(n26018) );
in01f01 g22228 ( .a(n26018), .o(n26019) );
na02f01 g22229 ( .a(n26019), .b(n26017), .o(n26020) );
no02f01 g22230 ( .a(n26009), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_28_), .o(n26021) );
no02f01 g22231 ( .a(n26021), .b(n26020), .o(n26022) );
in01f01 g22232 ( .a(n26022), .o(n26023) );
no02f01 g22233 ( .a(n26009), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_29_), .o(n26024) );
no02f01 g22234 ( .a(n26024), .b(n26023), .o(n26025) );
in01f01 g22235 ( .a(n26025), .o(n26026) );
no02f01 g22236 ( .a(n26009), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_30_), .o(n26027) );
na02f01 g22237 ( .a(n26009), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_30_), .o(n26028) );
in01f01 g22238 ( .a(n26028), .o(n26029) );
in01f01 g22239 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_26_), .o(n26030) );
in01f01 g22240 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_27_), .o(n26031) );
ao12f01 g22241 ( .a(n26002), .b(n26031), .c(n26030), .o(n26032) );
in01f01 g22242 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_25_), .o(n26033) );
in01f01 g22243 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_24_), .o(n26034) );
ao12f01 g22244 ( .a(n26002), .b(n26034), .c(n26033), .o(n26035) );
no02f01 g22245 ( .a(n26035), .b(n26032), .o(n26036) );
in01f01 g22246 ( .a(n26036), .o(n26037) );
in01f01 g22247 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_28_), .o(n26038) );
in01f01 g22248 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_29_), .o(n26039) );
ao12f01 g22249 ( .a(n26002), .b(n26039), .c(n26038), .o(n26040) );
no02f01 g22250 ( .a(n26040), .b(n26037), .o(n26041) );
in01f01 g22251 ( .a(n26041), .o(n26042) );
no02f01 g22252 ( .a(n26042), .b(n26029), .o(n26043) );
oa12f01 g22253 ( .a(n26043), .b(n26027), .c(n26026), .o(n26044) );
in01f01 g22254 ( .a(n26044), .o(n26045) );
no02f01 g22255 ( .a(n26009), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_31_), .o(n26046) );
na02f01 g22256 ( .a(n26009), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_31_), .o(n26047) );
in01f01 g22257 ( .a(n26047), .o(n26048) );
no02f01 g22258 ( .a(n26048), .b(n26046), .o(n26049) );
no02f01 g22259 ( .a(n26049), .b(n26045), .o(n26050) );
na02f01 g22260 ( .a(n26049), .b(n26045), .o(n26051) );
in01f01 g22261 ( .a(n26051), .o(n26052) );
no02f01 g22262 ( .a(n26052), .b(n26050), .o(n26053) );
no02f01 g22263 ( .a(n26053), .b(n25965), .o(n26054) );
in01f01 g22264 ( .a(n25964), .o(n26055) );
no02f01 g22265 ( .a(n26055), .b(n25962), .o(n26056) );
in01f01 g22266 ( .a(n26053), .o(n26057) );
no02f01 g22267 ( .a(n26057), .b(n26056), .o(n26058) );
no02f01 g22268 ( .a(n26058), .b(n26054), .o(n26059) );
no02f01 g22269 ( .a(n26009), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_24_), .o(n26060) );
no02f01 g22270 ( .a(n26060), .b(n26014), .o(n26061) );
no02f01 g22271 ( .a(n26002), .b(n26034), .o(n26062) );
no02f01 g22272 ( .a(n26062), .b(n26061), .o(n26063) );
no02f01 g22273 ( .a(n26002), .b(n26033), .o(n26064) );
no02f01 g22274 ( .a(n26009), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_25_), .o(n26065) );
no02f01 g22275 ( .a(n26065), .b(n26064), .o(n26066) );
na02f01 g22276 ( .a(n26066), .b(n26063), .o(n26067) );
in01f01 g22277 ( .a(n26067), .o(n26068) );
no02f01 g22278 ( .a(n26066), .b(n26063), .o(n26069) );
no02f01 g22279 ( .a(n26069), .b(n26068), .o(n26070) );
in01f01 g22280 ( .a(n26070), .o(n26071) );
in01f01 g22281 ( .a(n26014), .o(n26072) );
no02f01 g22282 ( .a(n26062), .b(n26060), .o(n26073) );
in01f01 g22283 ( .a(n26073), .o(n26074) );
na02f01 g22284 ( .a(n26074), .b(n26072), .o(n26075) );
in01f01 g22285 ( .a(n26075), .o(n26076) );
no02f01 g22286 ( .a(n26074), .b(n26072), .o(n26077) );
no02f01 g22287 ( .a(n26077), .b(n26076), .o(n26078) );
in01f01 g22288 ( .a(n26078), .o(n26079) );
ao12f01 g22289 ( .a(n26056), .b(n26079), .c(n26071), .o(n26080) );
in01f01 g22290 ( .a(n16785), .o(n26081) );
na02f01 g22291 ( .a(n26081), .b(n16771), .o(n26082) );
ao12f01 g22292 ( .a(n25985), .b(n25991), .c(n26082), .o(n26083) );
no02f01 g22293 ( .a(n25993), .b(n25977), .o(n26084) );
in01f01 g22294 ( .a(n26084), .o(n26085) );
no03f01 g22295 ( .a(n26085), .b(n26083), .c(n25995), .o(n26086) );
no02f01 g22296 ( .a(n16785), .b(n16831), .o(n26087) );
in01f01 g22297 ( .a(n25985), .o(n26088) );
oa12f01 g22298 ( .a(n26088), .b(n25990), .c(n26087), .o(n26089) );
ao12f01 g22299 ( .a(n26084), .b(n26089), .c(n25994), .o(n26090) );
no02f01 g22300 ( .a(n26090), .b(n26086), .o(n26091) );
na02f01 g22301 ( .a(n26091), .b(n25965), .o(n26092) );
in01f01 g22302 ( .a(n25961), .o(n26093) );
oa12f01 g22303 ( .a(n25941), .b(n17435), .c(n17474), .o(n26094) );
na02f01 g22304 ( .a(n26094), .b(n26093), .o(n26095) );
no02f01 g22305 ( .a(n26094), .b(n26093), .o(n26096) );
in01f01 g22306 ( .a(n26096), .o(n26097) );
no02f01 g22307 ( .a(n25990), .b(n26087), .o(n26098) );
no02f01 g22308 ( .a(n25995), .b(n25985), .o(n26099) );
in01f01 g22309 ( .a(n26099), .o(n26100) );
no02f01 g22310 ( .a(n26100), .b(n25990), .o(n26101) );
na02f01 g22311 ( .a(n26101), .b(n26082), .o(n26102) );
oa12f01 g22312 ( .a(n26102), .b(n26099), .c(n26098), .o(n26103) );
na03f01 g22313 ( .a(n26103), .b(n26097), .c(n26095), .o(n26104) );
no02f01 g22314 ( .a(n17791), .b(n17734), .o(n26105) );
ao12f01 g22315 ( .a(n16835), .b(n17476), .c(n17438), .o(n26106) );
no02f01 g22316 ( .a(n17724), .b(n26106), .o(n26107) );
ao12f01 g22317 ( .a(n26106), .b(n17727), .c(n17477), .o(n26108) );
ao12f01 g22318 ( .a(n26108), .b(n26107), .c(n26105), .o(n26109) );
ao12f01 g22319 ( .a(n26103), .b(n26097), .c(n26095), .o(n26110) );
oa12f01 g22320 ( .a(n26104), .b(n26110), .c(n26109), .o(n26111) );
no02f01 g22321 ( .a(n26091), .b(n25965), .o(n26112) );
oa12f01 g22322 ( .a(n26092), .b(n26112), .c(n26111), .o(n26113) );
no02f01 g22323 ( .a(n26002), .b(n26003), .o(n26114) );
no02f01 g22324 ( .a(n26009), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_21_), .o(n26115) );
no02f01 g22325 ( .a(n26115), .b(n26114), .o(n26116) );
in01f01 g22326 ( .a(n26116), .o(n26117) );
no02f01 g22327 ( .a(n26009), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_20_), .o(n26118) );
no02f01 g22328 ( .a(n26118), .b(n26000), .o(n26119) );
no02f01 g22329 ( .a(n26002), .b(n26004), .o(n26120) );
no02f01 g22330 ( .a(n26120), .b(n26119), .o(n26121) );
in01f01 g22331 ( .a(n26121), .o(n26122) );
no02f01 g22332 ( .a(n26122), .b(n26117), .o(n26123) );
no02f01 g22333 ( .a(n26121), .b(n26116), .o(n26124) );
no02f01 g22334 ( .a(n26124), .b(n26123), .o(n26125) );
in01f01 g22335 ( .a(n26125), .o(n26126) );
no02f01 g22336 ( .a(n26120), .b(n26118), .o(n26127) );
in01f01 g22337 ( .a(n26127), .o(n26128) );
no03f01 g22338 ( .a(n26128), .b(n25999), .c(n25988), .o(n26129) );
in01f01 g22339 ( .a(n26129), .o(n26130) );
oa12f01 g22340 ( .a(n26128), .b(n25999), .c(n25988), .o(n26131) );
na02f01 g22341 ( .a(n26131), .b(n26130), .o(n26132) );
ao12f01 g22342 ( .a(n26056), .b(n26132), .c(n26126), .o(n26133) );
no03f01 g22343 ( .a(n26012), .b(n25987), .c(n26082), .o(n26134) );
no02f01 g22344 ( .a(n26012), .b(n25998), .o(n26135) );
no02f01 g22345 ( .a(n26135), .b(n26134), .o(n26136) );
no02f01 g22346 ( .a(n26136), .b(n26010), .o(n26137) );
na02f01 g22347 ( .a(n26009), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_22_), .o(n26138) );
in01f01 g22348 ( .a(n26138), .o(n26139) );
no03f01 g22349 ( .a(n26139), .b(n26137), .c(n26005), .o(n26140) );
na02f01 g22350 ( .a(n26009), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_23_), .o(n26141) );
in01f01 g22351 ( .a(n26141), .o(n26142) );
no02f01 g22352 ( .a(n26142), .b(n26011), .o(n26143) );
na02f01 g22353 ( .a(n26143), .b(n26140), .o(n26144) );
no02f01 g22354 ( .a(n26143), .b(n26140), .o(n26145) );
in01f01 g22355 ( .a(n26145), .o(n26146) );
na02f01 g22356 ( .a(n26146), .b(n26144), .o(n26147) );
no02f01 g22357 ( .a(n26147), .b(n26056), .o(n26148) );
no02f01 g22358 ( .a(n26135), .b(n26005), .o(n26149) );
in01f01 g22359 ( .a(n26149), .o(n26150) );
no02f01 g22360 ( .a(n26150), .b(n26134), .o(n26151) );
no02f01 g22361 ( .a(n26139), .b(n26010), .o(n26152) );
in01f01 g22362 ( .a(n26134), .o(n26153) );
na03f01 g22363 ( .a(n26152), .b(n26149), .c(n26153), .o(n26154) );
oa12f01 g22364 ( .a(n26154), .b(n26152), .c(n26151), .o(n26155) );
no02f01 g22365 ( .a(n26155), .b(n26056), .o(n26156) );
no04f01 g22366 ( .a(n26156), .b(n26148), .c(n26133), .d(n26113), .o(n26157) );
in01f01 g22367 ( .a(n26132), .o(n26158) );
ao12f01 g22368 ( .a(n25965), .b(n26158), .c(n26125), .o(n26159) );
in01f01 g22369 ( .a(n26144), .o(n26160) );
no02f01 g22370 ( .a(n26145), .b(n26160), .o(n26161) );
in01f01 g22371 ( .a(n26155), .o(n26162) );
ao12f01 g22372 ( .a(n25965), .b(n26162), .c(n26161), .o(n26163) );
no02f01 g22373 ( .a(n26163), .b(n26159), .o(n26164) );
in01f01 g22374 ( .a(n26164), .o(n26165) );
no02f01 g22375 ( .a(n26165), .b(n26157), .o(n26166) );
no02f01 g22376 ( .a(n26166), .b(n26080), .o(n26167) );
no02f01 g22377 ( .a(n26002), .b(n26030), .o(n26168) );
no02f01 g22378 ( .a(n26168), .b(n26015), .o(n26169) );
in01f01 g22379 ( .a(n26016), .o(n26170) );
oa12f01 g22380 ( .a(n26170), .b(n26035), .c(n26072), .o(n26171) );
no02f01 g22381 ( .a(n26171), .b(n26169), .o(n26172) );
na02f01 g22382 ( .a(n26171), .b(n26169), .o(n26173) );
in01f01 g22383 ( .a(n26173), .o(n26174) );
no02f01 g22384 ( .a(n26174), .b(n26172), .o(n26175) );
in01f01 g22385 ( .a(n26175), .o(n26176) );
no02f01 g22386 ( .a(n26176), .b(n26056), .o(n26177) );
no03f01 g22387 ( .a(n26035), .b(n26168), .c(n26017), .o(n26178) );
in01f01 g22388 ( .a(n26178), .o(n26179) );
no02f01 g22389 ( .a(n26002), .b(n26031), .o(n26180) );
no02f01 g22390 ( .a(n26180), .b(n26018), .o(n26181) );
in01f01 g22391 ( .a(n26181), .o(n26182) );
no02f01 g22392 ( .a(n26182), .b(n26179), .o(n26183) );
no02f01 g22393 ( .a(n26181), .b(n26178), .o(n26184) );
no02f01 g22394 ( .a(n26184), .b(n26183), .o(n26185) );
in01f01 g22395 ( .a(n26185), .o(n26186) );
no02f01 g22396 ( .a(n26186), .b(n26056), .o(n26187) );
no02f01 g22397 ( .a(n26187), .b(n26177), .o(n26188) );
na02f01 g22398 ( .a(n26188), .b(n26167), .o(n26189) );
na02f01 g22399 ( .a(n26036), .b(n26020), .o(n26190) );
no02f01 g22400 ( .a(n26002), .b(n26038), .o(n26191) );
no02f01 g22401 ( .a(n26191), .b(n26021), .o(n26192) );
in01f01 g22402 ( .a(n26192), .o(n26193) );
na02f01 g22403 ( .a(n26193), .b(n26190), .o(n26194) );
no02f01 g22404 ( .a(n26193), .b(n26190), .o(n26195) );
in01f01 g22405 ( .a(n26195), .o(n26196) );
na02f01 g22406 ( .a(n26196), .b(n26194), .o(n26197) );
no02f01 g22407 ( .a(n26197), .b(n26056), .o(n26198) );
no02f01 g22408 ( .a(n26002), .b(n26039), .o(n26199) );
no02f01 g22409 ( .a(n26199), .b(n26024), .o(n26200) );
in01f01 g22410 ( .a(n26200), .o(n26201) );
no03f01 g22411 ( .a(n26191), .b(n26037), .c(n26022), .o(n26202) );
in01f01 g22412 ( .a(n26202), .o(n26203) );
no02f01 g22413 ( .a(n26203), .b(n26201), .o(n26204) );
no02f01 g22414 ( .a(n26202), .b(n26200), .o(n26205) );
no02f01 g22415 ( .a(n26205), .b(n26204), .o(n26206) );
in01f01 g22416 ( .a(n26206), .o(n26207) );
no02f01 g22417 ( .a(n26207), .b(n26056), .o(n26208) );
no02f01 g22418 ( .a(n26208), .b(n26198), .o(n26209) );
no02f01 g22419 ( .a(n26042), .b(n26025), .o(n26210) );
no02f01 g22420 ( .a(n26029), .b(n26027), .o(n26211) );
no02f01 g22421 ( .a(n26211), .b(n26210), .o(n26212) );
na02f01 g22422 ( .a(n26211), .b(n26210), .o(n26213) );
in01f01 g22423 ( .a(n26213), .o(n26214) );
no02f01 g22424 ( .a(n26214), .b(n26212), .o(n26215) );
in01f01 g22425 ( .a(n26215), .o(n26216) );
no02f01 g22426 ( .a(n26216), .b(n26056), .o(n26217) );
in01f01 g22427 ( .a(n26217), .o(n26218) );
na02f01 g22428 ( .a(n26218), .b(n26209), .o(n26219) );
ao12f01 g22429 ( .a(n25965), .b(n26078), .c(n26070), .o(n26220) );
ao12f01 g22430 ( .a(n25965), .b(n26185), .c(n26175), .o(n26221) );
no02f01 g22431 ( .a(n26221), .b(n26220), .o(n26222) );
in01f01 g22432 ( .a(n26222), .o(n26223) );
no02f01 g22433 ( .a(n26207), .b(n26197), .o(n26224) );
ao12f01 g22434 ( .a(n25965), .b(n26224), .c(n26215), .o(n26225) );
no02f01 g22435 ( .a(n26225), .b(n26223), .o(n26226) );
oa12f01 g22436 ( .a(n26226), .b(n26219), .c(n26189), .o(n26227) );
in01f01 g22437 ( .a(n26227), .o(n26228) );
no02f01 g22438 ( .a(n26228), .b(n26059), .o(n26229) );
na02f01 g22439 ( .a(n26228), .b(n26059), .o(n26230) );
in01f01 g22440 ( .a(n26230), .o(n26231) );
no02f01 g22441 ( .a(n26231), .b(n26229), .o(n26232) );
no02f01 g22442 ( .a(n26232), .b(n7682), .o(n26233) );
no02f01 g22443 ( .a(n26232), .b(n7712), .o(n26234) );
no02f01 g22444 ( .a(n26234), .b(n26233), .o(n26235) );
in01f01 g22445 ( .a(n26198), .o(n26236) );
ao12f01 g22446 ( .a(n26223), .b(n26188), .c(n26167), .o(n26237) );
in01f01 g22447 ( .a(n26194), .o(n26238) );
no02f01 g22448 ( .a(n26195), .b(n26238), .o(n26239) );
no02f01 g22449 ( .a(n26239), .b(n25965), .o(n26240) );
in01f01 g22450 ( .a(n26240), .o(n26241) );
na02f01 g22451 ( .a(n26241), .b(n26237), .o(n26242) );
no02f01 g22452 ( .a(n26206), .b(n25965), .o(n26243) );
no02f01 g22453 ( .a(n26243), .b(n26208), .o(n26244) );
in01f01 g22454 ( .a(n26244), .o(n26245) );
ao12f01 g22455 ( .a(n26245), .b(n26242), .c(n26236), .o(n26246) );
na02f01 g22456 ( .a(n26222), .b(n26189), .o(n26247) );
no02f01 g22457 ( .a(n26240), .b(n26247), .o(n26248) );
no03f01 g22458 ( .a(n26244), .b(n26248), .c(n26198), .o(n26249) );
no02f01 g22459 ( .a(n26249), .b(n26246), .o(n26250) );
no02f01 g22460 ( .a(n26250), .b(n7712), .o(n26251) );
no02f01 g22461 ( .a(n26240), .b(n26198), .o(n26252) );
no02f01 g22462 ( .a(n26252), .b(n26237), .o(n26253) );
na02f01 g22463 ( .a(n26252), .b(n26237), .o(n26254) );
in01f01 g22464 ( .a(n26254), .o(n26255) );
no02f01 g22465 ( .a(n26255), .b(n26253), .o(n26256) );
no02f01 g22466 ( .a(n26256), .b(n7712), .o(n26257) );
in01f01 g22467 ( .a(n26257), .o(n26258) );
in01f01 g22468 ( .a(n26177), .o(n26259) );
no02f01 g22469 ( .a(n26185), .b(n25965), .o(n26260) );
no02f01 g22470 ( .a(n26260), .b(n26187), .o(n26261) );
in01f01 g22471 ( .a(n26261), .o(n26262) );
no02f01 g22472 ( .a(n26175), .b(n25965), .o(n26263) );
in01f01 g22473 ( .a(n26263), .o(n26264) );
no02f01 g22474 ( .a(n26220), .b(n26167), .o(n26265) );
na02f01 g22475 ( .a(n26265), .b(n26264), .o(n26266) );
ao12f01 g22476 ( .a(n26262), .b(n26266), .c(n26259), .o(n26267) );
in01f01 g22477 ( .a(n26220), .o(n26268) );
oa12f01 g22478 ( .a(n26268), .b(n26166), .c(n26080), .o(n26269) );
no02f01 g22479 ( .a(n26269), .b(n26263), .o(n26270) );
no03f01 g22480 ( .a(n26270), .b(n26261), .c(n26177), .o(n26271) );
no02f01 g22481 ( .a(n26271), .b(n26267), .o(n26272) );
no02f01 g22482 ( .a(n26272), .b(n7712), .o(n26273) );
na03f01 g22483 ( .a(n26084), .b(n26089), .c(n25994), .o(n26274) );
oa12f01 g22484 ( .a(n26085), .b(n26083), .c(n25995), .o(n26275) );
na02f01 g22485 ( .a(n26275), .b(n26274), .o(n26276) );
na02f01 g22486 ( .a(n26276), .b(n26056), .o(n26277) );
na02f01 g22487 ( .a(n26277), .b(n26092), .o(n26278) );
no02f01 g22488 ( .a(n26278), .b(n26111), .o(n26279) );
no04f01 g22489 ( .a(n17724), .b(n17791), .c(n17734), .d(n26106), .o(n26280) );
in01f01 g22490 ( .a(n26095), .o(n26281) );
in01f01 g22491 ( .a(n26103), .o(n26282) );
oa12f01 g22492 ( .a(n26282), .b(n26096), .c(n26281), .o(n26283) );
oa12f01 g22493 ( .a(n26283), .b(n26108), .c(n26280), .o(n26284) );
no02f01 g22494 ( .a(n26276), .b(n26056), .o(n26285) );
no02f01 g22495 ( .a(n26112), .b(n26285), .o(n26286) );
ao12f01 g22496 ( .a(n26286), .b(n26284), .c(n26104), .o(n26287) );
oa12f01 g22497 ( .a(n7712), .b(n26287), .c(n26279), .o(n26288) );
na02f01 g22498 ( .a(n26283), .b(n26104), .o(n26289) );
no03f01 g22499 ( .a(n26289), .b(n26108), .c(n26280), .o(n26290) );
no03f01 g22500 ( .a(n26282), .b(n26096), .c(n26281), .o(n26291) );
no02f01 g22501 ( .a(n26110), .b(n26291), .o(n26292) );
no02f01 g22502 ( .a(n26292), .b(n26109), .o(n26293) );
oa12f01 g22503 ( .a(n7712), .b(n26293), .c(n26290), .o(n26294) );
na02f01 g22504 ( .a(n26294), .b(n26288), .o(n26295) );
na03f01 g22505 ( .a(n26107), .b(n17716), .c(n17498), .o(n26296) );
in01f01 g22506 ( .a(n26108), .o(n26297) );
ao12f01 g22507 ( .a(n26110), .b(n26297), .c(n26296), .o(n26298) );
no03f01 g22508 ( .a(n26112), .b(n26298), .c(n26291), .o(n26299) );
no02f01 g22509 ( .a(n26158), .b(n25965), .o(n26300) );
no02f01 g22510 ( .a(n26132), .b(n26056), .o(n26301) );
no02f01 g22511 ( .a(n26301), .b(n26300), .o(n26302) );
no03f01 g22512 ( .a(n26302), .b(n26299), .c(n26285), .o(n26303) );
na03f01 g22513 ( .a(n26277), .b(n26284), .c(n26104), .o(n26304) );
in01f01 g22514 ( .a(n26302), .o(n26305) );
ao12f01 g22515 ( .a(n26305), .b(n26304), .c(n26092), .o(n26306) );
oa12f01 g22516 ( .a(n7682), .b(n26306), .c(n26303), .o(n26307) );
na03f01 g22517 ( .a(n26286), .b(n26284), .c(n26104), .o(n26308) );
na02f01 g22518 ( .a(n26278), .b(n26111), .o(n26309) );
ao12f01 g22519 ( .a(n7712), .b(n26309), .c(n26308), .o(n26310) );
no02f01 g22520 ( .a(n17838), .b(n17796), .o(n26311) );
na02f01 g22521 ( .a(n17839), .b(n17826), .o(n26312) );
oa12f01 g22522 ( .a(n7682), .b(n26293), .c(n26290), .o(n26313) );
oa12f01 g22523 ( .a(n26313), .b(n26312), .c(n26311), .o(n26314) );
no02f01 g22524 ( .a(n26314), .b(n26310), .o(n26315) );
ao12f01 g22525 ( .a(n26295), .b(n26315), .c(n26307), .o(n26316) );
no02f01 g22526 ( .a(n26126), .b(n26056), .o(n26317) );
no02f01 g22527 ( .a(n26125), .b(n25965), .o(n26318) );
no02f01 g22528 ( .a(n26318), .b(n26317), .o(n26319) );
in01f01 g22529 ( .a(n26319), .o(n26320) );
no03f01 g22530 ( .a(n26301), .b(n26299), .c(n26285), .o(n26321) );
no03f01 g22531 ( .a(n26321), .b(n26320), .c(n26300), .o(n26322) );
in01f01 g22532 ( .a(n26300), .o(n26323) );
in01f01 g22533 ( .a(n26301), .o(n26324) );
na03f01 g22534 ( .a(n26324), .b(n26304), .c(n26092), .o(n26325) );
ao12f01 g22535 ( .a(n26319), .b(n26325), .c(n26323), .o(n26326) );
no02f01 g22536 ( .a(n26326), .b(n26322), .o(n26327) );
no02f01 g22537 ( .a(n26327), .b(n7712), .o(n26328) );
no02f01 g22538 ( .a(n26328), .b(n26316), .o(n26329) );
na03f01 g22539 ( .a(n26305), .b(n26304), .c(n26092), .o(n26330) );
oa12f01 g22540 ( .a(n26302), .b(n26299), .c(n26285), .o(n26331) );
na02f01 g22541 ( .a(n26331), .b(n26330), .o(n26332) );
na02f01 g22542 ( .a(n26332), .b(n7712), .o(n26333) );
na03f01 g22543 ( .a(n26325), .b(n26319), .c(n26323), .o(n26334) );
oa12f01 g22544 ( .a(n26320), .b(n26321), .c(n26300), .o(n26335) );
na02f01 g22545 ( .a(n26335), .b(n26334), .o(n26336) );
na02f01 g22546 ( .a(n26336), .b(n7712), .o(n26337) );
na02f01 g22547 ( .a(n26337), .b(n26333), .o(n26338) );
in01f01 g22548 ( .a(n26159), .o(n26339) );
oa12f01 g22549 ( .a(n26339), .b(n26133), .c(n26113), .o(n26340) );
no02f01 g22550 ( .a(n26162), .b(n25965), .o(n26341) );
no02f01 g22551 ( .a(n26341), .b(n26156), .o(n26342) );
in01f01 g22552 ( .a(n26342), .o(n26343) );
na02f01 g22553 ( .a(n26343), .b(n26340), .o(n26344) );
no02f01 g22554 ( .a(n26343), .b(n26340), .o(n26345) );
in01f01 g22555 ( .a(n26345), .o(n26346) );
na02f01 g22556 ( .a(n26346), .b(n26344), .o(n26347) );
na02f01 g22557 ( .a(n26347), .b(n7682), .o(n26348) );
oa12f01 g22558 ( .a(n26348), .b(n26338), .c(n26329), .o(n26349) );
no02f01 g22559 ( .a(n26161), .b(n25965), .o(n26350) );
no02f01 g22560 ( .a(n26350), .b(n26148), .o(n26351) );
no02f01 g22561 ( .a(n26340), .b(n26341), .o(n26352) );
no03f01 g22562 ( .a(n26352), .b(n26351), .c(n26156), .o(n26353) );
in01f01 g22563 ( .a(n26156), .o(n26354) );
in01f01 g22564 ( .a(n26351), .o(n26355) );
no02f01 g22565 ( .a(n26299), .b(n26285), .o(n26356) );
in01f01 g22566 ( .a(n26133), .o(n26357) );
ao12f01 g22567 ( .a(n26159), .b(n26357), .c(n26356), .o(n26358) );
oa12f01 g22568 ( .a(n26358), .b(n26162), .c(n25965), .o(n26359) );
ao12f01 g22569 ( .a(n26355), .b(n26359), .c(n26354), .o(n26360) );
no02f01 g22570 ( .a(n26360), .b(n26353), .o(n26361) );
no02f01 g22571 ( .a(n26361), .b(n7712), .o(n26362) );
no02f01 g22572 ( .a(n26156), .b(n26148), .o(n26363) );
na03f01 g22573 ( .a(n26363), .b(n26357), .c(n26356), .o(n26364) );
na02f01 g22574 ( .a(n26164), .b(n26364), .o(n26365) );
no02f01 g22575 ( .a(n26079), .b(n26056), .o(n26366) );
no02f01 g22576 ( .a(n26078), .b(n25965), .o(n26367) );
no02f01 g22577 ( .a(n26367), .b(n26366), .o(n26368) );
in01f01 g22578 ( .a(n26368), .o(n26369) );
na02f01 g22579 ( .a(n26369), .b(n26365), .o(n26370) );
in01f01 g22580 ( .a(n26370), .o(n26371) );
no02f01 g22581 ( .a(n26369), .b(n26365), .o(n26372) );
no02f01 g22582 ( .a(n26372), .b(n26371), .o(n26373) );
no02f01 g22583 ( .a(n26373), .b(n7712), .o(n26374) );
in01f01 g22584 ( .a(n26367), .o(n26375) );
no02f01 g22585 ( .a(n26071), .b(n26056), .o(n26376) );
no02f01 g22586 ( .a(n26070), .b(n25965), .o(n26377) );
no02f01 g22587 ( .a(n26377), .b(n26376), .o(n26378) );
in01f01 g22588 ( .a(n26366), .o(n26379) );
oa12f01 g22589 ( .a(n26379), .b(n26165), .c(n26157), .o(n26380) );
na03f01 g22590 ( .a(n26380), .b(n26378), .c(n26375), .o(n26381) );
in01f01 g22591 ( .a(n26378), .o(n26382) );
ao12f01 g22592 ( .a(n26366), .b(n26164), .c(n26364), .o(n26383) );
oa12f01 g22593 ( .a(n26382), .b(n26383), .c(n26367), .o(n26384) );
ao12f01 g22594 ( .a(n7712), .b(n26384), .c(n26381), .o(n26385) );
no04f01 g22595 ( .a(n26385), .b(n26374), .c(n26362), .d(n26349), .o(n26386) );
no02f01 g22596 ( .a(n26342), .b(n26358), .o(n26387) );
no02f01 g22597 ( .a(n26345), .b(n26387), .o(n26388) );
no02f01 g22598 ( .a(n26388), .b(n7682), .o(n26389) );
in01f01 g22599 ( .a(n26389), .o(n26390) );
na03f01 g22600 ( .a(n26359), .b(n26355), .c(n26354), .o(n26391) );
oa12f01 g22601 ( .a(n26351), .b(n26352), .c(n26156), .o(n26392) );
na02f01 g22602 ( .a(n26392), .b(n26391), .o(n26393) );
na02f01 g22603 ( .a(n26393), .b(n7712), .o(n26394) );
in01f01 g22604 ( .a(n26372), .o(n26395) );
na02f01 g22605 ( .a(n26395), .b(n26370), .o(n26396) );
na02f01 g22606 ( .a(n26396), .b(n7712), .o(n26397) );
no03f01 g22607 ( .a(n26383), .b(n26382), .c(n26367), .o(n26398) );
ao12f01 g22608 ( .a(n26378), .b(n26380), .c(n26375), .o(n26399) );
oa12f01 g22609 ( .a(n7712), .b(n26399), .c(n26398), .o(n26400) );
na04f01 g22610 ( .a(n26400), .b(n26397), .c(n26394), .d(n26390), .o(n26401) );
no02f01 g22611 ( .a(n26263), .b(n26177), .o(n26402) );
in01f01 g22612 ( .a(n26402), .o(n26403) );
na02f01 g22613 ( .a(n26403), .b(n26269), .o(n26404) );
in01f01 g22614 ( .a(n26404), .o(n26405) );
no02f01 g22615 ( .a(n26403), .b(n26269), .o(n26406) );
no02f01 g22616 ( .a(n26406), .b(n26405), .o(n26407) );
oa22f01 g22617 ( .a(n26407), .b(n7712), .c(n26401), .d(n26386), .o(n26408) );
oa12f01 g22618 ( .a(n26261), .b(n26270), .c(n26177), .o(n26409) );
in01f01 g22619 ( .a(n26271), .o(n26410) );
na02f01 g22620 ( .a(n26410), .b(n26409), .o(n26411) );
in01f01 g22621 ( .a(n26406), .o(n26412) );
na02f01 g22622 ( .a(n26412), .b(n26404), .o(n26413) );
oa12f01 g22623 ( .a(n7712), .b(n26413), .c(n26411), .o(n26414) );
oa12f01 g22624 ( .a(n26414), .b(n26408), .c(n26273), .o(n26415) );
ao12f01 g22625 ( .a(n7682), .b(n26256), .c(n26250), .o(n26416) );
ao12f01 g22626 ( .a(n26416), .b(n26415), .c(n26258), .o(n26417) );
no02f01 g22627 ( .a(n26417), .b(n26251), .o(n26418) );
no02f01 g22628 ( .a(n26215), .b(n25965), .o(n26419) );
no02f01 g22629 ( .a(n26419), .b(n26217), .o(n26420) );
in01f01 g22630 ( .a(n26420), .o(n26421) );
no02f01 g22631 ( .a(n26224), .b(n25965), .o(n26422) );
ao12f01 g22632 ( .a(n26422), .b(n26247), .c(n26209), .o(n26423) );
in01f01 g22633 ( .a(n26423), .o(n26424) );
no02f01 g22634 ( .a(n26424), .b(n26421), .o(n26425) );
in01f01 g22635 ( .a(n26425), .o(n26426) );
na02f01 g22636 ( .a(n26424), .b(n26421), .o(n26427) );
na02f01 g22637 ( .a(n26427), .b(n26426), .o(n26428) );
na02f01 g22638 ( .a(n26428), .b(n7682), .o(n26429) );
in01f01 g22639 ( .a(n26429), .o(n26430) );
no02f01 g22640 ( .a(n26430), .b(n26234), .o(n26431) );
na02f01 g22641 ( .a(n26431), .b(n26418), .o(n26432) );
na02f01 g22642 ( .a(n26428), .b(n7712), .o(n26433) );
in01f01 g22643 ( .a(n26433), .o(n26434) );
no02f01 g22644 ( .a(n26434), .b(n26233), .o(n26435) );
na03f01 g22645 ( .a(n26435), .b(n26432), .c(n26235), .o(n26436) );
in01f01 g22646 ( .a(n26436), .o(n26437) );
in01f01 g22647 ( .a(n26428), .o(n26438) );
no02f01 g22648 ( .a(n26232), .b(n7682), .o(n26439) );
no02f01 g22649 ( .a(n26439), .b(n26437), .o(n26440) );
in01f01 g22650 ( .a(n26440), .o(n26441) );
in01f01 g22651 ( .a(n17433), .o(n26442) );
ao12f01 g22652 ( .a(n_17093), .b(n26215), .c(n26206), .o(n26443) );
in01f01 g22653 ( .a(n26443), .o(n26444) );
no02f01 g22654 ( .a(n17846), .b(n17844), .o(n26445) );
na02f01 g22655 ( .a(n17723), .b(n_17093), .o(n26446) );
na02f01 g22656 ( .a(n26446), .b(n26445), .o(n26447) );
ao12f01 g22657 ( .a(n26447), .b(n16835), .c(n_17093), .o(n26448) );
oa12f01 g22658 ( .a(n26448), .b(n26282), .c(n7550), .o(n26449) );
ao12f01 g22659 ( .a(n26449), .b(n26276), .c(n_17093), .o(n26450) );
in01f01 g22660 ( .a(n26131), .o(n26451) );
no03f01 g22661 ( .a(n26451), .b(n26129), .c(n7550), .o(n26452) );
ao12f01 g22662 ( .a(n_17093), .b(n26131), .c(n26130), .o(n26453) );
no02f01 g22663 ( .a(n26453), .b(n26452), .o(n26454) );
oa12f01 g22664 ( .a(n7550), .b(n26090), .c(n26086), .o(n26455) );
na02f01 g22665 ( .a(n26455), .b(n26454), .o(n26456) );
oa12f01 g22666 ( .a(n7550), .b(n26456), .c(n26450), .o(n26457) );
na03f01 g22667 ( .a(n26131), .b(n26130), .c(n_17093), .o(n26458) );
oa12f01 g22668 ( .a(n7550), .b(n26451), .c(n26129), .o(n26459) );
na02f01 g22669 ( .a(n26459), .b(n26458), .o(n26460) );
oa12f01 g22670 ( .a(n7550), .b(n26103), .c(n16835), .o(n26461) );
in01f01 g22671 ( .a(n26461), .o(n26462) );
ao12f01 g22672 ( .a(n26462), .b(n26460), .c(n26450), .o(n26463) );
ao22f01 g22673 ( .a(n26463), .b(n26457), .c(n26126), .d(n_17093), .o(n26464) );
na02f01 g22674 ( .a(n26155), .b(n_17093), .o(n26465) );
na02f01 g22675 ( .a(n26147), .b(n_17093), .o(n26466) );
no02f01 g22676 ( .a(n26078), .b(n7550), .o(n26467) );
in01f01 g22677 ( .a(n26467), .o(n26468) );
na04f01 g22678 ( .a(n26468), .b(n26466), .c(n26465), .d(n26464), .o(n26469) );
ao12f01 g22679 ( .a(n_17093), .b(n26162), .c(n26125), .o(n26470) );
ao12f01 g22680 ( .a(n_17093), .b(n26161), .c(n26078), .o(n26471) );
no02f01 g22681 ( .a(n26471), .b(n26470), .o(n26472) );
na02f01 g22682 ( .a(n26472), .b(n26469), .o(n26473) );
oa12f01 g22683 ( .a(n_17093), .b(n26176), .c(n26071), .o(n26474) );
no02f01 g22684 ( .a(n26185), .b(n7550), .o(n26475) );
in01f01 g22685 ( .a(n26475), .o(n26476) );
na03f01 g22686 ( .a(n26476), .b(n26474), .c(n26473), .o(n26477) );
na02f01 g22687 ( .a(n26239), .b(n_17093), .o(n26478) );
na02f01 g22688 ( .a(n26197), .b(n7550), .o(n26479) );
na02f01 g22689 ( .a(n26479), .b(n26478), .o(n26480) );
no02f01 g22690 ( .a(n26185), .b(n_17093), .o(n26481) );
no02f01 g22691 ( .a(n26481), .b(n26480), .o(n26482) );
na02f01 g22692 ( .a(n26482), .b(n26477), .o(n26483) );
na02f01 g22693 ( .a(n26483), .b(n7550), .o(n26484) );
in01f01 g22694 ( .a(n26480), .o(n26485) );
ao12f01 g22695 ( .a(n_17093), .b(n26175), .c(n26070), .o(n26486) );
in01f01 g22696 ( .a(n26486), .o(n26487) );
oa12f01 g22697 ( .a(n26487), .b(n26485), .c(n26477), .o(n26488) );
in01f01 g22698 ( .a(n26488), .o(n26489) );
na02f01 g22699 ( .a(n26489), .b(n26484), .o(n26490) );
no02f01 g22700 ( .a(n26206), .b(n7550), .o(n26491) );
in01f01 g22701 ( .a(n26491), .o(n26492) );
na02f01 g22702 ( .a(n26492), .b(n26490), .o(n26493) );
no02f01 g22703 ( .a(n26215), .b(n7550), .o(n26494) );
oa12f01 g22704 ( .a(n26444), .b(n26494), .c(n26493), .o(n26495) );
oa12f01 g22705 ( .a(n7550), .b(n26495), .c(n26057), .o(n26496) );
no02f01 g22706 ( .a(n26494), .b(n26493), .o(n26497) );
na03f01 g22707 ( .a(n26497), .b(n26053), .c(n_17093), .o(n26498) );
na03f01 g22708 ( .a(n26498), .b(n26496), .c(n26053), .o(n26499) );
no02f01 g22709 ( .a(n26053), .b(n_17093), .o(n26500) );
in01f01 g22710 ( .a(n26500), .o(n26501) );
na02f01 g22711 ( .a(n26501), .b(n26499), .o(n26502) );
no02f01 g22712 ( .a(n26502), .b(n26442), .o(n26503) );
in01f01 g22713 ( .a(n26502), .o(n26504) );
no02f01 g22714 ( .a(n26504), .b(n17433), .o(n26505) );
no02f01 g22715 ( .a(n26505), .b(n26503), .o(n26506) );
in01f01 g22716 ( .a(n26506), .o(n26507) );
ao12f01 g22717 ( .a(n26504), .b(n17416), .c(n17401), .o(n26508) );
no02f01 g22718 ( .a(n26206), .b(n_17093), .o(n26509) );
ao12f01 g22719 ( .a(n26488), .b(n26483), .c(n7550), .o(n26510) );
no02f01 g22720 ( .a(n26491), .b(n26510), .o(n26511) );
no03f01 g22721 ( .a(n26511), .b(n26509), .c(n26216), .o(n26512) );
oa12f01 g22722 ( .a(n26216), .b(n26511), .c(n26509), .o(n26513) );
in01f01 g22723 ( .a(n26513), .o(n26514) );
no03f01 g22724 ( .a(n26514), .b(n26512), .c(n17200), .o(n26515) );
in01f01 g22725 ( .a(n26515), .o(n26516) );
no02f01 g22726 ( .a(n26491), .b(n26509), .o(n26517) );
na02f01 g22727 ( .a(n26517), .b(n26510), .o(n26518) );
in01f01 g22728 ( .a(n26518), .o(n26519) );
no02f01 g22729 ( .a(n26517), .b(n26510), .o(n26520) );
oa12f01 g22730 ( .a(n17260), .b(n26520), .c(n26519), .o(n26521) );
in01f01 g22731 ( .a(n26474), .o(n26522) );
no03f01 g22732 ( .a(n26486), .b(n26471), .c(n26470), .o(n26523) );
oa12f01 g22733 ( .a(n26523), .b(n26522), .c(n26469), .o(n26524) );
oa12f01 g22734 ( .a(n26476), .b(n26524), .c(n26481), .o(n26525) );
na02f01 g22735 ( .a(n26525), .b(n26239), .o(n26526) );
in01f01 g22736 ( .a(n26526), .o(n26527) );
no02f01 g22737 ( .a(n26525), .b(n26239), .o(n26528) );
no03f01 g22738 ( .a(n26528), .b(n26527), .c(n17214), .o(n26529) );
in01f01 g22739 ( .a(n26529), .o(n26530) );
no02f01 g22740 ( .a(n26070), .b(n_17093), .o(n26531) );
no02f01 g22741 ( .a(n26070), .b(n7550), .o(n26532) );
ao12f01 g22742 ( .a(n26532), .b(n26472), .c(n26469), .o(n26533) );
no03f01 g22743 ( .a(n26533), .b(n26531), .c(n26176), .o(n26534) );
oa12f01 g22744 ( .a(n26176), .b(n26533), .c(n26531), .o(n26535) );
in01f01 g22745 ( .a(n26535), .o(n26536) );
no03f01 g22746 ( .a(n26536), .b(n26534), .c(n17268), .o(n26537) );
in01f01 g22747 ( .a(n26537), .o(n26538) );
na02f01 g22748 ( .a(n26465), .b(n26464), .o(n26539) );
in01f01 g22749 ( .a(n26466), .o(n26540) );
ao12f01 g22750 ( .a(n26470), .b(n26147), .c(n7550), .o(n26541) );
oa12f01 g22751 ( .a(n26541), .b(n26540), .c(n26539), .o(n26542) );
na02f01 g22752 ( .a(n26542), .b(n26079), .o(n26543) );
no02f01 g22753 ( .a(n26542), .b(n26079), .o(n26544) );
in01f01 g22754 ( .a(n26544), .o(n26545) );
no02f01 g22755 ( .a(n17087), .b(n16969), .o(n26546) );
no02f01 g22756 ( .a(n17089), .b(n16960), .o(n26547) );
no02f01 g22757 ( .a(n26547), .b(n26546), .o(n26548) );
na02f01 g22758 ( .a(n26547), .b(n26546), .o(n26549) );
in01f01 g22759 ( .a(n26549), .o(n26550) );
no02f01 g22760 ( .a(n26550), .b(n26548), .o(n26551) );
na03f01 g22761 ( .a(n26551), .b(n26545), .c(n26543), .o(n26552) );
in01f01 g22762 ( .a(n26552), .o(n26553) );
in01f01 g22763 ( .a(n26470), .o(n26554) );
na03f01 g22764 ( .a(n26554), .b(n26539), .c(n26161), .o(n26555) );
in01f01 g22765 ( .a(n26555), .o(n26556) );
ao12f01 g22766 ( .a(n26161), .b(n26554), .c(n26539), .o(n26557) );
na02f01 g22767 ( .a(n17172), .b(n17145), .o(n26558) );
no02f01 g22768 ( .a(n17086), .b(n16969), .o(n26559) );
no02f01 g22769 ( .a(n26559), .b(n26558), .o(n26560) );
na02f01 g22770 ( .a(n26559), .b(n26558), .o(n26561) );
in01f01 g22771 ( .a(n26561), .o(n26562) );
no02f01 g22772 ( .a(n26562), .b(n26560), .o(n26563) );
in01f01 g22773 ( .a(n26563), .o(n26564) );
oa12f01 g22774 ( .a(n26564), .b(n26557), .c(n26556), .o(n26565) );
na02f01 g22775 ( .a(n17850), .b(n17848), .o(n26566) );
no02f01 g22776 ( .a(n17843), .b(n7550), .o(n26567) );
no02f01 g22777 ( .a(n26567), .b(n26566), .o(n26568) );
oa12f01 g22778 ( .a(n26568), .b(n17479), .c(n7550), .o(n26569) );
ao12f01 g22779 ( .a(n26569), .b(n26103), .c(n_17093), .o(n26570) );
oa12f01 g22780 ( .a(n26570), .b(n26091), .c(n7550), .o(n26571) );
no02f01 g22781 ( .a(n26091), .b(n_17093), .o(n26572) );
no02f01 g22782 ( .a(n26572), .b(n26460), .o(n26573) );
ao12f01 g22783 ( .a(n_17093), .b(n26573), .c(n26571), .o(n26574) );
oa12f01 g22784 ( .a(n26461), .b(n26454), .c(n26571), .o(n26575) );
oa22f01 g22785 ( .a(n26575), .b(n26574), .c(n26125), .d(n7550), .o(n26576) );
no02f01 g22786 ( .a(n26125), .b(n_17093), .o(n26577) );
in01f01 g22787 ( .a(n26577), .o(n26578) );
na03f01 g22788 ( .a(n26578), .b(n26576), .c(n26162), .o(n26579) );
oa12f01 g22789 ( .a(n26155), .b(n26577), .c(n26464), .o(n26580) );
no02f01 g22790 ( .a(n17081), .b(n16989), .o(n26581) );
no02f01 g22791 ( .a(n17083), .b(n16978), .o(n26582) );
no02f01 g22792 ( .a(n26582), .b(n26581), .o(n26583) );
na02f01 g22793 ( .a(n26582), .b(n26581), .o(n26584) );
in01f01 g22794 ( .a(n26584), .o(n26585) );
no02f01 g22795 ( .a(n26585), .b(n26583), .o(n26586) );
na03f01 g22796 ( .a(n26586), .b(n26580), .c(n26579), .o(n26587) );
ao12f01 g22797 ( .a(n26586), .b(n26580), .c(n26579), .o(n26588) );
no03f01 g22798 ( .a(n26575), .b(n26574), .c(n26126), .o(n26589) );
ao12f01 g22799 ( .a(n26125), .b(n26463), .c(n26457), .o(n26590) );
no02f01 g22800 ( .a(n17079), .b(n16998), .o(n26591) );
no02f01 g22801 ( .a(n17080), .b(n16989), .o(n26592) );
in01f01 g22802 ( .a(n26592), .o(n26593) );
no02f01 g22803 ( .a(n26593), .b(n26591), .o(n26594) );
na02f01 g22804 ( .a(n26593), .b(n26591), .o(n26595) );
in01f01 g22805 ( .a(n26595), .o(n26596) );
no02f01 g22806 ( .a(n26596), .b(n26594), .o(n26597) );
in01f01 g22807 ( .a(n26597), .o(n26598) );
oa12f01 g22808 ( .a(n26598), .b(n26590), .c(n26589), .o(n26599) );
no03f01 g22809 ( .a(n26598), .b(n26590), .c(n26589), .o(n26600) );
na02f01 g22810 ( .a(n26461), .b(n26455), .o(n26601) );
in01f01 g22811 ( .a(n26601), .o(n26602) );
na03f01 g22812 ( .a(n26602), .b(n26571), .c(n26158), .o(n26603) );
oa12f01 g22813 ( .a(n26132), .b(n26601), .c(n26450), .o(n26604) );
no02f01 g22814 ( .a(n17078), .b(n17011), .o(n26605) );
no02f01 g22815 ( .a(n17000), .b(n16998), .o(n26606) );
no02f01 g22816 ( .a(n26606), .b(n26605), .o(n26607) );
na02f01 g22817 ( .a(n26606), .b(n26605), .o(n26608) );
in01f01 g22818 ( .a(n26608), .o(n26609) );
no02f01 g22819 ( .a(n26609), .b(n26607), .o(n26610) );
ao12f01 g22820 ( .a(n26610), .b(n26604), .c(n26603), .o(n26611) );
no02f01 g22821 ( .a(n26570), .b(n26276), .o(n26612) );
no02f01 g22822 ( .a(n26449), .b(n26091), .o(n26613) );
no02f01 g22823 ( .a(n17075), .b(n17018), .o(n26614) );
no02f01 g22824 ( .a(n17077), .b(n17011), .o(n26615) );
in01f01 g22825 ( .a(n26615), .o(n26616) );
no02f01 g22826 ( .a(n26616), .b(n26614), .o(n26617) );
na02f01 g22827 ( .a(n26616), .b(n26614), .o(n26618) );
in01f01 g22828 ( .a(n26618), .o(n26619) );
no02f01 g22829 ( .a(n26619), .b(n26617), .o(n26620) );
in01f01 g22830 ( .a(n26620), .o(n26621) );
oa12f01 g22831 ( .a(n26621), .b(n26613), .c(n26612), .o(n26622) );
na02f01 g22832 ( .a(n26569), .b(n26282), .o(n26623) );
na02f01 g22833 ( .a(n26448), .b(n26103), .o(n26624) );
na02f01 g22834 ( .a(n17165), .b(n17151), .o(n26625) );
no02f01 g22835 ( .a(n17074), .b(n17018), .o(n26626) );
in01f01 g22836 ( .a(n26626), .o(n26627) );
no02f01 g22837 ( .a(n26627), .b(n26625), .o(n26628) );
na02f01 g22838 ( .a(n26627), .b(n26625), .o(n26629) );
in01f01 g22839 ( .a(n26629), .o(n26630) );
no02f01 g22840 ( .a(n26630), .b(n26628), .o(n26631) );
na03f01 g22841 ( .a(n26631), .b(n26624), .c(n26623), .o(n26632) );
no03f01 g22842 ( .a(n26567), .b(n26566), .c(n17479), .o(n26633) );
ao12f01 g22843 ( .a(n16835), .b(n26446), .c(n26445), .o(n26634) );
na02f01 g22844 ( .a(n17164), .b(n17152), .o(n26635) );
no02f01 g22845 ( .a(n17071), .b(n17027), .o(n26636) );
no02f01 g22846 ( .a(n26636), .b(n26635), .o(n26637) );
na02f01 g22847 ( .a(n26636), .b(n26635), .o(n26638) );
in01f01 g22848 ( .a(n26638), .o(n26639) );
no02f01 g22849 ( .a(n26639), .b(n26637), .o(n26640) );
in01f01 g22850 ( .a(n26640), .o(n26641) );
oa12f01 g22851 ( .a(n26641), .b(n26634), .c(n26633), .o(n26642) );
na03f01 g22852 ( .a(n17858), .b(n17851), .c(n17847), .o(n26643) );
oa12f01 g22853 ( .a(n17909), .b(n17903), .c(n17873), .o(n26644) );
no03f01 g22854 ( .a(n17909), .b(n17903), .c(n17873), .o(n26645) );
oa12f01 g22855 ( .a(n26644), .b(n17907), .c(n26645), .o(n26646) );
ao12f01 g22856 ( .a(n17859), .b(n26646), .c(n26643), .o(n26647) );
no03f01 g22857 ( .a(n26641), .b(n26634), .c(n26633), .o(n26648) );
oa12f01 g22858 ( .a(n26642), .b(n26648), .c(n26647), .o(n26649) );
ao12f01 g22859 ( .a(n26631), .b(n26624), .c(n26623), .o(n26650) );
ao12f01 g22860 ( .a(n26650), .b(n26649), .c(n26632), .o(n26651) );
no03f01 g22861 ( .a(n26621), .b(n26613), .c(n26612), .o(n26652) );
oa12f01 g22862 ( .a(n26622), .b(n26652), .c(n26651), .o(n26653) );
na03f01 g22863 ( .a(n26610), .b(n26604), .c(n26603), .o(n26654) );
ao12f01 g22864 ( .a(n26611), .b(n26654), .c(n26653), .o(n26655) );
oa12f01 g22865 ( .a(n26599), .b(n26655), .c(n26600), .o(n26656) );
oa12f01 g22866 ( .a(n26587), .b(n26656), .c(n26588), .o(n26657) );
no03f01 g22867 ( .a(n26564), .b(n26557), .c(n26556), .o(n26658) );
oa12f01 g22868 ( .a(n26565), .b(n26658), .c(n26657), .o(n26659) );
ao12f01 g22869 ( .a(n26551), .b(n26545), .c(n26543), .o(n26660) );
no02f01 g22870 ( .a(n26660), .b(n26659), .o(n26661) );
na03f01 g22871 ( .a(n26472), .b(n26469), .c(n26070), .o(n26662) );
na02f01 g22872 ( .a(n26473), .b(n26071), .o(n26663) );
na02f01 g22873 ( .a(n26663), .b(n26662), .o(n26664) );
no02f01 g22874 ( .a(n17090), .b(n16960), .o(n26665) );
no02f01 g22875 ( .a(n17092), .b(n16951), .o(n26666) );
in01f01 g22876 ( .a(n26666), .o(n26667) );
no02f01 g22877 ( .a(n26667), .b(n26665), .o(n26668) );
na02f01 g22878 ( .a(n26667), .b(n26665), .o(n26669) );
in01f01 g22879 ( .a(n26669), .o(n26670) );
no02f01 g22880 ( .a(n26670), .b(n26668), .o(n26671) );
in01f01 g22881 ( .a(n26671), .o(n26672) );
no02f01 g22882 ( .a(n26672), .b(n26664), .o(n26673) );
no03f01 g22883 ( .a(n26673), .b(n26661), .c(n26553), .o(n26674) );
oa12f01 g22884 ( .a(n17268), .b(n26536), .c(n26534), .o(n26675) );
na02f01 g22885 ( .a(n26672), .b(n26664), .o(n26676) );
na02f01 g22886 ( .a(n26676), .b(n26675), .o(n26677) );
oa12f01 g22887 ( .a(n26538), .b(n26677), .c(n26674), .o(n26678) );
no02f01 g22888 ( .a(n26524), .b(n26186), .o(n26679) );
na02f01 g22889 ( .a(n26524), .b(n26186), .o(n26680) );
in01f01 g22890 ( .a(n26680), .o(n26681) );
no02f01 g22891 ( .a(n26681), .b(n26679), .o(n26682) );
in01f01 g22892 ( .a(n26682), .o(n26683) );
no02f01 g22893 ( .a(n26683), .b(n17266), .o(n26684) );
in01f01 g22894 ( .a(n26528), .o(n26685) );
ao12f01 g22895 ( .a(n17263), .b(n26685), .c(n26526), .o(n26686) );
no02f01 g22896 ( .a(n26682), .b(n17219), .o(n26687) );
no02f01 g22897 ( .a(n26687), .b(n26686), .o(n26688) );
oa12f01 g22898 ( .a(n26688), .b(n26684), .c(n26678), .o(n26689) );
no03f01 g22899 ( .a(n26520), .b(n26519), .c(n17260), .o(n26690) );
in01f01 g22900 ( .a(n26690), .o(n26691) );
na03f01 g22901 ( .a(n26691), .b(n26689), .c(n26530), .o(n26692) );
in01f01 g22902 ( .a(n26512), .o(n26693) );
ao12f01 g22903 ( .a(n17251), .b(n26513), .c(n26693), .o(n26694) );
in01f01 g22904 ( .a(n26694), .o(n26695) );
na03f01 g22905 ( .a(n26695), .b(n26692), .c(n26521), .o(n26696) );
no02f01 g22906 ( .a(n26495), .b(n26057), .o(n26697) );
in01f01 g22907 ( .a(n26697), .o(n26698) );
na02f01 g22908 ( .a(n26495), .b(n26057), .o(n26699) );
na03f01 g22909 ( .a(n26699), .b(n26698), .c(n17236), .o(n26700) );
na03f01 g22910 ( .a(n26700), .b(n26696), .c(n26516), .o(n26701) );
in01f01 g22911 ( .a(n26699), .o(n26702) );
oa12f01 g22912 ( .a(n17570), .b(n26702), .c(n26697), .o(n26703) );
ao12f01 g22913 ( .a(n17629), .b(n26501), .c(n26499), .o(n26704) );
in01f01 g22914 ( .a(n26704), .o(n26705) );
na03f01 g22915 ( .a(n26705), .b(n26703), .c(n26701), .o(n26706) );
na03f01 g22916 ( .a(n26501), .b(n26499), .c(n17629), .o(n26707) );
na02f01 g22917 ( .a(n26504), .b(n17335), .o(n26708) );
no02f01 g22918 ( .a(n26502), .b(n17189), .o(n26709) );
no02f01 g22919 ( .a(n26502), .b(n17195), .o(n26710) );
no02f01 g22920 ( .a(n26710), .b(n26709), .o(n26711) );
na04f01 g22921 ( .a(n26711), .b(n26708), .c(n26707), .d(n26706), .o(n26712) );
ao12f01 g22922 ( .a(n17512), .b(n26502), .c(n17295), .o(n26713) );
na02f01 g22923 ( .a(n26713), .b(n26712), .o(n26714) );
ao12f01 g22924 ( .a(n26504), .b(n17440), .c(n17332), .o(n26715) );
in01f01 g22925 ( .a(n26715), .o(n26716) );
oa12f01 g22926 ( .a(n26716), .b(n26712), .c(n17325), .o(n26717) );
ao12f01 g22927 ( .a(n26717), .b(n26714), .c(n26502), .o(n26718) );
no02f01 g22928 ( .a(n17398), .b(n17499), .o(n26719) );
no02f01 g22929 ( .a(n26719), .b(n26502), .o(n26720) );
no02f01 g22930 ( .a(n26720), .b(n26718), .o(n26721) );
in01f01 g22931 ( .a(n17393), .o(n26722) );
no02f01 g22932 ( .a(n26502), .b(n26722), .o(n26723) );
no02f01 g22933 ( .a(n26502), .b(n17462), .o(n26724) );
no02f01 g22934 ( .a(n26724), .b(n26723), .o(n26725) );
na02f01 g22935 ( .a(n26725), .b(n26721), .o(n26726) );
ao12f01 g22936 ( .a(n26504), .b(n17398), .c(n17499), .o(n26727) );
ao12f01 g22937 ( .a(n26504), .b(n17393), .c(n17364), .o(n26728) );
no02f01 g22938 ( .a(n26728), .b(n26727), .o(n26729) );
na02f01 g22939 ( .a(n26729), .b(n26726), .o(n26730) );
no02f01 g22940 ( .a(n26502), .b(n17383), .o(n26731) );
no02f01 g22941 ( .a(n26502), .b(n17472), .o(n26732) );
no02f01 g22942 ( .a(n26732), .b(n26731), .o(n26733) );
ao12f01 g22943 ( .a(n26508), .b(n26733), .c(n26730), .o(n26734) );
in01f01 g22944 ( .a(n26734), .o(n26735) );
no02f01 g22945 ( .a(n26735), .b(n26507), .o(n26736) );
no02f01 g22946 ( .a(n26734), .b(n26506), .o(n26737) );
no02f01 g22947 ( .a(n26737), .b(n26736), .o(n26738) );
in01f01 g22948 ( .a(n26738), .o(n26739) );
no02f01 g22949 ( .a(n26739), .b(n26441), .o(n26740) );
no02f01 g22950 ( .a(n26738), .b(n26440), .o(n26741) );
no02f01 g22951 ( .a(n26741), .b(n26740), .o(n26742) );
in01f01 g22952 ( .a(n26439), .o(n26743) );
na02f01 g22953 ( .a(n26502), .b(n17295), .o(n26744) );
na03f01 g22954 ( .a(n26711), .b(n26707), .c(n26706), .o(n26745) );
na03f01 g22955 ( .a(n26745), .b(n26716), .c(n26744), .o(n26746) );
na02f01 g22956 ( .a(n26746), .b(n26708), .o(n26747) );
no02f01 g22957 ( .a(n26502), .b(n17512), .o(n26748) );
no02f01 g22958 ( .a(n26504), .b(n17325), .o(n26749) );
no02f01 g22959 ( .a(n26749), .b(n26748), .o(n26750) );
na02f01 g22960 ( .a(n26750), .b(n26747), .o(n26751) );
in01f01 g22961 ( .a(n26750), .o(n26752) );
na03f01 g22962 ( .a(n26752), .b(n26746), .c(n26708), .o(n26753) );
na02f01 g22963 ( .a(n26753), .b(n26751), .o(n26754) );
in01f01 g22964 ( .a(n26754), .o(n26755) );
na03f01 g22965 ( .a(n26755), .b(n26743), .c(n26436), .o(n26756) );
in01f01 g22966 ( .a(n26520), .o(n26757) );
ao12f01 g22967 ( .a(n17207), .b(n26757), .c(n26518), .o(n26758) );
in01f01 g22968 ( .a(n26557), .o(n26759) );
ao12f01 g22969 ( .a(n26563), .b(n26759), .c(n26555), .o(n26760) );
no03f01 g22970 ( .a(n26577), .b(n26464), .c(n26155), .o(n26761) );
ao12f01 g22971 ( .a(n26162), .b(n26578), .c(n26576), .o(n26762) );
in01f01 g22972 ( .a(n26586), .o(n26763) );
no03f01 g22973 ( .a(n26763), .b(n26762), .c(n26761), .o(n26764) );
oa12f01 g22974 ( .a(n26763), .b(n26762), .c(n26761), .o(n26765) );
na03f01 g22975 ( .a(n26463), .b(n26457), .c(n26125), .o(n26766) );
oa12f01 g22976 ( .a(n26126), .b(n26575), .c(n26574), .o(n26767) );
ao12f01 g22977 ( .a(n26597), .b(n26767), .c(n26766), .o(n26768) );
na03f01 g22978 ( .a(n26597), .b(n26767), .c(n26766), .o(n26769) );
no03f01 g22979 ( .a(n26601), .b(n26450), .c(n26132), .o(n26770) );
ao12f01 g22980 ( .a(n26158), .b(n26602), .c(n26571), .o(n26771) );
in01f01 g22981 ( .a(n26610), .o(n26772) );
oa12f01 g22982 ( .a(n26772), .b(n26771), .c(n26770), .o(n26773) );
na02f01 g22983 ( .a(n26449), .b(n26091), .o(n26774) );
na02f01 g22984 ( .a(n26570), .b(n26276), .o(n26775) );
ao12f01 g22985 ( .a(n26620), .b(n26775), .c(n26774), .o(n26776) );
no02f01 g22986 ( .a(n26448), .b(n26103), .o(n26777) );
no02f01 g22987 ( .a(n26569), .b(n26282), .o(n26778) );
in01f01 g22988 ( .a(n26631), .o(n26779) );
no03f01 g22989 ( .a(n26779), .b(n26778), .c(n26777), .o(n26780) );
na02f01 g22990 ( .a(n26568), .b(n16835), .o(n26781) );
na02f01 g22991 ( .a(n26447), .b(n17479), .o(n26782) );
ao12f01 g22992 ( .a(n26640), .b(n26782), .c(n26781), .o(n26783) );
oa12f01 g22993 ( .a(n17862), .b(n17861), .c(n17860), .o(n26784) );
oa12f01 g22994 ( .a(n26784), .b(n17889), .c(n17863), .o(n26785) );
na03f01 g22995 ( .a(n26640), .b(n26782), .c(n26781), .o(n26786) );
ao12f01 g22996 ( .a(n26783), .b(n26786), .c(n26785), .o(n26787) );
oa12f01 g22997 ( .a(n26779), .b(n26778), .c(n26777), .o(n26788) );
oa12f01 g22998 ( .a(n26788), .b(n26787), .c(n26780), .o(n26789) );
na03f01 g22999 ( .a(n26620), .b(n26775), .c(n26774), .o(n26790) );
ao12f01 g23000 ( .a(n26776), .b(n26790), .c(n26789), .o(n26791) );
no03f01 g23001 ( .a(n26772), .b(n26771), .c(n26770), .o(n26792) );
oa12f01 g23002 ( .a(n26773), .b(n26792), .c(n26791), .o(n26793) );
ao12f01 g23003 ( .a(n26768), .b(n26793), .c(n26769), .o(n26794) );
ao12f01 g23004 ( .a(n26764), .b(n26794), .c(n26765), .o(n26795) );
na03f01 g23005 ( .a(n26563), .b(n26759), .c(n26555), .o(n26796) );
ao12f01 g23006 ( .a(n26760), .b(n26796), .c(n26795), .o(n26797) );
in01f01 g23007 ( .a(n26543), .o(n26798) );
in01f01 g23008 ( .a(n26551), .o(n26799) );
oa12f01 g23009 ( .a(n26799), .b(n26544), .c(n26798), .o(n26800) );
na02f01 g23010 ( .a(n26800), .b(n26797), .o(n26801) );
in01f01 g23011 ( .a(n26673), .o(n26802) );
na03f01 g23012 ( .a(n26802), .b(n26801), .c(n26552), .o(n26803) );
in01f01 g23013 ( .a(n26534), .o(n26804) );
ao12f01 g23014 ( .a(n17225), .b(n26535), .c(n26804), .o(n26805) );
in01f01 g23015 ( .a(n26676), .o(n26806) );
no02f01 g23016 ( .a(n26806), .b(n26805), .o(n26807) );
ao12f01 g23017 ( .a(n26537), .b(n26807), .c(n26803), .o(n26808) );
in01f01 g23018 ( .a(n26684), .o(n26809) );
oa12f01 g23019 ( .a(n17214), .b(n26528), .c(n26527), .o(n26810) );
in01f01 g23020 ( .a(n26687), .o(n26811) );
na02f01 g23021 ( .a(n26811), .b(n26810), .o(n26812) );
ao12f01 g23022 ( .a(n26812), .b(n26809), .c(n26808), .o(n26813) );
no03f01 g23023 ( .a(n26690), .b(n26813), .c(n26529), .o(n26814) );
no03f01 g23024 ( .a(n26694), .b(n26814), .c(n26758), .o(n26815) );
no03f01 g23025 ( .a(n26702), .b(n26697), .c(n17570), .o(n26816) );
no03f01 g23026 ( .a(n26816), .b(n26815), .c(n26515), .o(n26817) );
ao12f01 g23027 ( .a(n17236), .b(n26699), .c(n26698), .o(n26818) );
no03f01 g23028 ( .a(n26704), .b(n26818), .c(n26817), .o(n26819) );
in01f01 g23029 ( .a(n26707), .o(n26820) );
na02f01 g23030 ( .a(n26502), .b(n17195), .o(n26821) );
in01f01 g23031 ( .a(n26821), .o(n26822) );
no02f01 g23032 ( .a(n26822), .b(n26710), .o(n26823) );
no03f01 g23033 ( .a(n26823), .b(n26820), .c(n26819), .o(n26824) );
in01f01 g23034 ( .a(n26710), .o(n26825) );
na02f01 g23035 ( .a(n26821), .b(n26825), .o(n26826) );
ao12f01 g23036 ( .a(n26826), .b(n26707), .c(n26706), .o(n26827) );
no02f01 g23037 ( .a(n26827), .b(n26824), .o(n26828) );
no03f01 g23038 ( .a(n26710), .b(n26820), .c(n26819), .o(n26829) );
in01f01 g23039 ( .a(n26709), .o(n26830) );
na02f01 g23040 ( .a(n26502), .b(n17189), .o(n26831) );
na02f01 g23041 ( .a(n26831), .b(n26830), .o(n26832) );
no03f01 g23042 ( .a(n26832), .b(n26829), .c(n26822), .o(n26833) );
na03f01 g23043 ( .a(n26825), .b(n26707), .c(n26706), .o(n26834) );
ao22f01 g23044 ( .a(n26831), .b(n26830), .c(n26834), .d(n26821), .o(n26835) );
no02f01 g23045 ( .a(n26835), .b(n26833), .o(n26836) );
no02f01 g23046 ( .a(n26836), .b(n26828), .o(n26837) );
in01f01 g23047 ( .a(n26837), .o(n26838) );
na03f01 g23048 ( .a(n26838), .b(n26743), .c(n26436), .o(n26839) );
na02f01 g23049 ( .a(n26745), .b(n26716), .o(n26840) );
na02f01 g23050 ( .a(n26744), .b(n26708), .o(n26841) );
na02f01 g23051 ( .a(n26841), .b(n26840), .o(n26842) );
na04f01 g23052 ( .a(n26745), .b(n26716), .c(n26744), .d(n26708), .o(n26843) );
na02f01 g23053 ( .a(n26843), .b(n26842), .o(n26844) );
in01f01 g23054 ( .a(n26844), .o(n26845) );
na03f01 g23055 ( .a(n26845), .b(n26743), .c(n26436), .o(n26846) );
na03f01 g23056 ( .a(n26846), .b(n26839), .c(n26756), .o(n26847) );
in01f01 g23057 ( .a(n26847), .o(n26848) );
oa12f01 g23058 ( .a(n26552), .b(n26660), .c(n26659), .o(n26849) );
oa12f01 g23059 ( .a(n26807), .b(n26673), .c(n26849), .o(n26850) );
ao12f01 g23060 ( .a(n26687), .b(n26850), .c(n26538), .o(n26851) );
no02f01 g23061 ( .a(n26686), .b(n26529), .o(n26852) );
oa12f01 g23062 ( .a(n26852), .b(n26851), .c(n26684), .o(n26853) );
ao12f01 g23063 ( .a(n26553), .b(n26800), .c(n26797), .o(n26854) );
ao12f01 g23064 ( .a(n26677), .b(n26802), .c(n26854), .o(n26855) );
oa12f01 g23065 ( .a(n26811), .b(n26855), .c(n26537), .o(n26856) );
in01f01 g23066 ( .a(n26852), .o(n26857) );
na03f01 g23067 ( .a(n26857), .b(n26856), .c(n26809), .o(n26858) );
na02f01 g23068 ( .a(n26858), .b(n26853), .o(n26859) );
no02f01 g23069 ( .a(n26250), .b(n7682), .o(n26860) );
no02f01 g23070 ( .a(n26860), .b(n26251), .o(n26861) );
no02f01 g23071 ( .a(n26256), .b(n7682), .o(n26862) );
oa12f01 g23072 ( .a(n26258), .b(n26862), .c(n26415), .o(n26863) );
na02f01 g23073 ( .a(n26863), .b(n26861), .o(n26864) );
in01f01 g23074 ( .a(n26861), .o(n26865) );
in01f01 g23075 ( .a(n26863), .o(n26866) );
na02f01 g23076 ( .a(n26866), .b(n26865), .o(n26867) );
na02f01 g23077 ( .a(n26867), .b(n26864), .o(n26868) );
no02f01 g23078 ( .a(n26868), .b(n26859), .o(n26869) );
in01f01 g23079 ( .a(n26869), .o(n26870) );
ao12f01 g23080 ( .a(n7712), .b(n26331), .c(n26330), .o(n26871) );
no03f01 g23081 ( .a(n26314), .b(n26310), .c(n26871), .o(n26872) );
oa22f01 g23082 ( .a(n26327), .b(n7712), .c(n26872), .d(n26295), .o(n26873) );
no02f01 g23083 ( .a(n26306), .b(n26303), .o(n26874) );
no02f01 g23084 ( .a(n26874), .b(n7682), .o(n26875) );
ao12f01 g23085 ( .a(n26875), .b(n26336), .c(n7712), .o(n26876) );
no02f01 g23086 ( .a(n26388), .b(n7712), .o(n26877) );
ao12f01 g23087 ( .a(n26877), .b(n26876), .c(n26873), .o(n26878) );
na02f01 g23088 ( .a(n26393), .b(n7682), .o(n26879) );
na02f01 g23089 ( .a(n26396), .b(n7682), .o(n26880) );
oa12f01 g23090 ( .a(n7682), .b(n26399), .c(n26398), .o(n26881) );
na04f01 g23091 ( .a(n26881), .b(n26880), .c(n26879), .d(n26878), .o(n26882) );
no02f01 g23092 ( .a(n26361), .b(n7682), .o(n26883) );
no02f01 g23093 ( .a(n26373), .b(n7682), .o(n26884) );
ao12f01 g23094 ( .a(n7682), .b(n26384), .c(n26381), .o(n26885) );
no04f01 g23095 ( .a(n26885), .b(n26884), .c(n26883), .d(n26389), .o(n26886) );
no02f01 g23096 ( .a(n26407), .b(n7712), .o(n26887) );
ao12f01 g23097 ( .a(n26887), .b(n26886), .c(n26882), .o(n26888) );
na02f01 g23098 ( .a(n26413), .b(n7712), .o(n26889) );
in01f01 g23099 ( .a(n26889), .o(n26890) );
no02f01 g23100 ( .a(n26890), .b(n26888), .o(n26891) );
no02f01 g23101 ( .a(n26272), .b(n7682), .o(n26892) );
no02f01 g23102 ( .a(n26892), .b(n26273), .o(n26893) );
no02f01 g23103 ( .a(n26893), .b(n26891), .o(n26894) );
na02f01 g23104 ( .a(n26893), .b(n26891), .o(n26895) );
in01f01 g23105 ( .a(n26895), .o(n26896) );
no02f01 g23106 ( .a(n26896), .b(n26894), .o(n26897) );
no02f01 g23107 ( .a(n26806), .b(n26674), .o(n26898) );
no02f01 g23108 ( .a(n26805), .b(n26537), .o(n26899) );
no02f01 g23109 ( .a(n26899), .b(n26898), .o(n26900) );
na02f01 g23110 ( .a(n26899), .b(n26898), .o(n26901) );
in01f01 g23111 ( .a(n26901), .o(n26902) );
no02f01 g23112 ( .a(n26902), .b(n26900), .o(n26903) );
no02f01 g23113 ( .a(n26903), .b(n26897), .o(n26904) );
na02f01 g23114 ( .a(n26886), .b(n26882), .o(n26905) );
no02f01 g23115 ( .a(n26890), .b(n26887), .o(n26906) );
in01f01 g23116 ( .a(n26906), .o(n26907) );
no02f01 g23117 ( .a(n26907), .b(n26905), .o(n26908) );
na02f01 g23118 ( .a(n26907), .b(n26905), .o(n26909) );
in01f01 g23119 ( .a(n26909), .o(n26910) );
no02f01 g23120 ( .a(n26910), .b(n26908), .o(n26911) );
no02f01 g23121 ( .a(n26806), .b(n26673), .o(n26912) );
no02f01 g23122 ( .a(n26912), .b(n26849), .o(n26913) );
na02f01 g23123 ( .a(n26912), .b(n26849), .o(n26914) );
in01f01 g23124 ( .a(n26914), .o(n26915) );
no02f01 g23125 ( .a(n26915), .b(n26913), .o(n26916) );
no02f01 g23126 ( .a(n26916), .b(n26911), .o(n26917) );
in01f01 g23127 ( .a(n26917), .o(n26918) );
na02f01 g23128 ( .a(n26879), .b(n26878), .o(n26919) );
no02f01 g23129 ( .a(n26374), .b(n26919), .o(n26920) );
na02f01 g23130 ( .a(n26394), .b(n26390), .o(n26921) );
no02f01 g23131 ( .a(n26884), .b(n26921), .o(n26922) );
in01f01 g23132 ( .a(n26922), .o(n26923) );
no02f01 g23133 ( .a(n26923), .b(n26920), .o(n26924) );
no02f01 g23134 ( .a(n26885), .b(n26385), .o(n26925) );
na02f01 g23135 ( .a(n26925), .b(n26922), .o(n26926) );
oa22f01 g23136 ( .a(n26926), .b(n26920), .c(n26925), .d(n26924), .o(n26927) );
no02f01 g23137 ( .a(n26660), .b(n26553), .o(n26928) );
no02f01 g23138 ( .a(n26928), .b(n26797), .o(n26929) );
na02f01 g23139 ( .a(n26928), .b(n26797), .o(n26930) );
in01f01 g23140 ( .a(n26930), .o(n26931) );
no02f01 g23141 ( .a(n26931), .b(n26929), .o(n26932) );
in01f01 g23142 ( .a(n26932), .o(n26933) );
no02f01 g23143 ( .a(n26933), .b(n26927), .o(n26934) );
in01f01 g23144 ( .a(n26934), .o(n26935) );
no02f01 g23145 ( .a(n26884), .b(n26374), .o(n26936) );
ao12f01 g23146 ( .a(n26921), .b(n26879), .c(n26878), .o(n26937) );
no02f01 g23147 ( .a(n26937), .b(n26936), .o(n26938) );
no02f01 g23148 ( .a(n26362), .b(n26349), .o(n26939) );
no04f01 g23149 ( .a(n26884), .b(n26921), .c(n26374), .d(n26939), .o(n26940) );
no02f01 g23150 ( .a(n26940), .b(n26938), .o(n26941) );
no03f01 g23151 ( .a(n26658), .b(n26795), .c(n26760), .o(n26942) );
ao12f01 g23152 ( .a(n26657), .b(n26796), .c(n26565), .o(n26943) );
no02f01 g23153 ( .a(n26943), .b(n26942), .o(n26944) );
no02f01 g23154 ( .a(n26944), .b(n26941), .o(n26945) );
in01f01 g23155 ( .a(n26945), .o(n26946) );
no02f01 g23156 ( .a(n26883), .b(n26362), .o(n26947) );
no02f01 g23157 ( .a(n26389), .b(n26878), .o(n26948) );
na02f01 g23158 ( .a(n26948), .b(n26947), .o(n26949) );
no02f01 g23159 ( .a(n26948), .b(n26947), .o(n26950) );
in01f01 g23160 ( .a(n26950), .o(n26951) );
no02f01 g23161 ( .a(n26588), .b(n26764), .o(n26952) );
no02f01 g23162 ( .a(n26952), .b(n26794), .o(n26953) );
na02f01 g23163 ( .a(n26952), .b(n26794), .o(n26954) );
in01f01 g23164 ( .a(n26954), .o(n26955) );
no02f01 g23165 ( .a(n26955), .b(n26953), .o(n26956) );
ao12f01 g23166 ( .a(n26956), .b(n26951), .c(n26949), .o(n26957) );
no02f01 g23167 ( .a(n26338), .b(n26329), .o(n26958) );
no02f01 g23168 ( .a(n26389), .b(n26877), .o(n26959) );
na02f01 g23169 ( .a(n26959), .b(n26958), .o(n26960) );
in01f01 g23170 ( .a(n26960), .o(n26961) );
no02f01 g23171 ( .a(n26959), .b(n26958), .o(n26962) );
no02f01 g23172 ( .a(n26600), .b(n26768), .o(n26963) );
no02f01 g23173 ( .a(n26963), .b(n26655), .o(n26964) );
na02f01 g23174 ( .a(n26963), .b(n26655), .o(n26965) );
in01f01 g23175 ( .a(n26965), .o(n26966) );
no02f01 g23176 ( .a(n26966), .b(n26964), .o(n26967) );
in01f01 g23177 ( .a(n26967), .o(n26968) );
oa12f01 g23178 ( .a(n26968), .b(n26962), .c(n26961), .o(n26969) );
na02f01 g23179 ( .a(n26336), .b(n7682), .o(n26970) );
na02f01 g23180 ( .a(n26337), .b(n26970), .o(n26971) );
na02f01 g23181 ( .a(n26333), .b(n26316), .o(n26972) );
na02f01 g23182 ( .a(n26972), .b(n26971), .o(n26973) );
no02f01 g23183 ( .a(n26327), .b(n7682), .o(n26974) );
no02f01 g23184 ( .a(n26974), .b(n26328), .o(n26975) );
na03f01 g23185 ( .a(n26975), .b(n26333), .c(n26316), .o(n26976) );
no02f01 g23186 ( .a(n26792), .b(n26611), .o(n26977) );
no02f01 g23187 ( .a(n26977), .b(n26791), .o(n26978) );
na02f01 g23188 ( .a(n26977), .b(n26791), .o(n26979) );
in01f01 g23189 ( .a(n26979), .o(n26980) );
no02f01 g23190 ( .a(n26980), .b(n26978), .o(n26981) );
na03f01 g23191 ( .a(n26981), .b(n26976), .c(n26973), .o(n26982) );
na02f01 g23192 ( .a(n26333), .b(n26307), .o(n26983) );
no03f01 g23193 ( .a(n26983), .b(n26315), .c(n26295), .o(n26984) );
no02f01 g23194 ( .a(n26875), .b(n26871), .o(n26985) );
no02f01 g23195 ( .a(n26315), .b(n26295), .o(n26986) );
no02f01 g23196 ( .a(n26986), .b(n26985), .o(n26987) );
no02f01 g23197 ( .a(n26652), .b(n26776), .o(n26988) );
no02f01 g23198 ( .a(n26988), .b(n26651), .o(n26989) );
na02f01 g23199 ( .a(n26988), .b(n26651), .o(n26990) );
in01f01 g23200 ( .a(n26990), .o(n26991) );
no02f01 g23201 ( .a(n26991), .b(n26989), .o(n26992) );
in01f01 g23202 ( .a(n26992), .o(n26993) );
oa12f01 g23203 ( .a(n26993), .b(n26987), .c(n26984), .o(n26994) );
na02f01 g23204 ( .a(n26292), .b(n26109), .o(n26995) );
oa12f01 g23205 ( .a(n26289), .b(n26108), .c(n26280), .o(n26996) );
ao12f01 g23206 ( .a(n7682), .b(n26996), .c(n26995), .o(n26997) );
no02f01 g23207 ( .a(n26312), .b(n26311), .o(n26998) );
ao12f01 g23208 ( .a(n7712), .b(n26996), .c(n26995), .o(n26999) );
no02f01 g23209 ( .a(n26999), .b(n26998), .o(n27000) );
oa12f01 g23210 ( .a(n7682), .b(n26287), .c(n26279), .o(n27001) );
na02f01 g23211 ( .a(n27001), .b(n26288), .o(n27002) );
oa12f01 g23212 ( .a(n27002), .b(n27000), .c(n26997), .o(n27003) );
ao12f01 g23213 ( .a(n7682), .b(n26309), .c(n26308), .o(n27004) );
no02f01 g23214 ( .a(n26310), .b(n27004), .o(n27005) );
na03f01 g23215 ( .a(n27005), .b(n26314), .c(n26294), .o(n27006) );
no02f01 g23216 ( .a(n26650), .b(n26780), .o(n27007) );
no02f01 g23217 ( .a(n27007), .b(n26787), .o(n27008) );
na02f01 g23218 ( .a(n27007), .b(n26787), .o(n27009) );
in01f01 g23219 ( .a(n27009), .o(n27010) );
no02f01 g23220 ( .a(n27010), .b(n27008), .o(n27011) );
ao12f01 g23221 ( .a(n27011), .b(n27006), .c(n27003), .o(n27012) );
na02f01 g23222 ( .a(n26313), .b(n26294), .o(n27013) );
no03f01 g23223 ( .a(n27013), .b(n26312), .c(n26311), .o(n27014) );
no02f01 g23224 ( .a(n26999), .b(n26997), .o(n27015) );
no02f01 g23225 ( .a(n27015), .b(n26998), .o(n27016) );
no03f01 g23226 ( .a(n26648), .b(n26785), .c(n26783), .o(n27017) );
ao12f01 g23227 ( .a(n26647), .b(n26786), .c(n26642), .o(n27018) );
no02f01 g23228 ( .a(n27018), .b(n27017), .o(n27019) );
in01f01 g23229 ( .a(n27019), .o(n27020) );
oa12f01 g23230 ( .a(n27020), .b(n27016), .c(n27014), .o(n27021) );
ao12f01 g23231 ( .a(n17941), .b(n17958), .c(n17898), .o(n27022) );
no03f01 g23232 ( .a(n27020), .b(n27016), .c(n27014), .o(n27023) );
oa12f01 g23233 ( .a(n27021), .b(n27023), .c(n27022), .o(n27024) );
na03f01 g23234 ( .a(n27011), .b(n27006), .c(n27003), .o(n27025) );
ao12f01 g23235 ( .a(n27012), .b(n27025), .c(n27024), .o(n27026) );
no03f01 g23236 ( .a(n26993), .b(n26987), .c(n26984), .o(n27027) );
oa12f01 g23237 ( .a(n26994), .b(n27027), .c(n27026), .o(n27028) );
ao12f01 g23238 ( .a(n26981), .b(n26976), .c(n26973), .o(n27029) );
oa12f01 g23239 ( .a(n26982), .b(n27029), .c(n27028), .o(n27030) );
no03f01 g23240 ( .a(n26968), .b(n26962), .c(n26961), .o(n27031) );
oa12f01 g23241 ( .a(n26969), .b(n27031), .c(n27030), .o(n27032) );
na03f01 g23242 ( .a(n26956), .b(n26951), .c(n26949), .o(n27033) );
ao12f01 g23243 ( .a(n26957), .b(n27033), .c(n27032), .o(n27034) );
na02f01 g23244 ( .a(n26944), .b(n26941), .o(n27035) );
in01f01 g23245 ( .a(n27035), .o(n27036) );
oa12f01 g23246 ( .a(n26946), .b(n27036), .c(n27034), .o(n27037) );
na02f01 g23247 ( .a(n26933), .b(n26927), .o(n27038) );
in01f01 g23248 ( .a(n27038), .o(n27039) );
oa12f01 g23249 ( .a(n26935), .b(n27039), .c(n27037), .o(n27040) );
na02f01 g23250 ( .a(n26916), .b(n26911), .o(n27041) );
in01f01 g23251 ( .a(n27041), .o(n27042) );
oa12f01 g23252 ( .a(n26918), .b(n27042), .c(n27040), .o(n27043) );
na02f01 g23253 ( .a(n26903), .b(n26897), .o(n27044) );
ao12f01 g23254 ( .a(n26904), .b(n27044), .c(n27043), .o(n27045) );
no02f01 g23255 ( .a(n26862), .b(n26257), .o(n27046) );
in01f01 g23256 ( .a(n27046), .o(n27047) );
no02f01 g23257 ( .a(n27047), .b(n26415), .o(n27048) );
na02f01 g23258 ( .a(n26411), .b(n7682), .o(n27049) );
oa12f01 g23259 ( .a(n26889), .b(n26272), .c(n7682), .o(n27050) );
ao12f01 g23260 ( .a(n27050), .b(n26888), .c(n27049), .o(n27051) );
no02f01 g23261 ( .a(n27046), .b(n27051), .o(n27052) );
no02f01 g23262 ( .a(n27052), .b(n27048), .o(n27053) );
in01f01 g23263 ( .a(n27053), .o(n27054) );
no02f01 g23264 ( .a(n26687), .b(n26684), .o(n27055) );
no02f01 g23265 ( .a(n27055), .b(n26678), .o(n27056) );
in01f01 g23266 ( .a(n27056), .o(n27057) );
na02f01 g23267 ( .a(n27055), .b(n26678), .o(n27058) );
na02f01 g23268 ( .a(n27058), .b(n27057), .o(n27059) );
no02f01 g23269 ( .a(n27059), .b(n27054), .o(n27060) );
na02f01 g23270 ( .a(n26868), .b(n26859), .o(n27061) );
in01f01 g23271 ( .a(n27058), .o(n27062) );
no02f01 g23272 ( .a(n27062), .b(n27056), .o(n27063) );
no02f01 g23273 ( .a(n27063), .b(n27053), .o(n27064) );
in01f01 g23274 ( .a(n27064), .o(n27065) );
na02f01 g23275 ( .a(n27065), .b(n27061), .o(n27066) );
in01f01 g23276 ( .a(n27066), .o(n27067) );
oa12f01 g23277 ( .a(n27067), .b(n27060), .c(n27045), .o(n27068) );
no02f01 g23278 ( .a(n26820), .b(n26704), .o(n27069) );
ao12f01 g23279 ( .a(n27069), .b(n26703), .c(n26701), .o(n27070) );
na02f01 g23280 ( .a(n26707), .b(n26705), .o(n27071) );
no03f01 g23281 ( .a(n27071), .b(n26818), .c(n26817), .o(n27072) );
no02f01 g23282 ( .a(n27072), .b(n27070), .o(n27073) );
no02f01 g23283 ( .a(n26818), .b(n26816), .o(n27074) );
no03f01 g23284 ( .a(n27074), .b(n26815), .c(n26515), .o(n27075) );
na02f01 g23285 ( .a(n26703), .b(n26700), .o(n27076) );
ao12f01 g23286 ( .a(n27076), .b(n26696), .c(n26516), .o(n27077) );
no02f01 g23287 ( .a(n27077), .b(n27075), .o(n27078) );
no02f01 g23288 ( .a(n27078), .b(n27073), .o(n27079) );
in01f01 g23289 ( .a(n27079), .o(n27080) );
na03f01 g23290 ( .a(n27080), .b(n26743), .c(n26436), .o(n27081) );
na02f01 g23291 ( .a(n26433), .b(n26429), .o(n27082) );
na02f01 g23292 ( .a(n27082), .b(n26418), .o(n27083) );
in01f01 g23293 ( .a(n26251), .o(n27084) );
no02f01 g23294 ( .a(n26860), .b(n26862), .o(n27085) );
oa12f01 g23295 ( .a(n27085), .b(n27051), .c(n26257), .o(n27086) );
na02f01 g23296 ( .a(n27086), .b(n27084), .o(n27087) );
in01f01 g23297 ( .a(n27082), .o(n27088) );
na02f01 g23298 ( .a(n27088), .b(n27087), .o(n27089) );
na02f01 g23299 ( .a(n27089), .b(n27083), .o(n27090) );
na02f01 g23300 ( .a(n26691), .b(n26521), .o(n27091) );
ao12f01 g23301 ( .a(n27091), .b(n26689), .c(n26530), .o(n27092) );
no02f01 g23302 ( .a(n26690), .b(n26758), .o(n27093) );
no03f01 g23303 ( .a(n27093), .b(n26813), .c(n26529), .o(n27094) );
no02f01 g23304 ( .a(n27094), .b(n27092), .o(n27095) );
in01f01 g23305 ( .a(n27095), .o(n27096) );
no02f01 g23306 ( .a(n27096), .b(n27090), .o(n27097) );
in01f01 g23307 ( .a(n27097), .o(n27098) );
no02f01 g23308 ( .a(n26694), .b(n26515), .o(n27099) );
ao12f01 g23309 ( .a(n27099), .b(n26692), .c(n26521), .o(n27100) );
in01f01 g23310 ( .a(n27099), .o(n27101) );
no03f01 g23311 ( .a(n27101), .b(n26814), .c(n26758), .o(n27102) );
no02f01 g23312 ( .a(n27102), .b(n27100), .o(n27103) );
na03f01 g23313 ( .a(n26429), .b(n27086), .c(n27084), .o(n27104) );
na03f01 g23314 ( .a(n27104), .b(n26433), .c(n26235), .o(n27105) );
in01f01 g23315 ( .a(n26235), .o(n27106) );
no03f01 g23316 ( .a(n26430), .b(n26417), .c(n26251), .o(n27107) );
oa12f01 g23317 ( .a(n27106), .b(n27107), .c(n26434), .o(n27108) );
na03f01 g23318 ( .a(n27108), .b(n27105), .c(n27103), .o(n27109) );
na03f01 g23319 ( .a(n27109), .b(n27098), .c(n27081), .o(n27110) );
in01f01 g23320 ( .a(n27110), .o(n27111) );
na04f01 g23321 ( .a(n27111), .b(n27068), .c(n26870), .d(n26848), .o(n27112) );
in01f01 g23322 ( .a(n27081), .o(n27113) );
ao12f01 g23323 ( .a(n27095), .b(n27089), .c(n27083), .o(n27114) );
ao12f01 g23324 ( .a(n27103), .b(n27108), .c(n27105), .o(n27115) );
oa12f01 g23325 ( .a(n27109), .b(n27115), .c(n27114), .o(n27116) );
ao22f01 g23326 ( .a(n27078), .b(n27073), .c(n26743), .d(n26436), .o(n27117) );
in01f01 g23327 ( .a(n27117), .o(n27118) );
ao12f01 g23328 ( .a(n27113), .b(n27118), .c(n27116), .o(n27119) );
ao22f01 g23329 ( .a(n26845), .b(n26755), .c(n26743), .d(n26436), .o(n27120) );
ao22f01 g23330 ( .a(n26836), .b(n26828), .c(n26743), .d(n26436), .o(n27121) );
no02f01 g23331 ( .a(n27121), .b(n27120), .o(n27122) );
in01f01 g23332 ( .a(n27122), .o(n27123) );
oa12f01 g23333 ( .a(n26848), .b(n27123), .c(n27119), .o(n27124) );
no02f01 g23334 ( .a(n26502), .b(n17349), .o(n27125) );
no02f01 g23335 ( .a(n26504), .b(n17398), .o(n27126) );
no02f01 g23336 ( .a(n27126), .b(n27125), .o(n27127) );
in01f01 g23337 ( .a(n27127), .o(n27128) );
no02f01 g23338 ( .a(n26504), .b(n17499), .o(n27129) );
in01f01 g23339 ( .a(n17499), .o(n27130) );
no02f01 g23340 ( .a(n26502), .b(n27130), .o(n27131) );
no02f01 g23341 ( .a(n27131), .b(n26718), .o(n27132) );
no03f01 g23342 ( .a(n27132), .b(n27129), .c(n27128), .o(n27133) );
oa12f01 g23343 ( .a(n27128), .b(n27132), .c(n27129), .o(n27134) );
in01f01 g23344 ( .a(n27134), .o(n27135) );
no02f01 g23345 ( .a(n27135), .b(n27133), .o(n27136) );
na02f01 g23346 ( .a(n26714), .b(n26502), .o(n27137) );
in01f01 g23347 ( .a(n26717), .o(n27138) );
na02f01 g23348 ( .a(n27138), .b(n27137), .o(n27139) );
no02f01 g23349 ( .a(n27131), .b(n27129), .o(n27140) );
in01f01 g23350 ( .a(n27140), .o(n27141) );
no02f01 g23351 ( .a(n27141), .b(n27139), .o(n27142) );
no02f01 g23352 ( .a(n27140), .b(n26718), .o(n27143) );
no02f01 g23353 ( .a(n27143), .b(n27142), .o(n27144) );
no02f01 g23354 ( .a(n27144), .b(n27136), .o(n27145) );
no02f01 g23355 ( .a(n27145), .b(n26441), .o(n27146) );
no02f01 g23356 ( .a(n26727), .b(n26721), .o(n27147) );
no02f01 g23357 ( .a(n26504), .b(n17364), .o(n27148) );
no02f01 g23358 ( .a(n27148), .b(n26724), .o(n27149) );
na02f01 g23359 ( .a(n27149), .b(n27147), .o(n27150) );
no02f01 g23360 ( .a(n27149), .b(n27147), .o(n27151) );
in01f01 g23361 ( .a(n27151), .o(n27152) );
na02f01 g23362 ( .a(n27152), .b(n27150), .o(n27153) );
no02f01 g23363 ( .a(n27153), .b(n26441), .o(n27154) );
no02f01 g23364 ( .a(n26504), .b(n17393), .o(n27155) );
no02f01 g23365 ( .a(n27155), .b(n26723), .o(n27156) );
no03f01 g23366 ( .a(n27148), .b(n26727), .c(n26721), .o(n27157) );
no03f01 g23367 ( .a(n27157), .b(n27156), .c(n26724), .o(n27158) );
oa12f01 g23368 ( .a(n27156), .b(n27157), .c(n26724), .o(n27159) );
in01f01 g23369 ( .a(n27159), .o(n27160) );
no02f01 g23370 ( .a(n27160), .b(n27158), .o(n27161) );
na02f01 g23371 ( .a(n27161), .b(n26440), .o(n27162) );
in01f01 g23372 ( .a(n27162), .o(n27163) );
no03f01 g23373 ( .a(n27163), .b(n27154), .c(n27146), .o(n27164) );
in01f01 g23374 ( .a(n27164), .o(n27165) );
ao12f01 g23375 ( .a(n27165), .b(n27124), .c(n27112), .o(n27166) );
ao12f01 g23376 ( .a(n26440), .b(n27144), .c(n27136), .o(n27167) );
in01f01 g23377 ( .a(n27150), .o(n27168) );
no02f01 g23378 ( .a(n27151), .b(n27168), .o(n27169) );
ao12f01 g23379 ( .a(n26440), .b(n27161), .c(n27169), .o(n27170) );
no02f01 g23380 ( .a(n27170), .b(n27167), .o(n27171) );
in01f01 g23381 ( .a(n27171), .o(n27172) );
in01f01 g23382 ( .a(n26731), .o(n27173) );
no02f01 g23383 ( .a(n26504), .b(n17416), .o(n27174) );
no02f01 g23384 ( .a(n27174), .b(n26732), .o(n27175) );
in01f01 g23385 ( .a(n27175), .o(n27176) );
no02f01 g23386 ( .a(n26504), .b(n17401), .o(n27177) );
in01f01 g23387 ( .a(n27177), .o(n27178) );
na03f01 g23388 ( .a(n27178), .b(n26729), .c(n26726), .o(n27179) );
ao12f01 g23389 ( .a(n27176), .b(n27179), .c(n27173), .o(n27180) );
na03f01 g23390 ( .a(n27179), .b(n27176), .c(n27173), .o(n27181) );
in01f01 g23391 ( .a(n27181), .o(n27182) );
no02f01 g23392 ( .a(n27182), .b(n27180), .o(n27183) );
no02f01 g23393 ( .a(n27177), .b(n26731), .o(n27184) );
in01f01 g23394 ( .a(n27184), .o(n27185) );
no02f01 g23395 ( .a(n27185), .b(n26730), .o(n27186) );
na02f01 g23396 ( .a(n27185), .b(n26730), .o(n27187) );
in01f01 g23397 ( .a(n27187), .o(n27188) );
no02f01 g23398 ( .a(n27188), .b(n27186), .o(n27189) );
ao12f01 g23399 ( .a(n26440), .b(n27189), .c(n27183), .o(n27190) );
no03f01 g23400 ( .a(n27190), .b(n27172), .c(n27166), .o(n27191) );
na02f01 g23401 ( .a(n27189), .b(n26440), .o(n27192) );
na02f01 g23402 ( .a(n27183), .b(n26440), .o(n27193) );
na02f01 g23403 ( .a(n27193), .b(n27192), .o(n27194) );
oa12f01 g23404 ( .a(n26742), .b(n27194), .c(n27191), .o(n27195) );
in01f01 g23405 ( .a(n26742), .o(n27196) );
in01f01 g23406 ( .a(n26904), .o(n27197) );
in01f01 g23407 ( .a(n26949), .o(n27198) );
in01f01 g23408 ( .a(n26956), .o(n27199) );
oa12f01 g23409 ( .a(n27199), .b(n26950), .c(n27198), .o(n27200) );
in01f01 g23410 ( .a(n26962), .o(n27201) );
ao12f01 g23411 ( .a(n26967), .b(n27201), .c(n26960), .o(n27202) );
ao12f01 g23412 ( .a(n26975), .b(n26333), .c(n26316), .o(n27203) );
no02f01 g23413 ( .a(n26972), .b(n26971), .o(n27204) );
in01f01 g23414 ( .a(n26981), .o(n27205) );
no03f01 g23415 ( .a(n27205), .b(n27204), .c(n27203), .o(n27206) );
na02f01 g23416 ( .a(n26986), .b(n26985), .o(n27207) );
oa12f01 g23417 ( .a(n26983), .b(n26315), .c(n26295), .o(n27208) );
ao12f01 g23418 ( .a(n26992), .b(n27208), .c(n27207), .o(n27209) );
ao12f01 g23419 ( .a(n27005), .b(n26314), .c(n26294), .o(n27210) );
no03f01 g23420 ( .a(n27002), .b(n27000), .c(n26997), .o(n27211) );
in01f01 g23421 ( .a(n27011), .o(n27212) );
oa12f01 g23422 ( .a(n27212), .b(n27211), .c(n27210), .o(n27213) );
in01f01 g23423 ( .a(n26311), .o(n27214) );
no02f01 g23424 ( .a(n17822), .b(n17795), .o(n27215) );
na03f01 g23425 ( .a(n27015), .b(n27215), .c(n27214), .o(n27216) );
oa12f01 g23426 ( .a(n27013), .b(n26312), .c(n26311), .o(n27217) );
ao12f01 g23427 ( .a(n27019), .b(n27217), .c(n27216), .o(n27218) );
oa12f01 g23428 ( .a(n17895), .b(n17939), .c(n17942), .o(n27219) );
na03f01 g23429 ( .a(n27019), .b(n27217), .c(n27216), .o(n27220) );
ao12f01 g23430 ( .a(n27218), .b(n27220), .c(n27219), .o(n27221) );
no03f01 g23431 ( .a(n27212), .b(n27211), .c(n27210), .o(n27222) );
oa12f01 g23432 ( .a(n27213), .b(n27222), .c(n27221), .o(n27223) );
na03f01 g23433 ( .a(n26992), .b(n27208), .c(n27207), .o(n27224) );
ao12f01 g23434 ( .a(n27209), .b(n27224), .c(n27223), .o(n27225) );
oa12f01 g23435 ( .a(n27205), .b(n27204), .c(n27203), .o(n27226) );
ao12f01 g23436 ( .a(n27206), .b(n27226), .c(n27225), .o(n27227) );
na03f01 g23437 ( .a(n26967), .b(n27201), .c(n26960), .o(n27228) );
ao12f01 g23438 ( .a(n27202), .b(n27228), .c(n27227), .o(n27229) );
no03f01 g23439 ( .a(n27199), .b(n26950), .c(n27198), .o(n27230) );
oa12f01 g23440 ( .a(n27200), .b(n27230), .c(n27229), .o(n27231) );
ao12f01 g23441 ( .a(n26945), .b(n27035), .c(n27231), .o(n27232) );
ao12f01 g23442 ( .a(n26934), .b(n27038), .c(n27232), .o(n27233) );
ao12f01 g23443 ( .a(n26917), .b(n27041), .c(n27233), .o(n27234) );
in01f01 g23444 ( .a(n27044), .o(n27235) );
oa12f01 g23445 ( .a(n27197), .b(n27235), .c(n27234), .o(n27236) );
in01f01 g23446 ( .a(n27060), .o(n27237) );
ao12f01 g23447 ( .a(n27066), .b(n27237), .c(n27236), .o(n27238) );
no04f01 g23448 ( .a(n27110), .b(n27238), .c(n26869), .d(n26847), .o(n27239) );
in01f01 g23449 ( .a(n27103), .o(n27240) );
no03f01 g23450 ( .a(n27107), .b(n26434), .c(n27106), .o(n27241) );
ao12f01 g23451 ( .a(n26235), .b(n27104), .c(n26433), .o(n27242) );
no03f01 g23452 ( .a(n27242), .b(n27241), .c(n27240), .o(n27243) );
na02f01 g23453 ( .a(n27096), .b(n27090), .o(n27244) );
oa12f01 g23454 ( .a(n27240), .b(n27242), .c(n27241), .o(n27245) );
ao12f01 g23455 ( .a(n27243), .b(n27245), .c(n27244), .o(n27246) );
oa12f01 g23456 ( .a(n27081), .b(n27117), .c(n27246), .o(n27247) );
ao12f01 g23457 ( .a(n26847), .b(n27122), .c(n27247), .o(n27248) );
oa12f01 g23458 ( .a(n27164), .b(n27248), .c(n27239), .o(n27249) );
in01f01 g23459 ( .a(n27190), .o(n27250) );
na03f01 g23460 ( .a(n27250), .b(n27171), .c(n27249), .o(n27251) );
in01f01 g23461 ( .a(n27194), .o(n27252) );
na03f01 g23462 ( .a(n27252), .b(n27251), .c(n27196), .o(n27253) );
na03f01 g23463 ( .a(n27253), .b(n27195), .c(n1821), .o(n27254) );
ao12f01 g23464 ( .a(n27196), .b(n27252), .c(n27251), .o(n27255) );
no03f01 g23465 ( .a(n27194), .b(n27191), .c(n26742), .o(n27256) );
oa12f01 g23466 ( .a(n8066), .b(n27256), .c(n27255), .o(n27257) );
na02f01 g23467 ( .a(n27257), .b(n27254), .o(n343) );
no02f01 g23468 ( .a(n16194), .b(n15090), .o(n27259) );
no02f01 g23469 ( .a(n16193), .b(n15087), .o(n27260) );
no02f01 g23470 ( .a(n27260), .b(n27259), .o(n27261) );
in01f01 g23471 ( .a(n27261), .o(n27262) );
no02f01 g23472 ( .a(n21600), .b(n21567), .o(n27263) );
in01f01 g23473 ( .a(n15155), .o(n27264) );
no02f01 g23474 ( .a(n16194), .b(n27264), .o(n27265) );
in01f01 g23475 ( .a(n27265), .o(n27266) );
na03f01 g23476 ( .a(n27266), .b(n27263), .c(n21560), .o(n27267) );
no02f01 g23477 ( .a(n15140), .b(n15123), .o(n27268) );
ao12f01 g23478 ( .a(n16193), .b(n27268), .c(n15155), .o(n27269) );
no02f01 g23479 ( .a(n27269), .b(n21564), .o(n27270) );
oa12f01 g23480 ( .a(n27270), .b(n27267), .c(n21483), .o(n27271) );
no02f01 g23481 ( .a(n27271), .b(n27262), .o(n27272) );
na02f01 g23482 ( .a(n27271), .b(n27262), .o(n27273) );
in01f01 g23483 ( .a(n27273), .o(n27274) );
no02f01 g23484 ( .a(n27274), .b(n27272), .o(n27275) );
no02f01 g23485 ( .a(n27275), .b(n15949), .o(n27276) );
no02f01 g23486 ( .a(n27275), .b(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .o(n27277) );
no02f01 g23487 ( .a(n27277), .b(n27276), .o(n27278) );
in01f01 g23488 ( .a(n27278), .o(n27279) );
oa12f01 g23489 ( .a(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .b(n21575), .c(n21548), .o(n27280) );
oa12f01 g23490 ( .a(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .b(n21605), .c(n21604), .o(n27281) );
na02f01 g23491 ( .a(n27281), .b(n27280), .o(n27282) );
no02f01 g23492 ( .a(n27268), .b(n16193), .o(n27283) );
in01f01 g23493 ( .a(n27283), .o(n27284) );
no02f01 g23494 ( .a(n16193), .b(n15155), .o(n27285) );
no02f01 g23495 ( .a(n27285), .b(n27265), .o(n27286) );
na02f01 g23496 ( .a(n27263), .b(n21566), .o(n27287) );
na03f01 g23497 ( .a(n27287), .b(n27286), .c(n27284), .o(n27288) );
in01f01 g23498 ( .a(n27288), .o(n27289) );
ao12f01 g23499 ( .a(n27286), .b(n27287), .c(n27284), .o(n27290) );
no02f01 g23500 ( .a(n27290), .b(n27289), .o(n27291) );
no02f01 g23501 ( .a(n27291), .b(n15949), .o(n27292) );
no02f01 g23502 ( .a(n27292), .b(n27282), .o(n27293) );
no02f01 g23503 ( .a(n27293), .b(n27279), .o(n27294) );
ao12f01 g23504 ( .a(n15949), .b(n21595), .c(n21589), .o(n27295) );
in01f01 g23505 ( .a(n21605), .o(n27296) );
ao12f01 g23506 ( .a(n15949), .b(n27296), .c(n21603), .o(n27297) );
no02f01 g23507 ( .a(n27297), .b(n27295), .o(n27298) );
in01f01 g23508 ( .a(n27290), .o(n27299) );
na02f01 g23509 ( .a(n27299), .b(n27288), .o(n27300) );
na02f01 g23510 ( .a(n27300), .b(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .o(n27301) );
na02f01 g23511 ( .a(n27301), .b(n27298), .o(n27302) );
no02f01 g23512 ( .a(n27302), .b(n27278), .o(n27303) );
no02f01 g23513 ( .a(n27303), .b(n27294), .o(n27304) );
no02f01 g23514 ( .a(n15892), .b(n15535), .o(n27305) );
no02f01 g23515 ( .a(n27305), .b(n15888), .o(n27306) );
na02f01 g23516 ( .a(n27305), .b(n15888), .o(n27307) );
in01f01 g23517 ( .a(n27307), .o(n27308) );
no02f01 g23518 ( .a(n27308), .b(n27306), .o(n27309) );
no02f01 g23519 ( .a(n27309), .b(n27304), .o(n27310) );
in01f01 g23520 ( .a(n27310), .o(n27311) );
no02f01 g23521 ( .a(n27291), .b(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .o(n27312) );
no02f01 g23522 ( .a(n27312), .b(n27292), .o(n27313) );
no02f01 g23523 ( .a(n27313), .b(n27282), .o(n27314) );
na02f01 g23524 ( .a(n27300), .b(n15949), .o(n27315) );
na02f01 g23525 ( .a(n27315), .b(n27301), .o(n27316) );
no02f01 g23526 ( .a(n27316), .b(n27298), .o(n27317) );
no02f01 g23527 ( .a(n15583), .b(n15870), .o(n27318) );
no02f01 g23528 ( .a(n27318), .b(n15582), .o(n27319) );
na02f01 g23529 ( .a(n27318), .b(n15582), .o(n27320) );
in01f01 g23530 ( .a(n27320), .o(n27321) );
no02f01 g23531 ( .a(n27321), .b(n27319), .o(n27322) );
in01f01 g23532 ( .a(n27322), .o(n27323) );
oa12f01 g23533 ( .a(n27323), .b(n27317), .c(n27314), .o(n27324) );
oa12f01 g23534 ( .a(n15949), .b(n21605), .c(n21604), .o(n27325) );
na03f01 g23535 ( .a(n27325), .b(n27281), .c(n27295), .o(n27326) );
ao12f01 g23536 ( .a(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .b(n27296), .c(n21603), .o(n27327) );
oa12f01 g23537 ( .a(n27280), .b(n27327), .c(n27297), .o(n27328) );
no02f01 g23538 ( .a(n15885), .b(n15560), .o(n27329) );
no02f01 g23539 ( .a(n27329), .b(n15884), .o(n27330) );
na02f01 g23540 ( .a(n27329), .b(n15884), .o(n27331) );
in01f01 g23541 ( .a(n27331), .o(n27332) );
no02f01 g23542 ( .a(n27332), .b(n27330), .o(n27333) );
ao12f01 g23543 ( .a(n27333), .b(n27328), .c(n27326), .o(n27334) );
ao12f01 g23544 ( .a(n21595), .b(n21548), .c(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .o(n27335) );
no03f01 g23545 ( .a(n21575), .b(n21589), .c(n15949), .o(n27336) );
no02f01 g23546 ( .a(n15883), .b(n15567), .o(n27337) );
no02f01 g23547 ( .a(n15579), .b(n15566), .o(n27338) );
no02f01 g23548 ( .a(n27338), .b(n27337), .o(n27339) );
no02f01 g23549 ( .a(n27339), .b(n15878), .o(n27340) );
na02f01 g23550 ( .a(n27339), .b(n15878), .o(n27341) );
in01f01 g23551 ( .a(n27341), .o(n27342) );
no02f01 g23552 ( .a(n27342), .b(n27340), .o(n27343) );
in01f01 g23553 ( .a(n27343), .o(n27344) );
no03f01 g23554 ( .a(n27344), .b(n27336), .c(n27335), .o(n27345) );
na02f01 g23555 ( .a(n21589), .b(n15949), .o(n27346) );
na02f01 g23556 ( .a(n21589), .b(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .o(n27347) );
no02f01 g23557 ( .a(n15569), .b(n15568), .o(n27348) );
no02f01 g23558 ( .a(n15573), .b(n27348), .o(n27349) );
na02f01 g23559 ( .a(n15573), .b(n27348), .o(n27350) );
in01f01 g23560 ( .a(n27350), .o(n27351) );
no02f01 g23561 ( .a(n27351), .b(n27349), .o(n27352) );
in01f01 g23562 ( .a(n27352), .o(n27353) );
na03f01 g23563 ( .a(n27353), .b(n27347), .c(n27346), .o(n27354) );
oa12f01 g23564 ( .a(n27344), .b(n27336), .c(n27335), .o(n27355) );
oa12f01 g23565 ( .a(n27355), .b(n27354), .c(n27345), .o(n27356) );
na03f01 g23566 ( .a(n27333), .b(n27328), .c(n27326), .o(n27357) );
ao12f01 g23567 ( .a(n27334), .b(n27357), .c(n27356), .o(n27358) );
no03f01 g23568 ( .a(n27323), .b(n27317), .c(n27314), .o(n27359) );
oa12f01 g23569 ( .a(n27324), .b(n27359), .c(n27358), .o(n27360) );
in01f01 g23570 ( .a(n27309), .o(n27361) );
no03f01 g23571 ( .a(n27361), .b(n27303), .c(n27294), .o(n27362) );
in01f01 g23572 ( .a(n27362), .o(n27363) );
na02f01 g23573 ( .a(n27363), .b(n27360), .o(n27364) );
no03f01 g23574 ( .a(n27293), .b(n27277), .c(n27276), .o(n27365) );
no03f01 g23575 ( .a(n27282), .b(n27275), .c(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .o(n27366) );
no02f01 g23576 ( .a(n27366), .b(n27365), .o(n27367) );
no02f01 g23577 ( .a(n15590), .b(n15525), .o(n27368) );
no02f01 g23578 ( .a(n27368), .b(n15586), .o(n27369) );
na02f01 g23579 ( .a(n27368), .b(n15586), .o(n27370) );
in01f01 g23580 ( .a(n27370), .o(n27371) );
no02f01 g23581 ( .a(n27371), .b(n27369), .o(n27372) );
no02f01 g23582 ( .a(n27372), .b(n27367), .o(n27373) );
in01f01 g23583 ( .a(n27373), .o(n27374) );
na03f01 g23584 ( .a(n27374), .b(n27364), .c(n27311), .o(n27375) );
na02f01 g23585 ( .a(n27372), .b(n27367), .o(n27376) );
no02f01 g23586 ( .a(n15607), .b(n15594), .o(n27377) );
no02f01 g23587 ( .a(n15591), .b(n15525), .o(n27378) );
no02f01 g23588 ( .a(n15611), .b(n15173), .o(n27379) );
no02f01 g23589 ( .a(n27379), .b(n27378), .o(n27380) );
no02f01 g23590 ( .a(n27380), .b(n27377), .o(n27381) );
no02f01 g23591 ( .a(n15610), .b(n15173), .o(n27382) );
no02f01 g23592 ( .a(n15600), .b(n15594), .o(n27383) );
no02f01 g23593 ( .a(n27383), .b(n27382), .o(n27384) );
no02f01 g23594 ( .a(n27384), .b(n27381), .o(n27385) );
na02f01 g23595 ( .a(n27384), .b(n27381), .o(n27386) );
in01f01 g23596 ( .a(n27386), .o(n27387) );
no02f01 g23597 ( .a(n27387), .b(n27385), .o(n27388) );
no04f01 g23598 ( .a(n27379), .b(n27377), .c(n15591), .d(n15525), .o(n27389) );
no02f01 g23599 ( .a(n27379), .b(n27377), .o(n27390) );
no02f01 g23600 ( .a(n27390), .b(n27378), .o(n27391) );
no02f01 g23601 ( .a(n27391), .b(n27389), .o(n27392) );
ao12f01 g23602 ( .a(n27367), .b(n27392), .c(n27388), .o(n27393) );
ao12f01 g23603 ( .a(n27393), .b(n27376), .c(n27375), .o(n27394) );
in01f01 g23604 ( .a(n27367), .o(n27395) );
in01f01 g23605 ( .a(n27392), .o(n27396) );
no02f01 g23606 ( .a(n27396), .b(n27395), .o(n27397) );
in01f01 g23607 ( .a(n27388), .o(n27398) );
no02f01 g23608 ( .a(n27398), .b(n27395), .o(n27399) );
no02f01 g23609 ( .a(n27399), .b(n27397), .o(n27400) );
in01f01 g23610 ( .a(n27400), .o(n27401) );
no02f01 g23611 ( .a(n15612), .b(n15609), .o(n27402) );
in01f01 g23612 ( .a(n27402), .o(n27403) );
no02f01 g23613 ( .a(n15903), .b(n27403), .o(n27404) );
no02f01 g23614 ( .a(n15621), .b(n15594), .o(n27405) );
no02f01 g23615 ( .a(n27405), .b(n15900), .o(n27406) );
in01f01 g23616 ( .a(n27406), .o(n27407) );
no03f01 g23617 ( .a(n27407), .b(n27404), .c(n15694), .o(n27408) );
no02f01 g23618 ( .a(n27404), .b(n15694), .o(n27409) );
no02f01 g23619 ( .a(n27406), .b(n27409), .o(n27410) );
no02f01 g23620 ( .a(n27410), .b(n27408), .o(n27411) );
na02f01 g23621 ( .a(n27411), .b(n27367), .o(n27412) );
na02f01 g23622 ( .a(n27404), .b(n15622), .o(n27413) );
no02f01 g23623 ( .a(n15694), .b(n27405), .o(n27414) );
na02f01 g23624 ( .a(n27414), .b(n27413), .o(n27415) );
in01f01 g23625 ( .a(n27415), .o(n27416) );
no02f01 g23626 ( .a(n15649), .b(n15594), .o(n27417) );
no02f01 g23627 ( .a(n27417), .b(n15905), .o(n27418) );
no02f01 g23628 ( .a(n27418), .b(n27416), .o(n27419) );
na02f01 g23629 ( .a(n27418), .b(n27416), .o(n27420) );
in01f01 g23630 ( .a(n27420), .o(n27421) );
no02f01 g23631 ( .a(n27421), .b(n27419), .o(n27422) );
na02f01 g23632 ( .a(n27422), .b(n27367), .o(n27423) );
no02f01 g23633 ( .a(n15638), .b(n15594), .o(n27424) );
no02f01 g23634 ( .a(n15902), .b(n15173), .o(n27425) );
no02f01 g23635 ( .a(n27425), .b(n27424), .o(n27426) );
in01f01 g23636 ( .a(n27426), .o(n27427) );
no02f01 g23637 ( .a(n27427), .b(n27402), .o(n27428) );
no02f01 g23638 ( .a(n27426), .b(n27403), .o(n27429) );
no02f01 g23639 ( .a(n27429), .b(n27428), .o(n27430) );
in01f01 g23640 ( .a(n27425), .o(n27431) );
ao12f01 g23641 ( .a(n27424), .b(n27431), .c(n27402), .o(n27432) );
no02f01 g23642 ( .a(n15633), .b(n15594), .o(n27433) );
no02f01 g23643 ( .a(n15901), .b(n15173), .o(n27434) );
no02f01 g23644 ( .a(n27434), .b(n27433), .o(n27435) );
no02f01 g23645 ( .a(n27435), .b(n27432), .o(n27436) );
na02f01 g23646 ( .a(n27435), .b(n27432), .o(n27437) );
in01f01 g23647 ( .a(n27437), .o(n27438) );
no02f01 g23648 ( .a(n27438), .b(n27436), .o(n27439) );
oa12f01 g23649 ( .a(n27367), .b(n27439), .c(n27430), .o(n27440) );
na03f01 g23650 ( .a(n27440), .b(n27423), .c(n27412), .o(n27441) );
no02f01 g23651 ( .a(n15651), .b(n27403), .o(n27442) );
in01f01 g23652 ( .a(n15695), .o(n27443) );
no02f01 g23653 ( .a(n27443), .b(n27442), .o(n27444) );
no02f01 g23654 ( .a(n15681), .b(n15594), .o(n27445) );
no02f01 g23655 ( .a(n15910), .b(n15173), .o(n27446) );
no02f01 g23656 ( .a(n27446), .b(n27445), .o(n27447) );
no02f01 g23657 ( .a(n27447), .b(n27444), .o(n27448) );
na02f01 g23658 ( .a(n27447), .b(n27444), .o(n27449) );
in01f01 g23659 ( .a(n27449), .o(n27450) );
no02f01 g23660 ( .a(n27450), .b(n27448), .o(n27451) );
na02f01 g23661 ( .a(n27451), .b(n27367), .o(n27452) );
in01f01 g23662 ( .a(n27452), .o(n27453) );
no02f01 g23663 ( .a(n27446), .b(n27444), .o(n27454) );
no02f01 g23664 ( .a(n27454), .b(n27445), .o(n27455) );
no02f01 g23665 ( .a(n15676), .b(n15594), .o(n27456) );
no02f01 g23666 ( .a(n15909), .b(n15173), .o(n27457) );
no02f01 g23667 ( .a(n27457), .b(n27456), .o(n27458) );
no02f01 g23668 ( .a(n27458), .b(n27455), .o(n27459) );
na02f01 g23669 ( .a(n27458), .b(n27455), .o(n27460) );
in01f01 g23670 ( .a(n27460), .o(n27461) );
no02f01 g23671 ( .a(n27461), .b(n27459), .o(n27462) );
na02f01 g23672 ( .a(n27462), .b(n27367), .o(n27463) );
in01f01 g23673 ( .a(n27463), .o(n27464) );
no02f01 g23674 ( .a(n27464), .b(n27453), .o(n27465) );
na02f01 g23675 ( .a(n15912), .b(n15173), .o(n27466) );
no02f01 g23676 ( .a(n15696), .b(n27443), .o(n27467) );
na02f01 g23677 ( .a(n15682), .b(n27442), .o(n27468) );
na02f01 g23678 ( .a(n27468), .b(n27467), .o(n27469) );
in01f01 g23679 ( .a(n27469), .o(n27470) );
ao12f01 g23680 ( .a(n15913), .b(n27470), .c(n27466), .o(n27471) );
in01f01 g23681 ( .a(n27471), .o(n27472) );
no02f01 g23682 ( .a(n15665), .b(n15594), .o(n27473) );
no02f01 g23683 ( .a(n27473), .b(n15908), .o(n27474) );
no02f01 g23684 ( .a(n27474), .b(n27472), .o(n27475) );
na02f01 g23685 ( .a(n27474), .b(n27472), .o(n27476) );
in01f01 g23686 ( .a(n27476), .o(n27477) );
no02f01 g23687 ( .a(n27477), .b(n27475), .o(n27478) );
na02f01 g23688 ( .a(n27478), .b(n27367), .o(n27479) );
na02f01 g23689 ( .a(n27466), .b(n15690), .o(n27480) );
in01f01 g23690 ( .a(n27480), .o(n27481) );
no02f01 g23691 ( .a(n27481), .b(n27470), .o(n27482) );
no02f01 g23692 ( .a(n27480), .b(n27469), .o(n27483) );
no02f01 g23693 ( .a(n27483), .b(n27482), .o(n27484) );
na02f01 g23694 ( .a(n27484), .b(n27367), .o(n27485) );
na03f01 g23695 ( .a(n27485), .b(n27479), .c(n27465), .o(n27486) );
no04f01 g23696 ( .a(n27486), .b(n27441), .c(n27401), .d(n27394), .o(n27487) );
ao12f01 g23697 ( .a(n27367), .b(n27439), .c(n27430), .o(n27488) );
ao12f01 g23698 ( .a(n27367), .b(n27422), .c(n27411), .o(n27489) );
no02f01 g23699 ( .a(n27489), .b(n27488), .o(n27490) );
ao12f01 g23700 ( .a(n27367), .b(n27462), .c(n27451), .o(n27491) );
ao12f01 g23701 ( .a(n27367), .b(n27484), .c(n27478), .o(n27492) );
no02f01 g23702 ( .a(n27492), .b(n27491), .o(n27493) );
na02f01 g23703 ( .a(n27493), .b(n27490), .o(n27494) );
no02f01 g23704 ( .a(n27494), .b(n27487), .o(n27495) );
in01f01 g23705 ( .a(n15742), .o(n27496) );
ao12f01 g23706 ( .a(n15837), .b(n27496), .c(n15917), .o(n27497) );
no02f01 g23707 ( .a(n15711), .b(n15594), .o(n27498) );
no02f01 g23708 ( .a(n27498), .b(n15713), .o(n27499) );
no02f01 g23709 ( .a(n27499), .b(n27497), .o(n27500) );
na02f01 g23710 ( .a(n27499), .b(n27497), .o(n27501) );
in01f01 g23711 ( .a(n27501), .o(n27502) );
no02f01 g23712 ( .a(n27502), .b(n27500), .o(n27503) );
in01f01 g23713 ( .a(n27503), .o(n27504) );
no02f01 g23714 ( .a(n27504), .b(n27395), .o(n27505) );
in01f01 g23715 ( .a(n27505), .o(n27506) );
no02f01 g23716 ( .a(n15740), .b(n15594), .o(n27507) );
no02f01 g23717 ( .a(n15741), .b(n15173), .o(n27508) );
in01f01 g23718 ( .a(n27508), .o(n27509) );
ao12f01 g23719 ( .a(n27507), .b(n27509), .c(n15917), .o(n27510) );
no02f01 g23720 ( .a(n15734), .b(n15594), .o(n27511) );
no02f01 g23721 ( .a(n15735), .b(n15173), .o(n27512) );
no02f01 g23722 ( .a(n27512), .b(n27511), .o(n27513) );
no02f01 g23723 ( .a(n27513), .b(n27510), .o(n27514) );
na02f01 g23724 ( .a(n27513), .b(n27510), .o(n27515) );
in01f01 g23725 ( .a(n27515), .o(n27516) );
no02f01 g23726 ( .a(n27516), .b(n27514), .o(n27517) );
no02f01 g23727 ( .a(n27508), .b(n27507), .o(n27518) );
no02f01 g23728 ( .a(n27518), .b(n15701), .o(n27519) );
na02f01 g23729 ( .a(n27518), .b(n15701), .o(n27520) );
in01f01 g23730 ( .a(n27520), .o(n27521) );
no02f01 g23731 ( .a(n27521), .b(n27519), .o(n27522) );
no02f01 g23732 ( .a(n27522), .b(n27517), .o(n27523) );
no02f01 g23733 ( .a(n27523), .b(n27395), .o(n27524) );
in01f01 g23734 ( .a(n27524), .o(n27525) );
no03f01 g23735 ( .a(n15742), .b(n15713), .c(n15701), .o(n27526) );
no02f01 g23736 ( .a(n15837), .b(n27498), .o(n27527) );
in01f01 g23737 ( .a(n27527), .o(n27528) );
no02f01 g23738 ( .a(n15721), .b(n15594), .o(n27529) );
no02f01 g23739 ( .a(n27529), .b(n15723), .o(n27530) );
in01f01 g23740 ( .a(n27530), .o(n27531) );
no03f01 g23741 ( .a(n27531), .b(n27528), .c(n27526), .o(n27532) );
no02f01 g23742 ( .a(n27528), .b(n27526), .o(n27533) );
no02f01 g23743 ( .a(n27530), .b(n27533), .o(n27534) );
no02f01 g23744 ( .a(n27534), .b(n27532), .o(n27535) );
in01f01 g23745 ( .a(n27535), .o(n27536) );
no02f01 g23746 ( .a(n27536), .b(n27395), .o(n27537) );
in01f01 g23747 ( .a(n27537), .o(n27538) );
na03f01 g23748 ( .a(n27538), .b(n27525), .c(n27506), .o(n27539) );
in01f01 g23749 ( .a(n15838), .o(n27540) );
no02f01 g23750 ( .a(n15774), .b(n15594), .o(n27541) );
no02f01 g23751 ( .a(n15775), .b(n15173), .o(n27542) );
no02f01 g23752 ( .a(n27542), .b(n27541), .o(n27543) );
in01f01 g23753 ( .a(n27543), .o(n27544) );
no03f01 g23754 ( .a(n27544), .b(n27540), .c(n16107), .o(n27545) );
no02f01 g23755 ( .a(n27540), .b(n16107), .o(n27546) );
no02f01 g23756 ( .a(n27543), .b(n27546), .o(n27547) );
no02f01 g23757 ( .a(n27547), .b(n27545), .o(n27548) );
in01f01 g23758 ( .a(n27548), .o(n27549) );
no02f01 g23759 ( .a(n27549), .b(n27395), .o(n27550) );
no02f01 g23760 ( .a(n27550), .b(n27539), .o(n27551) );
in01f01 g23761 ( .a(n27551), .o(n27552) );
no02f01 g23762 ( .a(n27542), .b(n27546), .o(n27553) );
no02f01 g23763 ( .a(n27553), .b(n27541), .o(n27554) );
no02f01 g23764 ( .a(n15768), .b(n15594), .o(n27555) );
no02f01 g23765 ( .a(n15769), .b(n15173), .o(n27556) );
no02f01 g23766 ( .a(n27556), .b(n27555), .o(n27557) );
no02f01 g23767 ( .a(n27557), .b(n27554), .o(n27558) );
na02f01 g23768 ( .a(n27557), .b(n27554), .o(n27559) );
in01f01 g23769 ( .a(n27559), .o(n27560) );
no02f01 g23770 ( .a(n27560), .b(n27558), .o(n27561) );
in01f01 g23771 ( .a(n27561), .o(n27562) );
no02f01 g23772 ( .a(n27562), .b(n27395), .o(n27563) );
in01f01 g23773 ( .a(n15776), .o(n27564) );
ao12f01 g23774 ( .a(n27540), .b(n27564), .c(n16107), .o(n27565) );
in01f01 g23775 ( .a(n27565), .o(n27566) );
no02f01 g23776 ( .a(n15756), .b(n15594), .o(n27567) );
no02f01 g23777 ( .a(n27567), .b(n15758), .o(n27568) );
in01f01 g23778 ( .a(n27568), .o(n27569) );
no03f01 g23779 ( .a(n27569), .b(n27566), .c(n15840), .o(n27570) );
ao12f01 g23780 ( .a(n27568), .b(n27565), .c(n15841), .o(n27571) );
no02f01 g23781 ( .a(n27571), .b(n27570), .o(n27572) );
in01f01 g23782 ( .a(n27572), .o(n27573) );
no02f01 g23783 ( .a(n27573), .b(n27395), .o(n27574) );
no02f01 g23784 ( .a(n27567), .b(n15840), .o(n27575) );
oa12f01 g23785 ( .a(n27575), .b(n27565), .c(n15758), .o(n27576) );
in01f01 g23786 ( .a(n27576), .o(n27577) );
no02f01 g23787 ( .a(n15786), .b(n15594), .o(n27578) );
no02f01 g23788 ( .a(n27578), .b(n15788), .o(n27579) );
no02f01 g23789 ( .a(n27579), .b(n27577), .o(n27580) );
na02f01 g23790 ( .a(n27579), .b(n27577), .o(n27581) );
in01f01 g23791 ( .a(n27581), .o(n27582) );
no02f01 g23792 ( .a(n27582), .b(n27580), .o(n27583) );
in01f01 g23793 ( .a(n27583), .o(n27584) );
no02f01 g23794 ( .a(n27584), .b(n27395), .o(n27585) );
no02f01 g23795 ( .a(n27585), .b(n27574), .o(n27586) );
in01f01 g23796 ( .a(n27586), .o(n27587) );
no04f01 g23797 ( .a(n27587), .b(n27563), .c(n27552), .d(n27495), .o(n27588) );
na02f01 g23798 ( .a(n15743), .b(n15917), .o(n27589) );
in01f01 g23799 ( .a(n15843), .o(n27590) );
oa12f01 g23800 ( .a(n27590), .b(n15926), .c(n27589), .o(n27591) );
no02f01 g23801 ( .a(n15817), .b(n15594), .o(n27592) );
no02f01 g23802 ( .a(n15818), .b(n15173), .o(n27593) );
no02f01 g23803 ( .a(n27593), .b(n27592), .o(n27594) );
in01f01 g23804 ( .a(n27594), .o(n27595) );
no02f01 g23805 ( .a(n27595), .b(n27591), .o(n27596) );
no02f01 g23806 ( .a(n27594), .b(n16108), .o(n27597) );
no02f01 g23807 ( .a(n27597), .b(n27596), .o(n27598) );
in01f01 g23808 ( .a(n27598), .o(n27599) );
no02f01 g23809 ( .a(n27599), .b(n27395), .o(n27600) );
in01f01 g23810 ( .a(n27593), .o(n27601) );
ao12f01 g23811 ( .a(n27592), .b(n27601), .c(n27591), .o(n27602) );
no02f01 g23812 ( .a(n15811), .b(n15594), .o(n27603) );
no02f01 g23813 ( .a(n15812), .b(n15173), .o(n27604) );
no02f01 g23814 ( .a(n27604), .b(n27603), .o(n27605) );
no02f01 g23815 ( .a(n27605), .b(n27602), .o(n27606) );
na02f01 g23816 ( .a(n27605), .b(n27602), .o(n27607) );
in01f01 g23817 ( .a(n27607), .o(n27608) );
no02f01 g23818 ( .a(n27608), .b(n27606), .o(n27609) );
in01f01 g23819 ( .a(n27609), .o(n27610) );
no02f01 g23820 ( .a(n27610), .b(n27395), .o(n27611) );
no02f01 g23821 ( .a(n27611), .b(n27600), .o(n27612) );
in01f01 g23822 ( .a(n15931), .o(n27613) );
ao12f01 g23823 ( .a(n27613), .b(n15927), .c(n16107), .o(n27614) );
no02f01 g23824 ( .a(n15929), .b(n15799), .o(n27615) );
no02f01 g23825 ( .a(n27615), .b(n27614), .o(n27616) );
na02f01 g23826 ( .a(n27615), .b(n27614), .o(n27617) );
in01f01 g23827 ( .a(n27617), .o(n27618) );
no02f01 g23828 ( .a(n27618), .b(n27616), .o(n27619) );
in01f01 g23829 ( .a(n27619), .o(n27620) );
no02f01 g23830 ( .a(n27620), .b(n27395), .o(n27621) );
no02f01 g23831 ( .a(n27395), .b(n15941), .o(n27622) );
no02f01 g23832 ( .a(n27622), .b(n27621), .o(n27623) );
na03f01 g23833 ( .a(n27623), .b(n27612), .c(n27588), .o(n27624) );
ao12f01 g23834 ( .a(n27367), .b(n27522), .c(n27517), .o(n27625) );
ao12f01 g23835 ( .a(n27367), .b(n27535), .c(n27503), .o(n27626) );
no02f01 g23836 ( .a(n27626), .b(n27625), .o(n27627) );
in01f01 g23837 ( .a(n27627), .o(n27628) );
ao12f01 g23838 ( .a(n27367), .b(n27561), .c(n27548), .o(n27629) );
no02f01 g23839 ( .a(n27629), .b(n27628), .o(n27630) );
in01f01 g23840 ( .a(n27630), .o(n27631) );
ao12f01 g23841 ( .a(n27367), .b(n27583), .c(n27572), .o(n27632) );
no02f01 g23842 ( .a(n27632), .b(n27631), .o(n27633) );
ao12f01 g23843 ( .a(n27367), .b(n27609), .c(n27598), .o(n27634) );
in01f01 g23844 ( .a(n27634), .o(n27635) );
na02f01 g23845 ( .a(n27635), .b(n27633), .o(n27636) );
ao12f01 g23846 ( .a(n27367), .b(n27619), .c(n15984), .o(n27637) );
no02f01 g23847 ( .a(n27637), .b(n27636), .o(n27638) );
no02f01 g23848 ( .a(n27367), .b(n15987), .o(n27639) );
no02f01 g23849 ( .a(n27395), .b(n15946), .o(n27640) );
no02f01 g23850 ( .a(n27640), .b(n27639), .o(n27641) );
na03f01 g23851 ( .a(n27641), .b(n27638), .c(n27624), .o(n27642) );
na02f01 g23852 ( .a(n27316), .b(n27298), .o(n27643) );
na02f01 g23853 ( .a(n27313), .b(n27282), .o(n27644) );
ao12f01 g23854 ( .a(n27322), .b(n27644), .c(n27643), .o(n27645) );
no03f01 g23855 ( .a(n27327), .b(n27297), .c(n27280), .o(n27646) );
ao12f01 g23856 ( .a(n27295), .b(n27325), .c(n27281), .o(n27647) );
in01f01 g23857 ( .a(n27333), .o(n27648) );
oa12f01 g23858 ( .a(n27648), .b(n27647), .c(n27646), .o(n27649) );
oa12f01 g23859 ( .a(n21575), .b(n21589), .c(n15949), .o(n27650) );
na03f01 g23860 ( .a(n21595), .b(n21548), .c(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .o(n27651) );
na03f01 g23861 ( .a(n27343), .b(n27651), .c(n27650), .o(n27652) );
no02f01 g23862 ( .a(n21548), .b(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .o(n27653) );
no02f01 g23863 ( .a(n21548), .b(n15949), .o(n27654) );
no03f01 g23864 ( .a(n27352), .b(n27654), .c(n27653), .o(n27655) );
ao12f01 g23865 ( .a(n27343), .b(n27651), .c(n27650), .o(n27656) );
ao12f01 g23866 ( .a(n27656), .b(n27655), .c(n27652), .o(n27657) );
no03f01 g23867 ( .a(n27648), .b(n27647), .c(n27646), .o(n27658) );
oa12f01 g23868 ( .a(n27649), .b(n27658), .c(n27657), .o(n27659) );
na03f01 g23869 ( .a(n27322), .b(n27644), .c(n27643), .o(n27660) );
ao12f01 g23870 ( .a(n27645), .b(n27660), .c(n27659), .o(n27661) );
no02f01 g23871 ( .a(n27362), .b(n27661), .o(n27662) );
no03f01 g23872 ( .a(n27373), .b(n27662), .c(n27310), .o(n27663) );
in01f01 g23873 ( .a(n27376), .o(n27664) );
in01f01 g23874 ( .a(n27393), .o(n27665) );
oa12f01 g23875 ( .a(n27665), .b(n27664), .c(n27663), .o(n27666) );
in01f01 g23876 ( .a(n27441), .o(n27667) );
in01f01 g23877 ( .a(n27486), .o(n27668) );
na04f01 g23878 ( .a(n27668), .b(n27667), .c(n27400), .d(n27666), .o(n27669) );
in01f01 g23879 ( .a(n27494), .o(n27670) );
na02f01 g23880 ( .a(n27670), .b(n27669), .o(n27671) );
in01f01 g23881 ( .a(n27563), .o(n27672) );
na04f01 g23882 ( .a(n27586), .b(n27672), .c(n27551), .d(n27671), .o(n27673) );
in01f01 g23883 ( .a(n27612), .o(n27674) );
in01f01 g23884 ( .a(n27623), .o(n27675) );
no03f01 g23885 ( .a(n27675), .b(n27674), .c(n27673), .o(n27676) );
in01f01 g23886 ( .a(n27638), .o(n27677) );
in01f01 g23887 ( .a(n27641), .o(n27678) );
oa12f01 g23888 ( .a(n27678), .b(n27677), .c(n27676), .o(n27679) );
na02f01 g23889 ( .a(n27679), .b(n27642), .o(n348) );
in01f01 g23890 ( .a(n_27014), .o(n27681) );
in01f01 g23891 ( .a(n_25834), .o(n27682) );
in01f01 g23892 ( .a(n_44722), .o(n27683) );
no02f01 g23893 ( .a(delay_xor_ln21_unr18_stage7_stallmux_q_3_), .b(n27683), .o(n27684) );
no02f01 g23894 ( .a(n27683), .b(delay_xor_ln21_unr18_stage7_stallmux_q_2_), .o(n27685) );
in01f01 g23895 ( .a(n27685), .o(n27686) );
no02f01 g23896 ( .a(n27683), .b(n_44695), .o(n27687) );
no02f01 g23897 ( .a(n_44422), .b(n27683), .o(n27688) );
no02f01 g23898 ( .a(n27688), .b(n27687), .o(n27689) );
na02f01 g23899 ( .a(n27689), .b(n27686), .o(n27690) );
no02f01 g23900 ( .a(n27690), .b(n27684), .o(n27691) );
no02f01 g23901 ( .a(delay_xor_ln21_unr18_stage7_stallmux_q_6_), .b(n27683), .o(n27692) );
no02f01 g23902 ( .a(delay_xor_ln21_unr18_stage7_stallmux_q_5_), .b(n27683), .o(n27693) );
no02f01 g23903 ( .a(n27683), .b(n_45202), .o(n27694) );
no03f01 g23904 ( .a(n27694), .b(n27693), .c(n27692), .o(n27695) );
na02f01 g23905 ( .a(n27695), .b(n27691), .o(n27696) );
no02f01 g23906 ( .a(delay_xor_ln21_unr18_stage7_stallmux_q_7_), .b(n27683), .o(n27697) );
no02f01 g23907 ( .a(n27697), .b(n27696), .o(n27698) );
in01f01 g23908 ( .a(n27698), .o(n27699) );
no02f01 g23909 ( .a(n27683), .b(delay_xor_ln21_unr18_stage7_stallmux_q_8_), .o(n27700) );
no02f01 g23910 ( .a(n27700), .b(n27699), .o(n27701) );
no02f01 g23911 ( .a(delay_xor_ln21_unr18_stage7_stallmux_q_11_), .b(n27683), .o(n27702) );
no02f01 g23912 ( .a(n27683), .b(delay_xor_ln21_unr18_stage7_stallmux_q_9_), .o(n27703) );
no02f01 g23913 ( .a(n27683), .b(delay_xor_ln21_unr18_stage7_stallmux_q_10_), .o(n27704) );
no03f01 g23914 ( .a(n27704), .b(n27703), .c(n27702), .o(n27705) );
na02f01 g23915 ( .a(n27705), .b(n27701), .o(n27706) );
no02f01 g23916 ( .a(n27683), .b(delay_xor_ln21_unr18_stage7_stallmux_q_12_), .o(n27707) );
no02f01 g23917 ( .a(n27707), .b(n27706), .o(n27708) );
in01f01 g23918 ( .a(n27708), .o(n27709) );
in01f01 g23919 ( .a(delay_xor_ln21_unr18_stage7_stallmux_q_12_), .o(n27710) );
ao12f01 g23920 ( .a(delay_xor_ln21_unr18_stage7_stallmux_q_13_), .b(n27683), .c(n27710), .o(n27711) );
in01f01 g23921 ( .a(delay_xor_ln21_unr18_stage7_stallmux_q_8_), .o(n27712) );
no03f01 g23922 ( .a(delay_xor_ln21_unr18_stage7_stallmux_q_11_), .b(delay_xor_ln21_unr18_stage7_stallmux_q_9_), .c(delay_xor_ln21_unr18_stage7_stallmux_q_10_), .o(n27713) );
ao12f01 g23923 ( .a(n_44722), .b(n27713), .c(n27712), .o(n27714) );
no02f01 g23924 ( .a(n27714), .b(n27711), .o(n27715) );
na02f01 g23925 ( .a(n27715), .b(n27709), .o(n27716) );
in01f01 g23926 ( .a(n27716), .o(n27717) );
in01f01 g23927 ( .a(delay_xor_ln21_unr18_stage7_stallmux_q_13_), .o(n27718) );
no02f01 g23928 ( .a(n_44722), .b(n27718), .o(n27719) );
no02f01 g23929 ( .a(n27719), .b(n27717), .o(n27720) );
in01f01 g23930 ( .a(n27720), .o(n27721) );
ao12f01 g23931 ( .a(n27720), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_28_), .c(delay_sub_ln21_0_unr17_stage7_stallmux_q_29_), .o(n27722) );
no02f01 g23932 ( .a(n27683), .b(delay_xor_ln21_unr18_stage7_stallmux_q_13_), .o(n27723) );
oa12f01 g23933 ( .a(n27708), .b(n27723), .c(n27719), .o(n27724) );
na02f01 g23934 ( .a(n27724), .b(n27716), .o(n27725) );
in01f01 g23935 ( .a(n27725), .o(n27726) );
no02f01 g23936 ( .a(n27726), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_13_), .o(n27727) );
in01f01 g23937 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_12_), .o(n27728) );
no02f01 g23938 ( .a(n_44722), .b(n27710), .o(n27729) );
no02f01 g23939 ( .a(n27729), .b(n27707), .o(n27730) );
in01f01 g23940 ( .a(n27730), .o(n27731) );
ao12f01 g23941 ( .a(n27731), .b(n27705), .c(n27701), .o(n27732) );
no02f01 g23942 ( .a(n27730), .b(n27706), .o(n27733) );
no03f01 g23943 ( .a(n27733), .b(n27732), .c(n27728), .o(n27734) );
in01f01 g23944 ( .a(n27696), .o(n27735) );
no03f01 g23945 ( .a(n27703), .b(n27700), .c(n27697), .o(n27736) );
na02f01 g23946 ( .a(n27736), .b(n27735), .o(n27737) );
in01f01 g23947 ( .a(n27737), .o(n27738) );
no02f01 g23948 ( .a(n27737), .b(n27704), .o(n27739) );
in01f01 g23949 ( .a(n27739), .o(n27740) );
na02f01 g23950 ( .a(delay_xor_ln21_unr18_stage7_stallmux_q_11_), .b(n27683), .o(n27741) );
in01f01 g23951 ( .a(n27741), .o(n27742) );
no02f01 g23952 ( .a(n27742), .b(n27702), .o(n27743) );
no02f01 g23953 ( .a(n27743), .b(n27704), .o(n27744) );
ao22f01 g23954 ( .a(n27744), .b(n27738), .c(n27743), .d(n27740), .o(n27745) );
no02f01 g23955 ( .a(n27745), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_11_), .o(n27746) );
in01f01 g23956 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_10_), .o(n27747) );
na02f01 g23957 ( .a(n27683), .b(delay_xor_ln21_unr18_stage7_stallmux_q_10_), .o(n27748) );
in01f01 g23958 ( .a(n27748), .o(n27749) );
no02f01 g23959 ( .a(n27749), .b(n27704), .o(n27750) );
in01f01 g23960 ( .a(n27750), .o(n27751) );
no02f01 g23961 ( .a(n27751), .b(n27738), .o(n27752) );
no02f01 g23962 ( .a(n27750), .b(n27737), .o(n27753) );
no03f01 g23963 ( .a(n27753), .b(n27752), .c(n27747), .o(n27754) );
na02f01 g23964 ( .a(n27683), .b(delay_xor_ln21_unr18_stage7_stallmux_q_9_), .o(n27755) );
in01f01 g23965 ( .a(n27755), .o(n27756) );
no02f01 g23966 ( .a(n27756), .b(n27703), .o(n27757) );
in01f01 g23967 ( .a(n27757), .o(n27758) );
no02f01 g23968 ( .a(n27758), .b(n27701), .o(n27759) );
na02f01 g23969 ( .a(n27758), .b(n27701), .o(n27760) );
in01f01 g23970 ( .a(n27760), .o(n27761) );
no02f01 g23971 ( .a(n27761), .b(n27759), .o(n27762) );
no02f01 g23972 ( .a(n27762), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_9_), .o(n27763) );
in01f01 g23973 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_8_), .o(n27764) );
no02f01 g23974 ( .a(n_44722), .b(n27712), .o(n27765) );
no02f01 g23975 ( .a(n27765), .b(n27700), .o(n27766) );
in01f01 g23976 ( .a(n27766), .o(n27767) );
no02f01 g23977 ( .a(n27767), .b(n27698), .o(n27768) );
no02f01 g23978 ( .a(n27766), .b(n27699), .o(n27769) );
no02f01 g23979 ( .a(n27769), .b(n27768), .o(n27770) );
in01f01 g23980 ( .a(n27770), .o(n27771) );
no02f01 g23981 ( .a(n27771), .b(n27764), .o(n27772) );
in01f01 g23982 ( .a(n27772), .o(n27773) );
na02f01 g23983 ( .a(delay_xor_ln21_unr18_stage7_stallmux_q_7_), .b(n27683), .o(n27774) );
in01f01 g23984 ( .a(n27774), .o(n27775) );
no02f01 g23985 ( .a(n27775), .b(n27697), .o(n27776) );
in01f01 g23986 ( .a(n27776), .o(n27777) );
no02f01 g23987 ( .a(n27777), .b(n27735), .o(n27778) );
no02f01 g23988 ( .a(n27776), .b(n27696), .o(n27779) );
no02f01 g23989 ( .a(n27779), .b(n27778), .o(n27780) );
no02f01 g23990 ( .a(n27780), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_7_), .o(n27781) );
in01f01 g23991 ( .a(n27781), .o(n27782) );
in01f01 g23992 ( .a(n27693), .o(n27783) );
na02f01 g23993 ( .a(delay_xor_ln21_unr18_stage7_stallmux_q_5_), .b(n27683), .o(n27784) );
na02f01 g23994 ( .a(n27784), .b(n27783), .o(n27785) );
no03f01 g23995 ( .a(n27694), .b(n27690), .c(n27684), .o(n27786) );
no02f01 g23996 ( .a(n27786), .b(n27785), .o(n27787) );
in01f01 g23997 ( .a(n27785), .o(n27788) );
in01f01 g23998 ( .a(n27786), .o(n27789) );
no02f01 g23999 ( .a(n27789), .b(n27788), .o(n27790) );
no02f01 g24000 ( .a(n27790), .b(n27787), .o(n27791) );
no02f01 g24001 ( .a(n27791), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_5_), .o(n27792) );
in01f01 g24002 ( .a(n27792), .o(n27793) );
na02f01 g24003 ( .a(delay_xor_ln21_unr18_stage7_stallmux_q_3_), .b(n27683), .o(n27794) );
in01f01 g24004 ( .a(n27794), .o(n27795) );
no02f01 g24005 ( .a(n27795), .b(n27684), .o(n27796) );
in01f01 g24006 ( .a(n27796), .o(n27797) );
ao12f01 g24007 ( .a(n27797), .b(n27689), .c(n27686), .o(n27798) );
no02f01 g24008 ( .a(n27796), .b(n27690), .o(n27799) );
no02f01 g24009 ( .a(n27799), .b(n27798), .o(n27800) );
no02f01 g24010 ( .a(n27800), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_3_), .o(n27801) );
in01f01 g24011 ( .a(n27801), .o(n27802) );
na02f01 g24012 ( .a(n27683), .b(delay_xor_ln21_unr18_stage7_stallmux_q_2_), .o(n27803) );
na02f01 g24013 ( .a(n27803), .b(n27686), .o(n27804) );
no02f01 g24014 ( .a(n27804), .b(n27689), .o(n27805) );
in01f01 g24015 ( .a(n_44695), .o(n27806) );
na02f01 g24016 ( .a(n_44722), .b(n27806), .o(n27807) );
in01f01 g24017 ( .a(n_44422), .o(n27808) );
na02f01 g24018 ( .a(n27808), .b(n_44722), .o(n27809) );
na02f01 g24019 ( .a(n27809), .b(n27807), .o(n27810) );
ao12f01 g24020 ( .a(n27810), .b(n27803), .c(n27686), .o(n27811) );
no02f01 g24021 ( .a(n27811), .b(n27805), .o(n27812) );
na02f01 g24022 ( .a(n27812), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_2_), .o(n27813) );
in01f01 g24023 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_1_), .o(n27814) );
na02f01 g24024 ( .a(n27809), .b(n27687), .o(n27815) );
no02f01 g24025 ( .a(n27808), .b(n_44722), .o(n27816) );
oa12f01 g24026 ( .a(n27807), .b(n27816), .c(n27688), .o(n27817) );
na02f01 g24027 ( .a(n27817), .b(n27815), .o(n27818) );
no02f01 g24028 ( .a(n27818), .b(n27814), .o(n27819) );
na02f01 g24029 ( .a(n27818), .b(n27814), .o(n27820) );
no02f01 g24030 ( .a(n_44722), .b(n_44695), .o(n27821) );
no02f01 g24031 ( .a(n27683), .b(n27806), .o(n27822) );
no02f01 g24032 ( .a(n27822), .b(n27821), .o(n27823) );
in01f01 g24033 ( .a(n27823), .o(n27824) );
no02f01 g24034 ( .a(n27824), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_0_), .o(n27825) );
in01f01 g24035 ( .a(n27825), .o(n27826) );
ao12f01 g24036 ( .a(n27819), .b(n27826), .c(n27820), .o(n27827) );
no02f01 g24037 ( .a(n27812), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_2_), .o(n27828) );
oa12f01 g24038 ( .a(n27813), .b(n27828), .c(n27827), .o(n27829) );
na02f01 g24039 ( .a(n27800), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_3_), .o(n27830) );
in01f01 g24040 ( .a(n27830), .o(n27831) );
oa12f01 g24041 ( .a(n27802), .b(n27831), .c(n27829), .o(n27832) );
in01f01 g24042 ( .a(n27694), .o(n27833) );
na02f01 g24043 ( .a(n27683), .b(n_45202), .o(n27834) );
na02f01 g24044 ( .a(n27834), .b(n27833), .o(n27835) );
no02f01 g24045 ( .a(n27835), .b(n27691), .o(n27836) );
na02f01 g24046 ( .a(n27835), .b(n27691), .o(n27837) );
in01f01 g24047 ( .a(n27837), .o(n27838) );
no02f01 g24048 ( .a(n27838), .b(n27836), .o(n27839) );
no02f01 g24049 ( .a(n27839), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_4_), .o(n27840) );
no02f01 g24050 ( .a(n27840), .b(n27832), .o(n27841) );
na02f01 g24051 ( .a(n27839), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_4_), .o(n27842) );
na02f01 g24052 ( .a(n27791), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_5_), .o(n27843) );
na02f01 g24053 ( .a(n27843), .b(n27842), .o(n27844) );
oa12f01 g24054 ( .a(n27793), .b(n27844), .c(n27841), .o(n27845) );
no02f01 g24055 ( .a(n27789), .b(n27693), .o(n27846) );
na02f01 g24056 ( .a(delay_xor_ln21_unr18_stage7_stallmux_q_6_), .b(n27683), .o(n27847) );
in01f01 g24057 ( .a(n27847), .o(n27848) );
no02f01 g24058 ( .a(n27848), .b(n27692), .o(n27849) );
in01f01 g24059 ( .a(n27849), .o(n27850) );
na02f01 g24060 ( .a(n27850), .b(n27846), .o(n27851) );
in01f01 g24061 ( .a(n27851), .o(n27852) );
no02f01 g24062 ( .a(n27850), .b(n27846), .o(n27853) );
no02f01 g24063 ( .a(n27853), .b(n27852), .o(n27854) );
no02f01 g24064 ( .a(n27854), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_6_), .o(n27855) );
na02f01 g24065 ( .a(n27780), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_7_), .o(n27856) );
in01f01 g24066 ( .a(n27856), .o(n27857) );
in01f01 g24067 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_6_), .o(n27858) );
no03f01 g24068 ( .a(n27853), .b(n27852), .c(n27858), .o(n27859) );
no02f01 g24069 ( .a(n27859), .b(n27857), .o(n27860) );
oa12f01 g24070 ( .a(n27860), .b(n27855), .c(n27845), .o(n27861) );
na02f01 g24071 ( .a(n27861), .b(n27782), .o(n27862) );
no02f01 g24072 ( .a(n27770), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_8_), .o(n27863) );
oa12f01 g24073 ( .a(n27773), .b(n27863), .c(n27862), .o(n27864) );
na02f01 g24074 ( .a(n27762), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_9_), .o(n27865) );
in01f01 g24075 ( .a(n27865), .o(n27866) );
no02f01 g24076 ( .a(n27866), .b(n27864), .o(n27867) );
no02f01 g24077 ( .a(n27867), .b(n27763), .o(n27868) );
in01f01 g24078 ( .a(n27868), .o(n27869) );
no02f01 g24079 ( .a(n27753), .b(n27752), .o(n27870) );
no02f01 g24080 ( .a(n27870), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_10_), .o(n27871) );
no02f01 g24081 ( .a(n27871), .b(n27869), .o(n27872) );
na02f01 g24082 ( .a(n27745), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_11_), .o(n27873) );
in01f01 g24083 ( .a(n27873), .o(n27874) );
no03f01 g24084 ( .a(n27874), .b(n27872), .c(n27754), .o(n27875) );
no02f01 g24085 ( .a(n27733), .b(n27732), .o(n27876) );
no02f01 g24086 ( .a(n27876), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_12_), .o(n27877) );
no03f01 g24087 ( .a(n27877), .b(n27875), .c(n27746), .o(n27878) );
na02f01 g24088 ( .a(n27726), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_13_), .o(n27879) );
in01f01 g24089 ( .a(n27879), .o(n27880) );
no03f01 g24090 ( .a(n27880), .b(n27878), .c(n27734), .o(n27881) );
in01f01 g24091 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_14_), .o(n27882) );
in01f01 g24092 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_15_), .o(n27883) );
ao12f01 g24093 ( .a(n27721), .b(n27883), .c(n27882), .o(n27884) );
in01f01 g24094 ( .a(n27884), .o(n27885) );
oa12f01 g24095 ( .a(n27885), .b(n27881), .c(n27727), .o(n27886) );
no02f01 g24096 ( .a(n27720), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_14_), .o(n27887) );
no02f01 g24097 ( .a(n27720), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_15_), .o(n27888) );
no02f01 g24098 ( .a(n27888), .b(n27887), .o(n27889) );
na02f01 g24099 ( .a(n27889), .b(n27886), .o(n27890) );
ao12f01 g24100 ( .a(n27720), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_17_), .c(delay_sub_ln21_0_unr17_stage7_stallmux_q_16_), .o(n27891) );
no02f01 g24101 ( .a(n27720), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_18_), .o(n27892) );
no02f01 g24102 ( .a(n27892), .b(n27891), .o(n27893) );
in01f01 g24103 ( .a(n27893), .o(n27894) );
no02f01 g24104 ( .a(n27720), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_19_), .o(n27895) );
no02f01 g24105 ( .a(n27895), .b(n27894), .o(n27896) );
in01f01 g24106 ( .a(n27896), .o(n27897) );
no02f01 g24107 ( .a(n27720), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_21_), .o(n27898) );
no02f01 g24108 ( .a(n27720), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_20_), .o(n27899) );
no03f01 g24109 ( .a(n27899), .b(n27898), .c(n27897), .o(n27900) );
in01f01 g24110 ( .a(n27900), .o(n27901) );
no02f01 g24111 ( .a(n27901), .b(n27890), .o(n27902) );
no02f01 g24112 ( .a(n27720), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_22_), .o(n27903) );
in01f01 g24113 ( .a(n27903), .o(n27904) );
na02f01 g24114 ( .a(n27904), .b(n27902), .o(n27905) );
no02f01 g24115 ( .a(n27720), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_23_), .o(n27906) );
no02f01 g24116 ( .a(n27906), .b(n27905), .o(n27907) );
no02f01 g24117 ( .a(n27720), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_24_), .o(n27908) );
in01f01 g24118 ( .a(n27908), .o(n27909) );
na02f01 g24119 ( .a(n27909), .b(n27907), .o(n27910) );
no02f01 g24120 ( .a(n27720), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_25_), .o(n27911) );
no02f01 g24121 ( .a(n27911), .b(n27910), .o(n27912) );
no02f01 g24122 ( .a(n27720), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_26_), .o(n27913) );
no02f01 g24123 ( .a(n27720), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_27_), .o(n27914) );
no02f01 g24124 ( .a(n27914), .b(n27913), .o(n27915) );
in01f01 g24125 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_18_), .o(n27916) );
in01f01 g24126 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_19_), .o(n27917) );
ao12f01 g24127 ( .a(n27721), .b(n27917), .c(n27916), .o(n27918) );
in01f01 g24128 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_16_), .o(n27919) );
in01f01 g24129 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_17_), .o(n27920) );
ao12f01 g24130 ( .a(n27721), .b(n27920), .c(n27919), .o(n27921) );
no02f01 g24131 ( .a(n27921), .b(n27918), .o(n27922) );
in01f01 g24132 ( .a(n27922), .o(n27923) );
in01f01 g24133 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_20_), .o(n27924) );
in01f01 g24134 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_21_), .o(n27925) );
ao12f01 g24135 ( .a(n27721), .b(n27925), .c(n27924), .o(n27926) );
no02f01 g24136 ( .a(n27926), .b(n27923), .o(n27927) );
in01f01 g24137 ( .a(n27927), .o(n27928) );
in01f01 g24138 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_23_), .o(n27929) );
in01f01 g24139 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_22_), .o(n27930) );
ao12f01 g24140 ( .a(n27721), .b(n27930), .c(n27929), .o(n27931) );
no02f01 g24141 ( .a(n27931), .b(n27928), .o(n27932) );
in01f01 g24142 ( .a(n27932), .o(n27933) );
in01f01 g24143 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_24_), .o(n27934) );
in01f01 g24144 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_25_), .o(n27935) );
ao12f01 g24145 ( .a(n27721), .b(n27935), .c(n27934), .o(n27936) );
no02f01 g24146 ( .a(n27936), .b(n27933), .o(n27937) );
in01f01 g24147 ( .a(n27937), .o(n27938) );
in01f01 g24148 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_26_), .o(n27939) );
in01f01 g24149 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_27_), .o(n27940) );
ao12f01 g24150 ( .a(n27721), .b(n27940), .c(n27939), .o(n27941) );
no02f01 g24151 ( .a(n27941), .b(n27938), .o(n27942) );
in01f01 g24152 ( .a(n27942), .o(n27943) );
ao12f01 g24153 ( .a(n27943), .b(n27915), .c(n27912), .o(n27944) );
in01f01 g24154 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_29_), .o(n27945) );
in01f01 g24155 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_28_), .o(n27946) );
ao12f01 g24156 ( .a(n27721), .b(n27946), .c(n27945), .o(n27947) );
in01f01 g24157 ( .a(n27947), .o(n27948) );
ao12f01 g24158 ( .a(n27722), .b(n27948), .c(n27944), .o(n27949) );
in01f01 g24159 ( .a(n27949), .o(n27950) );
na02f01 g24160 ( .a(n27944), .b(n27721), .o(n27951) );
in01f01 g24161 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_30_), .o(n27952) );
no02f01 g24162 ( .a(n27722), .b(n27952), .o(n27953) );
na02f01 g24163 ( .a(n27953), .b(n27951), .o(n27954) );
oa12f01 g24164 ( .a(n27954), .b(n27950), .c(n27721), .o(n27955) );
no02f01 g24165 ( .a(n27720), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_31_), .o(n27956) );
na02f01 g24166 ( .a(n27720), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_31_), .o(n27957) );
in01f01 g24167 ( .a(n27957), .o(n27958) );
no02f01 g24168 ( .a(n27958), .b(n27956), .o(n27959) );
in01f01 g24169 ( .a(n27959), .o(n27960) );
no02f01 g24170 ( .a(n27960), .b(n27955), .o(n27961) );
na02f01 g24171 ( .a(n27960), .b(n27955), .o(n27962) );
in01f01 g24172 ( .a(n27962), .o(n27963) );
no02f01 g24173 ( .a(n27963), .b(n27961), .o(n27964) );
no02f01 g24174 ( .a(n27964), .b(n27682), .o(n27965) );
no02f01 g24175 ( .a(n27721), .b(n27917), .o(n27966) );
no02f01 g24176 ( .a(n27966), .b(n27895), .o(n27967) );
in01f01 g24177 ( .a(n27967), .o(n27968) );
no02f01 g24178 ( .a(n27894), .b(n27890), .o(n27969) );
no02f01 g24179 ( .a(n27721), .b(n27916), .o(n27970) );
no02f01 g24180 ( .a(n27921), .b(n27970), .o(n27971) );
in01f01 g24181 ( .a(n27971), .o(n27972) );
no03f01 g24182 ( .a(n27972), .b(n27969), .c(n27968), .o(n27973) );
in01f01 g24183 ( .a(n27973), .o(n27974) );
oa12f01 g24184 ( .a(n27968), .b(n27972), .c(n27969), .o(n27975) );
ao12f01 g24185 ( .a(n27682), .b(n27975), .c(n27974), .o(n27976) );
na03f01 g24186 ( .a(n27896), .b(n27889), .c(n27886), .o(n27977) );
no02f01 g24187 ( .a(n27721), .b(n27924), .o(n27978) );
no02f01 g24188 ( .a(n27978), .b(n27899), .o(n27979) );
na03f01 g24189 ( .a(n27979), .b(n27977), .c(n27922), .o(n27980) );
in01f01 g24190 ( .a(n27980), .o(n27981) );
ao12f01 g24191 ( .a(n27979), .b(n27977), .c(n27922), .o(n27982) );
no02f01 g24192 ( .a(n27982), .b(n27981), .o(n27983) );
no02f01 g24193 ( .a(n27983), .b(n27682), .o(n27984) );
no02f01 g24194 ( .a(n27984), .b(n27976), .o(n27985) );
no02f01 g24195 ( .a(n27721), .b(n27925), .o(n27986) );
no02f01 g24196 ( .a(n27986), .b(n27898), .o(n27987) );
in01f01 g24197 ( .a(n27987), .o(n27988) );
no02f01 g24198 ( .a(n27977), .b(n27899), .o(n27989) );
no02f01 g24199 ( .a(n27978), .b(n27923), .o(n27990) );
in01f01 g24200 ( .a(n27990), .o(n27991) );
no03f01 g24201 ( .a(n27991), .b(n27989), .c(n27988), .o(n27992) );
in01f01 g24202 ( .a(n27992), .o(n27993) );
oa12f01 g24203 ( .a(n27988), .b(n27991), .c(n27989), .o(n27994) );
na02f01 g24204 ( .a(n27994), .b(n27993), .o(n27995) );
na02f01 g24205 ( .a(n27995), .b(n_25834), .o(n27996) );
no02f01 g24206 ( .a(n27721), .b(n27930), .o(n27997) );
no02f01 g24207 ( .a(n27997), .b(n27903), .o(n27998) );
no02f01 g24208 ( .a(n27928), .b(n27902), .o(n27999) );
na02f01 g24209 ( .a(n27999), .b(n27998), .o(n28000) );
in01f01 g24210 ( .a(n27998), .o(n28001) );
oa12f01 g24211 ( .a(n28001), .b(n27928), .c(n27902), .o(n28002) );
na02f01 g24212 ( .a(n28002), .b(n28000), .o(n28003) );
na02f01 g24213 ( .a(n28003), .b(n_25834), .o(n28004) );
na03f01 g24214 ( .a(n28004), .b(n27996), .c(n27985), .o(n28005) );
no02f01 g24215 ( .a(n27881), .b(n27727), .o(n28006) );
no02f01 g24216 ( .a(n27884), .b(n28006), .o(n28007) );
in01f01 g24217 ( .a(n27889), .o(n28008) );
no02f01 g24218 ( .a(n28008), .b(n28007), .o(n28009) );
na02f01 g24219 ( .a(n27900), .b(n28009), .o(n28010) );
no02f01 g24220 ( .a(n27903), .b(n28010), .o(n28011) );
no03f01 g24221 ( .a(n27997), .b(n27928), .c(n28011), .o(n28012) );
no02f01 g24222 ( .a(n27721), .b(n27929), .o(n28013) );
no02f01 g24223 ( .a(n28013), .b(n27906), .o(n28014) );
no02f01 g24224 ( .a(n28014), .b(n28012), .o(n28015) );
in01f01 g24225 ( .a(n28015), .o(n28016) );
na02f01 g24226 ( .a(n28014), .b(n28012), .o(n28017) );
na02f01 g24227 ( .a(n28017), .b(n28016), .o(n28018) );
ao12f01 g24228 ( .a(n28005), .b(n28018), .c(n_25834), .o(n28019) );
no02f01 g24229 ( .a(n27933), .b(n27907), .o(n28020) );
no02f01 g24230 ( .a(n27721), .b(n27934), .o(n28021) );
no02f01 g24231 ( .a(n28021), .b(n27908), .o(n28022) );
no02f01 g24232 ( .a(n28022), .b(n28020), .o(n28023) );
na02f01 g24233 ( .a(n28022), .b(n28020), .o(n28024) );
in01f01 g24234 ( .a(n28024), .o(n28025) );
no02f01 g24235 ( .a(n28025), .b(n28023), .o(n28026) );
oa12f01 g24236 ( .a(n28019), .b(n28026), .c(n27682), .o(n28027) );
no02f01 g24237 ( .a(n27721), .b(n27935), .o(n28028) );
no02f01 g24238 ( .a(n28028), .b(n27911), .o(n28029) );
in01f01 g24239 ( .a(n28029), .o(n28030) );
no02f01 g24240 ( .a(n28021), .b(n27933), .o(n28031) );
na02f01 g24241 ( .a(n28031), .b(n27910), .o(n28032) );
no02f01 g24242 ( .a(n28032), .b(n28030), .o(n28033) );
in01f01 g24243 ( .a(n28033), .o(n28034) );
na02f01 g24244 ( .a(n28032), .b(n28030), .o(n28035) );
na02f01 g24245 ( .a(n28035), .b(n28034), .o(n28036) );
ao12f01 g24246 ( .a(n28027), .b(n28036), .c(n_25834), .o(n28037) );
oa12f01 g24247 ( .a(n27937), .b(n27911), .c(n27910), .o(n28038) );
no02f01 g24248 ( .a(n27721), .b(n27939), .o(n28039) );
no02f01 g24249 ( .a(n28039), .b(n27913), .o(n28040) );
in01f01 g24250 ( .a(n28040), .o(n28041) );
na02f01 g24251 ( .a(n28041), .b(n28038), .o(n28042) );
in01f01 g24252 ( .a(n28042), .o(n28043) );
no02f01 g24253 ( .a(n28041), .b(n28038), .o(n28044) );
oa12f01 g24254 ( .a(n27682), .b(n28044), .c(n28043), .o(n28045) );
in01f01 g24255 ( .a(n28044), .o(n28046) );
na03f01 g24256 ( .a(n28046), .b(n28042), .c(n_25834), .o(n28047) );
na02f01 g24257 ( .a(n28036), .b(n27682), .o(n28048) );
na03f01 g24258 ( .a(n28048), .b(n28047), .c(n28045), .o(n28049) );
oa12f01 g24259 ( .a(n27682), .b(n28049), .c(n28037), .o(n28050) );
na02f01 g24260 ( .a(n28047), .b(n28045), .o(n28051) );
in01f01 g24261 ( .a(n28017), .o(n28052) );
no02f01 g24262 ( .a(n28052), .b(n28015), .o(n28053) );
ao12f01 g24263 ( .a(n_25834), .b(n28026), .c(n28053), .o(n28054) );
ao12f01 g24264 ( .a(n28054), .b(n28051), .c(n28037), .o(n28055) );
no02f01 g24265 ( .a(n27721), .b(n27940), .o(n28056) );
no02f01 g24266 ( .a(n28056), .b(n27914), .o(n28057) );
no02f01 g24267 ( .a(n28038), .b(n28039), .o(n28058) );
no02f01 g24268 ( .a(n28058), .b(n27913), .o(n28059) );
in01f01 g24269 ( .a(n28059), .o(n28060) );
no02f01 g24270 ( .a(n28060), .b(n28057), .o(n28061) );
in01f01 g24271 ( .a(n28057), .o(n28062) );
no02f01 g24272 ( .a(n28059), .b(n28062), .o(n28063) );
no02f01 g24273 ( .a(n28063), .b(n28061), .o(n28064) );
no02f01 g24274 ( .a(n27721), .b(n27946), .o(n28065) );
no02f01 g24275 ( .a(n27720), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_28_), .o(n28066) );
no02f01 g24276 ( .a(n28066), .b(n28065), .o(n28067) );
no02f01 g24277 ( .a(n28067), .b(n27944), .o(n28068) );
na02f01 g24278 ( .a(n28067), .b(n27944), .o(n28069) );
in01f01 g24279 ( .a(n28069), .o(n28070) );
no02f01 g24280 ( .a(n28070), .b(n28068), .o(n28071) );
ao12f01 g24281 ( .a(n27682), .b(n28071), .c(n28064), .o(n28072) );
ao12f01 g24282 ( .a(n28072), .b(n28055), .c(n28050), .o(n28073) );
in01f01 g24283 ( .a(n28073), .o(n28074) );
no02f01 g24284 ( .a(n27720), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_30_), .o(n28075) );
no02f01 g24285 ( .a(n27721), .b(n27952), .o(n28076) );
no02f01 g24286 ( .a(n28076), .b(n28075), .o(n28077) );
no02f01 g24287 ( .a(n28077), .b(n27950), .o(n28078) );
na02f01 g24288 ( .a(n28077), .b(n27950), .o(n28079) );
in01f01 g24289 ( .a(n28079), .o(n28080) );
no02f01 g24290 ( .a(n28080), .b(n28078), .o(n28081) );
in01f01 g24291 ( .a(n28065), .o(n28082) );
ao12f01 g24292 ( .a(n28066), .b(n28082), .c(n27944), .o(n28083) );
no02f01 g24293 ( .a(n27720), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_29_), .o(n28084) );
no02f01 g24294 ( .a(n27721), .b(n27945), .o(n28085) );
no02f01 g24295 ( .a(n28085), .b(n28084), .o(n28086) );
in01f01 g24296 ( .a(n28086), .o(n28087) );
na02f01 g24297 ( .a(n28087), .b(n28083), .o(n28088) );
no02f01 g24298 ( .a(n28087), .b(n28083), .o(n28089) );
in01f01 g24299 ( .a(n28089), .o(n28090) );
na02f01 g24300 ( .a(n28090), .b(n28088), .o(n28091) );
in01f01 g24301 ( .a(n28091), .o(n28092) );
ao12f01 g24302 ( .a(n27682), .b(n28092), .c(n28081), .o(n28093) );
no02f01 g24303 ( .a(n28093), .b(n28074), .o(n28094) );
ao12f01 g24304 ( .a(n_25834), .b(n28071), .c(n28064), .o(n28095) );
ao12f01 g24305 ( .a(n28095), .b(n28091), .c(n27682), .o(n28096) );
oa12f01 g24306 ( .a(n28096), .b(n28081), .c(n_25834), .o(n28097) );
no02f01 g24307 ( .a(n28097), .b(n28094), .o(n28098) );
in01f01 g24308 ( .a(n28098), .o(n28099) );
no02f01 g24309 ( .a(n27964), .b(n_25834), .o(n28100) );
in01f01 g24310 ( .a(n28100), .o(n28101) );
ao12f01 g24311 ( .a(n27965), .b(n28101), .c(n28099), .o(n28102) );
no02f01 g24312 ( .a(n27683), .b(delay_xor_ln22_unr18_stage7_stallmux_q_4_), .o(n28103) );
no02f01 g24313 ( .a(delay_xor_ln22_unr18_stage7_stallmux_q_3_), .b(n27683), .o(n28104) );
in01f01 g24314 ( .a(n28104), .o(n28105) );
no02f01 g24315 ( .a(delay_xor_ln22_unr18_stage7_stallmux_q_2_), .b(n27683), .o(n28106) );
in01f01 g24316 ( .a(delay_xor_ln22_unr18_stage7_stallmux_q_1_), .o(n28107) );
na02f01 g24317 ( .a(n28107), .b(n_44722), .o(n28108) );
in01f01 g24318 ( .a(delay_xor_ln22_unr18_stage7_stallmux_q_0_), .o(n28109) );
na02f01 g24319 ( .a(n_44722), .b(n28109), .o(n28110) );
na02f01 g24320 ( .a(n28110), .b(n28108), .o(n28111) );
no02f01 g24321 ( .a(n28111), .b(n28106), .o(n28112) );
na02f01 g24322 ( .a(n28112), .b(n28105), .o(n28113) );
no02f01 g24323 ( .a(n28113), .b(n28103), .o(n28114) );
no02f01 g24324 ( .a(n27683), .b(delay_xor_ln22_unr18_stage7_stallmux_q_5_), .o(n28115) );
in01f01 g24325 ( .a(n28115), .o(n28116) );
na02f01 g24326 ( .a(n28116), .b(n28114), .o(n28117) );
no02f01 g24327 ( .a(n27683), .b(delay_xor_ln22_unr18_stage7_stallmux_q_6_), .o(n28118) );
no02f01 g24328 ( .a(n28118), .b(n28117), .o(n28119) );
in01f01 g24329 ( .a(n28119), .o(n28120) );
no02f01 g24330 ( .a(n27683), .b(delay_xor_ln22_unr18_stage7_stallmux_q_7_), .o(n28121) );
no02f01 g24331 ( .a(delay_xor_ln22_unr18_stage7_stallmux_q_8_), .b(n27683), .o(n28122) );
no03f01 g24332 ( .a(n28122), .b(n28121), .c(n28120), .o(n28123) );
no02f01 g24333 ( .a(delay_xor_ln22_unr18_stage7_stallmux_q_9_), .b(n27683), .o(n28124) );
in01f01 g24334 ( .a(n28124), .o(n28125) );
na02f01 g24335 ( .a(n28125), .b(n28123), .o(n28126) );
no02f01 g24336 ( .a(delay_xor_ln22_unr18_stage7_stallmux_q_10_), .b(n27683), .o(n28127) );
no02f01 g24337 ( .a(n28127), .b(n28126), .o(n28128) );
in01f01 g24338 ( .a(n28128), .o(n28129) );
no02f01 g24339 ( .a(delay_xor_ln22_unr18_stage7_stallmux_q_11_), .b(n27683), .o(n28130) );
no02f01 g24340 ( .a(n28130), .b(n28129), .o(n28131) );
in01f01 g24341 ( .a(n28131), .o(n28132) );
no02f01 g24342 ( .a(n27683), .b(delay_xor_ln22_unr18_stage7_stallmux_q_12_), .o(n28133) );
no02f01 g24343 ( .a(n28133), .b(n28132), .o(n28134) );
in01f01 g24344 ( .a(delay_xor_ln22_unr18_stage7_stallmux_q_8_), .o(n28135) );
no03f01 g24345 ( .a(delay_xor_ln22_unr18_stage7_stallmux_q_11_), .b(delay_xor_ln22_unr18_stage7_stallmux_q_10_), .c(delay_xor_ln22_unr18_stage7_stallmux_q_9_), .o(n28136) );
ao12f01 g24346 ( .a(n_44722), .b(n28136), .c(n28135), .o(n28137) );
in01f01 g24347 ( .a(delay_xor_ln22_unr18_stage7_stallmux_q_12_), .o(n28138) );
ao12f01 g24348 ( .a(delay_xor_ln22_unr18_stage7_stallmux_q_13_), .b(n27683), .c(n28138), .o(n28139) );
no03f01 g24349 ( .a(n28139), .b(n28137), .c(n28134), .o(n28140) );
in01f01 g24350 ( .a(delay_xor_ln22_unr18_stage7_stallmux_q_13_), .o(n28141) );
no02f01 g24351 ( .a(n_44722), .b(n28141), .o(n28142) );
no02f01 g24352 ( .a(n28142), .b(n28140), .o(n28143) );
in01f01 g24353 ( .a(n28143), .o(n28144) );
ao12f01 g24354 ( .a(n28144), .b(delay_add_ln22_unr17_stage7_stallmux_q_28_), .c(delay_add_ln22_unr17_stage7_stallmux_q_29_), .o(n28145) );
no02f01 g24355 ( .a(n28144), .b(delay_add_ln22_unr17_stage7_stallmux_q_23_), .o(n28146) );
in01f01 g24356 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_13_), .o(n28147) );
in01f01 g24357 ( .a(n28134), .o(n28148) );
in01f01 g24358 ( .a(n28142), .o(n28149) );
no02f01 g24359 ( .a(n27683), .b(delay_xor_ln22_unr18_stage7_stallmux_q_13_), .o(n28150) );
in01f01 g24360 ( .a(n28150), .o(n28151) );
ao12f01 g24361 ( .a(n28148), .b(n28151), .c(n28149), .o(n28152) );
no02f01 g24362 ( .a(n28152), .b(n28140), .o(n28153) );
no02f01 g24363 ( .a(n28153), .b(n28147), .o(n28154) );
in01f01 g24364 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_12_), .o(n28155) );
no02f01 g24365 ( .a(n_44722), .b(n28138), .o(n28156) );
no02f01 g24366 ( .a(n28156), .b(n28133), .o(n28157) );
in01f01 g24367 ( .a(n28157), .o(n28158) );
no02f01 g24368 ( .a(n28158), .b(n28131), .o(n28159) );
na02f01 g24369 ( .a(n28158), .b(n28131), .o(n28160) );
in01f01 g24370 ( .a(n28160), .o(n28161) );
no02f01 g24371 ( .a(n28161), .b(n28159), .o(n28162) );
no02f01 g24372 ( .a(n28162), .b(n28155), .o(n28163) );
in01f01 g24373 ( .a(n28163), .o(n28164) );
na02f01 g24374 ( .a(delay_xor_ln22_unr18_stage7_stallmux_q_11_), .b(n27683), .o(n28165) );
in01f01 g24375 ( .a(n28165), .o(n28166) );
no02f01 g24376 ( .a(n28166), .b(n28130), .o(n28167) );
in01f01 g24377 ( .a(n28167), .o(n28168) );
no02f01 g24378 ( .a(n28168), .b(n28128), .o(n28169) );
in01f01 g24379 ( .a(n28169), .o(n28170) );
na02f01 g24380 ( .a(n28168), .b(n28128), .o(n28171) );
na02f01 g24381 ( .a(n28171), .b(n28170), .o(n28172) );
no02f01 g24382 ( .a(n28172), .b(delay_add_ln22_unr17_stage7_stallmux_q_11_), .o(n28173) );
in01f01 g24383 ( .a(n28173), .o(n28174) );
in01f01 g24384 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_10_), .o(n28175) );
na02f01 g24385 ( .a(delay_xor_ln22_unr18_stage7_stallmux_q_10_), .b(n27683), .o(n28176) );
in01f01 g24386 ( .a(n28176), .o(n28177) );
no02f01 g24387 ( .a(n28177), .b(n28127), .o(n28178) );
no02f01 g24388 ( .a(n28178), .b(n28126), .o(n28179) );
na02f01 g24389 ( .a(n28178), .b(n28126), .o(n28180) );
in01f01 g24390 ( .a(n28180), .o(n28181) );
no02f01 g24391 ( .a(n28181), .b(n28179), .o(n28182) );
no02f01 g24392 ( .a(n28182), .b(n28175), .o(n28183) );
in01f01 g24393 ( .a(n28183), .o(n28184) );
in01f01 g24394 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_9_), .o(n28185) );
na02f01 g24395 ( .a(delay_xor_ln22_unr18_stage7_stallmux_q_9_), .b(n27683), .o(n28186) );
na02f01 g24396 ( .a(n28186), .b(n28125), .o(n28187) );
no02f01 g24397 ( .a(n28187), .b(n28123), .o(n28188) );
in01f01 g24398 ( .a(n28188), .o(n28189) );
na02f01 g24399 ( .a(n28187), .b(n28123), .o(n28190) );
ao12f01 g24400 ( .a(n28185), .b(n28190), .c(n28189), .o(n28191) );
in01f01 g24401 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_8_), .o(n28192) );
no02f01 g24402 ( .a(n28121), .b(n28120), .o(n28193) );
no02f01 g24403 ( .a(n28135), .b(n_44722), .o(n28194) );
no02f01 g24404 ( .a(n28194), .b(n28122), .o(n28195) );
in01f01 g24405 ( .a(n28195), .o(n28196) );
no02f01 g24406 ( .a(n28196), .b(n28193), .o(n28197) );
na02f01 g24407 ( .a(n28196), .b(n28193), .o(n28198) );
in01f01 g24408 ( .a(n28198), .o(n28199) );
no02f01 g24409 ( .a(n28199), .b(n28197), .o(n28200) );
no02f01 g24410 ( .a(n28200), .b(n28192), .o(n28201) );
in01f01 g24411 ( .a(n28201), .o(n28202) );
na02f01 g24412 ( .a(n27683), .b(delay_xor_ln22_unr18_stage7_stallmux_q_7_), .o(n28203) );
in01f01 g24413 ( .a(n28203), .o(n28204) );
no02f01 g24414 ( .a(n28204), .b(n28121), .o(n28205) );
in01f01 g24415 ( .a(n28205), .o(n28206) );
na02f01 g24416 ( .a(n28206), .b(n28119), .o(n28207) );
no02f01 g24417 ( .a(n28206), .b(n28119), .o(n28208) );
in01f01 g24418 ( .a(n28208), .o(n28209) );
na02f01 g24419 ( .a(n28209), .b(n28207), .o(n28210) );
no02f01 g24420 ( .a(n28210), .b(delay_add_ln22_unr17_stage7_stallmux_q_7_), .o(n28211) );
in01f01 g24421 ( .a(n28211), .o(n28212) );
in01f01 g24422 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_6_), .o(n28213) );
na02f01 g24423 ( .a(n27683), .b(delay_xor_ln22_unr18_stage7_stallmux_q_6_), .o(n28214) );
in01f01 g24424 ( .a(n28214), .o(n28215) );
no02f01 g24425 ( .a(n28215), .b(n28118), .o(n28216) );
na02f01 g24426 ( .a(n28216), .b(n28117), .o(n28217) );
in01f01 g24427 ( .a(n28217), .o(n28218) );
no02f01 g24428 ( .a(n28216), .b(n28117), .o(n28219) );
no02f01 g24429 ( .a(n28219), .b(n28218), .o(n28220) );
no02f01 g24430 ( .a(n28220), .b(n28213), .o(n28221) );
in01f01 g24431 ( .a(n28221), .o(n28222) );
in01f01 g24432 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_5_), .o(n28223) );
na02f01 g24433 ( .a(n27683), .b(delay_xor_ln22_unr18_stage7_stallmux_q_5_), .o(n28224) );
na02f01 g24434 ( .a(n28224), .b(n28116), .o(n28225) );
na02f01 g24435 ( .a(n28225), .b(n28114), .o(n28226) );
no02f01 g24436 ( .a(n28225), .b(n28114), .o(n28227) );
in01f01 g24437 ( .a(n28227), .o(n28228) );
ao12f01 g24438 ( .a(n28223), .b(n28228), .c(n28226), .o(n28229) );
na02f01 g24439 ( .a(n27683), .b(delay_xor_ln22_unr18_stage7_stallmux_q_4_), .o(n28230) );
in01f01 g24440 ( .a(n28230), .o(n28231) );
no02f01 g24441 ( .a(n28231), .b(n28103), .o(n28232) );
na02f01 g24442 ( .a(n28232), .b(n28113), .o(n28233) );
no02f01 g24443 ( .a(n28232), .b(n28113), .o(n28234) );
in01f01 g24444 ( .a(n28234), .o(n28235) );
na02f01 g24445 ( .a(n28235), .b(n28233), .o(n28236) );
no02f01 g24446 ( .a(n28236), .b(delay_add_ln22_unr17_stage7_stallmux_q_4_), .o(n28237) );
na02f01 g24447 ( .a(delay_xor_ln22_unr18_stage7_stallmux_q_3_), .b(n27683), .o(n28238) );
na02f01 g24448 ( .a(n28238), .b(n28105), .o(n28239) );
in01f01 g24449 ( .a(n28239), .o(n28240) );
oa12f01 g24450 ( .a(n28240), .b(n28111), .c(n28106), .o(n28241) );
na02f01 g24451 ( .a(n28239), .b(n28112), .o(n28242) );
na02f01 g24452 ( .a(n28242), .b(n28241), .o(n28243) );
no02f01 g24453 ( .a(n28243), .b(delay_add_ln22_unr17_stage7_stallmux_q_3_), .o(n28244) );
no02f01 g24454 ( .a(delay_xor_ln22_unr18_stage7_stallmux_q_1_), .b(n27683), .o(n28245) );
no02f01 g24455 ( .a(n27683), .b(delay_xor_ln22_unr18_stage7_stallmux_q_0_), .o(n28246) );
no02f01 g24456 ( .a(n28246), .b(n28245), .o(n28247) );
in01f01 g24457 ( .a(delay_xor_ln22_unr18_stage7_stallmux_q_2_), .o(n28248) );
na02f01 g24458 ( .a(n28248), .b(n_44722), .o(n28249) );
na02f01 g24459 ( .a(delay_xor_ln22_unr18_stage7_stallmux_q_2_), .b(n27683), .o(n28250) );
na02f01 g24460 ( .a(n28250), .b(n28249), .o(n28251) );
na02f01 g24461 ( .a(n28251), .b(n28247), .o(n28252) );
na03f01 g24462 ( .a(n28250), .b(n28111), .c(n28249), .o(n28253) );
na02f01 g24463 ( .a(n28253), .b(n28252), .o(n28254) );
no02f01 g24464 ( .a(n28254), .b(delay_add_ln22_unr17_stage7_stallmux_q_2_), .o(n28255) );
in01f01 g24465 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_1_), .o(n28256) );
no02f01 g24466 ( .a(n_44722), .b(delay_xor_ln22_unr18_stage7_stallmux_q_0_), .o(n28257) );
no02f01 g24467 ( .a(n27683), .b(n28109), .o(n28258) );
no02f01 g24468 ( .a(n28258), .b(n28257), .o(n28259) );
na02f01 g24469 ( .a(n28259), .b(delay_add_ln22_unr17_stage7_stallmux_q_0_), .o(n28260) );
no02f01 g24470 ( .a(n28260), .b(n28256), .o(n28261) );
na03f01 g24471 ( .a(delay_xor_ln22_unr18_stage7_stallmux_q_1_), .b(n_44722), .c(n28109), .o(n28262) );
no02f01 g24472 ( .a(n28107), .b(n_44722), .o(n28263) );
oa12f01 g24473 ( .a(n28110), .b(n28263), .c(n28245), .o(n28264) );
na02f01 g24474 ( .a(n28264), .b(n28262), .o(n28265) );
na02f01 g24475 ( .a(n28260), .b(n28256), .o(n28266) );
ao12f01 g24476 ( .a(n28261), .b(n28266), .c(n28265), .o(n28267) );
na02f01 g24477 ( .a(n28254), .b(delay_add_ln22_unr17_stage7_stallmux_q_2_), .o(n28268) );
oa12f01 g24478 ( .a(n28268), .b(n28267), .c(n28255), .o(n28269) );
in01f01 g24479 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_3_), .o(n28270) );
ao12f01 g24480 ( .a(n28270), .b(n28242), .c(n28241), .o(n28271) );
no02f01 g24481 ( .a(n28271), .b(n28269), .o(n28272) );
no03f01 g24482 ( .a(n28272), .b(n28244), .c(n28237), .o(n28273) );
in01f01 g24483 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_4_), .o(n28274) );
ao12f01 g24484 ( .a(n28274), .b(n28235), .c(n28233), .o(n28275) );
no02f01 g24485 ( .a(n28275), .b(n28273), .o(n28276) );
in01f01 g24486 ( .a(n28226), .o(n28277) );
no03f01 g24487 ( .a(n28227), .b(n28277), .c(delay_add_ln22_unr17_stage7_stallmux_q_5_), .o(n28278) );
no02f01 g24488 ( .a(n28278), .b(n28276), .o(n28279) );
no03f01 g24489 ( .a(n28219), .b(n28218), .c(delay_add_ln22_unr17_stage7_stallmux_q_6_), .o(n28280) );
in01f01 g24490 ( .a(n28280), .o(n28281) );
oa12f01 g24491 ( .a(n28281), .b(n28279), .c(n28229), .o(n28282) );
in01f01 g24492 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_7_), .o(n28283) );
ao12f01 g24493 ( .a(n28283), .b(n28209), .c(n28207), .o(n28284) );
in01f01 g24494 ( .a(n28284), .o(n28285) );
na03f01 g24495 ( .a(n28285), .b(n28282), .c(n28222), .o(n28286) );
no03f01 g24496 ( .a(n28199), .b(n28197), .c(delay_add_ln22_unr17_stage7_stallmux_q_8_), .o(n28287) );
in01f01 g24497 ( .a(n28287), .o(n28288) );
na03f01 g24498 ( .a(n28288), .b(n28286), .c(n28212), .o(n28289) );
in01f01 g24499 ( .a(n28190), .o(n28290) );
no03f01 g24500 ( .a(n28290), .b(n28188), .c(delay_add_ln22_unr17_stage7_stallmux_q_9_), .o(n28291) );
ao12f01 g24501 ( .a(n28291), .b(n28289), .c(n28202), .o(n28292) );
no03f01 g24502 ( .a(n28181), .b(n28179), .c(delay_add_ln22_unr17_stage7_stallmux_q_10_), .o(n28293) );
in01f01 g24503 ( .a(n28293), .o(n28294) );
oa12f01 g24504 ( .a(n28294), .b(n28292), .c(n28191), .o(n28295) );
in01f01 g24505 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_11_), .o(n28296) );
ao12f01 g24506 ( .a(n28296), .b(n28171), .c(n28170), .o(n28297) );
in01f01 g24507 ( .a(n28297), .o(n28298) );
na03f01 g24508 ( .a(n28298), .b(n28295), .c(n28184), .o(n28299) );
no03f01 g24509 ( .a(n28161), .b(n28159), .c(delay_add_ln22_unr17_stage7_stallmux_q_12_), .o(n28300) );
in01f01 g24510 ( .a(n28300), .o(n28301) );
na03f01 g24511 ( .a(n28301), .b(n28299), .c(n28174), .o(n28302) );
no03f01 g24512 ( .a(n28152), .b(n28140), .c(delay_add_ln22_unr17_stage7_stallmux_q_13_), .o(n28303) );
ao12f01 g24513 ( .a(n28303), .b(n28302), .c(n28164), .o(n28304) );
in01f01 g24514 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_14_), .o(n28305) );
in01f01 g24515 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_15_), .o(n28306) );
ao12f01 g24516 ( .a(n28143), .b(n28306), .c(n28305), .o(n28307) );
no03f01 g24517 ( .a(n28307), .b(n28304), .c(n28154), .o(n28308) );
no02f01 g24518 ( .a(n28144), .b(delay_add_ln22_unr17_stage7_stallmux_q_15_), .o(n28309) );
no02f01 g24519 ( .a(n28144), .b(delay_add_ln22_unr17_stage7_stallmux_q_14_), .o(n28310) );
no02f01 g24520 ( .a(n28310), .b(n28309), .o(n28311) );
in01f01 g24521 ( .a(n28311), .o(n28312) );
in01f01 g24522 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_16_), .o(n28313) );
in01f01 g24523 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_17_), .o(n28314) );
no02f01 g24524 ( .a(n28314), .b(n28313), .o(n28315) );
no02f01 g24525 ( .a(n28315), .b(n28144), .o(n28316) );
no02f01 g24526 ( .a(n28144), .b(delay_add_ln22_unr17_stage7_stallmux_q_18_), .o(n28317) );
no02f01 g24527 ( .a(n28317), .b(n28316), .o(n28318) );
in01f01 g24528 ( .a(n28318), .o(n28319) );
no02f01 g24529 ( .a(n28144), .b(delay_add_ln22_unr17_stage7_stallmux_q_19_), .o(n28320) );
no04f01 g24530 ( .a(n28320), .b(n28319), .c(n28312), .d(n28308), .o(n28321) );
no02f01 g24531 ( .a(n28144), .b(delay_add_ln22_unr17_stage7_stallmux_q_20_), .o(n28322) );
in01f01 g24532 ( .a(n28322), .o(n28323) );
na02f01 g24533 ( .a(n28323), .b(n28321), .o(n28324) );
no02f01 g24534 ( .a(n28144), .b(delay_add_ln22_unr17_stage7_stallmux_q_21_), .o(n28325) );
no02f01 g24535 ( .a(n28325), .b(n28324), .o(n28326) );
no02f01 g24536 ( .a(n28144), .b(delay_add_ln22_unr17_stage7_stallmux_q_22_), .o(n28327) );
in01f01 g24537 ( .a(n28327), .o(n28328) );
na02f01 g24538 ( .a(n28328), .b(n28326), .o(n28329) );
no02f01 g24539 ( .a(n28329), .b(n28146), .o(n28330) );
no02f01 g24540 ( .a(n28144), .b(delay_add_ln22_unr17_stage7_stallmux_q_24_), .o(n28331) );
in01f01 g24541 ( .a(n28331), .o(n28332) );
na02f01 g24542 ( .a(n28332), .b(n28330), .o(n28333) );
no02f01 g24543 ( .a(n28144), .b(delay_add_ln22_unr17_stage7_stallmux_q_25_), .o(n28334) );
no02f01 g24544 ( .a(n28334), .b(n28333), .o(n28335) );
no02f01 g24545 ( .a(n28144), .b(delay_add_ln22_unr17_stage7_stallmux_q_27_), .o(n28336) );
no02f01 g24546 ( .a(n28144), .b(delay_add_ln22_unr17_stage7_stallmux_q_26_), .o(n28337) );
no02f01 g24547 ( .a(n28337), .b(n28336), .o(n28338) );
ao12f01 g24548 ( .a(n28143), .b(n28314), .c(n28313), .o(n28339) );
in01f01 g24549 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_18_), .o(n28340) );
no02f01 g24550 ( .a(n28143), .b(n28340), .o(n28341) );
no02f01 g24551 ( .a(n28341), .b(n28339), .o(n28342) );
in01f01 g24552 ( .a(n28342), .o(n28343) );
na02f01 g24553 ( .a(n28144), .b(delay_add_ln22_unr17_stage7_stallmux_q_19_), .o(n28344) );
in01f01 g24554 ( .a(n28344), .o(n28345) );
no02f01 g24555 ( .a(n28345), .b(n28343), .o(n28346) );
in01f01 g24556 ( .a(n28346), .o(n28347) );
in01f01 g24557 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_21_), .o(n28348) );
in01f01 g24558 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_20_), .o(n28349) );
ao12f01 g24559 ( .a(n28143), .b(n28349), .c(n28348), .o(n28350) );
no02f01 g24560 ( .a(n28350), .b(n28347), .o(n28351) );
in01f01 g24561 ( .a(n28351), .o(n28352) );
in01f01 g24562 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_22_), .o(n28353) );
in01f01 g24563 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_23_), .o(n28354) );
ao12f01 g24564 ( .a(n28143), .b(n28354), .c(n28353), .o(n28355) );
no02f01 g24565 ( .a(n28355), .b(n28352), .o(n28356) );
in01f01 g24566 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_24_), .o(n28357) );
in01f01 g24567 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_25_), .o(n28358) );
ao12f01 g24568 ( .a(n28143), .b(n28358), .c(n28357), .o(n28359) );
na02f01 g24569 ( .a(n28144), .b(delay_add_ln22_unr17_stage7_stallmux_q_27_), .o(n28360) );
in01f01 g24570 ( .a(n28360), .o(n28361) );
na02f01 g24571 ( .a(n28144), .b(delay_add_ln22_unr17_stage7_stallmux_q_26_), .o(n28362) );
in01f01 g24572 ( .a(n28362), .o(n28363) );
no03f01 g24573 ( .a(n28363), .b(n28361), .c(n28359), .o(n28364) );
na02f01 g24574 ( .a(n28364), .b(n28356), .o(n28365) );
ao12f01 g24575 ( .a(n28365), .b(n28338), .c(n28335), .o(n28366) );
in01f01 g24576 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_29_), .o(n28367) );
in01f01 g24577 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_28_), .o(n28368) );
ao12f01 g24578 ( .a(n28143), .b(n28368), .c(n28367), .o(n28369) );
in01f01 g24579 ( .a(n28369), .o(n28370) );
ao12f01 g24580 ( .a(n28145), .b(n28370), .c(n28366), .o(n28371) );
in01f01 g24581 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_30_), .o(n28372) );
no02f01 g24582 ( .a(n28143), .b(n28372), .o(n28373) );
no02f01 g24583 ( .a(n28144), .b(delay_add_ln22_unr17_stage7_stallmux_q_30_), .o(n28374) );
no02f01 g24584 ( .a(n28374), .b(n28373), .o(n28375) );
in01f01 g24585 ( .a(n28375), .o(n28376) );
no02f01 g24586 ( .a(n28376), .b(n28371), .o(n28377) );
na02f01 g24587 ( .a(n28376), .b(n28371), .o(n28378) );
in01f01 g24588 ( .a(n28378), .o(n28379) );
no02f01 g24589 ( .a(n28379), .b(n28377), .o(n28380) );
in01f01 g24590 ( .a(n28380), .o(n28381) );
no02f01 g24591 ( .a(n28381), .b(n28102), .o(n28382) );
in01f01 g24592 ( .a(n28102), .o(n28383) );
no02f01 g24593 ( .a(n28380), .b(n28383), .o(n28384) );
no02f01 g24594 ( .a(n28384), .b(n28382), .o(n28385) );
no02f01 g24595 ( .a(n28100), .b(n27965), .o(n28386) );
na02f01 g24596 ( .a(n28386), .b(n28098), .o(n28387) );
no02f01 g24597 ( .a(n28386), .b(n28098), .o(n28388) );
in01f01 g24598 ( .a(n28388), .o(n28389) );
na02f01 g24599 ( .a(n28389), .b(n28387), .o(n28390) );
in01f01 g24600 ( .a(n28299), .o(n28391) );
no02f01 g24601 ( .a(n28391), .b(n28173), .o(n28392) );
no02f01 g24602 ( .a(n28300), .b(n28163), .o(n28393) );
in01f01 g24603 ( .a(n28393), .o(n28394) );
no02f01 g24604 ( .a(n28394), .b(n28392), .o(n28395) );
na02f01 g24605 ( .a(n28394), .b(n28392), .o(n28396) );
in01f01 g24606 ( .a(n28396), .o(n28397) );
no02f01 g24607 ( .a(n28397), .b(n28395), .o(n28398) );
in01f01 g24608 ( .a(n28398), .o(n28399) );
na02f01 g24609 ( .a(n28399), .b(n28390), .o(n28400) );
in01f01 g24610 ( .a(n28302), .o(n28401) );
no02f01 g24611 ( .a(n28401), .b(n28163), .o(n28402) );
no02f01 g24612 ( .a(n28303), .b(n28154), .o(n28403) );
no02f01 g24613 ( .a(n28403), .b(n28402), .o(n28404) );
na02f01 g24614 ( .a(n28403), .b(n28402), .o(n28405) );
in01f01 g24615 ( .a(n28405), .o(n28406) );
no02f01 g24616 ( .a(n28406), .b(n28404), .o(n28407) );
in01f01 g24617 ( .a(n28407), .o(n28408) );
na02f01 g24618 ( .a(n28408), .b(n28102), .o(n28409) );
no02f01 g24619 ( .a(n28408), .b(n28102), .o(n28410) );
ao12f01 g24620 ( .a(n28410), .b(n28409), .c(n28400), .o(n28411) );
in01f01 g24621 ( .a(n28411), .o(n28412) );
in01f01 g24622 ( .a(n28410), .o(n28413) );
in01f01 g24623 ( .a(n28081), .o(n28414) );
na02f01 g24624 ( .a(n28091), .b(n_25834), .o(n28415) );
na02f01 g24625 ( .a(n28415), .b(n28073), .o(n28416) );
na02f01 g24626 ( .a(n28416), .b(n28096), .o(n28417) );
no02f01 g24627 ( .a(n28417), .b(n28414), .o(n28418) );
ao12f01 g24628 ( .a(n28081), .b(n28416), .c(n28096), .o(n28419) );
in01f01 g24629 ( .a(n28295), .o(n28420) );
no02f01 g24630 ( .a(n28297), .b(n28173), .o(n28421) );
in01f01 g24631 ( .a(n28421), .o(n28422) );
no03f01 g24632 ( .a(n28422), .b(n28420), .c(n28183), .o(n28423) );
ao12f01 g24633 ( .a(n28421), .b(n28295), .c(n28184), .o(n28424) );
no02f01 g24634 ( .a(n28424), .b(n28423), .o(n28425) );
in01f01 g24635 ( .a(n28425), .o(n28426) );
no03f01 g24636 ( .a(n28426), .b(n28419), .c(n28418), .o(n28427) );
in01f01 g24637 ( .a(n28427), .o(n28428) );
na02f01 g24638 ( .a(n28055), .b(n28050), .o(n28429) );
no02f01 g24639 ( .a(n28064), .b(n27682), .o(n28430) );
in01f01 g24640 ( .a(n28430), .o(n28431) );
na02f01 g24641 ( .a(n28431), .b(n28429), .o(n28432) );
no02f01 g24642 ( .a(n28064), .b(n_25834), .o(n28433) );
in01f01 g24643 ( .a(n28433), .o(n28434) );
ao12f01 g24644 ( .a(n28071), .b(n28434), .c(n28432), .o(n28435) );
in01f01 g24645 ( .a(n28071), .o(n28436) );
ao12f01 g24646 ( .a(n28430), .b(n28055), .c(n28050), .o(n28437) );
no03f01 g24647 ( .a(n28433), .b(n28437), .c(n28436), .o(n28438) );
in01f01 g24648 ( .a(n28289), .o(n28439) );
no02f01 g24649 ( .a(n28291), .b(n28191), .o(n28440) );
in01f01 g24650 ( .a(n28440), .o(n28441) );
no03f01 g24651 ( .a(n28441), .b(n28439), .c(n28201), .o(n28442) );
ao12f01 g24652 ( .a(n28440), .b(n28289), .c(n28202), .o(n28443) );
no02f01 g24653 ( .a(n28443), .b(n28442), .o(n28444) );
in01f01 g24654 ( .a(n28444), .o(n28445) );
oa12f01 g24655 ( .a(n28445), .b(n28438), .c(n28435), .o(n28446) );
no02f01 g24656 ( .a(n28433), .b(n28430), .o(n28447) );
ao12f01 g24657 ( .a(n28447), .b(n28055), .c(n28050), .o(n28448) );
in01f01 g24658 ( .a(n28448), .o(n28449) );
na03f01 g24659 ( .a(n28447), .b(n28055), .c(n28050), .o(n28450) );
in01f01 g24660 ( .a(n28286), .o(n28451) );
no02f01 g24661 ( .a(n28451), .b(n28211), .o(n28452) );
no02f01 g24662 ( .a(n28287), .b(n28201), .o(n28453) );
in01f01 g24663 ( .a(n28453), .o(n28454) );
no02f01 g24664 ( .a(n28454), .b(n28452), .o(n28455) );
na02f01 g24665 ( .a(n28454), .b(n28452), .o(n28456) );
in01f01 g24666 ( .a(n28456), .o(n28457) );
no02f01 g24667 ( .a(n28457), .b(n28455), .o(n28458) );
ao12f01 g24668 ( .a(n28458), .b(n28450), .c(n28449), .o(n28459) );
in01f01 g24669 ( .a(n28459), .o(n28460) );
no02f01 g24670 ( .a(n28044), .b(n28043), .o(n28461) );
in01f01 g24671 ( .a(n28461), .o(n28462) );
ao12f01 g24672 ( .a(n28054), .b(n28036), .c(n27682), .o(n28463) );
in01f01 g24673 ( .a(n28463), .o(n28464) );
oa12f01 g24674 ( .a(n28462), .b(n28464), .c(n28037), .o(n28465) );
in01f01 g24675 ( .a(n28465), .o(n28466) );
no03f01 g24676 ( .a(n28464), .b(n28462), .c(n28037), .o(n28467) );
in01f01 g24677 ( .a(n28282), .o(n28468) );
no02f01 g24678 ( .a(n28284), .b(n28211), .o(n28469) );
in01f01 g24679 ( .a(n28469), .o(n28470) );
no03f01 g24680 ( .a(n28470), .b(n28468), .c(n28221), .o(n28471) );
ao12f01 g24681 ( .a(n28469), .b(n28282), .c(n28222), .o(n28472) );
no02f01 g24682 ( .a(n28472), .b(n28471), .o(n28473) );
in01f01 g24683 ( .a(n28473), .o(n28474) );
no03f01 g24684 ( .a(n28474), .b(n28467), .c(n28466), .o(n28475) );
in01f01 g24685 ( .a(n28475), .o(n28476) );
in01f01 g24686 ( .a(n28036), .o(n28477) );
na02f01 g24687 ( .a(n28477), .b(n28027), .o(n28478) );
no02f01 g24688 ( .a(n28477), .b(n28027), .o(n28479) );
in01f01 g24689 ( .a(n28479), .o(n28480) );
no02f01 g24690 ( .a(n28280), .b(n28221), .o(n28481) );
in01f01 g24691 ( .a(n28481), .o(n28482) );
no03f01 g24692 ( .a(n28482), .b(n28279), .c(n28229), .o(n28483) );
no02f01 g24693 ( .a(n28279), .b(n28229), .o(n28484) );
no02f01 g24694 ( .a(n28481), .b(n28484), .o(n28485) );
no02f01 g24695 ( .a(n28485), .b(n28483), .o(n28486) );
ao12f01 g24696 ( .a(n28486), .b(n28480), .c(n28478), .o(n28487) );
in01f01 g24697 ( .a(n28487), .o(n28488) );
in01f01 g24698 ( .a(n27975), .o(n28489) );
oa12f01 g24699 ( .a(n_25834), .b(n28489), .c(n27973), .o(n28490) );
in01f01 g24700 ( .a(n27982), .o(n28491) );
na02f01 g24701 ( .a(n28491), .b(n27980), .o(n28492) );
na02f01 g24702 ( .a(n28492), .b(n_25834), .o(n28493) );
na02f01 g24703 ( .a(n28493), .b(n28490), .o(n28494) );
in01f01 g24704 ( .a(n27994), .o(n28495) );
no02f01 g24705 ( .a(n28495), .b(n27992), .o(n28496) );
no02f01 g24706 ( .a(n28496), .b(n27682), .o(n28497) );
in01f01 g24707 ( .a(n28004), .o(n28498) );
no03f01 g24708 ( .a(n28498), .b(n28497), .c(n28494), .o(n28499) );
no02f01 g24709 ( .a(n28018), .b(n28499), .o(n28500) );
in01f01 g24710 ( .a(n28500), .o(n28501) );
no02f01 g24711 ( .a(n28053), .b(n28005), .o(n28502) );
in01f01 g24712 ( .a(n28502), .o(n28503) );
no02f01 g24713 ( .a(n28272), .b(n28244), .o(n28504) );
no02f01 g24714 ( .a(n28275), .b(n28237), .o(n28505) );
in01f01 g24715 ( .a(n28505), .o(n28506) );
no02f01 g24716 ( .a(n28506), .b(n28504), .o(n28507) );
na02f01 g24717 ( .a(n28506), .b(n28504), .o(n28508) );
in01f01 g24718 ( .a(n28508), .o(n28509) );
no02f01 g24719 ( .a(n28509), .b(n28507), .o(n28510) );
ao12f01 g24720 ( .a(n28510), .b(n28503), .c(n28501), .o(n28511) );
in01f01 g24721 ( .a(n28511), .o(n28512) );
in01f01 g24722 ( .a(n28003), .o(n28513) );
oa12f01 g24723 ( .a(n28513), .b(n28497), .c(n28494), .o(n28514) );
na03f01 g24724 ( .a(n28003), .b(n27996), .c(n27985), .o(n28515) );
no02f01 g24725 ( .a(n28271), .b(n28244), .o(n28516) );
in01f01 g24726 ( .a(n28516), .o(n28517) );
no02f01 g24727 ( .a(n28517), .b(n28269), .o(n28518) );
na02f01 g24728 ( .a(n28517), .b(n28269), .o(n28519) );
in01f01 g24729 ( .a(n28519), .o(n28520) );
no02f01 g24730 ( .a(n28520), .b(n28518), .o(n28521) );
ao12f01 g24731 ( .a(n28521), .b(n28515), .c(n28514), .o(n28522) );
oa12f01 g24732 ( .a(n28496), .b(n27984), .c(n27976), .o(n28523) );
na03f01 g24733 ( .a(n27995), .b(n28493), .c(n28490), .o(n28524) );
na02f01 g24734 ( .a(n28524), .b(n28523), .o(n28525) );
in01f01 g24735 ( .a(n28268), .o(n28526) );
no02f01 g24736 ( .a(n28526), .b(n28255), .o(n28527) );
no02f01 g24737 ( .a(n28527), .b(n28267), .o(n28528) );
na02f01 g24738 ( .a(n28527), .b(n28267), .o(n28529) );
in01f01 g24739 ( .a(n28529), .o(n28530) );
no02f01 g24740 ( .a(n28530), .b(n28528), .o(n28531) );
in01f01 g24741 ( .a(n28531), .o(n28532) );
na02f01 g24742 ( .a(n28532), .b(n28525), .o(n28533) );
na02f01 g24743 ( .a(n27975), .b(n27974), .o(n28534) );
no03f01 g24744 ( .a(n28258), .b(n28257), .c(delay_add_ln22_unr17_stage7_stallmux_q_0_), .o(n28535) );
in01f01 g24745 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_0_), .o(n28536) );
no02f01 g24746 ( .a(n28259), .b(n28536), .o(n28537) );
no02f01 g24747 ( .a(n28537), .b(n28535), .o(n28538) );
in01f01 g24748 ( .a(n28538), .o(n28539) );
na02f01 g24749 ( .a(n28539), .b(n28534), .o(n28540) );
in01f01 g24750 ( .a(n28260), .o(n28541) );
no02f01 g24751 ( .a(n28265), .b(delay_add_ln22_unr17_stage7_stallmux_q_1_), .o(n28542) );
na02f01 g24752 ( .a(n28265), .b(delay_add_ln22_unr17_stage7_stallmux_q_1_), .o(n28543) );
in01f01 g24753 ( .a(n28543), .o(n28544) );
no03f01 g24754 ( .a(n28544), .b(n28542), .c(n28541), .o(n28545) );
in01f01 g24755 ( .a(n28542), .o(n28546) );
ao12f01 g24756 ( .a(n28260), .b(n28543), .c(n28546), .o(n28547) );
no02f01 g24757 ( .a(n28547), .b(n28545), .o(n28548) );
no02f01 g24758 ( .a(n28548), .b(n28540), .o(n28549) );
na02f01 g24759 ( .a(n28492), .b(n28490), .o(n28550) );
na02f01 g24760 ( .a(n27983), .b(n27976), .o(n28551) );
ao22f01 g24761 ( .a(n28551), .b(n28550), .c(n28548), .d(n28540), .o(n28552) );
oa22f01 g24762 ( .a(n28552), .b(n28549), .c(n28532), .d(n28525), .o(n28553) );
ao12f01 g24763 ( .a(n28003), .b(n27996), .c(n27985), .o(n28554) );
in01f01 g24764 ( .a(n28515), .o(n28555) );
in01f01 g24765 ( .a(n28521), .o(n28556) );
no03f01 g24766 ( .a(n28556), .b(n28555), .c(n28554), .o(n28557) );
ao12f01 g24767 ( .a(n28557), .b(n28553), .c(n28533), .o(n28558) );
in01f01 g24768 ( .a(n28510), .o(n28559) );
no03f01 g24769 ( .a(n28559), .b(n28502), .c(n28500), .o(n28560) );
in01f01 g24770 ( .a(n28560), .o(n28561) );
oa12f01 g24771 ( .a(n28561), .b(n28558), .c(n28522), .o(n28562) );
oa12f01 g24772 ( .a(n28499), .b(n28053), .c(n27682), .o(n28563) );
na02f01 g24773 ( .a(n28026), .b(n28563), .o(n28564) );
in01f01 g24774 ( .a(n28026), .o(n28565) );
na02f01 g24775 ( .a(n28565), .b(n28019), .o(n28566) );
na02f01 g24776 ( .a(n28566), .b(n28564), .o(n28567) );
no02f01 g24777 ( .a(n28278), .b(n28229), .o(n28568) );
no02f01 g24778 ( .a(n28568), .b(n28276), .o(n28569) );
na02f01 g24779 ( .a(n28568), .b(n28276), .o(n28570) );
in01f01 g24780 ( .a(n28570), .o(n28571) );
no02f01 g24781 ( .a(n28571), .b(n28569), .o(n28572) );
in01f01 g24782 ( .a(n28572), .o(n28573) );
na02f01 g24783 ( .a(n28573), .b(n28567), .o(n28574) );
na03f01 g24784 ( .a(n28574), .b(n28562), .c(n28512), .o(n28575) );
no02f01 g24785 ( .a(n28573), .b(n28567), .o(n28576) );
in01f01 g24786 ( .a(n28576), .o(n28577) );
na03f01 g24787 ( .a(n28486), .b(n28480), .c(n28478), .o(n28578) );
na03f01 g24788 ( .a(n28578), .b(n28577), .c(n28575), .o(n28579) );
oa12f01 g24789 ( .a(n28474), .b(n28467), .c(n28466), .o(n28580) );
na03f01 g24790 ( .a(n28580), .b(n28579), .c(n28488), .o(n28581) );
na03f01 g24791 ( .a(n28458), .b(n28450), .c(n28449), .o(n28582) );
na03f01 g24792 ( .a(n28582), .b(n28581), .c(n28476), .o(n28583) );
na03f01 g24793 ( .a(n28583), .b(n28460), .c(n28446), .o(n28584) );
no03f01 g24794 ( .a(n28445), .b(n28438), .c(n28435), .o(n28585) );
in01f01 g24795 ( .a(n28585), .o(n28586) );
no02f01 g24796 ( .a(n28095), .b(n28073), .o(n28587) );
in01f01 g24797 ( .a(n28587), .o(n28588) );
no02f01 g24798 ( .a(n28588), .b(n28091), .o(n28589) );
no02f01 g24799 ( .a(n28587), .b(n28092), .o(n28590) );
no02f01 g24800 ( .a(n28293), .b(n28183), .o(n28591) );
in01f01 g24801 ( .a(n28591), .o(n28592) );
no03f01 g24802 ( .a(n28592), .b(n28292), .c(n28191), .o(n28593) );
no02f01 g24803 ( .a(n28292), .b(n28191), .o(n28594) );
no02f01 g24804 ( .a(n28591), .b(n28594), .o(n28595) );
no02f01 g24805 ( .a(n28595), .b(n28593), .o(n28596) );
in01f01 g24806 ( .a(n28596), .o(n28597) );
no03f01 g24807 ( .a(n28597), .b(n28590), .c(n28589), .o(n28598) );
in01f01 g24808 ( .a(n28598), .o(n28599) );
na03f01 g24809 ( .a(n28599), .b(n28586), .c(n28584), .o(n28600) );
no02f01 g24810 ( .a(n28419), .b(n28418), .o(n28601) );
no02f01 g24811 ( .a(n28425), .b(n28601), .o(n28602) );
oa12f01 g24812 ( .a(n28597), .b(n28590), .c(n28589), .o(n28603) );
in01f01 g24813 ( .a(n28603), .o(n28604) );
no02f01 g24814 ( .a(n28604), .b(n28602), .o(n28605) );
na02f01 g24815 ( .a(n28605), .b(n28600), .o(n28606) );
no02f01 g24816 ( .a(n28399), .b(n28390), .o(n28607) );
in01f01 g24817 ( .a(n28607), .o(n28608) );
na04f01 g24818 ( .a(n28608), .b(n28606), .c(n28428), .d(n28413), .o(n28609) );
no02f01 g24819 ( .a(n28304), .b(n28154), .o(n28610) );
no02f01 g24820 ( .a(n28143), .b(n28305), .o(n28611) );
in01f01 g24821 ( .a(n28611), .o(n28612) );
ao12f01 g24822 ( .a(n28310), .b(n28612), .c(n28610), .o(n28613) );
no02f01 g24823 ( .a(n28143), .b(n28306), .o(n28614) );
no02f01 g24824 ( .a(n28614), .b(n28309), .o(n28615) );
in01f01 g24825 ( .a(n28615), .o(n28616) );
no02f01 g24826 ( .a(n28616), .b(n28613), .o(n28617) );
na02f01 g24827 ( .a(n28616), .b(n28613), .o(n28618) );
in01f01 g24828 ( .a(n28618), .o(n28619) );
no02f01 g24829 ( .a(n28619), .b(n28617), .o(n28620) );
no02f01 g24830 ( .a(n28310), .b(n28611), .o(n28621) );
no02f01 g24831 ( .a(n28621), .b(n28610), .o(n28622) );
na02f01 g24832 ( .a(n28621), .b(n28610), .o(n28623) );
in01f01 g24833 ( .a(n28623), .o(n28624) );
no02f01 g24834 ( .a(n28624), .b(n28622), .o(n28625) );
ao12f01 g24835 ( .a(n28383), .b(n28625), .c(n28620), .o(n28626) );
in01f01 g24836 ( .a(n28626), .o(n28627) );
na03f01 g24837 ( .a(n28627), .b(n28609), .c(n28412), .o(n28628) );
in01f01 g24838 ( .a(n28620), .o(n28629) );
no02f01 g24839 ( .a(n28629), .b(n28102), .o(n28630) );
in01f01 g24840 ( .a(n28625), .o(n28631) );
no02f01 g24841 ( .a(n28631), .b(n28102), .o(n28632) );
no02f01 g24842 ( .a(n28632), .b(n28630), .o(n28633) );
no02f01 g24843 ( .a(n28345), .b(n28320), .o(n28634) );
in01f01 g24844 ( .a(n28634), .o(n28635) );
no03f01 g24845 ( .a(n28319), .b(n28312), .c(n28308), .o(n28636) );
no03f01 g24846 ( .a(n28636), .b(n28635), .c(n28343), .o(n28637) );
in01f01 g24847 ( .a(n28637), .o(n28638) );
oa12f01 g24848 ( .a(n28635), .b(n28636), .c(n28343), .o(n28639) );
na02f01 g24849 ( .a(n28639), .b(n28638), .o(n28640) );
no02f01 g24850 ( .a(n28640), .b(n28102), .o(n28641) );
in01f01 g24851 ( .a(n28641), .o(n28642) );
no02f01 g24852 ( .a(n28312), .b(n28308), .o(n28643) );
no02f01 g24853 ( .a(n28143), .b(n28313), .o(n28644) );
no02f01 g24854 ( .a(n28144), .b(delay_add_ln22_unr17_stage7_stallmux_q_16_), .o(n28645) );
in01f01 g24855 ( .a(n28645), .o(n28646) );
ao12f01 g24856 ( .a(n28644), .b(n28646), .c(n28643), .o(n28647) );
in01f01 g24857 ( .a(n28647), .o(n28648) );
no02f01 g24858 ( .a(n28144), .b(delay_add_ln22_unr17_stage7_stallmux_q_17_), .o(n28649) );
no02f01 g24859 ( .a(n28143), .b(n28314), .o(n28650) );
no02f01 g24860 ( .a(n28650), .b(n28649), .o(n28651) );
in01f01 g24861 ( .a(n28651), .o(n28652) );
no02f01 g24862 ( .a(n28652), .b(n28648), .o(n28653) );
no02f01 g24863 ( .a(n28651), .b(n28647), .o(n28654) );
no02f01 g24864 ( .a(n28654), .b(n28653), .o(n28655) );
in01f01 g24865 ( .a(n28655), .o(n28656) );
in01f01 g24866 ( .a(n28643), .o(n28657) );
no02f01 g24867 ( .a(n28645), .b(n28644), .o(n28658) );
no02f01 g24868 ( .a(n28658), .b(n28657), .o(n28659) );
na02f01 g24869 ( .a(n28658), .b(n28657), .o(n28660) );
in01f01 g24870 ( .a(n28660), .o(n28661) );
no02f01 g24871 ( .a(n28661), .b(n28659), .o(n28662) );
in01f01 g24872 ( .a(n28662), .o(n28663) );
ao12f01 g24873 ( .a(n28102), .b(n28663), .c(n28656), .o(n28664) );
in01f01 g24874 ( .a(n28664), .o(n28665) );
in01f01 g24875 ( .a(n28316), .o(n28666) );
ao12f01 g24876 ( .a(n28339), .b(n28666), .c(n28643), .o(n28667) );
in01f01 g24877 ( .a(n28667), .o(n28668) );
no02f01 g24878 ( .a(n28341), .b(n28317), .o(n28669) );
in01f01 g24879 ( .a(n28669), .o(n28670) );
no02f01 g24880 ( .a(n28670), .b(n28668), .o(n28671) );
no02f01 g24881 ( .a(n28669), .b(n28667), .o(n28672) );
no02f01 g24882 ( .a(n28672), .b(n28671), .o(n28673) );
in01f01 g24883 ( .a(n28673), .o(n28674) );
no02f01 g24884 ( .a(n28674), .b(n28102), .o(n28675) );
in01f01 g24885 ( .a(n28675), .o(n28676) );
na04f01 g24886 ( .a(n28676), .b(n28665), .c(n28642), .d(n28633), .o(n28677) );
in01f01 g24887 ( .a(n28677), .o(n28678) );
ao12f01 g24888 ( .a(n28383), .b(n28662), .c(n28655), .o(n28679) );
in01f01 g24889 ( .a(n28639), .o(n28680) );
no02f01 g24890 ( .a(n28680), .b(n28637), .o(n28681) );
ao12f01 g24891 ( .a(n28383), .b(n28673), .c(n28681), .o(n28682) );
no02f01 g24892 ( .a(n28682), .b(n28679), .o(n28683) );
in01f01 g24893 ( .a(n28683), .o(n28684) );
ao12f01 g24894 ( .a(n28684), .b(n28678), .c(n28628), .o(n28685) );
no02f01 g24895 ( .a(n28320), .b(n28319), .o(n28686) );
na02f01 g24896 ( .a(n28686), .b(n28643), .o(n28687) );
no02f01 g24897 ( .a(n28143), .b(n28349), .o(n28688) );
no02f01 g24898 ( .a(n28688), .b(n28322), .o(n28689) );
na03f01 g24899 ( .a(n28689), .b(n28346), .c(n28687), .o(n28690) );
in01f01 g24900 ( .a(n28689), .o(n28691) );
oa12f01 g24901 ( .a(n28691), .b(n28347), .c(n28321), .o(n28692) );
na02f01 g24902 ( .a(n28692), .b(n28690), .o(n28693) );
no02f01 g24903 ( .a(n28693), .b(n28102), .o(n28694) );
no02f01 g24904 ( .a(n28688), .b(n28347), .o(n28695) );
no02f01 g24905 ( .a(n28143), .b(n28348), .o(n28696) );
no02f01 g24906 ( .a(n28696), .b(n28325), .o(n28697) );
na03f01 g24907 ( .a(n28697), .b(n28695), .c(n28324), .o(n28698) );
ao12f01 g24908 ( .a(n28697), .b(n28695), .c(n28324), .o(n28699) );
in01f01 g24909 ( .a(n28699), .o(n28700) );
na02f01 g24910 ( .a(n28700), .b(n28698), .o(n28701) );
no02f01 g24911 ( .a(n28701), .b(n28102), .o(n28702) );
no03f01 g24912 ( .a(n28702), .b(n28694), .c(n28685), .o(n28703) );
no02f01 g24913 ( .a(n28143), .b(n28354), .o(n28704) );
no02f01 g24914 ( .a(n28704), .b(n28146), .o(n28705) );
in01f01 g24915 ( .a(n28705), .o(n28706) );
no02f01 g24916 ( .a(n28143), .b(n28353), .o(n28707) );
no02f01 g24917 ( .a(n28707), .b(n28352), .o(n28708) );
na02f01 g24918 ( .a(n28708), .b(n28329), .o(n28709) );
na02f01 g24919 ( .a(n28709), .b(n28706), .o(n28710) );
no02f01 g24920 ( .a(n28709), .b(n28706), .o(n28711) );
in01f01 g24921 ( .a(n28711), .o(n28712) );
na02f01 g24922 ( .a(n28712), .b(n28710), .o(n28713) );
no02f01 g24923 ( .a(n28713), .b(n28102), .o(n28714) );
no02f01 g24924 ( .a(n28707), .b(n28327), .o(n28715) );
no02f01 g24925 ( .a(n28352), .b(n28326), .o(n28716) );
na02f01 g24926 ( .a(n28716), .b(n28715), .o(n28717) );
in01f01 g24927 ( .a(n28715), .o(n28718) );
no02f01 g24928 ( .a(n28322), .b(n28687), .o(n28719) );
in01f01 g24929 ( .a(n28325), .o(n28720) );
na02f01 g24930 ( .a(n28720), .b(n28719), .o(n28721) );
na02f01 g24931 ( .a(n28351), .b(n28721), .o(n28722) );
na02f01 g24932 ( .a(n28722), .b(n28718), .o(n28723) );
na02f01 g24933 ( .a(n28723), .b(n28717), .o(n28724) );
no02f01 g24934 ( .a(n28724), .b(n28102), .o(n28725) );
no02f01 g24935 ( .a(n28725), .b(n28714), .o(n28726) );
no03f01 g24936 ( .a(n28691), .b(n28347), .c(n28321), .o(n28727) );
ao12f01 g24937 ( .a(n28689), .b(n28346), .c(n28687), .o(n28728) );
no02f01 g24938 ( .a(n28728), .b(n28727), .o(n28729) );
in01f01 g24939 ( .a(n28698), .o(n28730) );
no02f01 g24940 ( .a(n28699), .b(n28730), .o(n28731) );
ao12f01 g24941 ( .a(n28383), .b(n28731), .c(n28729), .o(n28732) );
in01f01 g24942 ( .a(n28710), .o(n28733) );
no02f01 g24943 ( .a(n28711), .b(n28733), .o(n28734) );
no02f01 g24944 ( .a(n28722), .b(n28718), .o(n28735) );
no02f01 g24945 ( .a(n28716), .b(n28715), .o(n28736) );
no02f01 g24946 ( .a(n28736), .b(n28735), .o(n28737) );
ao12f01 g24947 ( .a(n28383), .b(n28737), .c(n28734), .o(n28738) );
no02f01 g24948 ( .a(n28738), .b(n28732), .o(n28739) );
in01f01 g24949 ( .a(n28739), .o(n28740) );
ao12f01 g24950 ( .a(n28740), .b(n28726), .c(n28703), .o(n28741) );
in01f01 g24951 ( .a(n28146), .o(n28742) );
no02f01 g24952 ( .a(n28327), .b(n28721), .o(n28743) );
na02f01 g24953 ( .a(n28743), .b(n28742), .o(n28744) );
na02f01 g24954 ( .a(n28356), .b(n28744), .o(n28745) );
no02f01 g24955 ( .a(n28143), .b(n28357), .o(n28746) );
no02f01 g24956 ( .a(n28746), .b(n28331), .o(n28747) );
in01f01 g24957 ( .a(n28747), .o(n28748) );
na02f01 g24958 ( .a(n28748), .b(n28745), .o(n28749) );
in01f01 g24959 ( .a(n28356), .o(n28750) );
no02f01 g24960 ( .a(n28750), .b(n28330), .o(n28751) );
na02f01 g24961 ( .a(n28747), .b(n28751), .o(n28752) );
na02f01 g24962 ( .a(n28752), .b(n28749), .o(n28753) );
no02f01 g24963 ( .a(n28753), .b(n28102), .o(n28754) );
no02f01 g24964 ( .a(n28746), .b(n28750), .o(n28755) );
na02f01 g24965 ( .a(n28755), .b(n28333), .o(n28756) );
no02f01 g24966 ( .a(n28143), .b(n28358), .o(n28757) );
no02f01 g24967 ( .a(n28757), .b(n28334), .o(n28758) );
in01f01 g24968 ( .a(n28758), .o(n28759) );
na02f01 g24969 ( .a(n28759), .b(n28756), .o(n28760) );
no02f01 g24970 ( .a(n28759), .b(n28756), .o(n28761) );
in01f01 g24971 ( .a(n28761), .o(n28762) );
na02f01 g24972 ( .a(n28762), .b(n28760), .o(n28763) );
no02f01 g24973 ( .a(n28763), .b(n28102), .o(n28764) );
no02f01 g24974 ( .a(n28764), .b(n28754), .o(n28765) );
in01f01 g24975 ( .a(n28765), .o(n28766) );
no02f01 g24976 ( .a(n28766), .b(n28741), .o(n28767) );
no02f01 g24977 ( .a(n28361), .b(n28336), .o(n28768) );
in01f01 g24978 ( .a(n28337), .o(n28769) );
no02f01 g24979 ( .a(n28359), .b(n28750), .o(n28770) );
oa12f01 g24980 ( .a(n28770), .b(n28334), .c(n28333), .o(n28771) );
oa12f01 g24981 ( .a(n28769), .b(n28771), .c(n28363), .o(n28772) );
na02f01 g24982 ( .a(n28772), .b(n28768), .o(n28773) );
no02f01 g24983 ( .a(n28772), .b(n28768), .o(n28774) );
in01f01 g24984 ( .a(n28774), .o(n28775) );
na02f01 g24985 ( .a(n28775), .b(n28773), .o(n28776) );
no02f01 g24986 ( .a(n28776), .b(n28102), .o(n28777) );
in01f01 g24987 ( .a(n28771), .o(n28778) );
no02f01 g24988 ( .a(n28363), .b(n28337), .o(n28779) );
no02f01 g24989 ( .a(n28779), .b(n28778), .o(n28780) );
in01f01 g24990 ( .a(n28780), .o(n28781) );
na02f01 g24991 ( .a(n28779), .b(n28778), .o(n28782) );
na02f01 g24992 ( .a(n28782), .b(n28781), .o(n28783) );
no02f01 g24993 ( .a(n28783), .b(n28102), .o(n28784) );
no02f01 g24994 ( .a(n28784), .b(n28777), .o(n28785) );
no02f01 g24995 ( .a(n28747), .b(n28751), .o(n28786) );
no02f01 g24996 ( .a(n28748), .b(n28745), .o(n28787) );
no02f01 g24997 ( .a(n28787), .b(n28786), .o(n28788) );
in01f01 g24998 ( .a(n28760), .o(n28789) );
no02f01 g24999 ( .a(n28761), .b(n28789), .o(n28790) );
ao12f01 g25000 ( .a(n28383), .b(n28790), .c(n28788), .o(n28791) );
in01f01 g25001 ( .a(n28773), .o(n28792) );
no02f01 g25002 ( .a(n28774), .b(n28792), .o(n28793) );
in01f01 g25003 ( .a(n28782), .o(n28794) );
no02f01 g25004 ( .a(n28794), .b(n28780), .o(n28795) );
ao12f01 g25005 ( .a(n28383), .b(n28795), .c(n28793), .o(n28796) );
no02f01 g25006 ( .a(n28796), .b(n28791), .o(n28797) );
in01f01 g25007 ( .a(n28797), .o(n28798) );
ao12f01 g25008 ( .a(n28798), .b(n28785), .c(n28767), .o(n28799) );
in01f01 g25009 ( .a(n28366), .o(n28800) );
no02f01 g25010 ( .a(n28143), .b(n28368), .o(n28801) );
no02f01 g25011 ( .a(n28144), .b(delay_add_ln22_unr17_stage7_stallmux_q_28_), .o(n28802) );
no02f01 g25012 ( .a(n28802), .b(n28801), .o(n28803) );
in01f01 g25013 ( .a(n28803), .o(n28804) );
no02f01 g25014 ( .a(n28804), .b(n28800), .o(n28805) );
no02f01 g25015 ( .a(n28803), .b(n28366), .o(n28806) );
no02f01 g25016 ( .a(n28806), .b(n28805), .o(n28807) );
in01f01 g25017 ( .a(n28807), .o(n28808) );
no02f01 g25018 ( .a(n28808), .b(n28102), .o(n28809) );
no02f01 g25019 ( .a(n28809), .b(n28799), .o(n28810) );
in01f01 g25020 ( .a(n28810), .o(n28811) );
no02f01 g25021 ( .a(n28144), .b(delay_add_ln22_unr17_stage7_stallmux_q_29_), .o(n28812) );
no02f01 g25022 ( .a(n28143), .b(n28367), .o(n28813) );
no02f01 g25023 ( .a(n28813), .b(n28812), .o(n28814) );
in01f01 g25024 ( .a(n28814), .o(n28815) );
no02f01 g25025 ( .a(n28802), .b(n28366), .o(n28816) );
no02f01 g25026 ( .a(n28816), .b(n28801), .o(n28817) );
in01f01 g25027 ( .a(n28817), .o(n28818) );
no02f01 g25028 ( .a(n28818), .b(n28815), .o(n28819) );
no02f01 g25029 ( .a(n28817), .b(n28814), .o(n28820) );
no02f01 g25030 ( .a(n28820), .b(n28819), .o(n28821) );
in01f01 g25031 ( .a(n28821), .o(n28822) );
no02f01 g25032 ( .a(n28822), .b(n28102), .o(n28823) );
no02f01 g25033 ( .a(n28823), .b(n28811), .o(n28824) );
no02f01 g25034 ( .a(n28807), .b(n28383), .o(n28825) );
no02f01 g25035 ( .a(n28821), .b(n28383), .o(n28826) );
no02f01 g25036 ( .a(n28826), .b(n28825), .o(n28827) );
in01f01 g25037 ( .a(n28827), .o(n28828) );
no02f01 g25038 ( .a(n28828), .b(n28824), .o(n28829) );
no02f01 g25039 ( .a(n28829), .b(n28385), .o(n28830) );
na02f01 g25040 ( .a(n28829), .b(n28385), .o(n28831) );
in01f01 g25041 ( .a(n28831), .o(n28832) );
no02f01 g25042 ( .a(n28832), .b(n28830), .o(n28833) );
no02f01 g25043 ( .a(n28833), .b(n27681), .o(n28834) );
oa12f01 g25044 ( .a(n28436), .b(n28433), .c(n28437), .o(n28835) );
na03f01 g25045 ( .a(n28434), .b(n28432), .c(n28071), .o(n28836) );
ao12f01 g25046 ( .a(n28444), .b(n28836), .c(n28835), .o(n28837) );
in01f01 g25047 ( .a(n28522), .o(n28838) );
ao12f01 g25048 ( .a(n27995), .b(n28493), .c(n28490), .o(n28839) );
no03f01 g25049 ( .a(n28496), .b(n27984), .c(n27976), .o(n28840) );
no02f01 g25050 ( .a(n28840), .b(n28839), .o(n28841) );
no02f01 g25051 ( .a(n28531), .b(n28841), .o(n28842) );
in01f01 g25052 ( .a(n28549), .o(n28843) );
no02f01 g25053 ( .a(n28489), .b(n27973), .o(n28844) );
no02f01 g25054 ( .a(n28538), .b(n28844), .o(n28845) );
in01f01 g25055 ( .a(n28548), .o(n28846) );
no02f01 g25056 ( .a(n27983), .b(n27976), .o(n28847) );
no02f01 g25057 ( .a(n28492), .b(n28490), .o(n28848) );
oa22f01 g25058 ( .a(n28848), .b(n28847), .c(n28846), .d(n28845), .o(n28849) );
ao22f01 g25059 ( .a(n28849), .b(n28843), .c(n28531), .d(n28841), .o(n28850) );
na03f01 g25060 ( .a(n28521), .b(n28515), .c(n28514), .o(n28851) );
oa12f01 g25061 ( .a(n28851), .b(n28850), .c(n28842), .o(n28852) );
ao12f01 g25062 ( .a(n28560), .b(n28852), .c(n28838), .o(n28853) );
no02f01 g25063 ( .a(n28565), .b(n28019), .o(n28854) );
no02f01 g25064 ( .a(n28026), .b(n28563), .o(n28855) );
no02f01 g25065 ( .a(n28855), .b(n28854), .o(n28856) );
no02f01 g25066 ( .a(n28572), .b(n28856), .o(n28857) );
no03f01 g25067 ( .a(n28857), .b(n28853), .c(n28511), .o(n28858) );
in01f01 g25068 ( .a(n28478), .o(n28859) );
in01f01 g25069 ( .a(n28486), .o(n28860) );
no03f01 g25070 ( .a(n28860), .b(n28479), .c(n28859), .o(n28861) );
no03f01 g25071 ( .a(n28861), .b(n28576), .c(n28858), .o(n28862) );
in01f01 g25072 ( .a(n28467), .o(n28863) );
ao12f01 g25073 ( .a(n28473), .b(n28863), .c(n28465), .o(n28864) );
no03f01 g25074 ( .a(n28864), .b(n28862), .c(n28487), .o(n28865) );
in01f01 g25075 ( .a(n28447), .o(n28866) );
no02f01 g25076 ( .a(n28866), .b(n28429), .o(n28867) );
in01f01 g25077 ( .a(n28458), .o(n28868) );
no03f01 g25078 ( .a(n28868), .b(n28867), .c(n28448), .o(n28869) );
no03f01 g25079 ( .a(n28869), .b(n28865), .c(n28475), .o(n28870) );
no03f01 g25080 ( .a(n28870), .b(n28459), .c(n28837), .o(n28871) );
no03f01 g25081 ( .a(n28598), .b(n28585), .c(n28871), .o(n28872) );
oa12f01 g25082 ( .a(n28603), .b(n28425), .c(n28601), .o(n28873) );
no02f01 g25083 ( .a(n28873), .b(n28872), .o(n28874) );
no04f01 g25084 ( .a(n28607), .b(n28874), .c(n28427), .d(n28410), .o(n28875) );
no03f01 g25085 ( .a(n28626), .b(n28875), .c(n28411), .o(n28876) );
oa12f01 g25086 ( .a(n28683), .b(n28677), .c(n28876), .o(n28877) );
in01f01 g25087 ( .a(n28694), .o(n28878) );
no02f01 g25088 ( .a(n28729), .b(n28383), .o(n28879) );
ao12f01 g25089 ( .a(n28879), .b(n28878), .c(n28877), .o(n28880) );
no02f01 g25090 ( .a(n28731), .b(n28383), .o(n28881) );
no02f01 g25091 ( .a(n28881), .b(n28702), .o(n28882) );
no02f01 g25092 ( .a(n28882), .b(n28880), .o(n28883) );
in01f01 g25093 ( .a(n28879), .o(n28884) );
oa12f01 g25094 ( .a(n28884), .b(n28694), .c(n28685), .o(n28885) );
in01f01 g25095 ( .a(n28882), .o(n28886) );
no02f01 g25096 ( .a(n28886), .b(n28885), .o(n28887) );
no02f01 g25097 ( .a(n28887), .b(n28883), .o(n28888) );
no02f01 g25098 ( .a(n28879), .b(n28694), .o(n28889) );
in01f01 g25099 ( .a(n28889), .o(n28890) );
no02f01 g25100 ( .a(n28890), .b(n28877), .o(n28891) );
no02f01 g25101 ( .a(n28889), .b(n28685), .o(n28892) );
no02f01 g25102 ( .a(n28892), .b(n28891), .o(n28893) );
ao12f01 g25103 ( .a(n27681), .b(n28893), .c(n28888), .o(n28894) );
in01f01 g25104 ( .a(n28702), .o(n28895) );
na03f01 g25105 ( .a(n28895), .b(n28878), .c(n28877), .o(n28896) );
in01f01 g25106 ( .a(n28732), .o(n28897) );
no02f01 g25107 ( .a(n28737), .b(n28383), .o(n28898) );
no02f01 g25108 ( .a(n28898), .b(n28725), .o(n28899) );
ao12f01 g25109 ( .a(n28899), .b(n28897), .c(n28896), .o(n28900) );
in01f01 g25110 ( .a(n28899), .o(n28901) );
no03f01 g25111 ( .a(n28901), .b(n28732), .c(n28703), .o(n28902) );
oa12f01 g25112 ( .a(n_27014), .b(n28902), .c(n28900), .o(n28903) );
in01f01 g25113 ( .a(n28903), .o(n28904) );
no02f01 g25114 ( .a(n28904), .b(n28894), .o(n28905) );
no03f01 g25115 ( .a(n28898), .b(n28732), .c(n28703), .o(n28906) );
no02f01 g25116 ( .a(n28734), .b(n28383), .o(n28907) );
no02f01 g25117 ( .a(n28907), .b(n28714), .o(n28908) );
no03f01 g25118 ( .a(n28908), .b(n28906), .c(n28725), .o(n28909) );
in01f01 g25119 ( .a(n28725), .o(n28910) );
in01f01 g25120 ( .a(n28898), .o(n28911) );
na03f01 g25121 ( .a(n28911), .b(n28897), .c(n28896), .o(n28912) );
in01f01 g25122 ( .a(n28908), .o(n28913) );
ao12f01 g25123 ( .a(n28913), .b(n28912), .c(n28910), .o(n28914) );
oa12f01 g25124 ( .a(n_27014), .b(n28914), .c(n28909), .o(n28915) );
oa12f01 g25125 ( .a(n27681), .b(n28914), .c(n28909), .o(n28916) );
in01f01 g25126 ( .a(n28916), .o(n28917) );
ao12f01 g25127 ( .a(n28917), .b(n28915), .c(n28905), .o(n28918) );
no02f01 g25128 ( .a(n28788), .b(n28383), .o(n28919) );
no02f01 g25129 ( .a(n28919), .b(n28754), .o(n28920) );
no02f01 g25130 ( .a(n28920), .b(n28741), .o(n28921) );
na02f01 g25131 ( .a(n28920), .b(n28741), .o(n28922) );
in01f01 g25132 ( .a(n28922), .o(n28923) );
no02f01 g25133 ( .a(n28923), .b(n28921), .o(n28924) );
no02f01 g25134 ( .a(n28924), .b(n27681), .o(n28925) );
no02f01 g25135 ( .a(n28925), .b(n28918), .o(n28926) );
no02f01 g25136 ( .a(n28790), .b(n28383), .o(n28927) );
no02f01 g25137 ( .a(n28927), .b(n28764), .o(n28928) );
in01f01 g25138 ( .a(n28928), .o(n28929) );
no02f01 g25139 ( .a(n28754), .b(n28741), .o(n28930) );
no03f01 g25140 ( .a(n28930), .b(n28929), .c(n28919), .o(n28931) );
in01f01 g25141 ( .a(n28931), .o(n28932) );
oa12f01 g25142 ( .a(n28929), .b(n28930), .c(n28919), .o(n28933) );
na02f01 g25143 ( .a(n28933), .b(n28932), .o(n28934) );
na02f01 g25144 ( .a(n28934), .b(n_27014), .o(n28935) );
no02f01 g25145 ( .a(n28795), .b(n28383), .o(n28936) );
no02f01 g25146 ( .a(n28936), .b(n28784), .o(n28937) );
no02f01 g25147 ( .a(n28791), .b(n28767), .o(n28938) );
no02f01 g25148 ( .a(n28938), .b(n28937), .o(n28939) );
in01f01 g25149 ( .a(n28937), .o(n28940) );
in01f01 g25150 ( .a(n28791), .o(n28941) );
oa12f01 g25151 ( .a(n28941), .b(n28766), .c(n28741), .o(n28942) );
no02f01 g25152 ( .a(n28942), .b(n28940), .o(n28943) );
no02f01 g25153 ( .a(n28943), .b(n28939), .o(n28944) );
no02f01 g25154 ( .a(n28944), .b(n27681), .o(n28945) );
in01f01 g25155 ( .a(n28945), .o(n28946) );
na03f01 g25156 ( .a(n28946), .b(n28935), .c(n28926), .o(n28947) );
in01f01 g25157 ( .a(n28784), .o(n28948) );
no02f01 g25158 ( .a(n28793), .b(n28383), .o(n28949) );
no02f01 g25159 ( .a(n28949), .b(n28777), .o(n28950) );
in01f01 g25160 ( .a(n28950), .o(n28951) );
in01f01 g25161 ( .a(n28936), .o(n28952) );
na02f01 g25162 ( .a(n28938), .b(n28952), .o(n28953) );
ao12f01 g25163 ( .a(n28951), .b(n28953), .c(n28948), .o(n28954) );
no02f01 g25164 ( .a(n28942), .b(n28936), .o(n28955) );
no03f01 g25165 ( .a(n28955), .b(n28950), .c(n28784), .o(n28956) );
no03f01 g25166 ( .a(n28956), .b(n28954), .c(n27681), .o(n28957) );
oa12f01 g25167 ( .a(n28950), .b(n28955), .c(n28784), .o(n28958) );
na03f01 g25168 ( .a(n28953), .b(n28951), .c(n28948), .o(n28959) );
ao12f01 g25169 ( .a(n_27014), .b(n28959), .c(n28958), .o(n28960) );
no02f01 g25170 ( .a(n28944), .b(n_27014), .o(n28961) );
no03f01 g25171 ( .a(n28961), .b(n28960), .c(n28957), .o(n28962) );
ao12f01 g25172 ( .a(n_27014), .b(n28962), .c(n28947), .o(n28963) );
no02f01 g25173 ( .a(n28960), .b(n28957), .o(n28964) );
in01f01 g25174 ( .a(n28924), .o(n28965) );
oa12f01 g25175 ( .a(n27681), .b(n28934), .c(n28965), .o(n28966) );
oa12f01 g25176 ( .a(n28966), .b(n28964), .c(n28947), .o(n28967) );
in01f01 g25177 ( .a(n28799), .o(n28968) );
no02f01 g25178 ( .a(n28825), .b(n28809), .o(n28969) );
in01f01 g25179 ( .a(n28969), .o(n28970) );
no02f01 g25180 ( .a(n28970), .b(n28968), .o(n28971) );
no02f01 g25181 ( .a(n28969), .b(n28799), .o(n28972) );
no02f01 g25182 ( .a(n28972), .b(n28971), .o(n28973) );
no02f01 g25183 ( .a(n28973), .b(n27681), .o(n28974) );
in01f01 g25184 ( .a(n28974), .o(n28975) );
oa12f01 g25185 ( .a(n28975), .b(n28967), .c(n28963), .o(n28976) );
no02f01 g25186 ( .a(n28825), .b(n28810), .o(n28977) );
no02f01 g25187 ( .a(n28826), .b(n28823), .o(n28978) );
no02f01 g25188 ( .a(n28978), .b(n28977), .o(n28979) );
na02f01 g25189 ( .a(n28978), .b(n28977), .o(n28980) );
in01f01 g25190 ( .a(n28980), .o(n28981) );
no02f01 g25191 ( .a(n28981), .b(n28979), .o(n28982) );
no02f01 g25192 ( .a(n28982), .b(n27681), .o(n28983) );
no03f01 g25193 ( .a(n28983), .b(n28976), .c(n28834), .o(n28984) );
ao12f01 g25194 ( .a(n_27014), .b(n28982), .c(n28973), .o(n28985) );
no02f01 g25195 ( .a(n28833), .b(n_27014), .o(n28986) );
no03f01 g25196 ( .a(n28986), .b(n28985), .c(n28984), .o(n28987) );
no02f01 g25197 ( .a(n28144), .b(delay_add_ln22_unr17_stage7_stallmux_q_31_), .o(n28988) );
na02f01 g25198 ( .a(n28144), .b(delay_add_ln22_unr17_stage7_stallmux_q_31_), .o(n28989) );
in01f01 g25199 ( .a(n28989), .o(n28990) );
no02f01 g25200 ( .a(n28990), .b(n28988), .o(n28991) );
in01f01 g25201 ( .a(n28991), .o(n28992) );
na02f01 g25202 ( .a(n28338), .b(n28335), .o(n28993) );
no03f01 g25203 ( .a(n28374), .b(n28993), .c(n28145), .o(n28994) );
no03f01 g25204 ( .a(n28373), .b(n28369), .c(n28365), .o(n28995) );
in01f01 g25205 ( .a(n28995), .o(n28996) );
no03f01 g25206 ( .a(n28996), .b(n28994), .c(n28992), .o(n28997) );
no02f01 g25207 ( .a(n28996), .b(n28994), .o(n28998) );
no02f01 g25208 ( .a(n28998), .b(n28991), .o(n28999) );
no02f01 g25209 ( .a(n28999), .b(n28997), .o(n29000) );
in01f01 g25210 ( .a(n29000), .o(n29001) );
no02f01 g25211 ( .a(n29001), .b(n28102), .o(n29002) );
no02f01 g25212 ( .a(n29000), .b(n28383), .o(n29003) );
no02f01 g25213 ( .a(n29003), .b(n29002), .o(n29004) );
na02f01 g25214 ( .a(n28829), .b(n28380), .o(n29005) );
ao22f01 g25215 ( .a(n29005), .b(n28102), .c(n28824), .d(n28381), .o(n29006) );
na02f01 g25216 ( .a(n29006), .b(n29004), .o(n29007) );
in01f01 g25217 ( .a(n29007), .o(n29008) );
no02f01 g25218 ( .a(n29006), .b(n29004), .o(n29009) );
no02f01 g25219 ( .a(n29009), .b(n29008), .o(n29010) );
no02f01 g25220 ( .a(n29010), .b(n_27014), .o(n29011) );
no02f01 g25221 ( .a(n29010), .b(n27681), .o(n29012) );
no02f01 g25222 ( .a(n29012), .b(n29011), .o(n29013) );
na02f01 g25223 ( .a(n29013), .b(n28987), .o(n29014) );
in01f01 g25224 ( .a(n28984), .o(n29015) );
no02f01 g25225 ( .a(n28986), .b(n28985), .o(n29016) );
na02f01 g25226 ( .a(n29016), .b(n29015), .o(n29017) );
in01f01 g25227 ( .a(n29009), .o(n29018) );
na02f01 g25228 ( .a(n29018), .b(n29007), .o(n29019) );
na02f01 g25229 ( .a(n29019), .b(n27681), .o(n29020) );
na02f01 g25230 ( .a(n29019), .b(n_27014), .o(n29021) );
na02f01 g25231 ( .a(n29021), .b(n29020), .o(n29022) );
na02f01 g25232 ( .a(n29022), .b(n29017), .o(n29023) );
no02f01 g25233 ( .a(n28807), .b(n27682), .o(n29024) );
in01f01 g25234 ( .a(n29024), .o(n29025) );
no02f01 g25235 ( .a(n28793), .b(n27682), .o(n29026) );
no02f01 g25236 ( .a(n28795), .b(n_25834), .o(n29027) );
no02f01 g25237 ( .a(n28731), .b(n27682), .o(n29028) );
ao12f01 g25238 ( .a(n27682), .b(n28729), .c(n28681), .o(n29029) );
no03f01 g25239 ( .a(n29029), .b(n29028), .c(n28724), .o(n29030) );
no02f01 g25240 ( .a(n29030), .b(n27682), .o(n29031) );
in01f01 g25241 ( .a(n29031), .o(n29032) );
oa12f01 g25242 ( .a(n_25834), .b(n28753), .c(n28713), .o(n29033) );
na02f01 g25243 ( .a(n29033), .b(n29032), .o(n29034) );
ao12f01 g25244 ( .a(n29034), .b(n28763), .c(n_25834), .o(n29035) );
na02f01 g25245 ( .a(n28783), .b(n_25834), .o(n29036) );
ao12f01 g25246 ( .a(n29027), .b(n29036), .c(n29035), .o(n29037) );
no02f01 g25247 ( .a(n29037), .b(n29026), .o(n29038) );
na02f01 g25248 ( .a(n29038), .b(n29025), .o(n29039) );
no02f01 g25249 ( .a(n29039), .b(n28821), .o(n29040) );
na02f01 g25250 ( .a(n28776), .b(n_25834), .o(n29041) );
na02f01 g25251 ( .a(n28783), .b(n27682), .o(n29042) );
ao12f01 g25252 ( .a(n27682), .b(n28788), .c(n28734), .o(n29043) );
no02f01 g25253 ( .a(n29043), .b(n29031), .o(n29044) );
oa12f01 g25254 ( .a(n29044), .b(n28790), .c(n27682), .o(n29045) );
no02f01 g25255 ( .a(n28795), .b(n27682), .o(n29046) );
oa12f01 g25256 ( .a(n29042), .b(n29046), .c(n29045), .o(n29047) );
na02f01 g25257 ( .a(n29047), .b(n29041), .o(n29048) );
no02f01 g25258 ( .a(n29048), .b(n29024), .o(n29049) );
no02f01 g25259 ( .a(n29049), .b(n28822), .o(n29050) );
no02f01 g25260 ( .a(n27871), .b(n27754), .o(n29051) );
in01f01 g25261 ( .a(n29051), .o(n29052) );
no02f01 g25262 ( .a(n29052), .b(n27868), .o(n29053) );
no02f01 g25263 ( .a(n29051), .b(n27869), .o(n29054) );
no02f01 g25264 ( .a(n29054), .b(n29053), .o(n29055) );
no03f01 g25265 ( .a(n29055), .b(n29050), .c(n29040), .o(n29056) );
na02f01 g25266 ( .a(n29038), .b(n28808), .o(n29057) );
na02f01 g25267 ( .a(n29048), .b(n28807), .o(n29058) );
no02f01 g25268 ( .a(n27866), .b(n27763), .o(n29059) );
in01f01 g25269 ( .a(n29059), .o(n29060) );
no02f01 g25270 ( .a(n29060), .b(n27864), .o(n29061) );
na02f01 g25271 ( .a(n29060), .b(n27864), .o(n29062) );
in01f01 g25272 ( .a(n29062), .o(n29063) );
no02f01 g25273 ( .a(n29063), .b(n29061), .o(n29064) );
in01f01 g25274 ( .a(n29064), .o(n29065) );
ao12f01 g25275 ( .a(n29065), .b(n29058), .c(n29057), .o(n29066) );
no02f01 g25276 ( .a(n28793), .b(n_25834), .o(n29067) );
no02f01 g25277 ( .a(n29067), .b(n29026), .o(n29068) );
no02f01 g25278 ( .a(n29068), .b(n29037), .o(n29069) );
na02f01 g25279 ( .a(n28776), .b(n27682), .o(n29070) );
na02f01 g25280 ( .a(n29070), .b(n29041), .o(n29071) );
no02f01 g25281 ( .a(n29071), .b(n29047), .o(n29072) );
no02f01 g25282 ( .a(n27863), .b(n27772), .o(n29073) );
in01f01 g25283 ( .a(n29073), .o(n29074) );
ao12f01 g25284 ( .a(n29074), .b(n27861), .c(n27782), .o(n29075) );
no02f01 g25285 ( .a(n29073), .b(n27862), .o(n29076) );
no02f01 g25286 ( .a(n29076), .b(n29075), .o(n29077) );
no03f01 g25287 ( .a(n29077), .b(n29072), .c(n29069), .o(n29078) );
in01f01 g25288 ( .a(n27859), .o(n29079) );
ao12f01 g25289 ( .a(n27855), .b(n29079), .c(n27845), .o(n29080) );
in01f01 g25290 ( .a(n29080), .o(n29081) );
no02f01 g25291 ( .a(n27857), .b(n27781), .o(n29082) );
no02f01 g25292 ( .a(n29082), .b(n29081), .o(n29083) );
na02f01 g25293 ( .a(n29082), .b(n29081), .o(n29084) );
in01f01 g25294 ( .a(n29084), .o(n29085) );
no02f01 g25295 ( .a(n29085), .b(n29083), .o(n29086) );
in01f01 g25296 ( .a(n29086), .o(n29087) );
na02f01 g25297 ( .a(n28701), .b(n_25834), .o(n29088) );
oa12f01 g25298 ( .a(n_25834), .b(n28693), .c(n28640), .o(n29089) );
na03f01 g25299 ( .a(n29089), .b(n29088), .c(n28737), .o(n29090) );
oa12f01 g25300 ( .a(n_25834), .b(n29090), .c(n28713), .o(n29091) );
no02f01 g25301 ( .a(n29091), .b(n28753), .o(n29092) );
ao12f01 g25302 ( .a(n27682), .b(n29030), .c(n28734), .o(n29093) );
no02f01 g25303 ( .a(n29093), .b(n28788), .o(n29094) );
in01f01 g25304 ( .a(n27842), .o(n29095) );
no02f01 g25305 ( .a(n29095), .b(n27841), .o(n29096) );
in01f01 g25306 ( .a(n27843), .o(n29097) );
no02f01 g25307 ( .a(n29097), .b(n27792), .o(n29098) );
no02f01 g25308 ( .a(n29098), .b(n29096), .o(n29099) );
na02f01 g25309 ( .a(n29098), .b(n29096), .o(n29100) );
in01f01 g25310 ( .a(n29100), .o(n29101) );
no02f01 g25311 ( .a(n29101), .b(n29099), .o(n29102) );
no03f01 g25312 ( .a(n29102), .b(n29094), .c(n29092), .o(n29103) );
oa12f01 g25313 ( .a(n28713), .b(n29030), .c(n27682), .o(n29104) );
na03f01 g25314 ( .a(n29090), .b(n28734), .c(n_25834), .o(n29105) );
in01f01 g25315 ( .a(n27832), .o(n29106) );
no03f01 g25316 ( .a(n29095), .b(n27840), .c(n29106), .o(n29107) );
in01f01 g25317 ( .a(n27840), .o(n29108) );
ao12f01 g25318 ( .a(n27832), .b(n27842), .c(n29108), .o(n29109) );
no02f01 g25319 ( .a(n29109), .b(n29107), .o(n29110) );
in01f01 g25320 ( .a(n29110), .o(n29111) );
na03f01 g25321 ( .a(n29111), .b(n29105), .c(n29104), .o(n29112) );
ao12f01 g25322 ( .a(n29111), .b(n29105), .c(n29104), .o(n29113) );
ao12f01 g25323 ( .a(n28724), .b(n29089), .c(n29088), .o(n29114) );
no03f01 g25324 ( .a(n29029), .b(n29028), .c(n28737), .o(n29115) );
in01f01 g25325 ( .a(n27829), .o(n29116) );
no02f01 g25326 ( .a(n27831), .b(n27801), .o(n29117) );
no02f01 g25327 ( .a(n29117), .b(n29116), .o(n29118) );
na02f01 g25328 ( .a(n29117), .b(n29116), .o(n29119) );
in01f01 g25329 ( .a(n29119), .o(n29120) );
no02f01 g25330 ( .a(n29120), .b(n29118), .o(n29121) );
no03f01 g25331 ( .a(n29121), .b(n29115), .c(n29114), .o(n29122) );
na02f01 g25332 ( .a(n29089), .b(n28701), .o(n29123) );
na02f01 g25333 ( .a(n29029), .b(n28731), .o(n29124) );
in01f01 g25334 ( .a(n27813), .o(n29125) );
in01f01 g25335 ( .a(n27827), .o(n29126) );
no03f01 g25336 ( .a(n27828), .b(n29126), .c(n29125), .o(n29127) );
in01f01 g25337 ( .a(n27828), .o(n29128) );
ao12f01 g25338 ( .a(n27827), .b(n29128), .c(n27813), .o(n29129) );
no02f01 g25339 ( .a(n29129), .b(n29127), .o(n29130) );
in01f01 g25340 ( .a(n29130), .o(n29131) );
na03f01 g25341 ( .a(n29131), .b(n29124), .c(n29123), .o(n29132) );
ao12f01 g25342 ( .a(n29131), .b(n29124), .c(n29123), .o(n29133) );
in01f01 g25343 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_0_), .o(n29134) );
no02f01 g25344 ( .a(n27824), .b(n29134), .o(n29135) );
no02f01 g25345 ( .a(n27823), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_0_), .o(n29136) );
no02f01 g25346 ( .a(n29136), .b(n29135), .o(n29137) );
no02f01 g25347 ( .a(n29137), .b(n28681), .o(n29138) );
in01f01 g25348 ( .a(n27820), .o(n29139) );
no03f01 g25349 ( .a(n27826), .b(n29139), .c(n27819), .o(n29140) );
in01f01 g25350 ( .a(n27819), .o(n29141) );
ao12f01 g25351 ( .a(n27825), .b(n27820), .c(n29141), .o(n29142) );
no02f01 g25352 ( .a(n29142), .b(n29140), .o(n29143) );
no02f01 g25353 ( .a(n29143), .b(n29138), .o(n29144) );
no03f01 g25354 ( .a(n28693), .b(n28681), .c(n27682), .o(n29145) );
ao12f01 g25355 ( .a(n28729), .b(n28640), .c(n_25834), .o(n29146) );
no02f01 g25356 ( .a(n29146), .b(n29145), .o(n29147) );
in01f01 g25357 ( .a(n29143), .o(n29148) );
no03f01 g25358 ( .a(n29148), .b(n29137), .c(n28681), .o(n29149) );
in01f01 g25359 ( .a(n29149), .o(n29150) );
ao12f01 g25360 ( .a(n29144), .b(n29150), .c(n29147), .o(n29151) );
oa12f01 g25361 ( .a(n29132), .b(n29151), .c(n29133), .o(n29152) );
oa12f01 g25362 ( .a(n29121), .b(n29115), .c(n29114), .o(n29153) );
ao12f01 g25363 ( .a(n29122), .b(n29153), .c(n29152), .o(n29154) );
oa12f01 g25364 ( .a(n29112), .b(n29154), .c(n29113), .o(n29155) );
oa12f01 g25365 ( .a(n29102), .b(n29094), .c(n29092), .o(n29156) );
ao12f01 g25366 ( .a(n29103), .b(n29156), .c(n29155), .o(n29157) );
oa12f01 g25367 ( .a(n28790), .b(n29043), .c(n29031), .o(n29158) );
na03f01 g25368 ( .a(n29033), .b(n29032), .c(n28763), .o(n29159) );
no02f01 g25369 ( .a(n27859), .b(n27855), .o(n29160) );
no02f01 g25370 ( .a(n29160), .b(n27845), .o(n29161) );
na02f01 g25371 ( .a(n29160), .b(n27845), .o(n29162) );
in01f01 g25372 ( .a(n29162), .o(n29163) );
no02f01 g25373 ( .a(n29163), .b(n29161), .o(n29164) );
in01f01 g25374 ( .a(n29164), .o(n29165) );
ao12f01 g25375 ( .a(n29165), .b(n29159), .c(n29158), .o(n29166) );
na03f01 g25376 ( .a(n29165), .b(n29159), .c(n29158), .o(n29167) );
oa12f01 g25377 ( .a(n29167), .b(n29166), .c(n29157), .o(n29168) );
no02f01 g25378 ( .a(n29046), .b(n29027), .o(n29169) );
no02f01 g25379 ( .a(n29169), .b(n29045), .o(n29170) );
na02f01 g25380 ( .a(n29036), .b(n29042), .o(n29171) );
no02f01 g25381 ( .a(n29171), .b(n29035), .o(n29172) );
no02f01 g25382 ( .a(n29172), .b(n29170), .o(n29173) );
ao12f01 g25383 ( .a(n28763), .b(n29033), .c(n29032), .o(n29174) );
no03f01 g25384 ( .a(n29043), .b(n29031), .c(n28790), .o(n29175) );
no03f01 g25385 ( .a(n29164), .b(n29175), .c(n29174), .o(n29176) );
no02f01 g25386 ( .a(n29176), .b(n29087), .o(n29177) );
oa12f01 g25387 ( .a(n29177), .b(n29166), .c(n29157), .o(n29178) );
ao22f01 g25388 ( .a(n29178), .b(n29173), .c(n29168), .d(n29087), .o(n29179) );
na02f01 g25389 ( .a(n29071), .b(n29047), .o(n29180) );
na02f01 g25390 ( .a(n29068), .b(n29037), .o(n29181) );
in01f01 g25391 ( .a(n29077), .o(n29182) );
ao12f01 g25392 ( .a(n29182), .b(n29181), .c(n29180), .o(n29183) );
no02f01 g25393 ( .a(n29183), .b(n29179), .o(n29184) );
no02f01 g25394 ( .a(n29048), .b(n28807), .o(n29185) );
no02f01 g25395 ( .a(n29038), .b(n28808), .o(n29186) );
no03f01 g25396 ( .a(n29064), .b(n29186), .c(n29185), .o(n29187) );
no03f01 g25397 ( .a(n29187), .b(n29184), .c(n29078), .o(n29188) );
oa12f01 g25398 ( .a(n29055), .b(n29050), .c(n29040), .o(n29189) );
in01f01 g25399 ( .a(n29189), .o(n29190) );
no03f01 g25400 ( .a(n29190), .b(n29188), .c(n29066), .o(n29191) );
no02f01 g25401 ( .a(n29191), .b(n29056), .o(n29192) );
oa12f01 g25402 ( .a(n29049), .b(n28821), .c(n27682), .o(n29193) );
na02f01 g25403 ( .a(n29193), .b(n28380), .o(n29194) );
ao12f01 g25404 ( .a(n29039), .b(n28822), .c(n_25834), .o(n29195) );
na02f01 g25405 ( .a(n29195), .b(n28381), .o(n29196) );
na02f01 g25406 ( .a(n29196), .b(n29194), .o(n29197) );
no02f01 g25407 ( .a(n27874), .b(n27746), .o(n29198) );
in01f01 g25408 ( .a(n29198), .o(n29199) );
no03f01 g25409 ( .a(n29199), .b(n27872), .c(n27754), .o(n29200) );
no02f01 g25410 ( .a(n27872), .b(n27754), .o(n29201) );
no02f01 g25411 ( .a(n29198), .b(n29201), .o(n29202) );
no02f01 g25412 ( .a(n29202), .b(n29200), .o(n29203) );
no02f01 g25413 ( .a(n29203), .b(n29197), .o(n29204) );
in01f01 g25414 ( .a(n29203), .o(n29205) );
ao12f01 g25415 ( .a(n29205), .b(n29196), .c(n29194), .o(n29206) );
no02f01 g25416 ( .a(n29206), .b(n29204), .o(n29207) );
no02f01 g25417 ( .a(n29207), .b(n29192), .o(n29208) );
na02f01 g25418 ( .a(n29207), .b(n29192), .o(n29209) );
in01f01 g25419 ( .a(n29209), .o(n29210) );
no02f01 g25420 ( .a(n29210), .b(n29208), .o(n29211) );
in01f01 g25421 ( .a(n29211), .o(n29212) );
ao12f01 g25422 ( .a(n29212), .b(n29023), .c(n29014), .o(n29213) );
no02f01 g25423 ( .a(n28983), .b(n28976), .o(n29214) );
no02f01 g25424 ( .a(n28986), .b(n28834), .o(n29215) );
in01f01 g25425 ( .a(n29215), .o(n29216) );
no03f01 g25426 ( .a(n29216), .b(n28985), .c(n29214), .o(n29217) );
no02f01 g25427 ( .a(n28985), .b(n29214), .o(n29218) );
no02f01 g25428 ( .a(n29218), .b(n29215), .o(n29219) );
in01f01 g25429 ( .a(n29066), .o(n29220) );
in01f01 g25430 ( .a(n29078), .o(n29221) );
in01f01 g25431 ( .a(n29103), .o(n29222) );
ao12f01 g25432 ( .a(n28734), .b(n29090), .c(n_25834), .o(n29223) );
no03f01 g25433 ( .a(n29030), .b(n28713), .c(n27682), .o(n29224) );
no03f01 g25434 ( .a(n29110), .b(n29224), .c(n29223), .o(n29225) );
oa12f01 g25435 ( .a(n29110), .b(n29224), .c(n29223), .o(n29226) );
oa12f01 g25436 ( .a(n28737), .b(n29029), .c(n29028), .o(n29227) );
na03f01 g25437 ( .a(n29089), .b(n29088), .c(n28724), .o(n29228) );
in01f01 g25438 ( .a(n29121), .o(n29229) );
na03f01 g25439 ( .a(n29229), .b(n29228), .c(n29227), .o(n29230) );
no02f01 g25440 ( .a(n29029), .b(n28731), .o(n29231) );
no02f01 g25441 ( .a(n29089), .b(n28701), .o(n29232) );
no03f01 g25442 ( .a(n29130), .b(n29232), .c(n29231), .o(n29233) );
oa12f01 g25443 ( .a(n29130), .b(n29232), .c(n29231), .o(n29234) );
in01f01 g25444 ( .a(n29144), .o(n29235) );
na03f01 g25445 ( .a(n28729), .b(n28640), .c(n_25834), .o(n29236) );
oa12f01 g25446 ( .a(n28693), .b(n28681), .c(n27682), .o(n29237) );
na02f01 g25447 ( .a(n29237), .b(n29236), .o(n29238) );
oa12f01 g25448 ( .a(n29235), .b(n29149), .c(n29238), .o(n29239) );
ao12f01 g25449 ( .a(n29233), .b(n29239), .c(n29234), .o(n29240) );
ao12f01 g25450 ( .a(n29229), .b(n29228), .c(n29227), .o(n29241) );
oa12f01 g25451 ( .a(n29230), .b(n29241), .c(n29240), .o(n29242) );
ao12f01 g25452 ( .a(n29225), .b(n29242), .c(n29226), .o(n29243) );
na02f01 g25453 ( .a(n29093), .b(n28788), .o(n29244) );
na02f01 g25454 ( .a(n29091), .b(n28753), .o(n29245) );
in01f01 g25455 ( .a(n29102), .o(n29246) );
ao12f01 g25456 ( .a(n29246), .b(n29245), .c(n29244), .o(n29247) );
oa12f01 g25457 ( .a(n29222), .b(n29247), .c(n29243), .o(n29248) );
in01f01 g25458 ( .a(n29166), .o(n29249) );
ao12f01 g25459 ( .a(n29176), .b(n29249), .c(n29248), .o(n29250) );
na02f01 g25460 ( .a(n29171), .b(n29035), .o(n29251) );
na02f01 g25461 ( .a(n29169), .b(n29045), .o(n29252) );
na02f01 g25462 ( .a(n29252), .b(n29251), .o(n29253) );
na02f01 g25463 ( .a(n29167), .b(n29086), .o(n29254) );
ao12f01 g25464 ( .a(n29254), .b(n29249), .c(n29248), .o(n29255) );
oa22f01 g25465 ( .a(n29255), .b(n29253), .c(n29250), .d(n29086), .o(n29256) );
oa12f01 g25466 ( .a(n29077), .b(n29072), .c(n29069), .o(n29257) );
na02f01 g25467 ( .a(n29257), .b(n29256), .o(n29258) );
na03f01 g25468 ( .a(n29065), .b(n29058), .c(n29057), .o(n29259) );
na03f01 g25469 ( .a(n29259), .b(n29258), .c(n29221), .o(n29260) );
na02f01 g25470 ( .a(n29260), .b(n29220), .o(n29261) );
no02f01 g25471 ( .a(n29190), .b(n29056), .o(n29262) );
no02f01 g25472 ( .a(n29262), .b(n29261), .o(n29263) );
na02f01 g25473 ( .a(n29262), .b(n29261), .o(n29264) );
in01f01 g25474 ( .a(n29264), .o(n29265) );
no02f01 g25475 ( .a(n29265), .b(n29263), .o(n29266) );
no03f01 g25476 ( .a(n29266), .b(n29219), .c(n29217), .o(n29267) );
no02f01 g25477 ( .a(n28973), .b(n_27014), .o(n29268) );
in01f01 g25478 ( .a(n29268), .o(n29269) );
no02f01 g25479 ( .a(n28982), .b(n_27014), .o(n29270) );
no02f01 g25480 ( .a(n29270), .b(n28983), .o(n29271) );
ao12f01 g25481 ( .a(n29271), .b(n29269), .c(n28976), .o(n29272) );
na03f01 g25482 ( .a(n29271), .b(n29269), .c(n28976), .o(n29273) );
in01f01 g25483 ( .a(n29273), .o(n29274) );
no02f01 g25484 ( .a(n29184), .b(n29078), .o(n29275) );
no02f01 g25485 ( .a(n29187), .b(n29066), .o(n29276) );
no02f01 g25486 ( .a(n29276), .b(n29275), .o(n29277) );
na02f01 g25487 ( .a(n29276), .b(n29275), .o(n29278) );
in01f01 g25488 ( .a(n29278), .o(n29279) );
no02f01 g25489 ( .a(n29279), .b(n29277), .o(n29280) );
no03f01 g25490 ( .a(n29280), .b(n29274), .c(n29272), .o(n29281) );
no02f01 g25491 ( .a(n29268), .b(n28974), .o(n29282) );
in01f01 g25492 ( .a(n29282), .o(n29283) );
oa12f01 g25493 ( .a(n29283), .b(n28967), .c(n28963), .o(n29284) );
in01f01 g25494 ( .a(n29284), .o(n29285) );
no03f01 g25495 ( .a(n29283), .b(n28967), .c(n28963), .o(n29286) );
no02f01 g25496 ( .a(n29183), .b(n29078), .o(n29287) );
no02f01 g25497 ( .a(n29287), .b(n29179), .o(n29288) );
na02f01 g25498 ( .a(n29287), .b(n29179), .o(n29289) );
in01f01 g25499 ( .a(n29289), .o(n29290) );
no02f01 g25500 ( .a(n29290), .b(n29288), .o(n29291) );
no03f01 g25501 ( .a(n29291), .b(n29286), .c(n29285), .o(n29292) );
na02f01 g25502 ( .a(n28886), .b(n28885), .o(n29293) );
na02f01 g25503 ( .a(n28882), .b(n28880), .o(n29294) );
na02f01 g25504 ( .a(n29294), .b(n29293), .o(n29295) );
in01f01 g25505 ( .a(n28893), .o(n29296) );
oa12f01 g25506 ( .a(n_27014), .b(n29296), .c(n29295), .o(n29297) );
na02f01 g25507 ( .a(n28903), .b(n29297), .o(n29298) );
in01f01 g25508 ( .a(n28915), .o(n29299) );
oa12f01 g25509 ( .a(n28916), .b(n29299), .c(n29298), .o(n29300) );
in01f01 g25510 ( .a(n28925), .o(n29301) );
na02f01 g25511 ( .a(n29301), .b(n29300), .o(n29302) );
in01f01 g25512 ( .a(n28935), .o(n29303) );
no03f01 g25513 ( .a(n28945), .b(n29303), .c(n29302), .o(n29304) );
in01f01 g25514 ( .a(n28961), .o(n29305) );
na02f01 g25515 ( .a(n28966), .b(n29305), .o(n29306) );
oa12f01 g25516 ( .a(n27681), .b(n28956), .c(n28954), .o(n29307) );
oa12f01 g25517 ( .a(n_27014), .b(n28956), .c(n28954), .o(n29308) );
na02f01 g25518 ( .a(n29308), .b(n29307), .o(n29309) );
oa12f01 g25519 ( .a(n29309), .b(n29306), .c(n29304), .o(n29310) );
in01f01 g25520 ( .a(n28966), .o(n29311) );
no02f01 g25521 ( .a(n29311), .b(n28961), .o(n29312) );
ao12f01 g25522 ( .a(n_27014), .b(n28959), .c(n28958), .o(n29313) );
ao12f01 g25523 ( .a(n27681), .b(n28959), .c(n28958), .o(n29314) );
no02f01 g25524 ( .a(n29314), .b(n29313), .o(n29315) );
na03f01 g25525 ( .a(n29315), .b(n29312), .c(n28947), .o(n29316) );
ao12f01 g25526 ( .a(n29166), .b(n29167), .c(n29157), .o(n29317) );
no02f01 g25527 ( .a(n29173), .b(n29087), .o(n29318) );
no02f01 g25528 ( .a(n29253), .b(n29086), .o(n29319) );
no02f01 g25529 ( .a(n29319), .b(n29318), .o(n29320) );
in01f01 g25530 ( .a(n29320), .o(n29321) );
no02f01 g25531 ( .a(n29321), .b(n29317), .o(n29322) );
na02f01 g25532 ( .a(n29321), .b(n29317), .o(n29323) );
in01f01 g25533 ( .a(n29323), .o(n29324) );
no02f01 g25534 ( .a(n29324), .b(n29322), .o(n29325) );
in01f01 g25535 ( .a(n29325), .o(n29326) );
ao12f01 g25536 ( .a(n29326), .b(n29316), .c(n29310), .o(n29327) );
na02f01 g25537 ( .a(n28934), .b(n27681), .o(n29328) );
na02f01 g25538 ( .a(n29328), .b(n28935), .o(n29329) );
na02f01 g25539 ( .a(n29329), .b(n28926), .o(n29330) );
no02f01 g25540 ( .a(n29329), .b(n28926), .o(n29331) );
in01f01 g25541 ( .a(n29331), .o(n29332) );
no03f01 g25542 ( .a(n29247), .b(n29155), .c(n29103), .o(n29333) );
ao12f01 g25543 ( .a(n29243), .b(n29156), .c(n29222), .o(n29334) );
no02f01 g25544 ( .a(n29334), .b(n29333), .o(n29335) );
in01f01 g25545 ( .a(n29335), .o(n29336) );
ao12f01 g25546 ( .a(n29336), .b(n29332), .c(n29330), .o(n29337) );
no02f01 g25547 ( .a(n28924), .b(n_27014), .o(n29338) );
no02f01 g25548 ( .a(n29338), .b(n28925), .o(n29339) );
no02f01 g25549 ( .a(n29339), .b(n28918), .o(n29340) );
no03f01 g25550 ( .a(n29338), .b(n28925), .c(n29300), .o(n29341) );
no03f01 g25551 ( .a(n29242), .b(n29113), .c(n29225), .o(n29342) );
ao12f01 g25552 ( .a(n29154), .b(n29226), .c(n29112), .o(n29343) );
no02f01 g25553 ( .a(n29343), .b(n29342), .o(n29344) );
no03f01 g25554 ( .a(n29344), .b(n29341), .c(n29340), .o(n29345) );
no03f01 g25555 ( .a(n29241), .b(n29152), .c(n29122), .o(n29346) );
ao12f01 g25556 ( .a(n29240), .b(n29153), .c(n29230), .o(n29347) );
no02f01 g25557 ( .a(n29347), .b(n29346), .o(n29348) );
in01f01 g25558 ( .a(n29348), .o(n29349) );
oa12f01 g25559 ( .a(n28905), .b(n28917), .c(n29299), .o(n29350) );
na03f01 g25560 ( .a(n28916), .b(n28915), .c(n29298), .o(n29351) );
na03f01 g25561 ( .a(n29351), .b(n29350), .c(n29349), .o(n29352) );
oa12f01 g25562 ( .a(n27681), .b(n28902), .c(n28900), .o(n29353) );
na02f01 g25563 ( .a(n29353), .b(n28903), .o(n29354) );
no02f01 g25564 ( .a(n29354), .b(n29297), .o(n29355) );
ao12f01 g25565 ( .a(n28894), .b(n29353), .c(n28903), .o(n29356) );
no03f01 g25566 ( .a(n29239), .b(n29133), .c(n29233), .o(n29357) );
ao12f01 g25567 ( .a(n29151), .b(n29234), .c(n29132), .o(n29358) );
no02f01 g25568 ( .a(n29358), .b(n29357), .o(n29359) );
no03f01 g25569 ( .a(n29359), .b(n29356), .c(n29355), .o(n29360) );
oa12f01 g25570 ( .a(n29359), .b(n29356), .c(n29355), .o(n29361) );
na03f01 g25571 ( .a(n29296), .b(n28888), .c(n_27014), .o(n29362) );
oa12f01 g25572 ( .a(n29295), .b(n28893), .c(n27681), .o(n29363) );
na02f01 g25573 ( .a(n29363), .b(n29362), .o(n29364) );
na02f01 g25574 ( .a(n28893), .b(n27681), .o(n29365) );
na02f01 g25575 ( .a(n28893), .b(n_27014), .o(n29366) );
no02f01 g25576 ( .a(n29137), .b(n28640), .o(n29367) );
in01f01 g25577 ( .a(n29137), .o(n29368) );
no02f01 g25578 ( .a(n29368), .b(n28681), .o(n29369) );
no02f01 g25579 ( .a(n29369), .b(n29367), .o(n29370) );
in01f01 g25580 ( .a(n29370), .o(n29371) );
na03f01 g25581 ( .a(n29371), .b(n29366), .c(n29365), .o(n29372) );
no02f01 g25582 ( .a(n29238), .b(n29143), .o(n29373) );
no02f01 g25583 ( .a(n29147), .b(n29148), .o(n29374) );
no02f01 g25584 ( .a(n29374), .b(n29373), .o(n29375) );
no02f01 g25585 ( .a(n29375), .b(n29138), .o(n29376) );
na02f01 g25586 ( .a(n29375), .b(n29138), .o(n29377) );
in01f01 g25587 ( .a(n29377), .o(n29378) );
no02f01 g25588 ( .a(n29378), .b(n29376), .o(n29379) );
in01f01 g25589 ( .a(n29379), .o(n29380) );
no02f01 g25590 ( .a(n29380), .b(n29372), .o(n29381) );
na02f01 g25591 ( .a(n29380), .b(n29372), .o(n29382) );
oa12f01 g25592 ( .a(n29382), .b(n29381), .c(n29364), .o(n29383) );
ao12f01 g25593 ( .a(n29360), .b(n29383), .c(n29361), .o(n29384) );
ao12f01 g25594 ( .a(n29349), .b(n29351), .c(n29350), .o(n29385) );
oa12f01 g25595 ( .a(n29352), .b(n29385), .c(n29384), .o(n29386) );
oa12f01 g25596 ( .a(n29344), .b(n29341), .c(n29340), .o(n29387) );
ao12f01 g25597 ( .a(n29345), .b(n29387), .c(n29386), .o(n29388) );
na03f01 g25598 ( .a(n29336), .b(n29332), .c(n29330), .o(n29389) );
ao12f01 g25599 ( .a(n29337), .b(n29389), .c(n29388), .o(n29390) );
no02f01 g25600 ( .a(n29303), .b(n29302), .o(n29391) );
no02f01 g25601 ( .a(n28961), .b(n28945), .o(n29392) );
in01f01 g25602 ( .a(n29392), .o(n29393) );
na02f01 g25603 ( .a(n29393), .b(n29391), .o(n29394) );
no02f01 g25604 ( .a(n29393), .b(n29391), .o(n29395) );
in01f01 g25605 ( .a(n29395), .o(n29396) );
no02f01 g25606 ( .a(n29176), .b(n29166), .o(n29397) );
no02f01 g25607 ( .a(n29397), .b(n29157), .o(n29398) );
na02f01 g25608 ( .a(n29397), .b(n29157), .o(n29399) );
in01f01 g25609 ( .a(n29399), .o(n29400) );
no02f01 g25610 ( .a(n29400), .b(n29398), .o(n29401) );
in01f01 g25611 ( .a(n29401), .o(n29402) );
ao12f01 g25612 ( .a(n29402), .b(n29396), .c(n29394), .o(n29403) );
in01f01 g25613 ( .a(n29403), .o(n29404) );
na03f01 g25614 ( .a(n29326), .b(n29316), .c(n29310), .o(n29405) );
na03f01 g25615 ( .a(n29402), .b(n29396), .c(n29394), .o(n29406) );
na02f01 g25616 ( .a(n29406), .b(n29405), .o(n29407) );
ao12f01 g25617 ( .a(n29407), .b(n29404), .c(n29390), .o(n29408) );
in01f01 g25618 ( .a(n29286), .o(n29409) );
in01f01 g25619 ( .a(n29291), .o(n29410) );
ao12f01 g25620 ( .a(n29410), .b(n29409), .c(n29284), .o(n29411) );
no03f01 g25621 ( .a(n29411), .b(n29408), .c(n29327), .o(n29412) );
no03f01 g25622 ( .a(n29412), .b(n29292), .c(n29281), .o(n29413) );
in01f01 g25623 ( .a(n29272), .o(n29414) );
in01f01 g25624 ( .a(n29280), .o(n29415) );
ao12f01 g25625 ( .a(n29415), .b(n29273), .c(n29414), .o(n29416) );
na02f01 g25626 ( .a(n29218), .b(n29215), .o(n29417) );
oa12f01 g25627 ( .a(n29216), .b(n28985), .c(n29214), .o(n29418) );
in01f01 g25628 ( .a(n29266), .o(n29419) );
ao12f01 g25629 ( .a(n29419), .b(n29418), .c(n29417), .o(n29420) );
no03f01 g25630 ( .a(n29420), .b(n29416), .c(n29413), .o(n29421) );
no02f01 g25631 ( .a(n29022), .b(n29017), .o(n29422) );
no02f01 g25632 ( .a(n29013), .b(n28987), .o(n29423) );
no03f01 g25633 ( .a(n29211), .b(n29423), .c(n29422), .o(n29424) );
no03f01 g25634 ( .a(n29424), .b(n29421), .c(n29267), .o(n29425) );
na02f01 g25635 ( .a(n29010), .b(n_27014), .o(n29426) );
na02f01 g25636 ( .a(n29019), .b(n27681), .o(n29427) );
na02f01 g25637 ( .a(n29427), .b(n29426), .o(n29428) );
no02f01 g25638 ( .a(n29017), .b(n_27014), .o(n29429) );
oa22f01 g25639 ( .a(n29429), .b(n29428), .c(n29015), .d(n27681), .o(n29430) );
ao12f01 g25640 ( .a(n27682), .b(n28821), .c(n28380), .o(n29431) );
no02f01 g25641 ( .a(n28381), .b(n_25834), .o(n29432) );
in01f01 g25642 ( .a(n29432), .o(n29433) );
oa12f01 g25643 ( .a(n29433), .b(n29431), .c(n29039), .o(n29434) );
no02f01 g25644 ( .a(n29000), .b(n27682), .o(n29435) );
no02f01 g25645 ( .a(n29000), .b(n_25834), .o(n29436) );
no02f01 g25646 ( .a(n29436), .b(n29435), .o(n29437) );
in01f01 g25647 ( .a(n29437), .o(n29438) );
no02f01 g25648 ( .a(n29438), .b(n29434), .o(n29439) );
na02f01 g25649 ( .a(n29438), .b(n29434), .o(n29440) );
in01f01 g25650 ( .a(n29440), .o(n29441) );
no02f01 g25651 ( .a(n29441), .b(n29439), .o(n29442) );
no02f01 g25652 ( .a(n27875), .b(n27746), .o(n29443) );
in01f01 g25653 ( .a(n29443), .o(n29444) );
no02f01 g25654 ( .a(n27877), .b(n27734), .o(n29445) );
no02f01 g25655 ( .a(n29445), .b(n29444), .o(n29446) );
na02f01 g25656 ( .a(n29445), .b(n29444), .o(n29447) );
in01f01 g25657 ( .a(n29447), .o(n29448) );
no02f01 g25658 ( .a(n29448), .b(n29446), .o(n29449) );
in01f01 g25659 ( .a(n29449), .o(n29450) );
no02f01 g25660 ( .a(n29450), .b(n29442), .o(n29451) );
no03f01 g25661 ( .a(n29449), .b(n29441), .c(n29439), .o(n29452) );
in01f01 g25662 ( .a(n29452), .o(n29453) );
in01f01 g25663 ( .a(n29056), .o(n29454) );
na03f01 g25664 ( .a(n29189), .b(n29260), .c(n29220), .o(n29455) );
ao12f01 g25665 ( .a(n29206), .b(n29455), .c(n29454), .o(n29456) );
no02f01 g25666 ( .a(n29456), .b(n29204), .o(n29457) );
ao12f01 g25667 ( .a(n29451), .b(n29457), .c(n29453), .o(n29458) );
in01f01 g25668 ( .a(n29436), .o(n29459) );
ao12f01 g25669 ( .a(n29435), .b(n29459), .c(n29434), .o(n29460) );
no02f01 g25670 ( .a(n27878), .b(n27734), .o(n29461) );
no02f01 g25671 ( .a(n27880), .b(n27727), .o(n29462) );
no02f01 g25672 ( .a(n29462), .b(n29461), .o(n29463) );
na02f01 g25673 ( .a(n29462), .b(n29461), .o(n29464) );
in01f01 g25674 ( .a(n29464), .o(n29465) );
no02f01 g25675 ( .a(n29465), .b(n29463), .o(n29466) );
na02f01 g25676 ( .a(n29466), .b(n29460), .o(n29467) );
in01f01 g25677 ( .a(n29467), .o(n29468) );
no02f01 g25678 ( .a(n29466), .b(n29460), .o(n29469) );
no02f01 g25679 ( .a(n29469), .b(n29468), .o(n29470) );
in01f01 g25680 ( .a(n29470), .o(n29471) );
no02f01 g25681 ( .a(n29471), .b(n29458), .o(n29472) );
na02f01 g25682 ( .a(n29471), .b(n29458), .o(n29473) );
in01f01 g25683 ( .a(n29473), .o(n29474) );
no02f01 g25684 ( .a(n29474), .b(n29472), .o(n29475) );
in01f01 g25685 ( .a(n29475), .o(n29476) );
no02f01 g25686 ( .a(n29452), .b(n29451), .o(n29477) );
no02f01 g25687 ( .a(n29477), .b(n29457), .o(n29478) );
na02f01 g25688 ( .a(n29477), .b(n29457), .o(n29479) );
in01f01 g25689 ( .a(n29479), .o(n29480) );
no02f01 g25690 ( .a(n29480), .b(n29478), .o(n29481) );
in01f01 g25691 ( .a(n29481), .o(n29482) );
ao12f01 g25692 ( .a(n29430), .b(n29482), .c(n29476), .o(n29483) );
oa12f01 g25693 ( .a(n29467), .b(n29469), .c(n29452), .o(n29484) );
in01f01 g25694 ( .a(n29484), .o(n29485) );
in01f01 g25695 ( .a(n29204), .o(n29486) );
in01f01 g25696 ( .a(n29206), .o(n29487) );
oa12f01 g25697 ( .a(n29487), .b(n29191), .c(n29056), .o(n29488) );
oa12f01 g25698 ( .a(n29467), .b(n29450), .c(n29442), .o(n29489) );
ao12f01 g25699 ( .a(n29489), .b(n29488), .c(n29486), .o(n29490) );
in01f01 g25700 ( .a(n29460), .o(n29491) );
no02f01 g25701 ( .a(n27721), .b(n27882), .o(n29492) );
no02f01 g25702 ( .a(n27887), .b(n29492), .o(n29493) );
in01f01 g25703 ( .a(n29493), .o(n29494) );
no02f01 g25704 ( .a(n29494), .b(n28006), .o(n29495) );
no03f01 g25705 ( .a(n29493), .b(n27881), .c(n27727), .o(n29496) );
no02f01 g25706 ( .a(n29496), .b(n29495), .o(n29497) );
in01f01 g25707 ( .a(n29497), .o(n29498) );
no02f01 g25708 ( .a(n29498), .b(n29491), .o(n29499) );
no02f01 g25709 ( .a(n29497), .b(n29460), .o(n29500) );
no02f01 g25710 ( .a(n29500), .b(n29499), .o(n29501) );
in01f01 g25711 ( .a(n29501), .o(n29502) );
no03f01 g25712 ( .a(n29502), .b(n29490), .c(n29485), .o(n29503) );
no02f01 g25713 ( .a(n29490), .b(n29485), .o(n29504) );
no02f01 g25714 ( .a(n29501), .b(n29504), .o(n29505) );
no02f01 g25715 ( .a(n29505), .b(n29503), .o(n29506) );
in01f01 g25716 ( .a(n29506), .o(n29507) );
in01f01 g25717 ( .a(n29500), .o(n29508) );
ao12f01 g25718 ( .a(n29499), .b(n29508), .c(n29504), .o(n29509) );
no02f01 g25719 ( .a(n29492), .b(n28006), .o(n29510) );
no02f01 g25720 ( .a(n29510), .b(n27887), .o(n29511) );
no02f01 g25721 ( .a(n27721), .b(n27883), .o(n29512) );
no02f01 g25722 ( .a(n29512), .b(n27888), .o(n29513) );
in01f01 g25723 ( .a(n29513), .o(n29514) );
no02f01 g25724 ( .a(n29514), .b(n29511), .o(n29515) );
na02f01 g25725 ( .a(n29514), .b(n29511), .o(n29516) );
in01f01 g25726 ( .a(n29516), .o(n29517) );
no02f01 g25727 ( .a(n29517), .b(n29515), .o(n29518) );
in01f01 g25728 ( .a(n29518), .o(n29519) );
no02f01 g25729 ( .a(n29519), .b(n29491), .o(n29520) );
no02f01 g25730 ( .a(n29518), .b(n29460), .o(n29521) );
no02f01 g25731 ( .a(n29521), .b(n29520), .o(n29522) );
in01f01 g25732 ( .a(n29522), .o(n29523) );
no02f01 g25733 ( .a(n29523), .b(n29509), .o(n29524) );
na02f01 g25734 ( .a(n29523), .b(n29509), .o(n29525) );
in01f01 g25735 ( .a(n29525), .o(n29526) );
no02f01 g25736 ( .a(n29526), .b(n29524), .o(n29527) );
in01f01 g25737 ( .a(n29527), .o(n29528) );
ao12f01 g25738 ( .a(n29430), .b(n29528), .c(n29507), .o(n29529) );
no04f01 g25739 ( .a(n29529), .b(n29483), .c(n29425), .d(n29213), .o(n29530) );
oa12f01 g25740 ( .a(n29430), .b(n29528), .c(n29507), .o(n29531) );
oa12f01 g25741 ( .a(n29430), .b(n29482), .c(n29476), .o(n29532) );
na02f01 g25742 ( .a(n29532), .b(n29531), .o(n29533) );
no02f01 g25743 ( .a(n27721), .b(n27919), .o(n29534) );
no02f01 g25744 ( .a(n27720), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_16_), .o(n29535) );
no02f01 g25745 ( .a(n29535), .b(n29534), .o(n29536) );
in01f01 g25746 ( .a(n29536), .o(n29537) );
no02f01 g25747 ( .a(n29537), .b(n28009), .o(n29538) );
no02f01 g25748 ( .a(n29536), .b(n27890), .o(n29539) );
no02f01 g25749 ( .a(n29539), .b(n29538), .o(n29540) );
no02f01 g25750 ( .a(n29540), .b(n29460), .o(n29541) );
oa12f01 g25751 ( .a(n29491), .b(n29519), .c(n29498), .o(n29542) );
in01f01 g25752 ( .a(n29542), .o(n29543) );
no03f01 g25753 ( .a(n29543), .b(n29490), .c(n29485), .o(n29544) );
no02f01 g25754 ( .a(n29520), .b(n29499), .o(n29545) );
in01f01 g25755 ( .a(n29545), .o(n29546) );
no02f01 g25756 ( .a(n29546), .b(n29544), .o(n29547) );
in01f01 g25757 ( .a(n29540), .o(n29548) );
no02f01 g25758 ( .a(n29548), .b(n29491), .o(n29549) );
in01f01 g25759 ( .a(n29549), .o(n29550) );
ao12f01 g25760 ( .a(n29541), .b(n29550), .c(n29547), .o(n29551) );
no02f01 g25761 ( .a(n29535), .b(n27890), .o(n29552) );
no02f01 g25762 ( .a(n29552), .b(n29534), .o(n29553) );
no02f01 g25763 ( .a(n27720), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_17_), .o(n29554) );
no02f01 g25764 ( .a(n27721), .b(n27920), .o(n29555) );
no02f01 g25765 ( .a(n29555), .b(n29554), .o(n29556) );
no02f01 g25766 ( .a(n29556), .b(n29553), .o(n29557) );
na02f01 g25767 ( .a(n29556), .b(n29553), .o(n29558) );
in01f01 g25768 ( .a(n29558), .o(n29559) );
no02f01 g25769 ( .a(n29559), .b(n29557), .o(n29560) );
in01f01 g25770 ( .a(n29560), .o(n29561) );
no02f01 g25771 ( .a(n29561), .b(n29491), .o(n29562) );
no02f01 g25772 ( .a(n29560), .b(n29460), .o(n29563) );
no02f01 g25773 ( .a(n29563), .b(n29562), .o(n29564) );
no02f01 g25774 ( .a(n29564), .b(n29551), .o(n29565) );
na02f01 g25775 ( .a(n29564), .b(n29551), .o(n29566) );
in01f01 g25776 ( .a(n29566), .o(n29567) );
no02f01 g25777 ( .a(n29567), .b(n29565), .o(n29568) );
no02f01 g25778 ( .a(n29549), .b(n29541), .o(n29569) );
in01f01 g25779 ( .a(n29569), .o(n29570) );
no02f01 g25780 ( .a(n29570), .b(n29547), .o(n29571) );
in01f01 g25781 ( .a(n29547), .o(n29572) );
no02f01 g25782 ( .a(n29569), .b(n29572), .o(n29573) );
no02f01 g25783 ( .a(n29573), .b(n29571), .o(n29574) );
no02f01 g25784 ( .a(n29574), .b(n29568), .o(n29575) );
no02f01 g25785 ( .a(n29575), .b(n29430), .o(n29576) );
in01f01 g25786 ( .a(n29576), .o(n29577) );
oa12f01 g25787 ( .a(n29577), .b(n29533), .c(n29530), .o(n29578) );
ao12f01 g25788 ( .a(n29491), .b(n29561), .c(n29548), .o(n29579) );
no02f01 g25789 ( .a(n29579), .b(n29572), .o(n29580) );
ao12f01 g25790 ( .a(n29460), .b(n29560), .c(n29540), .o(n29581) );
no02f01 g25791 ( .a(n27891), .b(n27890), .o(n29582) );
no02f01 g25792 ( .a(n29582), .b(n27921), .o(n29583) );
no02f01 g25793 ( .a(n27970), .b(n27892), .o(n29584) );
no02f01 g25794 ( .a(n29584), .b(n29583), .o(n29585) );
na02f01 g25795 ( .a(n29584), .b(n29583), .o(n29586) );
in01f01 g25796 ( .a(n29586), .o(n29587) );
no02f01 g25797 ( .a(n29587), .b(n29585), .o(n29588) );
in01f01 g25798 ( .a(n29588), .o(n29589) );
no02f01 g25799 ( .a(n29589), .b(n29491), .o(n29590) );
na02f01 g25800 ( .a(n29589), .b(n29491), .o(n29591) );
in01f01 g25801 ( .a(n29591), .o(n29592) );
no02f01 g25802 ( .a(n29592), .b(n29590), .o(n29593) );
in01f01 g25803 ( .a(n29593), .o(n29594) );
no03f01 g25804 ( .a(n29594), .b(n29581), .c(n29580), .o(n29595) );
no02f01 g25805 ( .a(n29581), .b(n29580), .o(n29596) );
no02f01 g25806 ( .a(n29593), .b(n29596), .o(n29597) );
no02f01 g25807 ( .a(n29597), .b(n29595), .o(n29598) );
in01f01 g25808 ( .a(n29598), .o(n29599) );
no02f01 g25809 ( .a(n29599), .b(n29430), .o(n29600) );
in01f01 g25810 ( .a(n29580), .o(n29601) );
no02f01 g25811 ( .a(n29592), .b(n29581), .o(n29602) );
oa12f01 g25812 ( .a(n29602), .b(n29590), .c(n29601), .o(n29603) );
no02f01 g25813 ( .a(n29491), .b(n28534), .o(n29604) );
no02f01 g25814 ( .a(n29460), .b(n28844), .o(n29605) );
no02f01 g25815 ( .a(n29605), .b(n29604), .o(n29606) );
in01f01 g25816 ( .a(n29606), .o(n29607) );
no02f01 g25817 ( .a(n29607), .b(n29603), .o(n29608) );
na02f01 g25818 ( .a(n29607), .b(n29603), .o(n29609) );
in01f01 g25819 ( .a(n29609), .o(n29610) );
no02f01 g25820 ( .a(n29610), .b(n29608), .o(n29611) );
in01f01 g25821 ( .a(n29611), .o(n29612) );
no02f01 g25822 ( .a(n29612), .b(n29430), .o(n29613) );
no02f01 g25823 ( .a(n29613), .b(n29600), .o(n29614) );
in01f01 g25824 ( .a(n29614), .o(n29615) );
no02f01 g25825 ( .a(n29615), .b(n29578), .o(n29616) );
no02f01 g25826 ( .a(n29491), .b(n28492), .o(n29617) );
no02f01 g25827 ( .a(n29460), .b(n27983), .o(n29618) );
no02f01 g25828 ( .a(n29618), .b(n29617), .o(n29619) );
no03f01 g25829 ( .a(n29604), .b(n29590), .c(n29579), .o(n29620) );
in01f01 g25830 ( .a(n29620), .o(n29621) );
no03f01 g25831 ( .a(n29621), .b(n29546), .c(n29544), .o(n29622) );
ao12f01 g25832 ( .a(n29460), .b(n29588), .c(n28844), .o(n29623) );
no02f01 g25833 ( .a(n29623), .b(n29581), .o(n29624) );
in01f01 g25834 ( .a(n29624), .o(n29625) );
no02f01 g25835 ( .a(n29625), .b(n29622), .o(n29626) );
na02f01 g25836 ( .a(n29626), .b(n29619), .o(n29627) );
in01f01 g25837 ( .a(n29619), .o(n29628) );
no02f01 g25838 ( .a(n29468), .b(n29451), .o(n29629) );
oa12f01 g25839 ( .a(n29629), .b(n29456), .c(n29204), .o(n29630) );
na03f01 g25840 ( .a(n29542), .b(n29630), .c(n29484), .o(n29631) );
na03f01 g25841 ( .a(n29620), .b(n29545), .c(n29631), .o(n29632) );
na02f01 g25842 ( .a(n29624), .b(n29632), .o(n29633) );
na02f01 g25843 ( .a(n29633), .b(n29628), .o(n29634) );
na02f01 g25844 ( .a(n29634), .b(n29627), .o(n29635) );
no02f01 g25845 ( .a(n29635), .b(n29430), .o(n29636) );
in01f01 g25846 ( .a(n29636), .o(n29637) );
na02f01 g25847 ( .a(n29637), .b(n29616), .o(n29638) );
in01f01 g25848 ( .a(n29430), .o(n29639) );
ao12f01 g25849 ( .a(n29639), .b(n29611), .c(n29598), .o(n29640) );
in01f01 g25850 ( .a(n29568), .o(n29641) );
in01f01 g25851 ( .a(n29574), .o(n29642) );
no02f01 g25852 ( .a(n29642), .b(n29641), .o(n29643) );
no02f01 g25853 ( .a(n29643), .b(n29639), .o(n29644) );
no02f01 g25854 ( .a(n29644), .b(n29640), .o(n29645) );
in01f01 g25855 ( .a(n29645), .o(n29646) );
no02f01 g25856 ( .a(n29633), .b(n29628), .o(n29647) );
no02f01 g25857 ( .a(n29626), .b(n29619), .o(n29648) );
no02f01 g25858 ( .a(n29648), .b(n29647), .o(n29649) );
no02f01 g25859 ( .a(n29649), .b(n29639), .o(n29650) );
no02f01 g25860 ( .a(n29650), .b(n29646), .o(n29651) );
in01f01 g25861 ( .a(n29618), .o(n29652) );
no02f01 g25862 ( .a(n29460), .b(n28496), .o(n29653) );
no02f01 g25863 ( .a(n29491), .b(n27995), .o(n29654) );
no02f01 g25864 ( .a(n29654), .b(n29653), .o(n29655) );
in01f01 g25865 ( .a(n29617), .o(n29656) );
oa12f01 g25866 ( .a(n29656), .b(n29625), .c(n29622), .o(n29657) );
na03f01 g25867 ( .a(n29657), .b(n29655), .c(n29652), .o(n29658) );
in01f01 g25868 ( .a(n29655), .o(n29659) );
ao12f01 g25869 ( .a(n29617), .b(n29624), .c(n29632), .o(n29660) );
oa12f01 g25870 ( .a(n29659), .b(n29660), .c(n29618), .o(n29661) );
na02f01 g25871 ( .a(n29661), .b(n29658), .o(n29662) );
no02f01 g25872 ( .a(n29662), .b(n29430), .o(n29663) );
no03f01 g25873 ( .a(n29660), .b(n29659), .c(n29618), .o(n29664) );
ao12f01 g25874 ( .a(n29655), .b(n29657), .c(n29652), .o(n29665) );
no02f01 g25875 ( .a(n29665), .b(n29664), .o(n29666) );
no02f01 g25876 ( .a(n29666), .b(n29639), .o(n29667) );
no02f01 g25877 ( .a(n29667), .b(n29663), .o(n29668) );
na03f01 g25878 ( .a(n29668), .b(n29651), .c(n29638), .o(n29669) );
in01f01 g25879 ( .a(n29213), .o(n29670) );
in01f01 g25880 ( .a(n29267), .o(n29671) );
na03f01 g25881 ( .a(n29415), .b(n29273), .c(n29414), .o(n29672) );
in01f01 g25882 ( .a(n29292), .o(n29673) );
in01f01 g25883 ( .a(n29327), .o(n29674) );
in01f01 g25884 ( .a(n29330), .o(n29675) );
oa12f01 g25885 ( .a(n29335), .b(n29331), .c(n29675), .o(n29676) );
in01f01 g25886 ( .a(n29345), .o(n29677) );
ao12f01 g25887 ( .a(n29298), .b(n28916), .c(n28915), .o(n29678) );
no03f01 g25888 ( .a(n28917), .b(n29299), .c(n28905), .o(n29679) );
no03f01 g25889 ( .a(n29679), .b(n29678), .c(n29348), .o(n29680) );
na03f01 g25890 ( .a(n29353), .b(n28903), .c(n28894), .o(n29681) );
na02f01 g25891 ( .a(n29354), .b(n29297), .o(n29682) );
in01f01 g25892 ( .a(n29359), .o(n29683) );
na03f01 g25893 ( .a(n29683), .b(n29682), .c(n29681), .o(n29684) );
ao12f01 g25894 ( .a(n29683), .b(n29682), .c(n29681), .o(n29685) );
no03f01 g25895 ( .a(n28893), .b(n29295), .c(n27681), .o(n29686) );
ao12f01 g25896 ( .a(n28888), .b(n29296), .c(n_27014), .o(n29687) );
no02f01 g25897 ( .a(n29687), .b(n29686), .o(n29688) );
in01f01 g25898 ( .a(n29381), .o(n29689) );
in01f01 g25899 ( .a(n29382), .o(n29690) );
ao12f01 g25900 ( .a(n29690), .b(n29689), .c(n29688), .o(n29691) );
oa12f01 g25901 ( .a(n29684), .b(n29691), .c(n29685), .o(n29692) );
oa12f01 g25902 ( .a(n29348), .b(n29679), .c(n29678), .o(n29693) );
ao12f01 g25903 ( .a(n29680), .b(n29693), .c(n29692), .o(n29694) );
oa12f01 g25904 ( .a(n29300), .b(n29338), .c(n28925), .o(n29695) );
na02f01 g25905 ( .a(n29339), .b(n28918), .o(n29696) );
in01f01 g25906 ( .a(n29344), .o(n29697) );
ao12f01 g25907 ( .a(n29697), .b(n29696), .c(n29695), .o(n29698) );
oa12f01 g25908 ( .a(n29677), .b(n29698), .c(n29694), .o(n29699) );
no03f01 g25909 ( .a(n29335), .b(n29331), .c(n29675), .o(n29700) );
oa12f01 g25910 ( .a(n29676), .b(n29700), .c(n29699), .o(n29701) );
ao12f01 g25911 ( .a(n29315), .b(n29312), .c(n28947), .o(n29702) );
no03f01 g25912 ( .a(n29309), .b(n29306), .c(n29304), .o(n29703) );
no03f01 g25913 ( .a(n29325), .b(n29703), .c(n29702), .o(n29704) );
in01f01 g25914 ( .a(n29394), .o(n29705) );
no03f01 g25915 ( .a(n29401), .b(n29395), .c(n29705), .o(n29706) );
no02f01 g25916 ( .a(n29706), .b(n29704), .o(n29707) );
oa12f01 g25917 ( .a(n29707), .b(n29403), .c(n29701), .o(n29708) );
oa12f01 g25918 ( .a(n29291), .b(n29286), .c(n29285), .o(n29709) );
na03f01 g25919 ( .a(n29709), .b(n29708), .c(n29674), .o(n29710) );
na03f01 g25920 ( .a(n29710), .b(n29673), .c(n29672), .o(n29711) );
in01f01 g25921 ( .a(n29416), .o(n29712) );
oa12f01 g25922 ( .a(n29266), .b(n29219), .c(n29217), .o(n29713) );
na03f01 g25923 ( .a(n29713), .b(n29712), .c(n29711), .o(n29714) );
na03f01 g25924 ( .a(n29212), .b(n29023), .c(n29014), .o(n29715) );
na03f01 g25925 ( .a(n29715), .b(n29714), .c(n29671), .o(n29716) );
in01f01 g25926 ( .a(n29483), .o(n29717) );
in01f01 g25927 ( .a(n29529), .o(n29718) );
na04f01 g25928 ( .a(n29718), .b(n29717), .c(n29716), .d(n29670), .o(n29719) );
in01f01 g25929 ( .a(n29533), .o(n29720) );
ao12f01 g25930 ( .a(n29576), .b(n29720), .c(n29719), .o(n29721) );
na02f01 g25931 ( .a(n29614), .b(n29721), .o(n29722) );
oa12f01 g25932 ( .a(n29651), .b(n29636), .c(n29722), .o(n29723) );
in01f01 g25933 ( .a(n29668), .o(n29724) );
na02f01 g25934 ( .a(n29724), .b(n29723), .o(n29725) );
na02f01 g25935 ( .a(n29725), .b(n29669), .o(n353) );
na03f01 g25936 ( .a(n27220), .b(n27022), .c(n27021), .o(n29727) );
oa12f01 g25937 ( .a(n27219), .b(n27023), .c(n27218), .o(n29728) );
na02f01 g25938 ( .a(n29728), .b(n29727), .o(n358) );
oa12f01 g25939 ( .a(n27627), .b(n27539), .c(n27495), .o(n29730) );
in01f01 g25940 ( .a(n29730), .o(n29731) );
no02f01 g25941 ( .a(n27548), .b(n27367), .o(n29732) );
no02f01 g25942 ( .a(n29732), .b(n27550), .o(n29733) );
na02f01 g25943 ( .a(n29733), .b(n29731), .o(n29734) );
in01f01 g25944 ( .a(n29733), .o(n29735) );
na02f01 g25945 ( .a(n29735), .b(n29730), .o(n29736) );
na02f01 g25946 ( .a(n29736), .b(n29734), .o(n363) );
no02f01 g25947 ( .a(n21065), .b(n18459), .o(n29738) );
ao12f01 g25948 ( .a(n18459), .b(n21092), .c(n21078), .o(n29739) );
no02f01 g25949 ( .a(n29739), .b(n29738), .o(n29740) );
na02f01 g25950 ( .a(n21047), .b(n18460), .o(n29741) );
na02f01 g25951 ( .a(n21047), .b(n18459), .o(n29742) );
oa12f01 g25952 ( .a(n18459), .b(n21064), .c(n21062), .o(n29743) );
na02f01 g25953 ( .a(n29743), .b(n29742), .o(n29744) );
ao12f01 g25954 ( .a(n29744), .b(n29741), .c(n29740), .o(n29745) );
in01f01 g25955 ( .a(n29745), .o(n29746) );
no02f01 g25956 ( .a(n21225), .b(n18460), .o(n29747) );
no02f01 g25957 ( .a(n21225), .b(n18459), .o(n29748) );
no03f01 g25958 ( .a(n29748), .b(n29747), .c(n29746), .o(n29749) );
no02f01 g25959 ( .a(n29748), .b(n29747), .o(n29750) );
no02f01 g25960 ( .a(n29750), .b(n29745), .o(n29751) );
no02f01 g25961 ( .a(n29751), .b(n29749), .o(n29752) );
no04f01 g25962 ( .a(n20052), .b(n19787), .c(n19778), .d(n19776), .o(n29753) );
ao22f01 g25963 ( .a(n19828), .b(n19788), .c(n20046), .d(n20045), .o(n29754) );
no02f01 g25964 ( .a(n29754), .b(n29753), .o(n29755) );
no02f01 g25965 ( .a(n29755), .b(n29752), .o(n29756) );
in01f01 g25966 ( .a(n29756), .o(n29757) );
in01f01 g25967 ( .a(n29740), .o(n29758) );
in01f01 g25968 ( .a(n29741), .o(n29759) );
in01f01 g25969 ( .a(n29742), .o(n29760) );
no02f01 g25970 ( .a(n29760), .b(n29759), .o(n29761) );
no02f01 g25971 ( .a(n29761), .b(n29758), .o(n29762) );
na02f01 g25972 ( .a(n29761), .b(n29758), .o(n29763) );
in01f01 g25973 ( .a(n29763), .o(n29764) );
no02f01 g25974 ( .a(n29764), .b(n29762), .o(n29765) );
no02f01 g25975 ( .a(n19826), .b(n19801), .o(n29766) );
no02f01 g25976 ( .a(n20051), .b(n19787), .o(n29767) );
no02f01 g25977 ( .a(n29767), .b(n29766), .o(n29768) );
na02f01 g25978 ( .a(n29767), .b(n29766), .o(n29769) );
in01f01 g25979 ( .a(n29769), .o(n29770) );
no02f01 g25980 ( .a(n29770), .b(n29768), .o(n29771) );
no02f01 g25981 ( .a(n29771), .b(n29765), .o(n29772) );
in01f01 g25982 ( .a(n29738), .o(n29773) );
na03f01 g25983 ( .a(n29743), .b(n29739), .c(n29773), .o(n29774) );
in01f01 g25984 ( .a(n29739), .o(n29775) );
in01f01 g25985 ( .a(n29743), .o(n29776) );
oa12f01 g25986 ( .a(n29775), .b(n29776), .c(n29738), .o(n29777) );
na02f01 g25987 ( .a(n29777), .b(n29774), .o(n29778) );
no02f01 g25988 ( .a(n20049), .b(n19817), .o(n29779) );
no02f01 g25989 ( .a(n19802), .b(n19801), .o(n29780) );
no02f01 g25990 ( .a(n29780), .b(n29779), .o(n29781) );
na02f01 g25991 ( .a(n29780), .b(n29779), .o(n29782) );
in01f01 g25992 ( .a(n29782), .o(n29783) );
no02f01 g25993 ( .a(n29783), .b(n29781), .o(n29784) );
in01f01 g25994 ( .a(n29784), .o(n29785) );
na02f01 g25995 ( .a(n29785), .b(n29778), .o(n29786) );
no03f01 g25996 ( .a(n21092), .b(n21079), .c(n18459), .o(n29787) );
in01f01 g25997 ( .a(n21092), .o(n29788) );
ao12f01 g25998 ( .a(n21078), .b(n29788), .c(n18460), .o(n29789) );
no02f01 g25999 ( .a(n29789), .b(n29787), .o(n29790) );
no02f01 g26000 ( .a(n19824), .b(n19819), .o(n29791) );
no02f01 g26001 ( .a(n20048), .b(n19816), .o(n29792) );
no02f01 g26002 ( .a(n29792), .b(n29791), .o(n29793) );
no02f01 g26003 ( .a(n29793), .b(n19807), .o(n29794) );
na02f01 g26004 ( .a(n29793), .b(n19807), .o(n29795) );
in01f01 g26005 ( .a(n29795), .o(n29796) );
no02f01 g26006 ( .a(n29796), .b(n29794), .o(n29797) );
na02f01 g26007 ( .a(n29797), .b(n29790), .o(n29798) );
na02f01 g26008 ( .a(n21092), .b(n18459), .o(n29799) );
no02f01 g26009 ( .a(n29788), .b(n18459), .o(n29800) );
in01f01 g26010 ( .a(n29800), .o(n29801) );
na02f01 g26011 ( .a(n29801), .b(n29799), .o(n29802) );
no02f01 g26012 ( .a(n19805), .b(n18919), .o(n29803) );
na02f01 g26013 ( .a(n19805), .b(n18919), .o(n29804) );
in01f01 g26014 ( .a(n29804), .o(n29805) );
no02f01 g26015 ( .a(n29805), .b(n29803), .o(n29806) );
no02f01 g26016 ( .a(n29806), .b(n29802), .o(n29807) );
no02f01 g26017 ( .a(n29797), .b(n29790), .o(n29808) );
ao12f01 g26018 ( .a(n29808), .b(n29807), .c(n29798), .o(n29809) );
no02f01 g26019 ( .a(n29785), .b(n29778), .o(n29810) );
oa12f01 g26020 ( .a(n29786), .b(n29810), .c(n29809), .o(n29811) );
na02f01 g26021 ( .a(n29771), .b(n29765), .o(n29812) );
ao12f01 g26022 ( .a(n29772), .b(n29812), .c(n29811), .o(n29813) );
na02f01 g26023 ( .a(n29755), .b(n29752), .o(n29814) );
in01f01 g26024 ( .a(n29814), .o(n29815) );
oa12f01 g26025 ( .a(n29757), .b(n29815), .c(n29813), .o(n29816) );
no02f01 g26026 ( .a(n29748), .b(n29745), .o(n29817) );
no02f01 g26027 ( .a(n29817), .b(n29747), .o(n29818) );
na02f01 g26028 ( .a(n21033), .b(n18459), .o(n29819) );
na02f01 g26029 ( .a(n21033), .b(n18460), .o(n29820) );
ao12f01 g26030 ( .a(n29818), .b(n29820), .c(n29819), .o(n29821) );
na03f01 g26031 ( .a(n29820), .b(n29819), .c(n29818), .o(n29822) );
in01f01 g26032 ( .a(n29822), .o(n29823) );
no02f01 g26033 ( .a(n29823), .b(n29821), .o(n29824) );
no04f01 g26034 ( .a(n20054), .b(n19829), .c(n19776), .d(n19763), .o(n29825) );
ao22f01 g26035 ( .a(n19830), .b(n19764), .c(n20053), .d(n20045), .o(n29826) );
no02f01 g26036 ( .a(n29826), .b(n29825), .o(n29827) );
no02f01 g26037 ( .a(n29827), .b(n29824), .o(n29828) );
na02f01 g26038 ( .a(n29827), .b(n29824), .o(n29829) );
in01f01 g26039 ( .a(n29829), .o(n29830) );
oa12f01 g26040 ( .a(n29816), .b(n29830), .c(n29828), .o(n29831) );
in01f01 g26041 ( .a(n29816), .o(n29832) );
in01f01 g26042 ( .a(n29828), .o(n29833) );
na03f01 g26043 ( .a(n29829), .b(n29833), .c(n29832), .o(n29834) );
na02f01 g26044 ( .a(n29834), .b(n29831), .o(n368) );
no02f01 g26045 ( .a(n27064), .b(n27060), .o(n29836) );
na02f01 g26046 ( .a(n29836), .b(n27045), .o(n29837) );
in01f01 g26047 ( .a(n29836), .o(n29838) );
na02f01 g26048 ( .a(n29838), .b(n27236), .o(n29839) );
na02f01 g26049 ( .a(n29839), .b(n29837), .o(n373) );
ao12f01 g26050 ( .a(n9228), .b(n9591), .c(n9231), .o(n29841) );
no02f01 g26051 ( .a(n29841), .b(n9591), .o(n29842) );
no03f01 g26052 ( .a(n4201), .b(n9231), .c(n9228), .o(n29843) );
no02f01 g26053 ( .a(n29843), .b(n29842), .o(n29844) );
na03f01 g26054 ( .a(n29844), .b(n9590), .c(n9589), .o(n29845) );
in01f01 g26055 ( .a(n29844), .o(n4098) );
oa12f01 g26056 ( .a(n4098), .b(n9646), .c(n9645), .o(n29847) );
na02f01 g26057 ( .a(n29847), .b(n29845), .o(n378) );
no03f01 g26058 ( .a(n18375), .b(n18373), .c(n18364), .o(n29849) );
na02f01 g26059 ( .a(n18367), .b(n18144), .o(n29850) );
no02f01 g26060 ( .a(n29850), .b(n29849), .o(n29851) );
no02f01 g26061 ( .a(n18147), .b(n18114), .o(n29852) );
no02f01 g26062 ( .a(n29852), .b(n29851), .o(n29853) );
na02f01 g26063 ( .a(n29852), .b(n29851), .o(n29854) );
in01f01 g26064 ( .a(n29854), .o(n29855) );
no03f01 g26065 ( .a(n29855), .b(n29853), .c(n18459), .o(n29856) );
in01f01 g26066 ( .a(n25662), .o(n29857) );
oa12f01 g26067 ( .a(n29857), .b(n25663), .c(n25652), .o(n29858) );
no02f01 g26068 ( .a(n29855), .b(n29853), .o(n29859) );
no02f01 g26069 ( .a(n29859), .b(n18460), .o(n29860) );
in01f01 g26070 ( .a(n29860), .o(n29861) );
ao12f01 g26071 ( .a(n29856), .b(n29861), .c(n29858), .o(n29862) );
in01f01 g26072 ( .a(n29862), .o(n29863) );
no02f01 g26073 ( .a(n18378), .b(n18149), .o(n29864) );
in01f01 g26074 ( .a(n29864), .o(n29865) );
no02f01 g26075 ( .a(n18451), .b(n18145), .o(n29866) );
no02f01 g26076 ( .a(n29866), .b(n18393), .o(n29867) );
in01f01 g26077 ( .a(n29867), .o(n29868) );
no02f01 g26078 ( .a(n29868), .b(n29865), .o(n29869) );
no02f01 g26079 ( .a(n29867), .b(n29864), .o(n29870) );
no02f01 g26080 ( .a(n29870), .b(n29869), .o(n29871) );
in01f01 g26081 ( .a(n29871), .o(n29872) );
no02f01 g26082 ( .a(n29872), .b(n18459), .o(n29873) );
no02f01 g26083 ( .a(n29871), .b(n18460), .o(n29874) );
no02f01 g26084 ( .a(n29874), .b(n29873), .o(n29875) );
na02f01 g26085 ( .a(n29875), .b(n29863), .o(n29876) );
in01f01 g26086 ( .a(n29875), .o(n29877) );
na02f01 g26087 ( .a(n29877), .b(n29862), .o(n29878) );
na02f01 g26088 ( .a(n29878), .b(n29876), .o(n383) );
no02f01 g26089 ( .a(n6932), .b(n6934), .o(n29880) );
no02f01 g26090 ( .a(n6933), .b(n5001), .o(n29881) );
no02f01 g26091 ( .a(n29881), .b(n29880), .o(n29882) );
na03f01 g26092 ( .a(n29882), .b(n6936), .c(n6923), .o(n29883) );
oa22f01 g26093 ( .a(n29881), .b(n29880), .c(n6935), .d(n6924), .o(n29884) );
na02f01 g26094 ( .a(n29884), .b(n29883), .o(n388) );
no02f01 g26095 ( .a(n24660), .b(n23151), .o(n29886) );
no02f01 g26096 ( .a(n24661), .b(n23150), .o(n29887) );
no02f01 g26097 ( .a(n29887), .b(n29886), .o(n29888) );
in01f01 g26098 ( .a(n29888), .o(n29889) );
ao12f01 g26099 ( .a(n24661), .b(n24945), .c(n23159), .o(n29890) );
in01f01 g26100 ( .a(n24664), .o(n29891) );
no03f01 g26101 ( .a(n24950), .b(n24940), .c(n24934), .o(n29892) );
oa12f01 g26102 ( .a(n24944), .b(n29892), .c(n29891), .o(n29893) );
in01f01 g26103 ( .a(n29893), .o(n29894) );
no03f01 g26104 ( .a(n29894), .b(n29890), .c(n29889), .o(n29895) );
in01f01 g26105 ( .a(n29890), .o(n29896) );
ao12f01 g26106 ( .a(n29888), .b(n29893), .c(n29896), .o(n29897) );
no02f01 g26107 ( .a(n29897), .b(n29895), .o(n29898) );
no02f01 g26108 ( .a(n29898), .b(n5529), .o(n29899) );
no02f01 g26109 ( .a(n25044), .b(n5527), .o(n29900) );
oa12f01 g26110 ( .a(n25177), .b(n25164), .c(n24663), .o(n29901) );
na03f01 g26111 ( .a(n25175), .b(n25174), .c(n25172), .o(n29902) );
ao12f01 g26112 ( .a(n5527), .b(n29902), .c(n29901), .o(n29903) );
no02f01 g26113 ( .a(n25157), .b(n5527), .o(n29904) );
oa12f01 g26114 ( .a(n5529), .b(n25144), .c(n25051), .o(n29905) );
oa12f01 g26115 ( .a(n25759), .b(n25217), .c(n5527), .o(n29906) );
ao12f01 g26116 ( .a(n25763), .b(n25293), .c(n5527), .o(n29907) );
ao22f01 g26117 ( .a(n29907), .b(n29906), .c(n25290), .d(n5529), .o(n29908) );
na02f01 g26118 ( .a(n29908), .b(n29905), .o(n29909) );
no03f01 g26119 ( .a(n29909), .b(n29904), .c(n29903), .o(n29910) );
ao12f01 g26120 ( .a(n5529), .b(n25541), .c(n25540), .o(n29911) );
oa12f01 g26121 ( .a(n5527), .b(n25144), .c(n25051), .o(n29912) );
na02f01 g26122 ( .a(n29912), .b(n25670), .o(n29913) );
ao12f01 g26123 ( .a(n5529), .b(n29902), .c(n29901), .o(n29914) );
no04f01 g26124 ( .a(n29914), .b(n29913), .c(n29911), .d(n29910), .o(n29915) );
in01f01 g26125 ( .a(n25169), .o(n29916) );
no02f01 g26126 ( .a(n29916), .b(n25167), .o(n29917) );
no02f01 g26127 ( .a(n29917), .b(n5527), .o(n29918) );
no02f01 g26128 ( .a(n29918), .b(n29915), .o(n29919) );
na02f01 g26129 ( .a(n25034), .b(n5529), .o(n29920) );
na02f01 g26130 ( .a(n29920), .b(n29919), .o(n29921) );
no02f01 g26131 ( .a(n29921), .b(n29900), .o(n29922) );
no02f01 g26132 ( .a(n24956), .b(n5527), .o(n29923) );
in01f01 g26133 ( .a(n29923), .o(n29924) );
no02f01 g26134 ( .a(n29917), .b(n5529), .o(n29925) );
in01f01 g26135 ( .a(n29925), .o(n29926) );
na02f01 g26136 ( .a(n25034), .b(n5527), .o(n29927) );
na02f01 g26137 ( .a(n29927), .b(n29926), .o(n29928) );
no02f01 g26138 ( .a(n25044), .b(n5529), .o(n29929) );
no02f01 g26139 ( .a(n29929), .b(n29928), .o(n29930) );
no02f01 g26140 ( .a(n24956), .b(n5529), .o(n29931) );
in01f01 g26141 ( .a(n29931), .o(n29932) );
na02f01 g26142 ( .a(n29932), .b(n29930), .o(n29933) );
ao12f01 g26143 ( .a(n29933), .b(n29924), .c(n29922), .o(n29934) );
no02f01 g26144 ( .a(n29898), .b(n5527), .o(n29935) );
in01f01 g26145 ( .a(n29935), .o(n29936) );
ao12f01 g26146 ( .a(n29899), .b(n29936), .c(n29934), .o(n29937) );
in01f01 g26147 ( .a(n29937), .o(n29938) );
no02f01 g26148 ( .a(n29938), .b(n24592), .o(n29939) );
no02f01 g26149 ( .a(n29937), .b(n24602), .o(n29940) );
no02f01 g26150 ( .a(n29940), .b(n29939), .o(n29941) );
no02f01 g26151 ( .a(n24547), .b(n24405), .o(n29942) );
no02f01 g26152 ( .a(n29942), .b(n29938), .o(n29943) );
in01f01 g26153 ( .a(n29943), .o(n29944) );
ao12f01 g26154 ( .a(n29937), .b(n24547), .c(n24405), .o(n29945) );
in01f01 g26155 ( .a(n29945), .o(n29946) );
oa12f01 g26156 ( .a(n29930), .b(n29921), .c(n29900), .o(n29947) );
no02f01 g26157 ( .a(n29931), .b(n29923), .o(n29948) );
in01f01 g26158 ( .a(n29948), .o(n29949) );
na02f01 g26159 ( .a(n29949), .b(n29947), .o(n29950) );
no02f01 g26160 ( .a(n29949), .b(n29947), .o(n29951) );
in01f01 g26161 ( .a(n29951), .o(n29952) );
na02f01 g26162 ( .a(n29952), .b(n29950), .o(n29953) );
na02f01 g26163 ( .a(n29953), .b(n24983), .o(n29954) );
no02f01 g26164 ( .a(n29929), .b(n29900), .o(n29955) );
ao12f01 g26165 ( .a(n29928), .b(n29920), .c(n29919), .o(n29956) );
no02f01 g26166 ( .a(n29956), .b(n29955), .o(n29957) );
na02f01 g26167 ( .a(n29956), .b(n29955), .o(n29958) );
in01f01 g26168 ( .a(n29958), .o(n29959) );
oa12f01 g26169 ( .a(n24978), .b(n29959), .c(n29957), .o(n29960) );
in01f01 g26170 ( .a(n29960), .o(n29961) );
in01f01 g26171 ( .a(n24431), .o(n29962) );
na02f01 g26172 ( .a(n29927), .b(n29920), .o(n29963) );
oa12f01 g26173 ( .a(n29963), .b(n29925), .c(n29919), .o(n29964) );
in01f01 g26174 ( .a(n29964), .o(n29965) );
no03f01 g26175 ( .a(n29963), .b(n29925), .c(n29919), .o(n29966) );
no03f01 g26176 ( .a(n29966), .b(n29965), .c(n29962), .o(n29967) );
oa12f01 g26177 ( .a(n5529), .b(n25178), .c(n25176), .o(n29968) );
na02f01 g26178 ( .a(n25542), .b(n5529), .o(n29969) );
na03f01 g26179 ( .a(n25143), .b(n25142), .c(n25138), .o(n29970) );
oa12f01 g26180 ( .a(n25050), .b(n24932), .c(n24923), .o(n29971) );
ao12f01 g26181 ( .a(n5527), .b(n29971), .c(n29970), .o(n29972) );
oa22f01 g26182 ( .a(n25712), .b(n25707), .c(n25212), .d(n5527), .o(n29973) );
no02f01 g26183 ( .a(n29973), .b(n29972), .o(n29974) );
na03f01 g26184 ( .a(n29974), .b(n29969), .c(n29968), .o(n29975) );
oa12f01 g26185 ( .a(n5527), .b(n25156), .c(n25152), .o(n29976) );
ao12f01 g26186 ( .a(n5529), .b(n29971), .c(n29970), .o(n29977) );
no02f01 g26187 ( .a(n29977), .b(n25716), .o(n29978) );
oa12f01 g26188 ( .a(n5527), .b(n25178), .c(n25176), .o(n29979) );
na04f01 g26189 ( .a(n29979), .b(n29978), .c(n29976), .d(n29975), .o(n29980) );
oa12f01 g26190 ( .a(n29980), .b(n29925), .c(n29918), .o(n29981) );
na02f01 g26191 ( .a(n25170), .b(n5529), .o(n29982) );
na03f01 g26192 ( .a(n29926), .b(n29982), .c(n29915), .o(n29983) );
ao12f01 g26193 ( .a(n24969), .b(n29983), .c(n29981), .o(n29984) );
na02f01 g26194 ( .a(n29979), .b(n29968), .o(n29985) );
na03f01 g26195 ( .a(n29978), .b(n29976), .c(n29909), .o(n29986) );
ao12f01 g26196 ( .a(n29985), .b(n29986), .c(n29969), .o(n29987) );
no02f01 g26197 ( .a(n29914), .b(n29903), .o(n29988) );
no03f01 g26198 ( .a(n29913), .b(n29911), .c(n29974), .o(n29989) );
no03f01 g26199 ( .a(n29989), .b(n29988), .c(n29904), .o(n29990) );
no03f01 g26200 ( .a(n29990), .b(n29987), .c(n24490), .o(n29991) );
ao22f01 g26201 ( .a(n29912), .b(n29905), .c(n29973), .d(n25670), .o(n29992) );
no04f01 g26202 ( .a(n29977), .b(n29908), .c(n29972), .d(n25716), .o(n29993) );
no03f01 g26203 ( .a(n29993), .b(n29992), .c(n25454), .o(n29994) );
in01f01 g26204 ( .a(n29994), .o(n29995) );
oa22f01 g26205 ( .a(n29977), .b(n29972), .c(n29908), .d(n25716), .o(n29996) );
na04f01 g26206 ( .a(n29912), .b(n29973), .c(n29905), .d(n25670), .o(n29997) );
ao12f01 g26207 ( .a(n24474), .b(n29997), .c(n29996), .o(n29998) );
no02f01 g26208 ( .a(n29998), .b(n25720), .o(n29999) );
oa12f01 g26209 ( .a(n29999), .b(n25922), .c(n25723), .o(n30000) );
na02f01 g26210 ( .a(n29978), .b(n29909), .o(n30001) );
oa12f01 g26211 ( .a(n30001), .b(n29911), .c(n29904), .o(n30002) );
no02f01 g26212 ( .a(n29913), .b(n29974), .o(n30003) );
na03f01 g26213 ( .a(n30003), .b(n29976), .c(n29969), .o(n30004) );
na03f01 g26214 ( .a(n30004), .b(n30002), .c(n25408), .o(n30005) );
na03f01 g26215 ( .a(n30005), .b(n30000), .c(n29995), .o(n30006) );
oa12f01 g26216 ( .a(n29988), .b(n29989), .c(n29904), .o(n30007) );
na03f01 g26217 ( .a(n29986), .b(n29985), .c(n29969), .o(n30008) );
ao12f01 g26218 ( .a(n24442), .b(n30008), .c(n30007), .o(n30009) );
ao12f01 g26219 ( .a(n25408), .b(n30004), .c(n30002), .o(n30010) );
no02f01 g26220 ( .a(n30010), .b(n30009), .o(n30011) );
ao12f01 g26221 ( .a(n29991), .b(n30011), .c(n30006), .o(n30012) );
na03f01 g26222 ( .a(n29983), .b(n29981), .c(n24969), .o(n30013) );
ao12f01 g26223 ( .a(n29984), .b(n30013), .c(n30012), .o(n30014) );
oa12f01 g26224 ( .a(n29962), .b(n29966), .c(n29965), .o(n30015) );
ao12f01 g26225 ( .a(n29967), .b(n30015), .c(n30014), .o(n30016) );
in01f01 g26226 ( .a(n29957), .o(n30017) );
na03f01 g26227 ( .a(n29958), .b(n30017), .c(n24427), .o(n30018) );
ao12f01 g26228 ( .a(n29961), .b(n30018), .c(n30016), .o(n30019) );
no02f01 g26229 ( .a(n29953), .b(n24983), .o(n30020) );
oa12f01 g26230 ( .a(n29954), .b(n30020), .c(n30019), .o(n30021) );
no02f01 g26231 ( .a(n29935), .b(n29899), .o(n30022) );
na02f01 g26232 ( .a(n30022), .b(n29934), .o(n30023) );
no02f01 g26233 ( .a(n30022), .b(n29934), .o(n30024) );
in01f01 g26234 ( .a(n30024), .o(n30025) );
na02f01 g26235 ( .a(n30025), .b(n30023), .o(n30026) );
no02f01 g26236 ( .a(n30026), .b(n24419), .o(n30027) );
in01f01 g26237 ( .a(n30027), .o(n30028) );
no02f01 g26238 ( .a(n24514), .b(n24513), .o(n30029) );
in01f01 g26239 ( .a(n30029), .o(n30030) );
no02f01 g26240 ( .a(n29938), .b(n30030), .o(n30031) );
in01f01 g26241 ( .a(n30031), .o(n30032) );
na03f01 g26242 ( .a(n30032), .b(n30028), .c(n30021), .o(n30033) );
no02f01 g26243 ( .a(n29937), .b(n30029), .o(n30034) );
ao12f01 g26244 ( .a(n24518), .b(n30025), .c(n30023), .o(n30035) );
oa12f01 g26245 ( .a(n30032), .b(n30035), .c(n30034), .o(n30036) );
na03f01 g26246 ( .a(n30036), .b(n30033), .c(n29946), .o(n30037) );
no02f01 g26247 ( .a(n29938), .b(n25016), .o(n30038) );
ao12f01 g26248 ( .a(n29938), .b(n24538), .c(n25005), .o(n30039) );
no02f01 g26249 ( .a(n29938), .b(n25003), .o(n30040) );
no03f01 g26250 ( .a(n30040), .b(n30039), .c(n30038), .o(n30041) );
na03f01 g26251 ( .a(n30041), .b(n30037), .c(n29944), .o(n30042) );
ao12f01 g26252 ( .a(n29937), .b(n24543), .c(n24563), .o(n30043) );
no02f01 g26253 ( .a(n29937), .b(n24561), .o(n30044) );
no02f01 g26254 ( .a(n30044), .b(n30043), .o(n30045) );
ao12f01 g26255 ( .a(n29937), .b(n30045), .c(n24598), .o(n30046) );
in01f01 g26256 ( .a(n30046), .o(n30047) );
na03f01 g26257 ( .a(n30047), .b(n30042), .c(n29941), .o(n30048) );
in01f01 g26258 ( .a(n29941), .o(n30049) );
in01f01 g26259 ( .a(n29950), .o(n30050) );
no02f01 g26260 ( .a(n29951), .b(n30050), .o(n30051) );
no02f01 g26261 ( .a(n30051), .b(n24504), .o(n30052) );
in01f01 g26262 ( .a(n29966), .o(n30053) );
na03f01 g26263 ( .a(n30053), .b(n29964), .c(n24431), .o(n30054) );
ao12f01 g26264 ( .a(n29915), .b(n29926), .c(n29982), .o(n30055) );
no03f01 g26265 ( .a(n29925), .b(n29918), .c(n29980), .o(n30056) );
oa12f01 g26266 ( .a(n24485), .b(n30056), .c(n30055), .o(n30057) );
in01f01 g26267 ( .a(n29991), .o(n30058) );
in01f01 g26268 ( .a(n25723), .o(n30059) );
na02f01 g26269 ( .a(n25764), .b(n25769), .o(n30060) );
na02f01 g26270 ( .a(n25765), .b(n25727), .o(n30061) );
na02f01 g26271 ( .a(n30061), .b(n30060), .o(n30062) );
na02f01 g26272 ( .a(n30062), .b(n24465), .o(n30063) );
in01f01 g26273 ( .a(n25777), .o(n30064) );
na02f01 g26274 ( .a(n25778), .b(n30064), .o(n30065) );
na03f01 g26275 ( .a(n25698), .b(n25798), .c(n25673), .o(n30066) );
na02f01 g26276 ( .a(n25796), .b(n25795), .o(n30067) );
na02f01 g26277 ( .a(n30067), .b(n30066), .o(n30068) );
oa22f01 g26278 ( .a(n25745), .b(n25691), .c(n25744), .d(n25741), .o(n30069) );
na04f01 g26279 ( .a(n25694), .b(n25693), .c(n25742), .d(n25688), .o(n30070) );
ao12f01 g26280 ( .a(n25807), .b(n30070), .c(n30069), .o(n30071) );
na03f01 g26281 ( .a(n25807), .b(n30070), .c(n30069), .o(n30072) );
no04f01 g26282 ( .a(n25744), .b(n25740), .c(n25686), .d(n25683), .o(n30073) );
ao22f01 g26283 ( .a(n25693), .b(n25687), .c(n25737), .d(n25734), .o(n30074) );
in01f01 g26284 ( .a(n25817), .o(n30075) );
oa12f01 g26285 ( .a(n30075), .b(n30074), .c(n30073), .o(n30076) );
ao12f01 g26286 ( .a(n25682), .b(n25685), .c(n25733), .o(n30077) );
no03f01 g26287 ( .a(n25736), .b(n25681), .c(n25680), .o(n30078) );
in01f01 g26288 ( .a(n25825), .o(n30079) );
oa12f01 g26289 ( .a(n30079), .b(n30078), .c(n30077), .o(n30080) );
no03f01 g26290 ( .a(n30079), .b(n30078), .c(n30077), .o(n30081) );
oa12f01 g26291 ( .a(n30080), .b(n25850), .c(n30081), .o(n30082) );
na03f01 g26292 ( .a(n25855), .b(n25684), .c(n25732), .o(n30083) );
oa12f01 g26293 ( .a(n25853), .b(n25735), .c(n25677), .o(n30084) );
na03f01 g26294 ( .a(n25859), .b(n30084), .c(n30083), .o(n30085) );
ao12f01 g26295 ( .a(n25859), .b(n30084), .c(n30083), .o(n30086) );
ao12f01 g26296 ( .a(n30086), .b(n30085), .c(n30082), .o(n30087) );
no03f01 g26297 ( .a(n30075), .b(n30074), .c(n30073), .o(n30088) );
oa12f01 g26298 ( .a(n30076), .b(n30088), .c(n30087), .o(n30089) );
ao12f01 g26299 ( .a(n30071), .b(n30089), .c(n30072), .o(n30090) );
no03f01 g26300 ( .a(n25889), .b(n25888), .c(n25887), .o(n30091) );
no02f01 g26301 ( .a(n30091), .b(n30090), .o(n30092) );
na02f01 g26302 ( .a(n25883), .b(n25890), .o(n30093) );
oa12f01 g26303 ( .a(n30068), .b(n30093), .c(n30092), .o(n30094) );
oa12f01 g26304 ( .a(n25884), .b(n25874), .c(n30092), .o(n30095) );
no02f01 g26305 ( .a(n25785), .b(n25784), .o(n30096) );
no02f01 g26306 ( .a(n25782), .b(n25781), .o(n30097) );
in01f01 g26307 ( .a(n25792), .o(n30098) );
no03f01 g26308 ( .a(n30098), .b(n30097), .c(n30096), .o(n30099) );
ao12f01 g26309 ( .a(n30099), .b(n30095), .c(n30094), .o(n30100) );
na03f01 g26310 ( .a(n25905), .b(n25910), .c(n25909), .o(n30101) );
oa12f01 g26311 ( .a(n30101), .b(n30100), .c(n25793), .o(n30102) );
in01f01 g26312 ( .a(n25911), .o(n30103) );
na03f01 g26313 ( .a(n25916), .b(n30103), .c(n30102), .o(n30104) );
ao12f01 g26314 ( .a(n25916), .b(n30103), .c(n30102), .o(n30105) );
ao12f01 g26315 ( .a(n30105), .b(n30104), .c(n30065), .o(n30106) );
no02f01 g26316 ( .a(n30062), .b(n24465), .o(n30107) );
oa12f01 g26317 ( .a(n30063), .b(n30107), .c(n30106), .o(n30108) );
oa12f01 g26318 ( .a(n24456), .b(n25722), .c(n25721), .o(n30109) );
oa12f01 g26319 ( .a(n25454), .b(n29993), .c(n29992), .o(n30110) );
na02f01 g26320 ( .a(n30110), .b(n30109), .o(n30111) );
ao12f01 g26321 ( .a(n30111), .b(n30108), .c(n30059), .o(n30112) );
ao12f01 g26322 ( .a(n30003), .b(n29976), .c(n29969), .o(n30113) );
no03f01 g26323 ( .a(n30001), .b(n29911), .c(n29904), .o(n30114) );
no03f01 g26324 ( .a(n30114), .b(n30113), .c(n24448), .o(n30115) );
no03f01 g26325 ( .a(n30115), .b(n30112), .c(n29994), .o(n30116) );
oa12f01 g26326 ( .a(n24490), .b(n29990), .c(n29987), .o(n30117) );
in01f01 g26327 ( .a(n30010), .o(n30118) );
na02f01 g26328 ( .a(n30118), .b(n30117), .o(n30119) );
oa12f01 g26329 ( .a(n30058), .b(n30119), .c(n30116), .o(n30120) );
no03f01 g26330 ( .a(n30056), .b(n30055), .c(n24485), .o(n30121) );
oa12f01 g26331 ( .a(n30057), .b(n30121), .c(n30120), .o(n30122) );
ao12f01 g26332 ( .a(n24431), .b(n30053), .c(n29964), .o(n30123) );
oa12f01 g26333 ( .a(n30054), .b(n30123), .c(n30122), .o(n30124) );
no03f01 g26334 ( .a(n29959), .b(n29957), .c(n24978), .o(n30125) );
oa12f01 g26335 ( .a(n29960), .b(n30125), .c(n30124), .o(n30126) );
na02f01 g26336 ( .a(n30051), .b(n24504), .o(n30127) );
ao12f01 g26337 ( .a(n30052), .b(n30127), .c(n30126), .o(n30128) );
no03f01 g26338 ( .a(n30031), .b(n30027), .c(n30128), .o(n30129) );
no02f01 g26339 ( .a(n30035), .b(n30034), .o(n30130) );
no02f01 g26340 ( .a(n30130), .b(n30031), .o(n30131) );
no03f01 g26341 ( .a(n30131), .b(n30129), .c(n29945), .o(n30132) );
in01f01 g26342 ( .a(n30041), .o(n30133) );
no03f01 g26343 ( .a(n30133), .b(n30132), .c(n29943), .o(n30134) );
oa12f01 g26344 ( .a(n30049), .b(n30046), .c(n30134), .o(n30135) );
na03f01 g26345 ( .a(n30135), .b(n30048), .c(n6037), .o(n30136) );
na02f01 g26346 ( .a(n30135), .b(n30048), .o(n3782) );
na02f01 g26347 ( .a(n3782), .b(n5873), .o(n30138) );
na02f01 g26348 ( .a(n30138), .b(n30136), .o(n393) );
no02f01 g26349 ( .a(n11845), .b(n11839), .o(n30140) );
no02f01 g26350 ( .a(n11862), .b(n11854), .o(n30141) );
na02f01 g26351 ( .a(n30141), .b(n30140), .o(n30142) );
in01f01 g26352 ( .a(n30141), .o(n30143) );
oa12f01 g26353 ( .a(n30143), .b(n11845), .c(n11839), .o(n30144) );
na02f01 g26354 ( .a(n30144), .b(n30142), .o(n398) );
in01f01 g26355 ( .a(n_44061), .o(n30146) );
no02f01 g26356 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_0_), .b(n30146), .o(n30147) );
no02f01 g26357 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_1_), .b(n30146), .o(n30148) );
no02f01 g26358 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_2_), .b(n30146), .o(n30149) );
no03f01 g26359 ( .a(n30149), .b(n30148), .c(n30147), .o(n30150) );
no02f01 g26360 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_3_), .b(n30146), .o(n30151) );
in01f01 g26361 ( .a(n30151), .o(n30152) );
na02f01 g26362 ( .a(n30152), .b(n30150), .o(n30153) );
no02f01 g26363 ( .a(n30146), .b(delay_xor_ln21_unr15_stage6_stallmux_q_5_), .o(n30154) );
no02f01 g26364 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_4_), .b(n30146), .o(n30155) );
no02f01 g26365 ( .a(n30155), .b(n30154), .o(n30156) );
in01f01 g26366 ( .a(n30156), .o(n30157) );
no02f01 g26367 ( .a(n30157), .b(n30153), .o(n30158) );
no02f01 g26368 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_6_), .b(n30146), .o(n30159) );
no02f01 g26369 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_7_), .b(n30146), .o(n30160) );
no02f01 g26370 ( .a(n30146), .b(delay_xor_ln21_unr15_stage6_stallmux_q_8_), .o(n30161) );
no03f01 g26371 ( .a(n30161), .b(n30160), .c(n30159), .o(n30162) );
na02f01 g26372 ( .a(n30162), .b(n30158), .o(n30163) );
no02f01 g26373 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_9_), .b(n30146), .o(n30164) );
no02f01 g26374 ( .a(n30164), .b(n30163), .o(n30165) );
no02f01 g26375 ( .a(n30146), .b(delay_xor_ln21_unr15_stage6_stallmux_q_12_), .o(n30166) );
no02f01 g26376 ( .a(n30146), .b(delay_xor_ln21_unr15_stage6_stallmux_q_10_), .o(n30167) );
no02f01 g26377 ( .a(n30146), .b(delay_xor_ln21_unr15_stage6_stallmux_q_11_), .o(n30168) );
no03f01 g26378 ( .a(n30168), .b(n30167), .c(n30166), .o(n30169) );
na02f01 g26379 ( .a(n30169), .b(n30165), .o(n30170) );
no02f01 g26380 ( .a(n30146), .b(delay_xor_ln21_unr15_stage6_stallmux_q_15_), .o(n30171) );
no02f01 g26381 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_13_), .b(n30146), .o(n30172) );
no02f01 g26382 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_14_), .b(n30146), .o(n30173) );
no02f01 g26383 ( .a(n30173), .b(n30172), .o(n30174) );
in01f01 g26384 ( .a(n30174), .o(n30175) );
no03f01 g26385 ( .a(n30175), .b(n30171), .c(n30170), .o(n30176) );
in01f01 g26386 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_16_), .o(n30177) );
no02f01 g26387 ( .a(n30177), .b(n_44061), .o(n30178) );
in01f01 g26388 ( .a(n30178), .o(n30179) );
no02f01 g26389 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_16_), .b(n30146), .o(n30180) );
ao12f01 g26390 ( .a(n30180), .b(n30179), .c(n30176), .o(n30181) );
in01f01 g26391 ( .a(n30181), .o(n30182) );
no02f01 g26392 ( .a(n30182), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_27_), .o(n30183) );
in01f01 g26393 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_27_), .o(n30184) );
no02f01 g26394 ( .a(n30181), .b(n30184), .o(n30185) );
no02f01 g26395 ( .a(n30185), .b(n30183), .o(n30186) );
no02f01 g26396 ( .a(n30182), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_26_), .o(n30187) );
in01f01 g26397 ( .a(n30187), .o(n30188) );
no02f01 g26398 ( .a(n30182), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_23_), .o(n30189) );
in01f01 g26399 ( .a(n30189), .o(n30190) );
no02f01 g26400 ( .a(n30182), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_21_), .o(n30191) );
no02f01 g26401 ( .a(n30182), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_17_), .o(n30192) );
in01f01 g26402 ( .a(n30192), .o(n30193) );
in01f01 g26403 ( .a(n30170), .o(n30194) );
in01f01 g26404 ( .a(n30172), .o(n30195) );
na02f01 g26405 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_13_), .b(n30146), .o(n30196) );
na02f01 g26406 ( .a(n30196), .b(n30195), .o(n30197) );
no02f01 g26407 ( .a(n30197), .b(n30194), .o(n30198) );
na02f01 g26408 ( .a(n30197), .b(n30194), .o(n30199) );
in01f01 g26409 ( .a(n30199), .o(n30200) );
no02f01 g26410 ( .a(n30200), .b(n30198), .o(n30201) );
no02f01 g26411 ( .a(n30201), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_13_), .o(n30202) );
in01f01 g26412 ( .a(n30202), .o(n30203) );
in01f01 g26413 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_12_), .o(n30204) );
in01f01 g26414 ( .a(n30159), .o(n30205) );
na02f01 g26415 ( .a(n30205), .b(n30158), .o(n30206) );
no02f01 g26416 ( .a(n30206), .b(n30160), .o(n30207) );
in01f01 g26417 ( .a(n30207), .o(n30208) );
no04f01 g26418 ( .a(n30208), .b(n30167), .c(n30164), .d(n30161), .o(n30209) );
in01f01 g26419 ( .a(n30209), .o(n30210) );
na02f01 g26420 ( .a(n30146), .b(delay_xor_ln21_unr15_stage6_stallmux_q_12_), .o(n30211) );
in01f01 g26421 ( .a(n30211), .o(n30212) );
no02f01 g26422 ( .a(n30212), .b(n30166), .o(n30213) );
no03f01 g26423 ( .a(n30213), .b(n30210), .c(n30168), .o(n30214) );
in01f01 g26424 ( .a(n30165), .o(n30215) );
no02f01 g26425 ( .a(n30167), .b(n30215), .o(n30216) );
in01f01 g26426 ( .a(n30216), .o(n30217) );
oa12f01 g26427 ( .a(n30213), .b(n30217), .c(n30168), .o(n30218) );
in01f01 g26428 ( .a(n30218), .o(n30219) );
no02f01 g26429 ( .a(n30219), .b(n30214), .o(n30220) );
in01f01 g26430 ( .a(n30220), .o(n30221) );
no02f01 g26431 ( .a(n30221), .b(n30204), .o(n30222) );
in01f01 g26432 ( .a(n30222), .o(n30223) );
na02f01 g26433 ( .a(n30146), .b(delay_xor_ln21_unr15_stage6_stallmux_q_11_), .o(n30224) );
in01f01 g26434 ( .a(n30224), .o(n30225) );
no02f01 g26435 ( .a(n30225), .b(n30168), .o(n30226) );
no02f01 g26436 ( .a(n30226), .b(n30217), .o(n30227) );
ao12f01 g26437 ( .a(n30227), .b(n30226), .c(n30210), .o(n30228) );
no02f01 g26438 ( .a(n30228), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_11_), .o(n30229) );
in01f01 g26439 ( .a(n30229), .o(n30230) );
in01f01 g26440 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_10_), .o(n30231) );
na02f01 g26441 ( .a(n30146), .b(delay_xor_ln21_unr15_stage6_stallmux_q_10_), .o(n30232) );
in01f01 g26442 ( .a(n30232), .o(n30233) );
no02f01 g26443 ( .a(n30233), .b(n30167), .o(n30234) );
no02f01 g26444 ( .a(n30234), .b(n30215), .o(n30235) );
na02f01 g26445 ( .a(n30234), .b(n30215), .o(n30236) );
in01f01 g26446 ( .a(n30236), .o(n30237) );
no02f01 g26447 ( .a(n30237), .b(n30235), .o(n30238) );
in01f01 g26448 ( .a(n30238), .o(n30239) );
no02f01 g26449 ( .a(n30239), .b(n30231), .o(n30240) );
in01f01 g26450 ( .a(n30240), .o(n30241) );
in01f01 g26451 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_8_), .o(n30242) );
na02f01 g26452 ( .a(n30146), .b(delay_xor_ln21_unr15_stage6_stallmux_q_8_), .o(n30243) );
in01f01 g26453 ( .a(n30243), .o(n30244) );
no02f01 g26454 ( .a(n30244), .b(n30161), .o(n30245) );
no03f01 g26455 ( .a(n30245), .b(n30160), .c(n30159), .o(n30246) );
ao22f01 g26456 ( .a(n30246), .b(n30158), .c(n30245), .d(n30208), .o(n30247) );
in01f01 g26457 ( .a(n30247), .o(n30248) );
no02f01 g26458 ( .a(n30248), .b(n30242), .o(n30249) );
in01f01 g26459 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_9_), .o(n30250) );
na02f01 g26460 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_9_), .b(n30146), .o(n30251) );
in01f01 g26461 ( .a(n30251), .o(n30252) );
no02f01 g26462 ( .a(n30252), .b(n30164), .o(n30253) );
in01f01 g26463 ( .a(n30253), .o(n30254) );
ao12f01 g26464 ( .a(n30254), .b(n30162), .c(n30158), .o(n30255) );
no02f01 g26465 ( .a(n30253), .b(n30163), .o(n30256) );
no02f01 g26466 ( .a(n30256), .b(n30255), .o(n30257) );
in01f01 g26467 ( .a(n30257), .o(n30258) );
no02f01 g26468 ( .a(n30258), .b(n30250), .o(n30259) );
no02f01 g26469 ( .a(n30259), .b(n30249), .o(n30260) );
no02f01 g26470 ( .a(n30257), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_9_), .o(n30261) );
no02f01 g26471 ( .a(n30261), .b(n30260), .o(n30262) );
na02f01 g26472 ( .a(n30146), .b(delay_xor_ln21_unr15_stage6_stallmux_q_5_), .o(n30263) );
in01f01 g26473 ( .a(n30263), .o(n30264) );
no02f01 g26474 ( .a(n30264), .b(n30154), .o(n30265) );
oa12f01 g26475 ( .a(n30265), .b(n30155), .c(n30153), .o(n30266) );
in01f01 g26476 ( .a(n30266), .o(n30267) );
no03f01 g26477 ( .a(n30265), .b(n30155), .c(n30153), .o(n30268) );
no02f01 g26478 ( .a(n30268), .b(n30267), .o(n30269) );
no02f01 g26479 ( .a(n30269), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_5_), .o(n30270) );
na02f01 g26480 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_3_), .b(n30146), .o(n30271) );
na02f01 g26481 ( .a(n30271), .b(n30152), .o(n30272) );
na02f01 g26482 ( .a(n30272), .b(n30150), .o(n30273) );
in01f01 g26483 ( .a(n30273), .o(n30274) );
no02f01 g26484 ( .a(n30272), .b(n30150), .o(n30275) );
no02f01 g26485 ( .a(n30275), .b(n30274), .o(n30276) );
no02f01 g26486 ( .a(n30276), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_3_), .o(n30277) );
in01f01 g26487 ( .a(n30277), .o(n30278) );
in01f01 g26488 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_2_), .o(n30279) );
no02f01 g26489 ( .a(n30148), .b(n30147), .o(n30280) );
in01f01 g26490 ( .a(n30280), .o(n30281) );
na02f01 g26491 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_2_), .b(n30146), .o(n30282) );
in01f01 g26492 ( .a(n30282), .o(n30283) );
no02f01 g26493 ( .a(n30283), .b(n30149), .o(n30284) );
na02f01 g26494 ( .a(n30284), .b(n30281), .o(n30285) );
no02f01 g26495 ( .a(n30284), .b(n30281), .o(n30286) );
in01f01 g26496 ( .a(n30286), .o(n30287) );
na02f01 g26497 ( .a(n30287), .b(n30285), .o(n30288) );
na02f01 g26498 ( .a(n30288), .b(n30279), .o(n30289) );
in01f01 g26499 ( .a(n30147), .o(n30290) );
in01f01 g26500 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_1_), .o(n30291) );
na02f01 g26501 ( .a(n30291), .b(n_44061), .o(n30292) );
na02f01 g26502 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_1_), .b(n30146), .o(n30293) );
na02f01 g26503 ( .a(n30293), .b(n30292), .o(n30294) );
no02f01 g26504 ( .a(n30294), .b(n30290), .o(n30295) );
ao12f01 g26505 ( .a(n30147), .b(n30293), .c(n30292), .o(n30296) );
no02f01 g26506 ( .a(n30296), .b(n30295), .o(n30297) );
na02f01 g26507 ( .a(n30297), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_1_), .o(n30298) );
no02f01 g26508 ( .a(n30297), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_1_), .o(n30299) );
na02f01 g26509 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_0_), .b(n_44061), .o(n30300) );
in01f01 g26510 ( .a(n30300), .o(n30301) );
no02f01 g26511 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_0_), .b(n_44061), .o(n30302) );
no02f01 g26512 ( .a(n30302), .b(n30301), .o(n30303) );
in01f01 g26513 ( .a(n30303), .o(n30304) );
no02f01 g26514 ( .a(n30304), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_0_), .o(n30305) );
oa12f01 g26515 ( .a(n30298), .b(n30305), .c(n30299), .o(n30306) );
no02f01 g26516 ( .a(n30288), .b(n30279), .o(n30307) );
ao12f01 g26517 ( .a(n30307), .b(n30306), .c(n30289), .o(n30308) );
in01f01 g26518 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_3_), .o(n30309) );
no03f01 g26519 ( .a(n30275), .b(n30274), .c(n30309), .o(n30310) );
in01f01 g26520 ( .a(n30310), .o(n30311) );
na02f01 g26521 ( .a(n30311), .b(n30308), .o(n30312) );
na02f01 g26522 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_4_), .b(n30146), .o(n30313) );
in01f01 g26523 ( .a(n30313), .o(n30314) );
no02f01 g26524 ( .a(n30314), .b(n30155), .o(n30315) );
no02f01 g26525 ( .a(n30315), .b(n30153), .o(n30316) );
na02f01 g26526 ( .a(n30315), .b(n30153), .o(n30317) );
in01f01 g26527 ( .a(n30317), .o(n30318) );
no02f01 g26528 ( .a(n30318), .b(n30316), .o(n30319) );
no02f01 g26529 ( .a(n30319), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_4_), .o(n30320) );
in01f01 g26530 ( .a(n30320), .o(n30321) );
na03f01 g26531 ( .a(n30321), .b(n30312), .c(n30278), .o(n30322) );
in01f01 g26532 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_4_), .o(n30323) );
no03f01 g26533 ( .a(n30318), .b(n30316), .c(n30323), .o(n30324) );
in01f01 g26534 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_5_), .o(n30325) );
no03f01 g26535 ( .a(n30268), .b(n30267), .c(n30325), .o(n30326) );
no02f01 g26536 ( .a(n30326), .b(n30324), .o(n30327) );
ao12f01 g26537 ( .a(n30270), .b(n30327), .c(n30322), .o(n30328) );
na02f01 g26538 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_6_), .b(n30146), .o(n30329) );
na02f01 g26539 ( .a(n30329), .b(n30205), .o(n30330) );
in01f01 g26540 ( .a(n30330), .o(n30331) );
no03f01 g26541 ( .a(n30331), .b(n30157), .c(n30153), .o(n30332) );
no02f01 g26542 ( .a(n30330), .b(n30158), .o(n30333) );
no02f01 g26543 ( .a(n30333), .b(n30332), .o(n30334) );
no02f01 g26544 ( .a(n30334), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_6_), .o(n30335) );
in01f01 g26545 ( .a(n30335), .o(n30336) );
na02f01 g26546 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_7_), .b(n30146), .o(n30337) );
in01f01 g26547 ( .a(n30337), .o(n30338) );
no02f01 g26548 ( .a(n30338), .b(n30160), .o(n30339) );
na02f01 g26549 ( .a(n30339), .b(n30206), .o(n30340) );
in01f01 g26550 ( .a(n30340), .o(n30341) );
no02f01 g26551 ( .a(n30339), .b(n30206), .o(n30342) );
no02f01 g26552 ( .a(n30342), .b(n30341), .o(n30343) );
na02f01 g26553 ( .a(n30343), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_7_), .o(n30344) );
na02f01 g26554 ( .a(n30334), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_6_), .o(n30345) );
na02f01 g26555 ( .a(n30345), .b(n30344), .o(n30346) );
ao12f01 g26556 ( .a(n30346), .b(n30336), .c(n30328), .o(n30347) );
no02f01 g26557 ( .a(n30343), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_7_), .o(n30348) );
no02f01 g26558 ( .a(n30247), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_8_), .o(n30349) );
no02f01 g26559 ( .a(n30349), .b(n30261), .o(n30350) );
in01f01 g26560 ( .a(n30350), .o(n30351) );
no03f01 g26561 ( .a(n30351), .b(n30348), .c(n30347), .o(n30352) );
no02f01 g26562 ( .a(n30238), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_10_), .o(n30353) );
in01f01 g26563 ( .a(n30353), .o(n30354) );
oa12f01 g26564 ( .a(n30354), .b(n30352), .c(n30262), .o(n30355) );
na02f01 g26565 ( .a(n30228), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_11_), .o(n30356) );
na03f01 g26566 ( .a(n30356), .b(n30355), .c(n30241), .o(n30357) );
no02f01 g26567 ( .a(n30220), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_12_), .o(n30358) );
in01f01 g26568 ( .a(n30358), .o(n30359) );
na03f01 g26569 ( .a(n30359), .b(n30357), .c(n30230), .o(n30360) );
na02f01 g26570 ( .a(n30201), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_13_), .o(n30361) );
na03f01 g26571 ( .a(n30361), .b(n30360), .c(n30223), .o(n30362) );
no02f01 g26572 ( .a(n30172), .b(n30170), .o(n30363) );
in01f01 g26573 ( .a(n30173), .o(n30364) );
na02f01 g26574 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_14_), .b(n30146), .o(n30365) );
na02f01 g26575 ( .a(n30365), .b(n30364), .o(n30366) );
no02f01 g26576 ( .a(n30366), .b(n30363), .o(n30367) );
na02f01 g26577 ( .a(n30366), .b(n30363), .o(n30368) );
in01f01 g26578 ( .a(n30368), .o(n30369) );
no02f01 g26579 ( .a(n30369), .b(n30367), .o(n30370) );
no02f01 g26580 ( .a(n30370), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_14_), .o(n30371) );
in01f01 g26581 ( .a(n30371), .o(n30372) );
na03f01 g26582 ( .a(n30372), .b(n30362), .c(n30203), .o(n30373) );
in01f01 g26583 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_15_), .o(n30374) );
na02f01 g26584 ( .a(n30363), .b(n30364), .o(n30375) );
in01f01 g26585 ( .a(n30171), .o(n30376) );
na02f01 g26586 ( .a(n30146), .b(delay_xor_ln21_unr15_stage6_stallmux_q_15_), .o(n30377) );
na02f01 g26587 ( .a(n30377), .b(n30376), .o(n30378) );
in01f01 g26588 ( .a(n30378), .o(n30379) );
no02f01 g26589 ( .a(n30379), .b(n30175), .o(n30380) );
ao22f01 g26590 ( .a(n30380), .b(n30194), .c(n30379), .d(n30375), .o(n30381) );
in01f01 g26591 ( .a(n30381), .o(n30382) );
no02f01 g26592 ( .a(n30382), .b(n30374), .o(n30383) );
na02f01 g26593 ( .a(n30370), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_14_), .o(n30384) );
in01f01 g26594 ( .a(n30384), .o(n30385) );
no02f01 g26595 ( .a(n30385), .b(n30383), .o(n30386) );
no02f01 g26596 ( .a(n30381), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_15_), .o(n30387) );
ao12f01 g26597 ( .a(n30387), .b(n30386), .c(n30373), .o(n30388) );
in01f01 g26598 ( .a(n30176), .o(n30389) );
no02f01 g26599 ( .a(n30180), .b(n30178), .o(n30390) );
no03f01 g26600 ( .a(n30390), .b(n30375), .c(n30171), .o(n30391) );
ao12f01 g26601 ( .a(n30391), .b(n30390), .c(n30389), .o(n30392) );
no02f01 g26602 ( .a(n30392), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_16_), .o(n30393) );
in01f01 g26603 ( .a(n30393), .o(n30394) );
na03f01 g26604 ( .a(n30394), .b(n30388), .c(n30193), .o(n30395) );
no02f01 g26605 ( .a(n30182), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_18_), .o(n30396) );
no02f01 g26606 ( .a(n30396), .b(n30395), .o(n30397) );
no02f01 g26607 ( .a(n30182), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_19_), .o(n30398) );
in01f01 g26608 ( .a(n30398), .o(n30399) );
na02f01 g26609 ( .a(n30399), .b(n30397), .o(n30400) );
no02f01 g26610 ( .a(n30182), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_20_), .o(n30401) );
no03f01 g26611 ( .a(n30401), .b(n30400), .c(n30191), .o(n30402) );
in01f01 g26612 ( .a(n30402), .o(n30403) );
no02f01 g26613 ( .a(n30182), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_22_), .o(n30404) );
no02f01 g26614 ( .a(n30404), .b(n30403), .o(n30405) );
na02f01 g26615 ( .a(n30405), .b(n30190), .o(n30406) );
no02f01 g26616 ( .a(n30182), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_24_), .o(n30407) );
no02f01 g26617 ( .a(n30407), .b(n30406), .o(n30408) );
no02f01 g26618 ( .a(n30182), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_25_), .o(n30409) );
in01f01 g26619 ( .a(n30409), .o(n30410) );
na02f01 g26620 ( .a(n30410), .b(n30408), .o(n30411) );
in01f01 g26621 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_18_), .o(n30412) );
in01f01 g26622 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_19_), .o(n30413) );
ao12f01 g26623 ( .a(n30181), .b(n30413), .c(n30412), .o(n30414) );
in01f01 g26624 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_17_), .o(n30415) );
na02f01 g26625 ( .a(n30392), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_16_), .o(n30416) );
ao12f01 g26626 ( .a(n30181), .b(n30416), .c(n30415), .o(n30417) );
no02f01 g26627 ( .a(n30417), .b(n30414), .o(n30418) );
in01f01 g26628 ( .a(n30418), .o(n30419) );
in01f01 g26629 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_21_), .o(n30420) );
in01f01 g26630 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_20_), .o(n30421) );
ao12f01 g26631 ( .a(n30181), .b(n30421), .c(n30420), .o(n30422) );
no02f01 g26632 ( .a(n30422), .b(n30419), .o(n30423) );
in01f01 g26633 ( .a(n30423), .o(n30424) );
in01f01 g26634 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_23_), .o(n30425) );
in01f01 g26635 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_22_), .o(n30426) );
ao12f01 g26636 ( .a(n30181), .b(n30426), .c(n30425), .o(n30427) );
no02f01 g26637 ( .a(n30427), .b(n30424), .o(n30428) );
in01f01 g26638 ( .a(n30428), .o(n30429) );
in01f01 g26639 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_24_), .o(n30430) );
in01f01 g26640 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_25_), .o(n30431) );
ao12f01 g26641 ( .a(n30181), .b(n30431), .c(n30430), .o(n30432) );
no02f01 g26642 ( .a(n30432), .b(n30429), .o(n30433) );
na02f01 g26643 ( .a(n30433), .b(n30411), .o(n30434) );
in01f01 g26644 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_26_), .o(n30435) );
no02f01 g26645 ( .a(n30181), .b(n30435), .o(n30436) );
oa12f01 g26646 ( .a(n30188), .b(n30436), .c(n30434), .o(n30437) );
na02f01 g26647 ( .a(n30437), .b(n30186), .o(n30438) );
no02f01 g26648 ( .a(n30437), .b(n30186), .o(n30439) );
in01f01 g26649 ( .a(n30439), .o(n30440) );
na02f01 g26650 ( .a(n30440), .b(n30438), .o(n30441) );
na02f01 g26651 ( .a(n30441), .b(delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n30442) );
in01f01 g26652 ( .a(delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n30443) );
in01f01 g26653 ( .a(n30417), .o(n30444) );
no02f01 g26654 ( .a(n30181), .b(n30412), .o(n30445) );
no02f01 g26655 ( .a(n30445), .b(n30396), .o(n30446) );
na03f01 g26656 ( .a(n30446), .b(n30444), .c(n30395), .o(n30447) );
ao12f01 g26657 ( .a(n30446), .b(n30444), .c(n30395), .o(n30448) );
in01f01 g26658 ( .a(n30448), .o(n30449) );
na02f01 g26659 ( .a(n30449), .b(n30447), .o(n30450) );
na02f01 g26660 ( .a(n30450), .b(delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n30451) );
na02f01 g26661 ( .a(n30394), .b(n30388), .o(n30452) );
no02f01 g26662 ( .a(n30181), .b(n30415), .o(n30453) );
no02f01 g26663 ( .a(n30453), .b(n30192), .o(n30454) );
ao12f01 g26664 ( .a(n30454), .b(n30416), .c(n30452), .o(n30455) );
in01f01 g26665 ( .a(n30455), .o(n30456) );
in01f01 g26666 ( .a(n30416), .o(n30457) );
in01f01 g26667 ( .a(n30454), .o(n30458) );
no02f01 g26668 ( .a(n30458), .b(n30457), .o(n30459) );
na02f01 g26669 ( .a(n30459), .b(n30452), .o(n30460) );
no02f01 g26670 ( .a(n30457), .b(n30393), .o(n30461) );
in01f01 g26671 ( .a(n30461), .o(n30462) );
na02f01 g26672 ( .a(n30462), .b(n30388), .o(n30463) );
in01f01 g26673 ( .a(n30463), .o(n30464) );
no02f01 g26674 ( .a(n30462), .b(n30388), .o(n30465) );
oa12f01 g26675 ( .a(delay_sub_ln23_0_unr15_stage6_stallmux_q), .b(n30465), .c(n30464), .o(n30466) );
na03f01 g26676 ( .a(n30466), .b(n30460), .c(n30456), .o(n30467) );
na02f01 g26677 ( .a(n30467), .b(delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n30468) );
no02f01 g26678 ( .a(n30181), .b(n30413), .o(n30469) );
no02f01 g26679 ( .a(n30469), .b(n30398), .o(n30470) );
in01f01 g26680 ( .a(n30470), .o(n30471) );
no02f01 g26681 ( .a(n30417), .b(n30445), .o(n30472) );
in01f01 g26682 ( .a(n30472), .o(n30473) );
no03f01 g26683 ( .a(n30473), .b(n30471), .c(n30397), .o(n30474) );
oa12f01 g26684 ( .a(n30471), .b(n30473), .c(n30397), .o(n30475) );
in01f01 g26685 ( .a(n30475), .o(n30476) );
no02f01 g26686 ( .a(n30476), .b(n30474), .o(n30477) );
na03f01 g26687 ( .a(n30477), .b(n30468), .c(n30451), .o(n30478) );
no02f01 g26688 ( .a(n30181), .b(n30421), .o(n30479) );
no02f01 g26689 ( .a(n30479), .b(n30401), .o(n30480) );
in01f01 g26690 ( .a(n30480), .o(n30481) );
na02f01 g26691 ( .a(n30418), .b(n30400), .o(n30482) );
no02f01 g26692 ( .a(n30482), .b(n30481), .o(n30483) );
in01f01 g26693 ( .a(n30483), .o(n30484) );
na02f01 g26694 ( .a(n30482), .b(n30481), .o(n30485) );
na02f01 g26695 ( .a(n30485), .b(n30484), .o(n30486) );
oa12f01 g26696 ( .a(delay_sub_ln23_0_unr15_stage6_stallmux_q), .b(n30486), .c(n30478), .o(n30487) );
no02f01 g26697 ( .a(n30181), .b(n30420), .o(n30488) );
no02f01 g26698 ( .a(n30488), .b(n30191), .o(n30489) );
no02f01 g26699 ( .a(n30401), .b(n30400), .o(n30490) );
in01f01 g26700 ( .a(n30479), .o(n30491) );
na02f01 g26701 ( .a(n30491), .b(n30418), .o(n30492) );
no02f01 g26702 ( .a(n30492), .b(n30490), .o(n30493) );
na02f01 g26703 ( .a(n30493), .b(n30489), .o(n30494) );
in01f01 g26704 ( .a(n30489), .o(n30495) );
oa12f01 g26705 ( .a(n30495), .b(n30492), .c(n30490), .o(n30496) );
na02f01 g26706 ( .a(n30496), .b(n30494), .o(n30497) );
na02f01 g26707 ( .a(n30497), .b(delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n30498) );
na02f01 g26708 ( .a(n30498), .b(n30487), .o(n30499) );
no02f01 g26709 ( .a(n30424), .b(n30402), .o(n30500) );
no02f01 g26710 ( .a(n30181), .b(n30426), .o(n30501) );
no02f01 g26711 ( .a(n30501), .b(n30404), .o(n30502) );
no02f01 g26712 ( .a(n30502), .b(n30500), .o(n30503) );
na02f01 g26713 ( .a(n30502), .b(n30500), .o(n30504) );
in01f01 g26714 ( .a(n30504), .o(n30505) );
no02f01 g26715 ( .a(n30505), .b(n30503), .o(n30506) );
in01f01 g26716 ( .a(n30506), .o(n30507) );
ao12f01 g26717 ( .a(n30499), .b(n30507), .c(delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n30508) );
no02f01 g26718 ( .a(n30181), .b(n30425), .o(n30509) );
no02f01 g26719 ( .a(n30509), .b(n30189), .o(n30510) );
in01f01 g26720 ( .a(n30510), .o(n30511) );
no03f01 g26721 ( .a(n30501), .b(n30424), .c(n30405), .o(n30512) );
in01f01 g26722 ( .a(n30512), .o(n30513) );
no02f01 g26723 ( .a(n30513), .b(n30511), .o(n30514) );
no02f01 g26724 ( .a(n30512), .b(n30510), .o(n30515) );
no02f01 g26725 ( .a(n30515), .b(n30514), .o(n30516) );
na02f01 g26726 ( .a(n30516), .b(n30508), .o(n30517) );
no02f01 g26727 ( .a(n30181), .b(n30430), .o(n30518) );
no02f01 g26728 ( .a(n30518), .b(n30407), .o(n30519) );
in01f01 g26729 ( .a(n30519), .o(n30520) );
na02f01 g26730 ( .a(n30428), .b(n30406), .o(n30521) );
no02f01 g26731 ( .a(n30521), .b(n30520), .o(n30522) );
na02f01 g26732 ( .a(n30521), .b(n30520), .o(n30523) );
in01f01 g26733 ( .a(n30523), .o(n30524) );
no02f01 g26734 ( .a(n30524), .b(n30522), .o(n30525) );
in01f01 g26735 ( .a(n30525), .o(n30526) );
oa12f01 g26736 ( .a(delay_sub_ln23_0_unr15_stage6_stallmux_q), .b(n30526), .c(n30517), .o(n30527) );
no02f01 g26737 ( .a(n30181), .b(n30431), .o(n30528) );
no02f01 g26738 ( .a(n30528), .b(n30409), .o(n30529) );
in01f01 g26739 ( .a(n30529), .o(n30530) );
no03f01 g26740 ( .a(n30518), .b(n30429), .c(n30408), .o(n30531) );
in01f01 g26741 ( .a(n30531), .o(n30532) );
no02f01 g26742 ( .a(n30532), .b(n30530), .o(n30533) );
no02f01 g26743 ( .a(n30531), .b(n30529), .o(n30534) );
no02f01 g26744 ( .a(n30534), .b(n30533), .o(n30535) );
oa12f01 g26745 ( .a(n30527), .b(n30535), .c(n30443), .o(n30536) );
no02f01 g26746 ( .a(n30436), .b(n30187), .o(n30537) );
in01f01 g26747 ( .a(n30537), .o(n30538) );
no02f01 g26748 ( .a(n30538), .b(n30434), .o(n30539) );
na02f01 g26749 ( .a(n30538), .b(n30434), .o(n30540) );
in01f01 g26750 ( .a(n30540), .o(n30541) );
no02f01 g26751 ( .a(n30541), .b(n30539), .o(n30542) );
in01f01 g26752 ( .a(n30542), .o(n30543) );
ao12f01 g26753 ( .a(n30536), .b(n30543), .c(delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n30544) );
na02f01 g26754 ( .a(n30544), .b(n30442), .o(n30545) );
in01f01 g26755 ( .a(n30545), .o(n30546) );
no02f01 g26756 ( .a(n30187), .b(n30183), .o(n30547) );
in01f01 g26757 ( .a(n30547), .o(n30548) );
no02f01 g26758 ( .a(n30548), .b(n30411), .o(n30549) );
in01f01 g26759 ( .a(n30549), .o(n30550) );
no02f01 g26760 ( .a(n30182), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_28_), .o(n30551) );
no02f01 g26761 ( .a(n30551), .b(n30550), .o(n30552) );
ao12f01 g26762 ( .a(n30181), .b(n30435), .c(n30184), .o(n30553) );
no02f01 g26763 ( .a(n30553), .b(n30432), .o(n30554) );
na02f01 g26764 ( .a(n30554), .b(n30428), .o(n30555) );
in01f01 g26765 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_28_), .o(n30556) );
no02f01 g26766 ( .a(n30181), .b(n30556), .o(n30557) );
no02f01 g26767 ( .a(n30557), .b(n30555), .o(n30558) );
in01f01 g26768 ( .a(n30558), .o(n30559) );
no02f01 g26769 ( .a(n30559), .b(n30552), .o(n30560) );
no02f01 g26770 ( .a(n30182), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_29_), .o(n30561) );
in01f01 g26771 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_29_), .o(n30562) );
no02f01 g26772 ( .a(n30181), .b(n30562), .o(n30563) );
no02f01 g26773 ( .a(n30563), .b(n30561), .o(n30564) );
no02f01 g26774 ( .a(n30564), .b(n30560), .o(n30565) );
in01f01 g26775 ( .a(n30565), .o(n30566) );
na02f01 g26776 ( .a(n30564), .b(n30560), .o(n30567) );
na02f01 g26777 ( .a(n30567), .b(n30566), .o(n30568) );
no02f01 g26778 ( .a(n30555), .b(n30549), .o(n30569) );
no02f01 g26779 ( .a(n30557), .b(n30551), .o(n30570) );
no02f01 g26780 ( .a(n30570), .b(n30569), .o(n30571) );
na02f01 g26781 ( .a(n30570), .b(n30569), .o(n30572) );
in01f01 g26782 ( .a(n30572), .o(n30573) );
no02f01 g26783 ( .a(n30573), .b(n30571), .o(n30574) );
in01f01 g26784 ( .a(n30574), .o(n30575) );
oa12f01 g26785 ( .a(delay_sub_ln23_0_unr15_stage6_stallmux_q), .b(n30575), .c(n30568), .o(n30576) );
na02f01 g26786 ( .a(n30576), .b(n30546), .o(n30577) );
no03f01 g26787 ( .a(n30561), .b(n30551), .c(n30550), .o(n30578) );
in01f01 g26788 ( .a(n30578), .o(n30579) );
ao12f01 g26789 ( .a(n30181), .b(n30562), .c(n30556), .o(n30580) );
no02f01 g26790 ( .a(n30580), .b(n30555), .o(n30581) );
in01f01 g26791 ( .a(n30581), .o(n30582) );
no02f01 g26792 ( .a(n30582), .b(n30578), .o(n30583) );
in01f01 g26793 ( .a(n30583), .o(n30584) );
no02f01 g26794 ( .a(n30182), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_30_), .o(n30585) );
na02f01 g26795 ( .a(n30182), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_30_), .o(n30586) );
in01f01 g26796 ( .a(n30586), .o(n30587) );
no02f01 g26797 ( .a(n30587), .b(n30585), .o(n30588) );
in01f01 g26798 ( .a(n30588), .o(n30589) );
no02f01 g26799 ( .a(n30589), .b(n30582), .o(n30590) );
ao22f01 g26800 ( .a(n30590), .b(n30579), .c(n30589), .d(n30584), .o(n30591) );
no02f01 g26801 ( .a(n30591), .b(delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n30592) );
in01f01 g26802 ( .a(n30591), .o(n30593) );
no02f01 g26803 ( .a(n30593), .b(n30443), .o(n30594) );
no02f01 g26804 ( .a(n30594), .b(n30592), .o(n30595) );
in01f01 g26805 ( .a(n30567), .o(n30596) );
no02f01 g26806 ( .a(n30596), .b(n30565), .o(n30597) );
ao12f01 g26807 ( .a(delay_sub_ln23_0_unr15_stage6_stallmux_q), .b(n30574), .c(n30597), .o(n30598) );
in01f01 g26808 ( .a(n30598), .o(n30599) );
oa12f01 g26809 ( .a(n30599), .b(n30595), .c(n30577), .o(n30600) );
na02f01 g26810 ( .a(n30600), .b(delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n30601) );
na02f01 g26811 ( .a(n30599), .b(n30577), .o(n30602) );
no02f01 g26812 ( .a(n30593), .b(delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n30603) );
in01f01 g26813 ( .a(n30603), .o(n30604) );
no02f01 g26814 ( .a(n30604), .b(n30602), .o(n30605) );
no02f01 g26815 ( .a(n30182), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_31_), .o(n30606) );
na02f01 g26816 ( .a(n30182), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_31_), .o(n30607) );
in01f01 g26817 ( .a(n30607), .o(n30608) );
no02f01 g26818 ( .a(n30608), .b(n30606), .o(n30609) );
in01f01 g26819 ( .a(n30609), .o(n30610) );
no02f01 g26820 ( .a(n30587), .b(n30582), .o(n30611) );
oa12f01 g26821 ( .a(n30611), .b(n30585), .c(n30579), .o(n30612) );
no02f01 g26822 ( .a(n30612), .b(n30610), .o(n30613) );
na02f01 g26823 ( .a(n30612), .b(n30610), .o(n30614) );
in01f01 g26824 ( .a(n30614), .o(n30615) );
no02f01 g26825 ( .a(n30615), .b(n30613), .o(n30616) );
na02f01 g26826 ( .a(n30616), .b(delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n30617) );
in01f01 g26827 ( .a(n30613), .o(n30618) );
na02f01 g26828 ( .a(n30614), .b(n30618), .o(n30619) );
na02f01 g26829 ( .a(n30619), .b(n30443), .o(n30620) );
na02f01 g26830 ( .a(n30620), .b(n30617), .o(n30621) );
oa12f01 g26831 ( .a(n30601), .b(n30621), .c(n30605), .o(n30622) );
in01f01 g26832 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_16_), .o(n30623) );
no02f01 g26833 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_2_), .b(n30146), .o(n30624) );
in01f01 g26834 ( .a(n30624), .o(n30625) );
no02f01 g26835 ( .a(n_45204), .b(n30146), .o(n30626) );
no02f01 g26836 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_0_), .b(n30146), .o(n30627) );
no02f01 g26837 ( .a(n30627), .b(n30626), .o(n30628) );
na02f01 g26838 ( .a(n30628), .b(n30625), .o(n30629) );
in01f01 g26839 ( .a(n30629), .o(n30630) );
no02f01 g26840 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_3_), .b(n30146), .o(n30631) );
no02f01 g26841 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_5_), .b(n30146), .o(n30632) );
no02f01 g26842 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_4_), .b(n30146), .o(n30633) );
no03f01 g26843 ( .a(n30633), .b(n30632), .c(n30631), .o(n30634) );
na02f01 g26844 ( .a(n30634), .b(n30630), .o(n30635) );
in01f01 g26845 ( .a(n30635), .o(n30636) );
no02f01 g26846 ( .a(n30146), .b(delay_xor_ln22_unr15_stage6_stallmux_q_7_), .o(n30637) );
no02f01 g26847 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_6_), .b(n30146), .o(n30638) );
no02f01 g26848 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_8_), .b(n30146), .o(n30639) );
no03f01 g26849 ( .a(n30639), .b(n30638), .c(n30637), .o(n30640) );
na02f01 g26850 ( .a(n30640), .b(n30636), .o(n30641) );
in01f01 g26851 ( .a(n30641), .o(n30642) );
no02f01 g26852 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_9_), .b(n30146), .o(n30643) );
no02f01 g26853 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_11_), .b(n30146), .o(n30644) );
no02f01 g26854 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_10_), .b(n30146), .o(n30645) );
no03f01 g26855 ( .a(n30645), .b(n30644), .c(n30643), .o(n30646) );
na02f01 g26856 ( .a(n30646), .b(n30642), .o(n30647) );
in01f01 g26857 ( .a(n30647), .o(n30648) );
no02f01 g26858 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_12_), .b(n30146), .o(n30649) );
no02f01 g26859 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_13_), .b(n30146), .o(n30650) );
no02f01 g26860 ( .a(n30650), .b(n30649), .o(n30651) );
na02f01 g26861 ( .a(n30651), .b(n30648), .o(n30652) );
no02f01 g26862 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_14_), .b(n30146), .o(n30653) );
no02f01 g26863 ( .a(n30653), .b(n30652), .o(n30654) );
in01f01 g26864 ( .a(n30654), .o(n30655) );
no02f01 g26865 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_15_), .b(n30146), .o(n30656) );
no02f01 g26866 ( .a(n30656), .b(n30655), .o(n30657) );
in01f01 g26867 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_16_), .o(n30658) );
no02f01 g26868 ( .a(n_44061), .b(n30658), .o(n30659) );
no02f01 g26869 ( .a(n30146), .b(delay_xor_ln22_unr15_stage6_stallmux_q_16_), .o(n30660) );
no02f01 g26870 ( .a(n30660), .b(n30659), .o(n30661) );
in01f01 g26871 ( .a(n30661), .o(n30662) );
no02f01 g26872 ( .a(n30662), .b(n30657), .o(n30663) );
no03f01 g26873 ( .a(n30661), .b(n30656), .c(n30655), .o(n30664) );
no02f01 g26874 ( .a(n30664), .b(n30663), .o(n30665) );
no02f01 g26875 ( .a(n30665), .b(n30623), .o(n30666) );
in01f01 g26876 ( .a(n30666), .o(n30667) );
in01f01 g26877 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_15_), .o(n30668) );
na02f01 g26878 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_15_), .b(n30146), .o(n30669) );
in01f01 g26879 ( .a(n30669), .o(n30670) );
no02f01 g26880 ( .a(n30670), .b(n30656), .o(n30671) );
in01f01 g26881 ( .a(n30671), .o(n30672) );
no02f01 g26882 ( .a(n30672), .b(n30654), .o(n30673) );
no02f01 g26883 ( .a(n30671), .b(n30655), .o(n30674) );
no02f01 g26884 ( .a(n30674), .b(n30673), .o(n30675) );
no02f01 g26885 ( .a(n30675), .b(n30668), .o(n30676) );
in01f01 g26886 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_14_), .o(n30677) );
na02f01 g26887 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_14_), .b(n30146), .o(n30678) );
in01f01 g26888 ( .a(n30678), .o(n30679) );
no02f01 g26889 ( .a(n30679), .b(n30653), .o(n30680) );
in01f01 g26890 ( .a(n30680), .o(n30681) );
ao12f01 g26891 ( .a(n30681), .b(n30651), .c(n30648), .o(n30682) );
no02f01 g26892 ( .a(n30680), .b(n30652), .o(n30683) );
no02f01 g26893 ( .a(n30683), .b(n30682), .o(n30684) );
no02f01 g26894 ( .a(n30684), .b(n30677), .o(n30685) );
in01f01 g26895 ( .a(n30685), .o(n30686) );
na02f01 g26896 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_13_), .b(n30146), .o(n30687) );
in01f01 g26897 ( .a(n30687), .o(n30688) );
no02f01 g26898 ( .a(n30688), .b(n30650), .o(n30689) );
in01f01 g26899 ( .a(n30649), .o(n30690) );
na02f01 g26900 ( .a(n30690), .b(n30648), .o(n30691) );
no02f01 g26901 ( .a(n30638), .b(n30635), .o(n30692) );
in01f01 g26902 ( .a(n30692), .o(n30693) );
no02f01 g26903 ( .a(n30693), .b(n30637), .o(n30694) );
no03f01 g26904 ( .a(n30645), .b(n30643), .c(n30639), .o(n30695) );
na02f01 g26905 ( .a(n30695), .b(n30694), .o(n30696) );
in01f01 g26906 ( .a(n30696), .o(n30697) );
no03f01 g26907 ( .a(n30689), .b(n30649), .c(n30644), .o(n30698) );
ao22f01 g26908 ( .a(n30698), .b(n30697), .c(n30691), .d(n30689), .o(n30699) );
in01f01 g26909 ( .a(n30699), .o(n30700) );
no02f01 g26910 ( .a(n30700), .b(delay_add_ln22_unr14_stage6_stallmux_q_13_), .o(n30701) );
in01f01 g26911 ( .a(n30701), .o(n30702) );
na02f01 g26912 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_11_), .b(n30146), .o(n30703) );
in01f01 g26913 ( .a(n30703), .o(n30704) );
no02f01 g26914 ( .a(n30704), .b(n30644), .o(n30705) );
no04f01 g26915 ( .a(n30705), .b(n30645), .c(n30643), .d(n30641), .o(n30706) );
ao12f01 g26916 ( .a(n30706), .b(n30705), .c(n30696), .o(n30707) );
in01f01 g26917 ( .a(n30707), .o(n30708) );
no02f01 g26918 ( .a(n30708), .b(delay_add_ln22_unr14_stage6_stallmux_q_11_), .o(n30709) );
in01f01 g26919 ( .a(n30709), .o(n30710) );
in01f01 g26920 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_10_), .o(n30711) );
na02f01 g26921 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_10_), .b(n30146), .o(n30712) );
in01f01 g26922 ( .a(n30712), .o(n30713) );
no02f01 g26923 ( .a(n30713), .b(n30645), .o(n30714) );
no02f01 g26924 ( .a(n30714), .b(n30643), .o(n30715) );
no02f01 g26925 ( .a(n30643), .b(n30641), .o(n30716) );
in01f01 g26926 ( .a(n30716), .o(n30717) );
ao22f01 g26927 ( .a(n30717), .b(n30714), .c(n30715), .d(n30642), .o(n30718) );
no02f01 g26928 ( .a(n30718), .b(n30711), .o(n30719) );
in01f01 g26929 ( .a(n30719), .o(n30720) );
in01f01 g26930 ( .a(n30637), .o(n30721) );
na02f01 g26931 ( .a(n30146), .b(delay_xor_ln22_unr15_stage6_stallmux_q_7_), .o(n30722) );
na02f01 g26932 ( .a(n30722), .b(n30721), .o(n30723) );
in01f01 g26933 ( .a(n30638), .o(n30724) );
na02f01 g26934 ( .a(n30723), .b(n30724), .o(n30725) );
oa22f01 g26935 ( .a(n30725), .b(n30635), .c(n30723), .d(n30692), .o(n30726) );
no02f01 g26936 ( .a(n30726), .b(delay_add_ln22_unr14_stage6_stallmux_q_7_), .o(n30727) );
in01f01 g26937 ( .a(n30727), .o(n30728) );
in01f01 g26938 ( .a(n30633), .o(n30729) );
no02f01 g26939 ( .a(n30631), .b(n30629), .o(n30730) );
na02f01 g26940 ( .a(n30730), .b(n30729), .o(n30731) );
na02f01 g26941 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_5_), .b(n30146), .o(n30732) );
in01f01 g26942 ( .a(n30732), .o(n30733) );
no02f01 g26943 ( .a(n30733), .b(n30632), .o(n30734) );
na02f01 g26944 ( .a(n30734), .b(n30731), .o(n30735) );
in01f01 g26945 ( .a(n30734), .o(n30736) );
na03f01 g26946 ( .a(n30736), .b(n30730), .c(n30729), .o(n30737) );
na02f01 g26947 ( .a(n30737), .b(n30735), .o(n30738) );
no02f01 g26948 ( .a(n30738), .b(delay_add_ln22_unr14_stage6_stallmux_q_5_), .o(n30739) );
in01f01 g26949 ( .a(n30631), .o(n30740) );
na02f01 g26950 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_3_), .b(n30146), .o(n30741) );
na03f01 g26951 ( .a(n30741), .b(n30740), .c(n30629), .o(n30742) );
na02f01 g26952 ( .a(n30741), .b(n30740), .o(n30743) );
na02f01 g26953 ( .a(n30743), .b(n30630), .o(n30744) );
na02f01 g26954 ( .a(n30744), .b(n30742), .o(n30745) );
no02f01 g26955 ( .a(n30745), .b(delay_add_ln22_unr14_stage6_stallmux_q_3_), .o(n30746) );
in01f01 g26956 ( .a(n30746), .o(n30747) );
na02f01 g26957 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_2_), .b(n30146), .o(n30748) );
na02f01 g26958 ( .a(n30748), .b(n30625), .o(n30749) );
na02f01 g26959 ( .a(n30749), .b(n30628), .o(n30750) );
no02f01 g26960 ( .a(n30749), .b(n30628), .o(n30751) );
in01f01 g26961 ( .a(n30751), .o(n30752) );
na02f01 g26962 ( .a(n30752), .b(n30750), .o(n30753) );
na02f01 g26963 ( .a(n30753), .b(delay_add_ln22_unr14_stage6_stallmux_q_2_), .o(n30754) );
in01f01 g26964 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_1_), .o(n30755) );
in01f01 g26965 ( .a(n30627), .o(n30756) );
in01f01 g26966 ( .a(n_45204), .o(n30757) );
na02f01 g26967 ( .a(n30757), .b(n_44061), .o(n30758) );
na02f01 g26968 ( .a(n_45204), .b(n30146), .o(n30759) );
na02f01 g26969 ( .a(n30759), .b(n30758), .o(n30760) );
no02f01 g26970 ( .a(n30760), .b(n30756), .o(n30761) );
ao12f01 g26971 ( .a(n30627), .b(n30759), .c(n30758), .o(n30762) );
no02f01 g26972 ( .a(n30762), .b(n30761), .o(n30763) );
no02f01 g26973 ( .a(n30763), .b(n30755), .o(n30764) );
na02f01 g26974 ( .a(n30763), .b(n30755), .o(n30765) );
in01f01 g26975 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_0_), .o(n30766) );
in01f01 g26976 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_0_), .o(n30767) );
no02f01 g26977 ( .a(n30767), .b(n30146), .o(n30768) );
no02f01 g26978 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_0_), .b(n_44061), .o(n30769) );
no02f01 g26979 ( .a(n30769), .b(n30768), .o(n30770) );
in01f01 g26980 ( .a(n30770), .o(n30771) );
no02f01 g26981 ( .a(n30771), .b(n30766), .o(n30772) );
ao12f01 g26982 ( .a(n30764), .b(n30772), .c(n30765), .o(n30773) );
no02f01 g26983 ( .a(n30753), .b(delay_add_ln22_unr14_stage6_stallmux_q_2_), .o(n30774) );
oa12f01 g26984 ( .a(n30754), .b(n30774), .c(n30773), .o(n30775) );
na02f01 g26985 ( .a(n30745), .b(delay_add_ln22_unr14_stage6_stallmux_q_3_), .o(n30776) );
in01f01 g26986 ( .a(n30776), .o(n30777) );
oa12f01 g26987 ( .a(n30747), .b(n30777), .c(n30775), .o(n30778) );
in01f01 g26988 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_4_), .o(n30779) );
na02f01 g26989 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_4_), .b(n30146), .o(n30780) );
na02f01 g26990 ( .a(n30780), .b(n30729), .o(n30781) );
no02f01 g26991 ( .a(n30781), .b(n30730), .o(n30782) );
na02f01 g26992 ( .a(n30781), .b(n30730), .o(n30783) );
in01f01 g26993 ( .a(n30783), .o(n30784) );
no02f01 g26994 ( .a(n30784), .b(n30782), .o(n30785) );
na02f01 g26995 ( .a(n30785), .b(n30779), .o(n30786) );
in01f01 g26996 ( .a(n30786), .o(n30787) );
no02f01 g26997 ( .a(n30787), .b(n30778), .o(n30788) );
in01f01 g26998 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_5_), .o(n30789) );
ao12f01 g26999 ( .a(n30789), .b(n30737), .c(n30735), .o(n30790) );
no02f01 g27000 ( .a(n30785), .b(n30779), .o(n30791) );
no02f01 g27001 ( .a(n30791), .b(n30790), .o(n30792) );
in01f01 g27002 ( .a(n30792), .o(n30793) );
no02f01 g27003 ( .a(n30793), .b(n30788), .o(n30794) );
na02f01 g27004 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_6_), .b(n30146), .o(n30795) );
na02f01 g27005 ( .a(n30795), .b(n30724), .o(n30796) );
in01f01 g27006 ( .a(n30796), .o(n30797) );
no02f01 g27007 ( .a(n30797), .b(n30635), .o(n30798) );
no02f01 g27008 ( .a(n30796), .b(n30636), .o(n30799) );
no02f01 g27009 ( .a(n30799), .b(n30798), .o(n30800) );
in01f01 g27010 ( .a(n30800), .o(n30801) );
no02f01 g27011 ( .a(n30801), .b(delay_add_ln22_unr14_stage6_stallmux_q_6_), .o(n30802) );
no03f01 g27012 ( .a(n30802), .b(n30794), .c(n30739), .o(n30803) );
na02f01 g27013 ( .a(n30801), .b(delay_add_ln22_unr14_stage6_stallmux_q_6_), .o(n30804) );
in01f01 g27014 ( .a(n30804), .o(n30805) );
na02f01 g27015 ( .a(n30726), .b(delay_add_ln22_unr14_stage6_stallmux_q_7_), .o(n30806) );
in01f01 g27016 ( .a(n30806), .o(n30807) );
no02f01 g27017 ( .a(n30807), .b(n30805), .o(n30808) );
in01f01 g27018 ( .a(n30808), .o(n30809) );
oa12f01 g27019 ( .a(n30728), .b(n30809), .c(n30803), .o(n30810) );
in01f01 g27020 ( .a(n30694), .o(n30811) );
na02f01 g27021 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_8_), .b(n30146), .o(n30812) );
in01f01 g27022 ( .a(n30812), .o(n30813) );
no02f01 g27023 ( .a(n30813), .b(n30639), .o(n30814) );
no03f01 g27024 ( .a(n30814), .b(n30638), .c(n30637), .o(n30815) );
ao22f01 g27025 ( .a(n30815), .b(n30636), .c(n30814), .d(n30811), .o(n30816) );
in01f01 g27026 ( .a(n30816), .o(n30817) );
no02f01 g27027 ( .a(n30817), .b(delay_add_ln22_unr14_stage6_stallmux_q_8_), .o(n30818) );
in01f01 g27028 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_9_), .o(n30819) );
na02f01 g27029 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_9_), .b(n30146), .o(n30820) );
in01f01 g27030 ( .a(n30820), .o(n30821) );
no02f01 g27031 ( .a(n30821), .b(n30643), .o(n30822) );
no02f01 g27032 ( .a(n30822), .b(n30641), .o(n30823) );
na02f01 g27033 ( .a(n30822), .b(n30641), .o(n30824) );
in01f01 g27034 ( .a(n30824), .o(n30825) );
no02f01 g27035 ( .a(n30825), .b(n30823), .o(n30826) );
no02f01 g27036 ( .a(n30826), .b(n30819), .o(n30827) );
na02f01 g27037 ( .a(n30817), .b(delay_add_ln22_unr14_stage6_stallmux_q_8_), .o(n30828) );
in01f01 g27038 ( .a(n30828), .o(n30829) );
no02f01 g27039 ( .a(n30829), .b(n30827), .o(n30830) );
oa12f01 g27040 ( .a(n30830), .b(n30818), .c(n30810), .o(n30831) );
na02f01 g27041 ( .a(n30718), .b(n30711), .o(n30832) );
in01f01 g27042 ( .a(n30832), .o(n30833) );
na02f01 g27043 ( .a(n30826), .b(n30819), .o(n30834) );
in01f01 g27044 ( .a(n30834), .o(n30835) );
no02f01 g27045 ( .a(n30835), .b(n30833), .o(n30836) );
na02f01 g27046 ( .a(n30836), .b(n30831), .o(n30837) );
na02f01 g27047 ( .a(n30837), .b(n30720), .o(n30838) );
na02f01 g27048 ( .a(n30708), .b(delay_add_ln22_unr14_stage6_stallmux_q_11_), .o(n30839) );
in01f01 g27049 ( .a(n30839), .o(n30840) );
oa12f01 g27050 ( .a(n30710), .b(n30840), .c(n30838), .o(n30841) );
na02f01 g27051 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_12_), .b(n30146), .o(n30842) );
na02f01 g27052 ( .a(n30842), .b(n30690), .o(n30843) );
no02f01 g27053 ( .a(n30843), .b(n30648), .o(n30844) );
na02f01 g27054 ( .a(n30843), .b(n30648), .o(n30845) );
in01f01 g27055 ( .a(n30845), .o(n30846) );
no02f01 g27056 ( .a(n30846), .b(n30844), .o(n30847) );
in01f01 g27057 ( .a(n30847), .o(n30848) );
no02f01 g27058 ( .a(n30848), .b(delay_add_ln22_unr14_stage6_stallmux_q_12_), .o(n30849) );
na02f01 g27059 ( .a(n30700), .b(delay_add_ln22_unr14_stage6_stallmux_q_13_), .o(n30850) );
in01f01 g27060 ( .a(n30850), .o(n30851) );
na02f01 g27061 ( .a(n30848), .b(delay_add_ln22_unr14_stage6_stallmux_q_12_), .o(n30852) );
in01f01 g27062 ( .a(n30852), .o(n30853) );
no02f01 g27063 ( .a(n30853), .b(n30851), .o(n30854) );
oa12f01 g27064 ( .a(n30854), .b(n30849), .c(n30841), .o(n30855) );
na02f01 g27065 ( .a(n30684), .b(n30677), .o(n30856) );
na03f01 g27066 ( .a(n30856), .b(n30855), .c(n30702), .o(n30857) );
na02f01 g27067 ( .a(n30675), .b(n30668), .o(n30858) );
in01f01 g27068 ( .a(n30858), .o(n30859) );
ao12f01 g27069 ( .a(n30859), .b(n30857), .c(n30686), .o(n30860) );
na02f01 g27070 ( .a(n30665), .b(n30623), .o(n30861) );
oa12f01 g27071 ( .a(n30861), .b(n30860), .c(n30676), .o(n30862) );
in01f01 g27072 ( .a(n30659), .o(n30863) );
ao12f01 g27073 ( .a(n30660), .b(n30863), .c(n30657), .o(n30864) );
no02f01 g27074 ( .a(n30864), .b(delay_add_ln22_unr14_stage6_stallmux_q_17_), .o(n30865) );
na02f01 g27075 ( .a(n30864), .b(delay_add_ln22_unr14_stage6_stallmux_q_17_), .o(n30866) );
in01f01 g27076 ( .a(n30866), .o(n30867) );
no02f01 g27077 ( .a(n30867), .b(n30865), .o(n30868) );
na03f01 g27078 ( .a(n30868), .b(n30862), .c(n30667), .o(n30869) );
na02f01 g27079 ( .a(n30862), .b(n30667), .o(n30870) );
in01f01 g27080 ( .a(n30868), .o(n30871) );
na02f01 g27081 ( .a(n30871), .b(n30870), .o(n30872) );
na02f01 g27082 ( .a(n30872), .b(n30869), .o(n30873) );
no02f01 g27083 ( .a(n30860), .b(n30676), .o(n30874) );
in01f01 g27084 ( .a(n30861), .o(n30875) );
no02f01 g27085 ( .a(n30875), .b(n30666), .o(n30876) );
na02f01 g27086 ( .a(n30876), .b(n30874), .o(n30877) );
in01f01 g27087 ( .a(n30676), .o(n30878) );
na02f01 g27088 ( .a(n30857), .b(n30686), .o(n30879) );
na02f01 g27089 ( .a(n30858), .b(n30879), .o(n30880) );
na02f01 g27090 ( .a(n30880), .b(n30878), .o(n30881) );
in01f01 g27091 ( .a(n30876), .o(n30882) );
na02f01 g27092 ( .a(n30882), .b(n30881), .o(n30883) );
na02f01 g27093 ( .a(n30883), .b(n30877), .o(n30884) );
no02f01 g27094 ( .a(n30884), .b(n30873), .o(n30885) );
no02f01 g27095 ( .a(n30885), .b(n30622), .o(n30886) );
no02f01 g27096 ( .a(n30865), .b(n30875), .o(n30887) );
oa12f01 g27097 ( .a(n30887), .b(n30860), .c(n30676), .o(n30888) );
ao12f01 g27098 ( .a(n30865), .b(n30866), .c(n30667), .o(n30889) );
in01f01 g27099 ( .a(n30889), .o(n30890) );
in01f01 g27100 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_18_), .o(n30891) );
in01f01 g27101 ( .a(n30864), .o(n30892) );
no02f01 g27102 ( .a(n30892), .b(n30891), .o(n30893) );
no02f01 g27103 ( .a(n30864), .b(delay_add_ln22_unr14_stage6_stallmux_q_18_), .o(n30894) );
no02f01 g27104 ( .a(n30894), .b(n30893), .o(n30895) );
na03f01 g27105 ( .a(n30895), .b(n30890), .c(n30888), .o(n30896) );
in01f01 g27106 ( .a(n30896), .o(n30897) );
ao12f01 g27107 ( .a(n30895), .b(n30890), .c(n30888), .o(n30898) );
no02f01 g27108 ( .a(n30898), .b(n30897), .o(n30899) );
in01f01 g27109 ( .a(n30893), .o(n30900) );
na02f01 g27110 ( .a(n30890), .b(n30888), .o(n30901) );
in01f01 g27111 ( .a(n30894), .o(n30902) );
na02f01 g27112 ( .a(n30902), .b(n30901), .o(n30903) );
in01f01 g27113 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_19_), .o(n30904) );
no02f01 g27114 ( .a(n30892), .b(n30904), .o(n30905) );
no02f01 g27115 ( .a(n30864), .b(delay_add_ln22_unr14_stage6_stallmux_q_19_), .o(n30906) );
no02f01 g27116 ( .a(n30906), .b(n30905), .o(n30907) );
na03f01 g27117 ( .a(n30907), .b(n30903), .c(n30900), .o(n30908) );
in01f01 g27118 ( .a(n30908), .o(n30909) );
ao12f01 g27119 ( .a(n30907), .b(n30903), .c(n30900), .o(n30910) );
no02f01 g27120 ( .a(n30910), .b(n30909), .o(n30911) );
ao12f01 g27121 ( .a(n30622), .b(n30911), .c(n30899), .o(n30912) );
no02f01 g27122 ( .a(n30912), .b(n30886), .o(n30913) );
in01f01 g27123 ( .a(n30913), .o(n30914) );
no02f01 g27124 ( .a(n30905), .b(n30893), .o(n30915) );
na03f01 g27125 ( .a(n30915), .b(n30890), .c(n30888), .o(n30916) );
ao12f01 g27126 ( .a(n30864), .b(delay_add_ln22_unr14_stage6_stallmux_q_18_), .c(delay_add_ln22_unr14_stage6_stallmux_q_19_), .o(n30917) );
in01f01 g27127 ( .a(n30917), .o(n30918) );
na02f01 g27128 ( .a(n30918), .b(n30916), .o(n30919) );
in01f01 g27129 ( .a(n30919), .o(n30920) );
no02f01 g27130 ( .a(n30864), .b(delay_add_ln22_unr14_stage6_stallmux_q_20_), .o(n30921) );
in01f01 g27131 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_20_), .o(n30922) );
no02f01 g27132 ( .a(n30892), .b(n30922), .o(n30923) );
no02f01 g27133 ( .a(n30923), .b(n30921), .o(n30924) );
in01f01 g27134 ( .a(n30924), .o(n30925) );
no02f01 g27135 ( .a(n30925), .b(n30920), .o(n30926) );
no02f01 g27136 ( .a(n30924), .b(n30919), .o(n30927) );
no02f01 g27137 ( .a(n30927), .b(n30926), .o(n30928) );
no02f01 g27138 ( .a(n30928), .b(n30622), .o(n30929) );
in01f01 g27139 ( .a(n30923), .o(n30930) );
no02f01 g27140 ( .a(n30864), .b(delay_add_ln22_unr14_stage6_stallmux_q_21_), .o(n30931) );
in01f01 g27141 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_21_), .o(n30932) );
no02f01 g27142 ( .a(n30892), .b(n30932), .o(n30933) );
no02f01 g27143 ( .a(n30933), .b(n30931), .o(n30934) );
in01f01 g27144 ( .a(n30921), .o(n30935) );
na02f01 g27145 ( .a(n30935), .b(n30920), .o(n30936) );
na03f01 g27146 ( .a(n30936), .b(n30934), .c(n30930), .o(n30937) );
in01f01 g27147 ( .a(n30937), .o(n30938) );
ao12f01 g27148 ( .a(n30934), .b(n30936), .c(n30930), .o(n30939) );
no02f01 g27149 ( .a(n30939), .b(n30938), .o(n30940) );
no02f01 g27150 ( .a(n30940), .b(n30622), .o(n30941) );
no03f01 g27151 ( .a(n30941), .b(n30929), .c(n30914), .o(n30942) );
no02f01 g27152 ( .a(n30864), .b(delay_add_ln22_unr14_stage6_stallmux_q_22_), .o(n30943) );
na02f01 g27153 ( .a(n30864), .b(delay_add_ln22_unr14_stage6_stallmux_q_22_), .o(n30944) );
in01f01 g27154 ( .a(n30944), .o(n30945) );
no02f01 g27155 ( .a(n30945), .b(n30943), .o(n30946) );
ao12f01 g27156 ( .a(n30892), .b(n30922), .c(n30932), .o(n30947) );
in01f01 g27157 ( .a(n30947), .o(n30948) );
no02f01 g27158 ( .a(n30931), .b(n30921), .o(n30949) );
in01f01 g27159 ( .a(n30949), .o(n30950) );
oa12f01 g27160 ( .a(n30948), .b(n30950), .c(n30919), .o(n30951) );
in01f01 g27161 ( .a(n30951), .o(n30952) );
na02f01 g27162 ( .a(n30952), .b(n30946), .o(n30953) );
in01f01 g27163 ( .a(n30946), .o(n30954) );
na02f01 g27164 ( .a(n30951), .b(n30954), .o(n30955) );
na02f01 g27165 ( .a(n30955), .b(n30953), .o(n30956) );
in01f01 g27166 ( .a(n30956), .o(n30957) );
no02f01 g27167 ( .a(n30947), .b(n30945), .o(n30958) );
in01f01 g27168 ( .a(n30958), .o(n30959) );
no03f01 g27169 ( .a(n30950), .b(n30943), .c(n30919), .o(n30960) );
no02f01 g27170 ( .a(n30864), .b(delay_add_ln22_unr14_stage6_stallmux_q_23_), .o(n30961) );
na02f01 g27171 ( .a(n30864), .b(delay_add_ln22_unr14_stage6_stallmux_q_23_), .o(n30962) );
in01f01 g27172 ( .a(n30962), .o(n30963) );
no02f01 g27173 ( .a(n30963), .b(n30961), .o(n30964) );
in01f01 g27174 ( .a(n30964), .o(n30965) );
oa12f01 g27175 ( .a(n30965), .b(n30960), .c(n30959), .o(n30966) );
in01f01 g27176 ( .a(n30966), .o(n30967) );
no03f01 g27177 ( .a(n30965), .b(n30960), .c(n30959), .o(n30968) );
no02f01 g27178 ( .a(n30968), .b(n30967), .o(n30969) );
ao12f01 g27179 ( .a(n30622), .b(n30969), .c(n30957), .o(n30970) );
in01f01 g27180 ( .a(n30970), .o(n30971) );
na02f01 g27181 ( .a(n30971), .b(n30942), .o(n30972) );
na02f01 g27182 ( .a(n30575), .b(n30443), .o(n30973) );
na02f01 g27183 ( .a(n30575), .b(delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n30974) );
na03f01 g27184 ( .a(n30974), .b(n30544), .c(n30442), .o(n30975) );
ao12f01 g27185 ( .a(n30597), .b(n30975), .c(n30973), .o(n30976) );
na03f01 g27186 ( .a(n30975), .b(n30973), .c(n30597), .o(n30977) );
in01f01 g27187 ( .a(n30977), .o(n30978) );
no02f01 g27188 ( .a(n30849), .b(n30841), .o(n30979) );
no02f01 g27189 ( .a(n30853), .b(n30979), .o(n30980) );
no02f01 g27190 ( .a(n30851), .b(n30701), .o(n30981) );
no02f01 g27191 ( .a(n30981), .b(n30980), .o(n30982) );
na02f01 g27192 ( .a(n30981), .b(n30980), .o(n30983) );
in01f01 g27193 ( .a(n30983), .o(n30984) );
no02f01 g27194 ( .a(n30984), .b(n30982), .o(n30985) );
in01f01 g27195 ( .a(n30985), .o(n30986) );
no03f01 g27196 ( .a(n30986), .b(n30978), .c(n30976), .o(n30987) );
in01f01 g27197 ( .a(n30987), .o(n30988) );
na02f01 g27198 ( .a(n30544), .b(n30441), .o(n30989) );
no02f01 g27199 ( .a(n30544), .b(n30441), .o(n30990) );
in01f01 g27200 ( .a(n30990), .o(n30991) );
na02f01 g27201 ( .a(n30991), .b(n30989), .o(n30992) );
in01f01 g27202 ( .a(n30838), .o(n30993) );
no02f01 g27203 ( .a(n30840), .b(n30709), .o(n30994) );
no02f01 g27204 ( .a(n30994), .b(n30993), .o(n30995) );
na02f01 g27205 ( .a(n30994), .b(n30993), .o(n30996) );
in01f01 g27206 ( .a(n30996), .o(n30997) );
no02f01 g27207 ( .a(n30997), .b(n30995), .o(n30998) );
in01f01 g27208 ( .a(n30998), .o(n30999) );
no02f01 g27209 ( .a(n30999), .b(n30992), .o(n31000) );
no02f01 g27210 ( .a(n30542), .b(n30536), .o(n31001) );
in01f01 g27211 ( .a(n31001), .o(n31002) );
na02f01 g27212 ( .a(n30542), .b(n30536), .o(n31003) );
no02f01 g27213 ( .a(n30833), .b(n30719), .o(n31004) );
in01f01 g27214 ( .a(n31004), .o(n31005) );
ao12f01 g27215 ( .a(n31005), .b(n30834), .c(n30831), .o(n31006) );
na02f01 g27216 ( .a(n30834), .b(n30831), .o(n31007) );
no02f01 g27217 ( .a(n31004), .b(n31007), .o(n31008) );
no02f01 g27218 ( .a(n31008), .b(n31006), .o(n31009) );
ao12f01 g27219 ( .a(n31009), .b(n31003), .c(n31002), .o(n31010) );
in01f01 g27220 ( .a(n30535), .o(n31011) );
no02f01 g27221 ( .a(n31011), .b(n30527), .o(n31012) );
na02f01 g27222 ( .a(n31011), .b(n30527), .o(n31013) );
in01f01 g27223 ( .a(n31013), .o(n31014) );
no02f01 g27224 ( .a(n30818), .b(n30810), .o(n31015) );
no02f01 g27225 ( .a(n30829), .b(n31015), .o(n31016) );
no02f01 g27226 ( .a(n30835), .b(n30827), .o(n31017) );
no02f01 g27227 ( .a(n31017), .b(n31016), .o(n31018) );
na02f01 g27228 ( .a(n31017), .b(n31016), .o(n31019) );
in01f01 g27229 ( .a(n31019), .o(n31020) );
no02f01 g27230 ( .a(n31020), .b(n31018), .o(n31021) );
in01f01 g27231 ( .a(n31021), .o(n31022) );
no03f01 g27232 ( .a(n31022), .b(n31014), .c(n31012), .o(n31023) );
na03f01 g27233 ( .a(n30525), .b(n30517), .c(delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n31024) );
ao12f01 g27234 ( .a(n30525), .b(n30517), .c(delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n31025) );
in01f01 g27235 ( .a(n31025), .o(n31026) );
in01f01 g27236 ( .a(n30810), .o(n31027) );
no02f01 g27237 ( .a(n30829), .b(n30818), .o(n31028) );
in01f01 g27238 ( .a(n31028), .o(n31029) );
no02f01 g27239 ( .a(n31029), .b(n31027), .o(n31030) );
no02f01 g27240 ( .a(n31028), .b(n30810), .o(n31031) );
no02f01 g27241 ( .a(n31031), .b(n31030), .o(n31032) );
ao12f01 g27242 ( .a(n31032), .b(n31026), .c(n31024), .o(n31033) );
in01f01 g27243 ( .a(n30516), .o(n31034) );
no02f01 g27244 ( .a(n31034), .b(n30508), .o(n31035) );
in01f01 g27245 ( .a(n30508), .o(n31036) );
no02f01 g27246 ( .a(n30516), .b(n31036), .o(n31037) );
no02f01 g27247 ( .a(n30805), .b(n30803), .o(n31038) );
no02f01 g27248 ( .a(n30807), .b(n30727), .o(n31039) );
no02f01 g27249 ( .a(n31039), .b(n31038), .o(n31040) );
na02f01 g27250 ( .a(n31039), .b(n31038), .o(n31041) );
in01f01 g27251 ( .a(n31041), .o(n31042) );
no02f01 g27252 ( .a(n31042), .b(n31040), .o(n31043) );
in01f01 g27253 ( .a(n31043), .o(n31044) );
no03f01 g27254 ( .a(n31044), .b(n31037), .c(n31035), .o(n31045) );
na02f01 g27255 ( .a(n30506), .b(n30499), .o(n31046) );
no02f01 g27256 ( .a(n30506), .b(n30499), .o(n31047) );
in01f01 g27257 ( .a(n31047), .o(n31048) );
no02f01 g27258 ( .a(n30794), .b(n30739), .o(n31049) );
in01f01 g27259 ( .a(n31049), .o(n31050) );
no02f01 g27260 ( .a(n30805), .b(n30802), .o(n31051) );
no02f01 g27261 ( .a(n31051), .b(n31050), .o(n31052) );
na02f01 g27262 ( .a(n31051), .b(n31050), .o(n31053) );
in01f01 g27263 ( .a(n31053), .o(n31054) );
no02f01 g27264 ( .a(n31054), .b(n31052), .o(n31055) );
ao12f01 g27265 ( .a(n31055), .b(n31048), .c(n31046), .o(n31056) );
no02f01 g27266 ( .a(n30497), .b(n30487), .o(n31057) );
in01f01 g27267 ( .a(n30447), .o(n31058) );
no02f01 g27268 ( .a(n30448), .b(n31058), .o(n31059) );
no02f01 g27269 ( .a(n31059), .b(n30443), .o(n31060) );
in01f01 g27270 ( .a(n30460), .o(n31061) );
in01f01 g27271 ( .a(n30465), .o(n31062) );
ao12f01 g27272 ( .a(n30443), .b(n31062), .c(n30463), .o(n31063) );
no03f01 g27273 ( .a(n31063), .b(n31061), .c(n30455), .o(n31064) );
no02f01 g27274 ( .a(n31064), .b(n30443), .o(n31065) );
in01f01 g27275 ( .a(n30474), .o(n31066) );
na02f01 g27276 ( .a(n30475), .b(n31066), .o(n31067) );
no03f01 g27277 ( .a(n31067), .b(n31065), .c(n31060), .o(n31068) );
in01f01 g27278 ( .a(n30485), .o(n31069) );
no02f01 g27279 ( .a(n31069), .b(n30483), .o(n31070) );
ao12f01 g27280 ( .a(n30443), .b(n31070), .c(n31068), .o(n31071) );
in01f01 g27281 ( .a(n30497), .o(n31072) );
no02f01 g27282 ( .a(n31072), .b(n31071), .o(n31073) );
no02f01 g27283 ( .a(n30790), .b(n30739), .o(n31074) );
in01f01 g27284 ( .a(n31074), .o(n31075) );
no03f01 g27285 ( .a(n31075), .b(n30791), .c(n30788), .o(n31076) );
no02f01 g27286 ( .a(n30791), .b(n30788), .o(n31077) );
no02f01 g27287 ( .a(n31074), .b(n31077), .o(n31078) );
no02f01 g27288 ( .a(n31078), .b(n31076), .o(n31079) );
in01f01 g27289 ( .a(n31079), .o(n31080) );
no03f01 g27290 ( .a(n31080), .b(n31073), .c(n31057), .o(n31081) );
ao12f01 g27291 ( .a(n31070), .b(n30478), .c(delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n31082) );
in01f01 g27292 ( .a(n31082), .o(n31083) );
na03f01 g27293 ( .a(n31070), .b(n30478), .c(delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n31084) );
in01f01 g27294 ( .a(n30778), .o(n31085) );
no02f01 g27295 ( .a(n30791), .b(n30787), .o(n31086) );
in01f01 g27296 ( .a(n31086), .o(n31087) );
no02f01 g27297 ( .a(n31087), .b(n31085), .o(n31088) );
no02f01 g27298 ( .a(n31086), .b(n30778), .o(n31089) );
no02f01 g27299 ( .a(n31089), .b(n31088), .o(n31090) );
ao12f01 g27300 ( .a(n31090), .b(n31084), .c(n31083), .o(n31091) );
no03f01 g27301 ( .a(n30486), .b(n31068), .c(n30443), .o(n31092) );
in01f01 g27302 ( .a(n31090), .o(n31093) );
no03f01 g27303 ( .a(n31093), .b(n31092), .c(n31082), .o(n31094) );
oa12f01 g27304 ( .a(n30477), .b(n31065), .c(n31060), .o(n31095) );
no03f01 g27305 ( .a(n30477), .b(n31065), .c(n31060), .o(n31096) );
in01f01 g27306 ( .a(n31096), .o(n31097) );
no03f01 g27307 ( .a(n30777), .b(n30775), .c(n30746), .o(n31098) );
in01f01 g27308 ( .a(n30775), .o(n31099) );
ao12f01 g27309 ( .a(n31099), .b(n30776), .c(n30747), .o(n31100) );
no02f01 g27310 ( .a(n31100), .b(n31098), .o(n31101) );
ao12f01 g27311 ( .a(n31101), .b(n31097), .c(n31095), .o(n31102) );
ao12f01 g27312 ( .a(n31059), .b(n30467), .c(delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n31103) );
no03f01 g27313 ( .a(n31064), .b(n30450), .c(n30443), .o(n31104) );
in01f01 g27314 ( .a(n30754), .o(n31105) );
in01f01 g27315 ( .a(n30773), .o(n31106) );
no03f01 g27316 ( .a(n30774), .b(n31106), .c(n31105), .o(n31107) );
in01f01 g27317 ( .a(n30774), .o(n31108) );
ao12f01 g27318 ( .a(n30773), .b(n31108), .c(n30754), .o(n31109) );
no02f01 g27319 ( .a(n31109), .b(n31107), .o(n31110) );
in01f01 g27320 ( .a(n31110), .o(n31111) );
oa12f01 g27321 ( .a(n31111), .b(n31104), .c(n31103), .o(n31112) );
no03f01 g27322 ( .a(n31111), .b(n31104), .c(n31103), .o(n31113) );
no02f01 g27323 ( .a(n30465), .b(n30464), .o(n31114) );
no02f01 g27324 ( .a(n30771), .b(delay_add_ln22_unr14_stage6_stallmux_q_0_), .o(n31115) );
no02f01 g27325 ( .a(n30770), .b(n30766), .o(n31116) );
no02f01 g27326 ( .a(n31116), .b(n31115), .o(n31117) );
no02f01 g27327 ( .a(n31117), .b(n31114), .o(n31118) );
in01f01 g27328 ( .a(n31118), .o(n31119) );
in01f01 g27329 ( .a(n30765), .o(n31120) );
no03f01 g27330 ( .a(n30772), .b(n31120), .c(n30764), .o(n31121) );
in01f01 g27331 ( .a(n30764), .o(n31122) );
in01f01 g27332 ( .a(n30772), .o(n31123) );
ao12f01 g27333 ( .a(n31123), .b(n30765), .c(n31122), .o(n31124) );
no02f01 g27334 ( .a(n31124), .b(n31121), .o(n31125) );
no02f01 g27335 ( .a(n31125), .b(n31119), .o(n31126) );
in01f01 g27336 ( .a(n31125), .o(n31127) );
no02f01 g27337 ( .a(n31127), .b(n31118), .o(n31128) );
in01f01 g27338 ( .a(n31128), .o(n31129) );
no02f01 g27339 ( .a(n31061), .b(n30455), .o(n31130) );
na02f01 g27340 ( .a(n31063), .b(n31130), .o(n31131) );
oa12f01 g27341 ( .a(n30466), .b(n31061), .c(n30455), .o(n31132) );
na02f01 g27342 ( .a(n31132), .b(n31131), .o(n31133) );
ao12f01 g27343 ( .a(n31126), .b(n31133), .c(n31129), .o(n31134) );
oa12f01 g27344 ( .a(n31112), .b(n31134), .c(n31113), .o(n31135) );
na03f01 g27345 ( .a(n31101), .b(n31097), .c(n31095), .o(n31136) );
ao12f01 g27346 ( .a(n31102), .b(n31136), .c(n31135), .o(n31137) );
no02f01 g27347 ( .a(n31137), .b(n31094), .o(n31138) );
na02f01 g27348 ( .a(n31072), .b(n31071), .o(n31139) );
na02f01 g27349 ( .a(n30497), .b(n30487), .o(n31140) );
ao12f01 g27350 ( .a(n31079), .b(n31140), .c(n31139), .o(n31141) );
no03f01 g27351 ( .a(n31141), .b(n31138), .c(n31091), .o(n31142) );
in01f01 g27352 ( .a(n31046), .o(n31143) );
in01f01 g27353 ( .a(n31055), .o(n31144) );
no03f01 g27354 ( .a(n31144), .b(n31047), .c(n31143), .o(n31145) );
no03f01 g27355 ( .a(n31145), .b(n31142), .c(n31081), .o(n31146) );
na02f01 g27356 ( .a(n30516), .b(n31036), .o(n31147) );
na02f01 g27357 ( .a(n31034), .b(n30508), .o(n31148) );
ao12f01 g27358 ( .a(n31043), .b(n31148), .c(n31147), .o(n31149) );
no03f01 g27359 ( .a(n31149), .b(n31146), .c(n31056), .o(n31150) );
in01f01 g27360 ( .a(n31024), .o(n31151) );
in01f01 g27361 ( .a(n31032), .o(n31152) );
no03f01 g27362 ( .a(n31152), .b(n31025), .c(n31151), .o(n31153) );
no03f01 g27363 ( .a(n31153), .b(n31150), .c(n31045), .o(n31154) );
in01f01 g27364 ( .a(n31012), .o(n31155) );
ao12f01 g27365 ( .a(n31021), .b(n31013), .c(n31155), .o(n31156) );
no03f01 g27366 ( .a(n31156), .b(n31154), .c(n31033), .o(n31157) );
in01f01 g27367 ( .a(n31003), .o(n31158) );
in01f01 g27368 ( .a(n31009), .o(n31159) );
no03f01 g27369 ( .a(n31159), .b(n31158), .c(n31001), .o(n31160) );
no03f01 g27370 ( .a(n31160), .b(n31157), .c(n31023), .o(n31161) );
ao12f01 g27371 ( .a(n30998), .b(n30991), .c(n30989), .o(n31162) );
no03f01 g27372 ( .a(n31162), .b(n31161), .c(n31010), .o(n31163) );
na02f01 g27373 ( .a(n30574), .b(n30545), .o(n31164) );
no02f01 g27374 ( .a(n30574), .b(n30545), .o(n31165) );
in01f01 g27375 ( .a(n31165), .o(n31166) );
na02f01 g27376 ( .a(n31166), .b(n31164), .o(n31167) );
no02f01 g27377 ( .a(n30853), .b(n30849), .o(n31168) );
no02f01 g27378 ( .a(n31168), .b(n30841), .o(n31169) );
na02f01 g27379 ( .a(n31168), .b(n30841), .o(n31170) );
in01f01 g27380 ( .a(n31170), .o(n31171) );
no02f01 g27381 ( .a(n31171), .b(n31169), .o(n31172) );
in01f01 g27382 ( .a(n31172), .o(n31173) );
no02f01 g27383 ( .a(n31173), .b(n31167), .o(n31174) );
no03f01 g27384 ( .a(n31174), .b(n31163), .c(n31000), .o(n31175) );
oa12f01 g27385 ( .a(n30986), .b(n30978), .c(n30976), .o(n31176) );
na02f01 g27386 ( .a(n31173), .b(n31167), .o(n31177) );
na02f01 g27387 ( .a(n31177), .b(n31176), .o(n31178) );
oa12f01 g27388 ( .a(n30988), .b(n31178), .c(n31175), .o(n31179) );
na02f01 g27389 ( .a(n30602), .b(n30593), .o(n31180) );
na03f01 g27390 ( .a(n30599), .b(n30591), .c(n30577), .o(n31181) );
na02f01 g27391 ( .a(n31181), .b(n31180), .o(n31182) );
na02f01 g27392 ( .a(n30855), .b(n30702), .o(n31183) );
in01f01 g27393 ( .a(n30856), .o(n31184) );
no02f01 g27394 ( .a(n31184), .b(n30685), .o(n31185) );
no02f01 g27395 ( .a(n31185), .b(n31183), .o(n31186) );
na02f01 g27396 ( .a(n31185), .b(n31183), .o(n31187) );
in01f01 g27397 ( .a(n31187), .o(n31188) );
no02f01 g27398 ( .a(n31188), .b(n31186), .o(n31189) );
in01f01 g27399 ( .a(n31189), .o(n31190) );
no02f01 g27400 ( .a(n31190), .b(n31182), .o(n31191) );
na02f01 g27401 ( .a(n30593), .b(delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n31192) );
na03f01 g27402 ( .a(n31192), .b(n30576), .c(n30546), .o(n31193) );
in01f01 g27403 ( .a(n31193), .o(n31194) );
ao12f01 g27404 ( .a(n30598), .b(n30593), .c(n30443), .o(n31195) );
in01f01 g27405 ( .a(n31195), .o(n31196) );
na02f01 g27406 ( .a(n30619), .b(n30443), .o(n31197) );
na02f01 g27407 ( .a(n30619), .b(delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n31198) );
na02f01 g27408 ( .a(n31198), .b(n31197), .o(n31199) );
oa12f01 g27409 ( .a(n31199), .b(n31196), .c(n31194), .o(n31200) );
no02f01 g27410 ( .a(n30616), .b(delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n31201) );
no02f01 g27411 ( .a(n30616), .b(n30443), .o(n31202) );
no02f01 g27412 ( .a(n31202), .b(n31201), .o(n31203) );
na03f01 g27413 ( .a(n31203), .b(n31195), .c(n31193), .o(n31204) );
no02f01 g27414 ( .a(n30859), .b(n30676), .o(n31205) );
in01f01 g27415 ( .a(n31205), .o(n31206) );
no02f01 g27416 ( .a(n31206), .b(n30879), .o(n31207) );
na02f01 g27417 ( .a(n31206), .b(n30879), .o(n31208) );
in01f01 g27418 ( .a(n31208), .o(n31209) );
no02f01 g27419 ( .a(n31209), .b(n31207), .o(n31210) );
ao12f01 g27420 ( .a(n31210), .b(n31204), .c(n31200), .o(n31211) );
ao12f01 g27421 ( .a(n31189), .b(n31181), .c(n31180), .o(n31212) );
no02f01 g27422 ( .a(n31212), .b(n31211), .o(n31213) );
oa12f01 g27423 ( .a(n31213), .b(n31191), .c(n31179), .o(n31214) );
ao12f01 g27424 ( .a(n31203), .b(n31195), .c(n31193), .o(n31215) );
no03f01 g27425 ( .a(n31199), .b(n31196), .c(n31194), .o(n31216) );
in01f01 g27426 ( .a(n31210), .o(n31217) );
no03f01 g27427 ( .a(n31217), .b(n31216), .c(n31215), .o(n31218) );
in01f01 g27428 ( .a(n31218), .o(n31219) );
no02f01 g27429 ( .a(n30882), .b(n30881), .o(n31220) );
no02f01 g27430 ( .a(n30876), .b(n30874), .o(n31221) );
no02f01 g27431 ( .a(n31221), .b(n31220), .o(n31222) );
na02f01 g27432 ( .a(n31222), .b(n30622), .o(n31223) );
in01f01 g27433 ( .a(n30869), .o(n31224) );
ao12f01 g27434 ( .a(n30868), .b(n30862), .c(n30667), .o(n31225) );
no02f01 g27435 ( .a(n31225), .b(n31224), .o(n31226) );
na02f01 g27436 ( .a(n31226), .b(n30622), .o(n31227) );
na02f01 g27437 ( .a(n31227), .b(n31223), .o(n31228) );
in01f01 g27438 ( .a(n31228), .o(n31229) );
in01f01 g27439 ( .a(n30622), .o(n31230) );
in01f01 g27440 ( .a(n30895), .o(n31231) );
na02f01 g27441 ( .a(n31231), .b(n30901), .o(n31232) );
na02f01 g27442 ( .a(n31232), .b(n30896), .o(n31233) );
no02f01 g27443 ( .a(n31233), .b(n31230), .o(n31234) );
in01f01 g27444 ( .a(n31234), .o(n31235) );
na04f01 g27445 ( .a(n31235), .b(n31229), .c(n31219), .d(n31214), .o(n31236) );
in01f01 g27446 ( .a(n30911), .o(n31237) );
no02f01 g27447 ( .a(n31237), .b(n31230), .o(n31238) );
no02f01 g27448 ( .a(n31238), .b(n31236), .o(n31239) );
no02f01 g27449 ( .a(n30956), .b(n31230), .o(n31240) );
in01f01 g27450 ( .a(n31240), .o(n31241) );
in01f01 g27451 ( .a(n30968), .o(n31242) );
na02f01 g27452 ( .a(n31242), .b(n30966), .o(n31243) );
no02f01 g27453 ( .a(n31243), .b(n31230), .o(n31244) );
in01f01 g27454 ( .a(n30928), .o(n31245) );
in01f01 g27455 ( .a(n30939), .o(n31246) );
na02f01 g27456 ( .a(n31246), .b(n30937), .o(n31247) );
ao12f01 g27457 ( .a(n31230), .b(n31247), .c(n31245), .o(n31248) );
no02f01 g27458 ( .a(n31248), .b(n31244), .o(n31249) );
na02f01 g27459 ( .a(n31249), .b(n31241), .o(n31250) );
in01f01 g27460 ( .a(n31250), .o(n31251) );
ao12f01 g27461 ( .a(n30972), .b(n31251), .c(n31239), .o(n31252) );
in01f01 g27462 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_26_), .o(n31253) );
no02f01 g27463 ( .a(n30892), .b(n31253), .o(n31254) );
no02f01 g27464 ( .a(n30864), .b(delay_add_ln22_unr14_stage6_stallmux_q_26_), .o(n31255) );
no02f01 g27465 ( .a(n31255), .b(n31254), .o(n31256) );
in01f01 g27466 ( .a(n31256), .o(n31257) );
no03f01 g27467 ( .a(n30961), .b(n30950), .c(n30943), .o(n31258) );
in01f01 g27468 ( .a(n31258), .o(n31259) );
no02f01 g27469 ( .a(n30963), .b(n30959), .o(n31260) );
oa12f01 g27470 ( .a(n31260), .b(n31259), .c(n30919), .o(n31261) );
in01f01 g27471 ( .a(n31261), .o(n31262) );
ao12f01 g27472 ( .a(n30864), .b(delay_add_ln22_unr14_stage6_stallmux_q_25_), .c(delay_add_ln22_unr14_stage6_stallmux_q_24_), .o(n31263) );
no02f01 g27473 ( .a(n31263), .b(n31262), .o(n31264) );
in01f01 g27474 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_24_), .o(n31265) );
in01f01 g27475 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_25_), .o(n31266) );
ao12f01 g27476 ( .a(n30892), .b(n31266), .c(n31265), .o(n31267) );
no02f01 g27477 ( .a(n31267), .b(n31264), .o(n31268) );
in01f01 g27478 ( .a(n31268), .o(n31269) );
no02f01 g27479 ( .a(n31269), .b(n31257), .o(n31270) );
no02f01 g27480 ( .a(n31268), .b(n31256), .o(n31271) );
no02f01 g27481 ( .a(n31271), .b(n31270), .o(n31272) );
in01f01 g27482 ( .a(n31272), .o(n31273) );
no02f01 g27483 ( .a(n31273), .b(n31230), .o(n31274) );
in01f01 g27484 ( .a(n31274), .o(n31275) );
no02f01 g27485 ( .a(n30864), .b(delay_add_ln22_unr14_stage6_stallmux_q_27_), .o(n31276) );
in01f01 g27486 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_27_), .o(n31277) );
no02f01 g27487 ( .a(n30892), .b(n31277), .o(n31278) );
no02f01 g27488 ( .a(n31278), .b(n31276), .o(n31279) );
no03f01 g27489 ( .a(n31263), .b(n31262), .c(n31255), .o(n31280) );
no03f01 g27490 ( .a(n31280), .b(n31267), .c(n31254), .o(n31281) );
na02f01 g27491 ( .a(n31281), .b(n31279), .o(n31282) );
in01f01 g27492 ( .a(n31282), .o(n31283) );
no02f01 g27493 ( .a(n31281), .b(n31279), .o(n31284) );
no02f01 g27494 ( .a(n31284), .b(n31283), .o(n31285) );
in01f01 g27495 ( .a(n31285), .o(n31286) );
no02f01 g27496 ( .a(n31286), .b(n31230), .o(n31287) );
no02f01 g27497 ( .a(n30864), .b(delay_add_ln22_unr14_stage6_stallmux_q_25_), .o(n31288) );
no02f01 g27498 ( .a(n30892), .b(n31266), .o(n31289) );
no02f01 g27499 ( .a(n31289), .b(n31288), .o(n31290) );
no02f01 g27500 ( .a(n30892), .b(n31265), .o(n31291) );
no02f01 g27501 ( .a(n30864), .b(delay_add_ln22_unr14_stage6_stallmux_q_24_), .o(n31292) );
in01f01 g27502 ( .a(n31292), .o(n31293) );
ao12f01 g27503 ( .a(n31291), .b(n31293), .c(n31261), .o(n31294) );
no02f01 g27504 ( .a(n31294), .b(n31290), .o(n31295) );
na02f01 g27505 ( .a(n31294), .b(n31290), .o(n31296) );
in01f01 g27506 ( .a(n31296), .o(n31297) );
no02f01 g27507 ( .a(n31297), .b(n31295), .o(n31298) );
in01f01 g27508 ( .a(n31298), .o(n31299) );
no02f01 g27509 ( .a(n31292), .b(n31291), .o(n31300) );
no02f01 g27510 ( .a(n31300), .b(n31262), .o(n31301) );
na02f01 g27511 ( .a(n31300), .b(n31262), .o(n31302) );
in01f01 g27512 ( .a(n31302), .o(n31303) );
no02f01 g27513 ( .a(n31303), .b(n31301), .o(n31304) );
in01f01 g27514 ( .a(n31304), .o(n31305) );
ao12f01 g27515 ( .a(n31230), .b(n31305), .c(n31299), .o(n31306) );
no02f01 g27516 ( .a(n31306), .b(n31287), .o(n31307) );
na02f01 g27517 ( .a(n31307), .b(n31275), .o(n31308) );
no02f01 g27518 ( .a(n30864), .b(delay_add_ln22_unr14_stage6_stallmux_q_28_), .o(n31309) );
in01f01 g27519 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_28_), .o(n31310) );
no02f01 g27520 ( .a(n30892), .b(n31310), .o(n31311) );
no02f01 g27521 ( .a(n31311), .b(n31309), .o(n31312) );
in01f01 g27522 ( .a(n31312), .o(n31313) );
no03f01 g27523 ( .a(n31276), .b(n31263), .c(n31255), .o(n31314) );
in01f01 g27524 ( .a(n31314), .o(n31315) );
no02f01 g27525 ( .a(n31315), .b(n31262), .o(n31316) );
ao12f01 g27526 ( .a(n30892), .b(n31253), .c(n31277), .o(n31317) );
no02f01 g27527 ( .a(n31317), .b(n31267), .o(n31318) );
in01f01 g27528 ( .a(n31318), .o(n31319) );
no03f01 g27529 ( .a(n31319), .b(n31316), .c(n31313), .o(n31320) );
no02f01 g27530 ( .a(n31319), .b(n31316), .o(n31321) );
no02f01 g27531 ( .a(n31321), .b(n31312), .o(n31322) );
no02f01 g27532 ( .a(n31322), .b(n31320), .o(n31323) );
in01f01 g27533 ( .a(n31323), .o(n31324) );
no02f01 g27534 ( .a(n30864), .b(delay_add_ln22_unr14_stage6_stallmux_q_29_), .o(n31325) );
in01f01 g27535 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_29_), .o(n31326) );
no02f01 g27536 ( .a(n30892), .b(n31326), .o(n31327) );
no02f01 g27537 ( .a(n31327), .b(n31325), .o(n31328) );
no03f01 g27538 ( .a(n31319), .b(n31311), .c(n31261), .o(n31329) );
no03f01 g27539 ( .a(n31329), .b(n31315), .c(n31309), .o(n31330) );
in01f01 g27540 ( .a(n31330), .o(n31331) );
no02f01 g27541 ( .a(n31331), .b(n31328), .o(n31332) );
na02f01 g27542 ( .a(n31331), .b(n31328), .o(n31333) );
in01f01 g27543 ( .a(n31333), .o(n31334) );
no02f01 g27544 ( .a(n31334), .b(n31332), .o(n31335) );
in01f01 g27545 ( .a(n31335), .o(n31336) );
ao12f01 g27546 ( .a(n31230), .b(n31336), .c(n31324), .o(n31337) );
no02f01 g27547 ( .a(n30864), .b(delay_add_ln22_unr14_stage6_stallmux_q_30_), .o(n31338) );
in01f01 g27548 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_30_), .o(n31339) );
no02f01 g27549 ( .a(n30892), .b(n31339), .o(n31340) );
no02f01 g27550 ( .a(n31340), .b(n31338), .o(n31341) );
in01f01 g27551 ( .a(n31341), .o(n31342) );
ao12f01 g27552 ( .a(n30892), .b(n31310), .c(n31326), .o(n31343) );
no03f01 g27553 ( .a(n31343), .b(n31319), .c(n31261), .o(n31344) );
no02f01 g27554 ( .a(n31325), .b(n31309), .o(n31345) );
in01f01 g27555 ( .a(n31345), .o(n31346) );
no03f01 g27556 ( .a(n31346), .b(n31344), .c(n31315), .o(n31347) );
no02f01 g27557 ( .a(n31347), .b(n31342), .o(n31348) );
na02f01 g27558 ( .a(n31347), .b(n31342), .o(n31349) );
in01f01 g27559 ( .a(n31349), .o(n31350) );
no02f01 g27560 ( .a(n31350), .b(n31348), .o(n31351) );
in01f01 g27561 ( .a(n31351), .o(n31352) );
no02f01 g27562 ( .a(n31352), .b(n31230), .o(n31353) );
no04f01 g27563 ( .a(n31353), .b(n31337), .c(n31308), .d(n31252), .o(n31354) );
ao12f01 g27564 ( .a(n30622), .b(n31304), .c(n31298), .o(n31355) );
ao12f01 g27565 ( .a(n30622), .b(n31285), .c(n31272), .o(n31356) );
no02f01 g27566 ( .a(n31356), .b(n31355), .o(n31357) );
in01f01 g27567 ( .a(n31357), .o(n31358) );
no02f01 g27568 ( .a(n31336), .b(n31324), .o(n31359) );
ao12f01 g27569 ( .a(n30622), .b(n31359), .c(n31351), .o(n31360) );
no03f01 g27570 ( .a(n31360), .b(n31358), .c(n31354), .o(n31361) );
no02f01 g27571 ( .a(n30864), .b(delay_add_ln22_unr14_stage6_stallmux_q_31_), .o(n31362) );
na02f01 g27572 ( .a(n30864), .b(delay_add_ln22_unr14_stage6_stallmux_q_31_), .o(n31363) );
in01f01 g27573 ( .a(n31363), .o(n31364) );
no02f01 g27574 ( .a(n31364), .b(n31362), .o(n31365) );
in01f01 g27575 ( .a(n31365), .o(n31366) );
no04f01 g27576 ( .a(n31346), .b(n31338), .c(n31315), .d(n31262), .o(n31367) );
oa12f01 g27577 ( .a(n30864), .b(n31343), .c(delay_add_ln22_unr14_stage6_stallmux_q_30_), .o(n31368) );
na02f01 g27578 ( .a(n31368), .b(n31318), .o(n31369) );
no03f01 g27579 ( .a(n31369), .b(n31367), .c(n31366), .o(n31370) );
no02f01 g27580 ( .a(n31369), .b(n31367), .o(n31371) );
no02f01 g27581 ( .a(n31371), .b(n31365), .o(n31372) );
no02f01 g27582 ( .a(n31372), .b(n31370), .o(n31373) );
in01f01 g27583 ( .a(n31373), .o(n31374) );
no02f01 g27584 ( .a(n31374), .b(n31230), .o(n31375) );
no02f01 g27585 ( .a(n31373), .b(n30622), .o(n31376) );
no02f01 g27586 ( .a(n31376), .b(n31375), .o(n31377) );
no02f01 g27587 ( .a(n31377), .b(n31361), .o(n31378) );
na02f01 g27588 ( .a(n31377), .b(n31361), .o(n31379) );
in01f01 g27589 ( .a(n31379), .o(n31380) );
no02f01 g27590 ( .a(n31380), .b(n31378), .o(n31381) );
no02f01 g27591 ( .a(n30969), .b(n30622), .o(n31382) );
no02f01 g27592 ( .a(n31382), .b(n31244), .o(n31383) );
no02f01 g27593 ( .a(n30957), .b(n30622), .o(n31384) );
in01f01 g27594 ( .a(n31384), .o(n31385) );
in01f01 g27595 ( .a(n30942), .o(n31386) );
in01f01 g27596 ( .a(n31248), .o(n31387) );
ao12f01 g27597 ( .a(n31386), .b(n31387), .c(n31239), .o(n31388) );
na02f01 g27598 ( .a(n31388), .b(n31385), .o(n31389) );
na02f01 g27599 ( .a(n31389), .b(n31241), .o(n31390) );
na02f01 g27600 ( .a(n31390), .b(n31383), .o(n31391) );
in01f01 g27601 ( .a(n31383), .o(n31392) );
na03f01 g27602 ( .a(n31389), .b(n31392), .c(n31241), .o(n31393) );
ao12f01 g27603 ( .a(n6075), .b(n31393), .c(n31391), .o(n31394) );
no02f01 g27604 ( .a(n31245), .b(n31230), .o(n31395) );
no02f01 g27605 ( .a(n31395), .b(n30929), .o(n31396) );
in01f01 g27606 ( .a(n31396), .o(n31397) );
no03f01 g27607 ( .a(n31397), .b(n31239), .c(n30914), .o(n31398) );
no02f01 g27608 ( .a(n31239), .b(n30914), .o(n31399) );
no02f01 g27609 ( .a(n31396), .b(n31399), .o(n31400) );
no02f01 g27610 ( .a(n31400), .b(n31398), .o(n31401) );
no02f01 g27611 ( .a(n31401), .b(n6075), .o(n31402) );
in01f01 g27612 ( .a(n30886), .o(n31403) );
na03f01 g27613 ( .a(n31229), .b(n31219), .c(n31214), .o(n31404) );
no02f01 g27614 ( .a(n30899), .b(n30622), .o(n31405) );
no02f01 g27615 ( .a(n31234), .b(n31405), .o(n31406) );
na03f01 g27616 ( .a(n31406), .b(n31404), .c(n31403), .o(n31407) );
in01f01 g27617 ( .a(n31000), .o(n31408) );
in01f01 g27618 ( .a(n31010), .o(n31409) );
in01f01 g27619 ( .a(n31023), .o(n31410) );
in01f01 g27620 ( .a(n31033), .o(n31411) );
in01f01 g27621 ( .a(n31045), .o(n31412) );
in01f01 g27622 ( .a(n31056), .o(n31413) );
in01f01 g27623 ( .a(n31081), .o(n31414) );
in01f01 g27624 ( .a(n31091), .o(n31415) );
na02f01 g27625 ( .a(n31084), .b(n31083), .o(n31416) );
oa12f01 g27626 ( .a(n30450), .b(n31064), .c(n30443), .o(n31417) );
na03f01 g27627 ( .a(n30467), .b(n31059), .c(delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n31418) );
ao12f01 g27628 ( .a(n31110), .b(n31418), .c(n31417), .o(n31419) );
na03f01 g27629 ( .a(n31110), .b(n31418), .c(n31417), .o(n31420) );
in01f01 g27630 ( .a(n31126), .o(n31421) );
no03f01 g27631 ( .a(n30466), .b(n31061), .c(n30455), .o(n31422) );
in01f01 g27632 ( .a(n31132), .o(n31423) );
no02f01 g27633 ( .a(n31423), .b(n31422), .o(n31424) );
oa12f01 g27634 ( .a(n31421), .b(n31424), .c(n31128), .o(n31425) );
ao12f01 g27635 ( .a(n31419), .b(n31425), .c(n31420), .o(n31426) );
in01f01 g27636 ( .a(n31095), .o(n31427) );
in01f01 g27637 ( .a(n31101), .o(n31428) );
no03f01 g27638 ( .a(n31428), .b(n31096), .c(n31427), .o(n31429) );
no02f01 g27639 ( .a(n31429), .b(n31426), .o(n31430) );
oa22f01 g27640 ( .a(n31430), .b(n31102), .c(n31093), .d(n31416), .o(n31431) );
oa12f01 g27641 ( .a(n31080), .b(n31073), .c(n31057), .o(n31432) );
na03f01 g27642 ( .a(n31432), .b(n31431), .c(n31415), .o(n31433) );
na03f01 g27643 ( .a(n31055), .b(n31048), .c(n31046), .o(n31434) );
na03f01 g27644 ( .a(n31434), .b(n31433), .c(n31414), .o(n31435) );
oa12f01 g27645 ( .a(n31044), .b(n31037), .c(n31035), .o(n31436) );
na03f01 g27646 ( .a(n31436), .b(n31435), .c(n31413), .o(n31437) );
na03f01 g27647 ( .a(n31032), .b(n31026), .c(n31024), .o(n31438) );
na03f01 g27648 ( .a(n31438), .b(n31437), .c(n31412), .o(n31439) );
oa12f01 g27649 ( .a(n31022), .b(n31014), .c(n31012), .o(n31440) );
na03f01 g27650 ( .a(n31440), .b(n31439), .c(n31411), .o(n31441) );
na03f01 g27651 ( .a(n31009), .b(n31003), .c(n31002), .o(n31442) );
na03f01 g27652 ( .a(n31442), .b(n31441), .c(n31410), .o(n31443) );
na02f01 g27653 ( .a(n30999), .b(n30992), .o(n31444) );
na03f01 g27654 ( .a(n31444), .b(n31443), .c(n31409), .o(n31445) );
in01f01 g27655 ( .a(n31164), .o(n31446) );
no02f01 g27656 ( .a(n31165), .b(n31446), .o(n31447) );
na02f01 g27657 ( .a(n31172), .b(n31447), .o(n31448) );
na03f01 g27658 ( .a(n31448), .b(n31445), .c(n31408), .o(n31449) );
in01f01 g27659 ( .a(n30976), .o(n31450) );
ao12f01 g27660 ( .a(n30985), .b(n30977), .c(n31450), .o(n31451) );
no02f01 g27661 ( .a(n31172), .b(n31447), .o(n31452) );
no02f01 g27662 ( .a(n31452), .b(n31451), .o(n31453) );
ao12f01 g27663 ( .a(n30987), .b(n31453), .c(n31449), .o(n31454) );
in01f01 g27664 ( .a(n31191), .o(n31455) );
oa12f01 g27665 ( .a(n31217), .b(n31216), .c(n31215), .o(n31456) );
in01f01 g27666 ( .a(n31212), .o(n31457) );
na02f01 g27667 ( .a(n31457), .b(n31456), .o(n31458) );
ao12f01 g27668 ( .a(n31458), .b(n31455), .c(n31454), .o(n31459) );
no03f01 g27669 ( .a(n31228), .b(n31218), .c(n31459), .o(n31460) );
in01f01 g27670 ( .a(n31406), .o(n31461) );
oa12f01 g27671 ( .a(n31461), .b(n31460), .c(n30886), .o(n31462) );
na02f01 g27672 ( .a(n31462), .b(n31407), .o(n31463) );
na02f01 g27673 ( .a(n30873), .b(n31230), .o(n31464) );
na02f01 g27674 ( .a(n31464), .b(n31227), .o(n31465) );
in01f01 g27675 ( .a(n31465), .o(n31466) );
no02f01 g27676 ( .a(n31222), .b(n30622), .o(n31467) );
in01f01 g27677 ( .a(n31467), .o(n31468) );
na03f01 g27678 ( .a(n31223), .b(n31219), .c(n31214), .o(n31469) );
na03f01 g27679 ( .a(n31469), .b(n31468), .c(n31466), .o(n31470) );
in01f01 g27680 ( .a(n31223), .o(n31471) );
no03f01 g27681 ( .a(n31471), .b(n31218), .c(n31459), .o(n31472) );
oa12f01 g27682 ( .a(n31465), .b(n31472), .c(n31467), .o(n31473) );
na02f01 g27683 ( .a(n31473), .b(n31470), .o(n31474) );
oa12f01 g27684 ( .a(n_22641), .b(n31474), .c(n31463), .o(n31475) );
no02f01 g27685 ( .a(n31405), .b(n30886), .o(n31476) );
no02f01 g27686 ( .a(n30911), .b(n30622), .o(n31477) );
no02f01 g27687 ( .a(n31477), .b(n31238), .o(n31478) );
ao12f01 g27688 ( .a(n31478), .b(n31476), .c(n31236), .o(n31479) );
na03f01 g27689 ( .a(n31478), .b(n31476), .c(n31236), .o(n31480) );
in01f01 g27690 ( .a(n31480), .o(n31481) );
oa12f01 g27691 ( .a(n_22641), .b(n31481), .c(n31479), .o(n31482) );
na02f01 g27692 ( .a(n31482), .b(n31475), .o(n31483) );
no02f01 g27693 ( .a(n31483), .b(n31402), .o(n31484) );
no02f01 g27694 ( .a(n31481), .b(n31479), .o(n31485) );
ao12f01 g27695 ( .a(n_22641), .b(n31485), .c(n31401), .o(n31486) );
no02f01 g27696 ( .a(n31486), .b(n31484), .o(n31487) );
in01f01 g27697 ( .a(n30929), .o(n31488) );
in01f01 g27698 ( .a(n31395), .o(n31489) );
oa12f01 g27699 ( .a(n31489), .b(n31239), .c(n30914), .o(n31490) );
no02f01 g27700 ( .a(n31247), .b(n31230), .o(n31491) );
no02f01 g27701 ( .a(n31491), .b(n30941), .o(n31492) );
na03f01 g27702 ( .a(n31492), .b(n31490), .c(n31488), .o(n31493) );
ao12f01 g27703 ( .a(n31492), .b(n31490), .c(n31488), .o(n31494) );
in01f01 g27704 ( .a(n31494), .o(n31495) );
ao12f01 g27705 ( .a(n6075), .b(n31495), .c(n31493), .o(n31496) );
in01f01 g27706 ( .a(n31388), .o(n31497) );
no02f01 g27707 ( .a(n31240), .b(n31384), .o(n31498) );
in01f01 g27708 ( .a(n31498), .o(n31499) );
no02f01 g27709 ( .a(n31499), .b(n31497), .o(n31500) );
no02f01 g27710 ( .a(n31498), .b(n31388), .o(n31501) );
no02f01 g27711 ( .a(n31501), .b(n31500), .o(n31502) );
no02f01 g27712 ( .a(n31502), .b(n6075), .o(n31503) );
no04f01 g27713 ( .a(n31503), .b(n31496), .c(n31487), .d(n31394), .o(n31504) );
no02f01 g27714 ( .a(n31304), .b(n30622), .o(n31505) );
no02f01 g27715 ( .a(n31305), .b(n31230), .o(n31506) );
no02f01 g27716 ( .a(n31506), .b(n31505), .o(n31507) );
no02f01 g27717 ( .a(n31507), .b(n31252), .o(n31508) );
na02f01 g27718 ( .a(n31507), .b(n31252), .o(n31509) );
in01f01 g27719 ( .a(n31509), .o(n31510) );
no02f01 g27720 ( .a(n31510), .b(n31508), .o(n31511) );
no02f01 g27721 ( .a(n31511), .b(n6075), .o(n31512) );
in01f01 g27722 ( .a(n31512), .o(n31513) );
in01f01 g27723 ( .a(n31493), .o(n31514) );
no02f01 g27724 ( .a(n31494), .b(n31514), .o(n31515) );
ao12f01 g27725 ( .a(n_22641), .b(n31502), .c(n31515), .o(n31516) );
in01f01 g27726 ( .a(n31516), .o(n31517) );
na02f01 g27727 ( .a(n31393), .b(n31391), .o(n31518) );
in01f01 g27728 ( .a(n31511), .o(n31519) );
oa12f01 g27729 ( .a(n6075), .b(n31519), .c(n31518), .o(n31520) );
na02f01 g27730 ( .a(n31520), .b(n31517), .o(n31521) );
ao12f01 g27731 ( .a(n31521), .b(n31513), .c(n31504), .o(n31522) );
no02f01 g27732 ( .a(n31299), .b(n31230), .o(n31523) );
no02f01 g27733 ( .a(n31298), .b(n30622), .o(n31524) );
no02f01 g27734 ( .a(n31524), .b(n31523), .o(n31525) );
in01f01 g27735 ( .a(n31525), .o(n31526) );
in01f01 g27736 ( .a(n31505), .o(n31527) );
oa12f01 g27737 ( .a(n31527), .b(n31506), .c(n31252), .o(n31528) );
no02f01 g27738 ( .a(n31528), .b(n31526), .o(n31529) );
na02f01 g27739 ( .a(n31528), .b(n31526), .o(n31530) );
in01f01 g27740 ( .a(n31530), .o(n31531) );
no02f01 g27741 ( .a(n31531), .b(n31529), .o(n31532) );
no02f01 g27742 ( .a(n31532), .b(n6075), .o(n31533) );
no02f01 g27743 ( .a(n31533), .b(n31522), .o(n31534) );
no02f01 g27744 ( .a(n31272), .b(n30622), .o(n31535) );
no02f01 g27745 ( .a(n31535), .b(n31274), .o(n31536) );
in01f01 g27746 ( .a(n31536), .o(n31537) );
in01f01 g27747 ( .a(n30972), .o(n31538) );
no02f01 g27748 ( .a(n31306), .b(n31250), .o(n31539) );
na02f01 g27749 ( .a(n31539), .b(n31239), .o(n31540) );
na02f01 g27750 ( .a(n31540), .b(n31538), .o(n31541) );
no03f01 g27751 ( .a(n31541), .b(n31537), .c(n31355), .o(n31542) );
no02f01 g27752 ( .a(n31541), .b(n31355), .o(n31543) );
no02f01 g27753 ( .a(n31543), .b(n31536), .o(n31544) );
no02f01 g27754 ( .a(n31544), .b(n31542), .o(n31545) );
no02f01 g27755 ( .a(n31545), .b(n6075), .o(n31546) );
in01f01 g27756 ( .a(n31546), .o(n31547) );
na02f01 g27757 ( .a(n31541), .b(n31275), .o(n31548) );
no02f01 g27758 ( .a(n31535), .b(n31355), .o(n31549) );
na02f01 g27759 ( .a(n31549), .b(n31548), .o(n31550) );
no02f01 g27760 ( .a(n31285), .b(n30622), .o(n31551) );
no02f01 g27761 ( .a(n31551), .b(n31287), .o(n31552) );
in01f01 g27762 ( .a(n31552), .o(n31553) );
no02f01 g27763 ( .a(n31553), .b(n31550), .o(n31554) );
na02f01 g27764 ( .a(n31553), .b(n31550), .o(n31555) );
in01f01 g27765 ( .a(n31555), .o(n31556) );
no02f01 g27766 ( .a(n31556), .b(n31554), .o(n31557) );
no02f01 g27767 ( .a(n31557), .b(n6075), .o(n31558) );
in01f01 g27768 ( .a(n31558), .o(n31559) );
na03f01 g27769 ( .a(n31559), .b(n31547), .c(n31534), .o(n31560) );
oa12f01 g27770 ( .a(n31357), .b(n31308), .c(n31252), .o(n31561) );
no02f01 g27771 ( .a(n31324), .b(n31230), .o(n31562) );
no02f01 g27772 ( .a(n31323), .b(n30622), .o(n31563) );
no02f01 g27773 ( .a(n31563), .b(n31562), .o(n31564) );
in01f01 g27774 ( .a(n31564), .o(n31565) );
no02f01 g27775 ( .a(n31565), .b(n31561), .o(n31566) );
in01f01 g27776 ( .a(n31561), .o(n31567) );
no02f01 g27777 ( .a(n31564), .b(n31567), .o(n31568) );
no02f01 g27778 ( .a(n31568), .b(n31566), .o(n31569) );
no02f01 g27779 ( .a(n31569), .b(n6075), .o(n31570) );
no02f01 g27780 ( .a(n31570), .b(n31560), .o(n31571) );
ao12f01 g27781 ( .a(n_22641), .b(n31545), .c(n31532), .o(n31572) );
ao12f01 g27782 ( .a(n_22641), .b(n31569), .c(n31557), .o(n31573) );
no02f01 g27783 ( .a(n31573), .b(n31572), .o(n31574) );
in01f01 g27784 ( .a(n31574), .o(n31575) );
no02f01 g27785 ( .a(n31575), .b(n31571), .o(n31576) );
in01f01 g27786 ( .a(n31562), .o(n31577) );
ao12f01 g27787 ( .a(n31563), .b(n31577), .c(n31561), .o(n31578) );
in01f01 g27788 ( .a(n31578), .o(n31579) );
no02f01 g27789 ( .a(n31336), .b(n31230), .o(n31580) );
no02f01 g27790 ( .a(n31335), .b(n30622), .o(n31581) );
no02f01 g27791 ( .a(n31581), .b(n31580), .o(n31582) );
in01f01 g27792 ( .a(n31582), .o(n31583) );
no02f01 g27793 ( .a(n31583), .b(n31579), .o(n31584) );
no02f01 g27794 ( .a(n31582), .b(n31578), .o(n31585) );
no02f01 g27795 ( .a(n31585), .b(n31584), .o(n31586) );
no02f01 g27796 ( .a(n31351), .b(n30622), .o(n31587) );
no02f01 g27797 ( .a(n31587), .b(n31353), .o(n31588) );
in01f01 g27798 ( .a(n31588), .o(n31589) );
in01f01 g27799 ( .a(n31337), .o(n31590) );
no02f01 g27800 ( .a(n31359), .b(n30622), .o(n31591) );
ao12f01 g27801 ( .a(n31591), .b(n31561), .c(n31590), .o(n31592) );
in01f01 g27802 ( .a(n31592), .o(n31593) );
no02f01 g27803 ( .a(n31593), .b(n31589), .o(n31594) );
no02f01 g27804 ( .a(n31592), .b(n31588), .o(n31595) );
no02f01 g27805 ( .a(n31595), .b(n31594), .o(n31596) );
ao12f01 g27806 ( .a(n6075), .b(n31596), .c(n31586), .o(n31597) );
no02f01 g27807 ( .a(n31597), .b(n31576), .o(n31598) );
ao12f01 g27808 ( .a(n_22641), .b(n31596), .c(n31586), .o(n31599) );
no02f01 g27809 ( .a(n31381), .b(n_22641), .o(n31600) );
no02f01 g27810 ( .a(n31381), .b(n6075), .o(n31601) );
no02f01 g27811 ( .a(n31381), .b(n_22641), .o(n31602) );
in01f01 g27812 ( .a(n31599), .o(n31603) );
ao12f01 g27813 ( .a(n_22641), .b(n31603), .c(n31381), .o(n31604) );
no04f01 g27814 ( .a(n31604), .b(n31598), .c(n31602), .d(n31601), .o(n31605) );
no02f01 g27815 ( .a(n31605), .b(n31600), .o(n31606) );
in01f01 g27816 ( .a(n31606), .o(n31607) );
na02f01 g27817 ( .a(n31233), .b(delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n31608) );
ao12f01 g27818 ( .a(n30443), .b(n30872), .c(n30869), .o(n31609) );
no02f01 g27819 ( .a(n31222), .b(n30443), .o(n31610) );
no02f01 g27820 ( .a(n31610), .b(n31609), .o(n31611) );
na02f01 g27821 ( .a(n31611), .b(n31608), .o(n31612) );
oa12f01 g27822 ( .a(n30443), .b(n30910), .c(n30909), .o(n31613) );
in01f01 g27823 ( .a(n30910), .o(n31614) );
na03f01 g27824 ( .a(n31614), .b(n30908), .c(delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n31615) );
ao12f01 g27825 ( .a(n31612), .b(n31615), .c(n31613), .o(n31616) );
no02f01 g27826 ( .a(n31233), .b(n30443), .o(n31617) );
no02f01 g27827 ( .a(n30899), .b(delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n31618) );
no02f01 g27828 ( .a(n31618), .b(n31617), .o(n31619) );
na04f01 g27829 ( .a(n31615), .b(n31613), .c(n31612), .d(n31619), .o(n31620) );
ao12f01 g27830 ( .a(n31616), .b(n31620), .c(n30443), .o(n31621) );
ao12f01 g27831 ( .a(n30443), .b(n30940), .c(n30928), .o(n31622) );
na02f01 g27832 ( .a(n30956), .b(delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n31623) );
in01f01 g27833 ( .a(n31623), .o(n31624) );
no03f01 g27834 ( .a(n31624), .b(n31622), .c(n31621), .o(n31625) );
no02f01 g27835 ( .a(n31243), .b(n30443), .o(n31626) );
no02f01 g27836 ( .a(n30969), .b(delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n31627) );
no02f01 g27837 ( .a(n31627), .b(n31626), .o(n31628) );
na02f01 g27838 ( .a(n30956), .b(n30443), .o(n31629) );
na02f01 g27839 ( .a(n31629), .b(n31628), .o(n31630) );
oa12f01 g27840 ( .a(n30443), .b(n31630), .c(n31625), .o(n31631) );
na02f01 g27841 ( .a(n30969), .b(delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n31632) );
na02f01 g27842 ( .a(n31243), .b(n30443), .o(n31633) );
na02f01 g27843 ( .a(n31633), .b(n31632), .o(n31634) );
ao12f01 g27844 ( .a(delay_sub_ln23_0_unr15_stage6_stallmux_q), .b(n30940), .c(n30928), .o(n31635) );
ao12f01 g27845 ( .a(n31635), .b(n31634), .c(n31625), .o(n31636) );
na02f01 g27846 ( .a(n31636), .b(n31631), .o(n31637) );
ao12f01 g27847 ( .a(n30443), .b(n31304), .c(n31298), .o(n31638) );
no02f01 g27848 ( .a(n31272), .b(n30443), .o(n31639) );
no02f01 g27849 ( .a(n31639), .b(n31638), .o(n31640) );
na02f01 g27850 ( .a(n31640), .b(n31637), .o(n31641) );
no02f01 g27851 ( .a(n31285), .b(n30443), .o(n31642) );
no02f01 g27852 ( .a(n31642), .b(n31641), .o(n31643) );
ao12f01 g27853 ( .a(delay_sub_ln23_0_unr15_stage6_stallmux_q), .b(n31304), .c(n31298), .o(n31644) );
ao12f01 g27854 ( .a(delay_sub_ln23_0_unr15_stage6_stallmux_q), .b(n31285), .c(n31272), .o(n31645) );
no02f01 g27855 ( .a(n31645), .b(n31644), .o(n31646) );
in01f01 g27856 ( .a(n31646), .o(n31647) );
no02f01 g27857 ( .a(n31647), .b(n31643), .o(n31648) );
ao12f01 g27858 ( .a(n30443), .b(n31335), .c(n31323), .o(n31649) );
no02f01 g27859 ( .a(n31649), .b(n31648), .o(n31650) );
in01f01 g27860 ( .a(n31650), .o(n31651) );
no02f01 g27861 ( .a(n31335), .b(delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n31652) );
no02f01 g27862 ( .a(n31336), .b(n30443), .o(n31653) );
no02f01 g27863 ( .a(n31323), .b(delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n31654) );
no03f01 g27864 ( .a(n31654), .b(n31653), .c(n31652), .o(n31655) );
no03f01 g27865 ( .a(n31651), .b(n31352), .c(n30443), .o(n31656) );
no02f01 g27866 ( .a(n31655), .b(delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n31657) );
no03f01 g27867 ( .a(n31657), .b(n31352), .c(delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n31658) );
no02f01 g27868 ( .a(n31373), .b(delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n31659) );
no02f01 g27869 ( .a(n31374), .b(n30443), .o(n31660) );
no02f01 g27870 ( .a(n31660), .b(n31659), .o(n31661) );
in01f01 g27871 ( .a(n31661), .o(n31662) );
ao12f01 g27872 ( .a(n31662), .b(n31658), .c(n31651), .o(n31663) );
no02f01 g27873 ( .a(n31663), .b(n31656), .o(n31664) );
no02f01 g27874 ( .a(n31664), .b(n30525), .o(n31665) );
in01f01 g27875 ( .a(n31664), .o(n31666) );
no02f01 g27876 ( .a(n31666), .b(n30526), .o(n31667) );
no02f01 g27877 ( .a(n31667), .b(n31665), .o(n31668) );
in01f01 g27878 ( .a(n31668), .o(n31669) );
ao12f01 g27879 ( .a(n31664), .b(n31114), .c(n31130), .o(n31670) );
ao12f01 g27880 ( .a(n31664), .b(n30477), .c(n31059), .o(n31671) );
no02f01 g27881 ( .a(n31671), .b(n31670), .o(n31672) );
in01f01 g27882 ( .a(n31672), .o(n31673) );
no02f01 g27883 ( .a(n31373), .b(n30443), .o(n31674) );
no02f01 g27884 ( .a(n31373), .b(delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n31675) );
no02f01 g27885 ( .a(n31675), .b(n31674), .o(n31676) );
no02f01 g27886 ( .a(n31351), .b(n30443), .o(n31677) );
in01f01 g27887 ( .a(n31643), .o(n31678) );
no02f01 g27888 ( .a(n31657), .b(n31647), .o(n31679) );
oa12f01 g27889 ( .a(n31679), .b(n31649), .c(n31678), .o(n31680) );
ao12f01 g27890 ( .a(n31680), .b(n31352), .c(n30443), .o(n31681) );
no03f01 g27891 ( .a(n31681), .b(n31677), .c(n31676), .o(n31682) );
in01f01 g27892 ( .a(n31676), .o(n31683) );
ao12f01 g27893 ( .a(n31681), .b(n31352), .c(delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n31684) );
no02f01 g27894 ( .a(n31684), .b(n31683), .o(n31685) );
no02f01 g27895 ( .a(n31685), .b(n31682), .o(n31686) );
in01f01 g27896 ( .a(n30362), .o(n31687) );
no02f01 g27897 ( .a(n31687), .b(n30202), .o(n31688) );
in01f01 g27898 ( .a(n31688), .o(n31689) );
ao12f01 g27899 ( .a(n30371), .b(n30384), .c(n31689), .o(n31690) );
in01f01 g27900 ( .a(n31690), .o(n31691) );
no02f01 g27901 ( .a(n30387), .b(n30383), .o(n31692) );
no02f01 g27902 ( .a(n31692), .b(n31691), .o(n31693) );
na02f01 g27903 ( .a(n31692), .b(n31691), .o(n31694) );
in01f01 g27904 ( .a(n31694), .o(n31695) );
no02f01 g27905 ( .a(n31695), .b(n31693), .o(n31696) );
in01f01 g27906 ( .a(n31696), .o(n31697) );
no02f01 g27907 ( .a(n31697), .b(n31686), .o(n31698) );
no02f01 g27908 ( .a(n31323), .b(n30443), .o(n31699) );
in01f01 g27909 ( .a(n31699), .o(n31700) );
no02f01 g27910 ( .a(n31654), .b(n31647), .o(n31701) );
in01f01 g27911 ( .a(n31701), .o(n31702) );
ao12f01 g27912 ( .a(n31702), .b(n31700), .c(n31643), .o(n31703) );
na02f01 g27913 ( .a(n31703), .b(n31335), .o(n31704) );
in01f01 g27914 ( .a(n31704), .o(n31705) );
no02f01 g27915 ( .a(n31703), .b(n31335), .o(n31706) );
in01f01 g27916 ( .a(n30360), .o(n31707) );
in01f01 g27917 ( .a(n30361), .o(n31708) );
no02f01 g27918 ( .a(n31708), .b(n30202), .o(n31709) );
in01f01 g27919 ( .a(n31709), .o(n31710) );
no03f01 g27920 ( .a(n31710), .b(n31707), .c(n30222), .o(n31711) );
ao12f01 g27921 ( .a(n31709), .b(n30360), .c(n30223), .o(n31712) );
no02f01 g27922 ( .a(n31712), .b(n31711), .o(n31713) );
no03f01 g27923 ( .a(n31713), .b(n31706), .c(n31705), .o(n31714) );
in01f01 g27924 ( .a(n30357), .o(n31715) );
no02f01 g27925 ( .a(n31715), .b(n30229), .o(n31716) );
no02f01 g27926 ( .a(n30358), .b(n30222), .o(n31717) );
in01f01 g27927 ( .a(n31717), .o(n31718) );
no02f01 g27928 ( .a(n31718), .b(n31716), .o(n31719) );
na02f01 g27929 ( .a(n31718), .b(n31716), .o(n31720) );
in01f01 g27930 ( .a(n31720), .o(n31721) );
no02f01 g27931 ( .a(n31721), .b(n31719), .o(n31722) );
no02f01 g27932 ( .a(n31654), .b(n31699), .o(n31723) );
na02f01 g27933 ( .a(n31723), .b(n31648), .o(n31724) );
no02f01 g27934 ( .a(n31723), .b(n31648), .o(n31725) );
in01f01 g27935 ( .a(n31725), .o(n31726) );
na02f01 g27936 ( .a(n31726), .b(n31724), .o(n31727) );
no02f01 g27937 ( .a(n31727), .b(n31722), .o(n31728) );
oa12f01 g27938 ( .a(n31713), .b(n31706), .c(n31705), .o(n31729) );
oa12f01 g27939 ( .a(n31729), .b(n31728), .c(n31714), .o(n31730) );
no02f01 g27940 ( .a(n31285), .b(delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n31731) );
no02f01 g27941 ( .a(n31731), .b(n31642), .o(n31732) );
in01f01 g27942 ( .a(n31732), .o(n31733) );
no02f01 g27943 ( .a(n31272), .b(delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n31734) );
no02f01 g27944 ( .a(n31734), .b(n31644), .o(n31735) );
na02f01 g27945 ( .a(n31735), .b(n31641), .o(n31736) );
no02f01 g27946 ( .a(n31736), .b(n31733), .o(n31737) );
ao12f01 g27947 ( .a(n31732), .b(n31735), .c(n31641), .o(n31738) );
no02f01 g27948 ( .a(n31738), .b(n31737), .o(n31739) );
in01f01 g27949 ( .a(n30355), .o(n31740) );
in01f01 g27950 ( .a(n30356), .o(n31741) );
no02f01 g27951 ( .a(n31741), .b(n30229), .o(n31742) );
in01f01 g27952 ( .a(n31742), .o(n31743) );
no03f01 g27953 ( .a(n31743), .b(n31740), .c(n30240), .o(n31744) );
ao12f01 g27954 ( .a(n31742), .b(n30355), .c(n30241), .o(n31745) );
no02f01 g27955 ( .a(n31745), .b(n31744), .o(n31746) );
in01f01 g27956 ( .a(n31746), .o(n31747) );
no02f01 g27957 ( .a(n31747), .b(n31739), .o(n31748) );
in01f01 g27958 ( .a(n31748), .o(n31749) );
no02f01 g27959 ( .a(n31734), .b(n31639), .o(n31750) );
in01f01 g27960 ( .a(n31638), .o(n31751) );
ao12f01 g27961 ( .a(n31644), .b(n31751), .c(n31637), .o(n31752) );
na02f01 g27962 ( .a(n31752), .b(n31750), .o(n31753) );
no02f01 g27963 ( .a(n31752), .b(n31750), .o(n31754) );
in01f01 g27964 ( .a(n31754), .o(n31755) );
na02f01 g27965 ( .a(n31755), .b(n31753), .o(n31756) );
no02f01 g27966 ( .a(n30353), .b(n30240), .o(n31757) );
in01f01 g27967 ( .a(n31757), .o(n31758) );
no03f01 g27968 ( .a(n31758), .b(n30352), .c(n30262), .o(n31759) );
no02f01 g27969 ( .a(n30352), .b(n30262), .o(n31760) );
no02f01 g27970 ( .a(n31757), .b(n31760), .o(n31761) );
no02f01 g27971 ( .a(n31761), .b(n31759), .o(n31762) );
no02f01 g27972 ( .a(n31762), .b(n31756), .o(n31763) );
in01f01 g27973 ( .a(n31763), .o(n31764) );
no02f01 g27974 ( .a(n31304), .b(delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n31765) );
in01f01 g27975 ( .a(n31765), .o(n31766) );
in01f01 g27976 ( .a(n31616), .o(n31767) );
oa12f01 g27977 ( .a(delay_sub_ln23_0_unr15_stage6_stallmux_q), .b(n31225), .c(n31224), .o(n31768) );
na02f01 g27978 ( .a(n30884), .b(delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n31769) );
na02f01 g27979 ( .a(n31769), .b(n31768), .o(n31770) );
oa12f01 g27980 ( .a(n31619), .b(n31770), .c(delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n31771) );
oa12f01 g27981 ( .a(n30443), .b(n31771), .c(n31237), .o(n31772) );
na02f01 g27982 ( .a(n31772), .b(n31767), .o(n31773) );
oa12f01 g27983 ( .a(delay_sub_ln23_0_unr15_stage6_stallmux_q), .b(n31247), .c(n31245), .o(n31774) );
na03f01 g27984 ( .a(n31623), .b(n31774), .c(n31773), .o(n31775) );
ao12f01 g27985 ( .a(n31634), .b(n30956), .c(n30443), .o(n31776) );
ao12f01 g27986 ( .a(delay_sub_ln23_0_unr15_stage6_stallmux_q), .b(n31776), .c(n31775), .o(n31777) );
in01f01 g27987 ( .a(n31635), .o(n31778) );
oa12f01 g27988 ( .a(n31778), .b(n31628), .c(n31775), .o(n31779) );
oa22f01 g27989 ( .a(n31779), .b(n31777), .c(n31304), .d(n30443), .o(n31780) );
na03f01 g27990 ( .a(n31780), .b(n31766), .c(n31298), .o(n31781) );
ao22f01 g27991 ( .a(n31636), .b(n31631), .c(n31305), .d(delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n31782) );
oa12f01 g27992 ( .a(n31299), .b(n31782), .c(n31765), .o(n31783) );
no02f01 g27993 ( .a(n30348), .b(n30347), .o(n31784) );
in01f01 g27994 ( .a(n30349), .o(n31785) );
ao12f01 g27995 ( .a(n30249), .b(n31785), .c(n31784), .o(n31786) );
in01f01 g27996 ( .a(n31786), .o(n31787) );
no02f01 g27997 ( .a(n30261), .b(n30259), .o(n31788) );
in01f01 g27998 ( .a(n31788), .o(n31789) );
no02f01 g27999 ( .a(n31789), .b(n31787), .o(n31790) );
no02f01 g28000 ( .a(n31788), .b(n31786), .o(n31791) );
no02f01 g28001 ( .a(n31791), .b(n31790), .o(n31792) );
in01f01 g28002 ( .a(n31792), .o(n31793) );
ao12f01 g28003 ( .a(n31793), .b(n31783), .c(n31781), .o(n31794) );
in01f01 g28004 ( .a(n31794), .o(n31795) );
na02f01 g28005 ( .a(n31778), .b(n31629), .o(n31796) );
no02f01 g28006 ( .a(n31796), .b(n31625), .o(n31797) );
no02f01 g28007 ( .a(n31797), .b(n30969), .o(n31798) );
no02f01 g28008 ( .a(n31796), .b(n31243), .o(n31799) );
ao12f01 g28009 ( .a(n31798), .b(n31799), .c(n31775), .o(n31800) );
in01f01 g28010 ( .a(n30328), .o(n31801) );
ao12f01 g28011 ( .a(n30335), .b(n30345), .c(n31801), .o(n31802) );
in01f01 g28012 ( .a(n30348), .o(n31803) );
na02f01 g28013 ( .a(n31803), .b(n30344), .o(n31804) );
no02f01 g28014 ( .a(n31804), .b(n31802), .o(n31805) );
na02f01 g28015 ( .a(n31804), .b(n31802), .o(n31806) );
in01f01 g28016 ( .a(n31806), .o(n31807) );
no02f01 g28017 ( .a(n31807), .b(n31805), .o(n31808) );
in01f01 g28018 ( .a(n31808), .o(n31809) );
no02f01 g28019 ( .a(n30928), .b(delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n31810) );
in01f01 g28020 ( .a(n31810), .o(n31811) );
na02f01 g28021 ( .a(n30899), .b(delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n31812) );
na02f01 g28022 ( .a(n31233), .b(n30443), .o(n31813) );
na02f01 g28023 ( .a(n31813), .b(n31812), .o(n31814) );
ao12f01 g28024 ( .a(n31814), .b(n31611), .c(n30443), .o(n31815) );
ao12f01 g28025 ( .a(delay_sub_ln23_0_unr15_stage6_stallmux_q), .b(n31815), .c(n30911), .o(n31816) );
oa22f01 g28026 ( .a(n31816), .b(n31616), .c(n30928), .d(n30443), .o(n31817) );
ao12f01 g28027 ( .a(n30940), .b(n31817), .c(n31811), .o(n31818) );
ao22f01 g28028 ( .a(n31772), .b(n31767), .c(n31245), .d(delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n31819) );
no03f01 g28029 ( .a(n31819), .b(n31810), .c(n31247), .o(n31820) );
in01f01 g28030 ( .a(n30322), .o(n31821) );
no02f01 g28031 ( .a(n30326), .b(n30270), .o(n31822) );
in01f01 g28032 ( .a(n31822), .o(n31823) );
no03f01 g28033 ( .a(n31823), .b(n30324), .c(n31821), .o(n31824) );
in01f01 g28034 ( .a(n30324), .o(n31825) );
ao12f01 g28035 ( .a(n31822), .b(n31825), .c(n30322), .o(n31826) );
no02f01 g28036 ( .a(n31826), .b(n31824), .o(n31827) );
no03f01 g28037 ( .a(n31827), .b(n31820), .c(n31818), .o(n31828) );
oa12f01 g28038 ( .a(n31827), .b(n31820), .c(n31818), .o(n31829) );
na03f01 g28039 ( .a(n31772), .b(n31767), .c(n30928), .o(n31830) );
oa12f01 g28040 ( .a(n31245), .b(n31816), .c(n31616), .o(n31831) );
in01f01 g28041 ( .a(n30312), .o(n31832) );
no02f01 g28042 ( .a(n31832), .b(n30277), .o(n31833) );
no02f01 g28043 ( .a(n30324), .b(n30320), .o(n31834) );
in01f01 g28044 ( .a(n31834), .o(n31835) );
no02f01 g28045 ( .a(n31835), .b(n31833), .o(n31836) );
na02f01 g28046 ( .a(n31835), .b(n31833), .o(n31837) );
in01f01 g28047 ( .a(n31837), .o(n31838) );
no02f01 g28048 ( .a(n31838), .b(n31836), .o(n31839) );
in01f01 g28049 ( .a(n31839), .o(n31840) );
ao12f01 g28050 ( .a(n31840), .b(n31831), .c(n31830), .o(n31841) );
in01f01 g28051 ( .a(n31612), .o(n31842) );
no02f01 g28052 ( .a(n31842), .b(n31237), .o(n31843) );
no02f01 g28053 ( .a(n31612), .b(n30911), .o(n31844) );
no02f01 g28054 ( .a(n31844), .b(n31843), .o(n31845) );
in01f01 g28055 ( .a(n30298), .o(n31846) );
in01f01 g28056 ( .a(n30305), .o(n31847) );
no03f01 g28057 ( .a(n31847), .b(n30299), .c(n31846), .o(n31848) );
in01f01 g28058 ( .a(n30299), .o(n31849) );
ao12f01 g28059 ( .a(n30305), .b(n31849), .c(n30298), .o(n31850) );
no02f01 g28060 ( .a(n31850), .b(n31848), .o(n31851) );
in01f01 g28061 ( .a(n31851), .o(n31852) );
in01f01 g28062 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_0_), .o(n31853) );
no02f01 g28063 ( .a(n30304), .b(n31853), .o(n31854) );
no02f01 g28064 ( .a(n30303), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_0_), .o(n31855) );
no02f01 g28065 ( .a(n31855), .b(n31854), .o(n31856) );
in01f01 g28066 ( .a(n31856), .o(n31857) );
na02f01 g28067 ( .a(n31857), .b(n30884), .o(n31858) );
na02f01 g28068 ( .a(n31858), .b(n31852), .o(n31859) );
no02f01 g28069 ( .a(n31858), .b(n31852), .o(n31860) );
na02f01 g28070 ( .a(n31610), .b(n31226), .o(n31861) );
na02f01 g28071 ( .a(n31769), .b(n30873), .o(n31862) );
na02f01 g28072 ( .a(n31862), .b(n31861), .o(n31863) );
oa12f01 g28073 ( .a(n31859), .b(n31863), .c(n31860), .o(n31864) );
no03f01 g28074 ( .a(n31610), .b(n31609), .c(n30899), .o(n31865) );
ao12f01 g28075 ( .a(n31233), .b(n31769), .c(n31768), .o(n31866) );
in01f01 g28076 ( .a(n30289), .o(n31867) );
no03f01 g28077 ( .a(n30307), .b(n30306), .c(n31867), .o(n31868) );
in01f01 g28078 ( .a(n30306), .o(n31869) );
in01f01 g28079 ( .a(n30307), .o(n31870) );
ao12f01 g28080 ( .a(n31869), .b(n31870), .c(n30289), .o(n31871) );
no02f01 g28081 ( .a(n31871), .b(n31868), .o(n31872) );
oa12f01 g28082 ( .a(n31872), .b(n31866), .c(n31865), .o(n31873) );
no03f01 g28083 ( .a(n31872), .b(n31866), .c(n31865), .o(n31874) );
ao12f01 g28084 ( .a(n31874), .b(n31873), .c(n31864), .o(n31875) );
in01f01 g28085 ( .a(n30308), .o(n31876) );
no02f01 g28086 ( .a(n30310), .b(n30277), .o(n31877) );
in01f01 g28087 ( .a(n31877), .o(n31878) );
no02f01 g28088 ( .a(n31878), .b(n31876), .o(n31879) );
no02f01 g28089 ( .a(n31877), .b(n30308), .o(n31880) );
no02f01 g28090 ( .a(n31880), .b(n31879), .o(n31881) );
na02f01 g28091 ( .a(n31881), .b(n31875), .o(n31882) );
no02f01 g28092 ( .a(n31881), .b(n31875), .o(n31883) );
ao12f01 g28093 ( .a(n31883), .b(n31882), .c(n31845), .o(n31884) );
na03f01 g28094 ( .a(n31840), .b(n31831), .c(n31830), .o(n31885) );
oa12f01 g28095 ( .a(n31885), .b(n31884), .c(n31841), .o(n31886) );
ao12f01 g28096 ( .a(n31828), .b(n31886), .c(n31829), .o(n31887) );
no02f01 g28097 ( .a(n31622), .b(n31621), .o(n31888) );
oa12f01 g28098 ( .a(n30956), .b(n31635), .c(n31888), .o(n31889) );
na02f01 g28099 ( .a(n31774), .b(n31773), .o(n31890) );
na03f01 g28100 ( .a(n31778), .b(n31890), .c(n30957), .o(n31891) );
in01f01 g28101 ( .a(n30345), .o(n31892) );
no02f01 g28102 ( .a(n31892), .b(n30335), .o(n31893) );
no02f01 g28103 ( .a(n31893), .b(n31801), .o(n31894) );
na02f01 g28104 ( .a(n31893), .b(n31801), .o(n31895) );
in01f01 g28105 ( .a(n31895), .o(n31896) );
no02f01 g28106 ( .a(n31896), .b(n31894), .o(n31897) );
in01f01 g28107 ( .a(n31897), .o(n31898) );
ao12f01 g28108 ( .a(n31898), .b(n31891), .c(n31889), .o(n31899) );
ao12f01 g28109 ( .a(n30957), .b(n31778), .c(n31890), .o(n31900) );
no03f01 g28110 ( .a(n31635), .b(n31888), .c(n30956), .o(n31901) );
no03f01 g28111 ( .a(n31897), .b(n31901), .c(n31900), .o(n31902) );
no02f01 g28112 ( .a(n31902), .b(n31809), .o(n31903) );
oa12f01 g28113 ( .a(n31903), .b(n31899), .c(n31887), .o(n31904) );
na03f01 g28114 ( .a(n31898), .b(n31891), .c(n31889), .o(n31905) );
oa12f01 g28115 ( .a(n31905), .b(n31899), .c(n31887), .o(n31906) );
ao22f01 g28116 ( .a(n31906), .b(n31809), .c(n31904), .d(n31800), .o(n31907) );
no02f01 g28117 ( .a(n31637), .b(n31305), .o(n31908) );
no02f01 g28118 ( .a(n31779), .b(n31777), .o(n31909) );
no02f01 g28119 ( .a(n31909), .b(n31304), .o(n31910) );
no02f01 g28120 ( .a(n31910), .b(n31908), .o(n31911) );
in01f01 g28121 ( .a(n31784), .o(n31912) );
no02f01 g28122 ( .a(n30349), .b(n30249), .o(n31913) );
no02f01 g28123 ( .a(n31913), .b(n31912), .o(n31914) );
na02f01 g28124 ( .a(n31913), .b(n31912), .o(n31915) );
in01f01 g28125 ( .a(n31915), .o(n31916) );
no02f01 g28126 ( .a(n31916), .b(n31914), .o(n31917) );
in01f01 g28127 ( .a(n31917), .o(n31918) );
no02f01 g28128 ( .a(n31918), .b(n31911), .o(n31919) );
no03f01 g28129 ( .a(n31917), .b(n31910), .c(n31908), .o(n31920) );
no03f01 g28130 ( .a(n31782), .b(n31765), .c(n31299), .o(n31921) );
ao12f01 g28131 ( .a(n31298), .b(n31780), .c(n31766), .o(n31922) );
no03f01 g28132 ( .a(n31792), .b(n31922), .c(n31921), .o(n31923) );
no02f01 g28133 ( .a(n31923), .b(n31920), .o(n31924) );
oa12f01 g28134 ( .a(n31924), .b(n31919), .c(n31907), .o(n31925) );
in01f01 g28135 ( .a(n31762), .o(n31926) );
ao12f01 g28136 ( .a(n31926), .b(n31755), .c(n31753), .o(n31927) );
in01f01 g28137 ( .a(n31927), .o(n31928) );
na03f01 g28138 ( .a(n31928), .b(n31925), .c(n31795), .o(n31929) );
na02f01 g28139 ( .a(n31747), .b(n31739), .o(n31930) );
na03f01 g28140 ( .a(n31930), .b(n31929), .c(n31764), .o(n31931) );
in01f01 g28141 ( .a(n31706), .o(n31932) );
in01f01 g28142 ( .a(n31713), .o(n31933) );
ao12f01 g28143 ( .a(n31933), .b(n31932), .c(n31704), .o(n31934) );
in01f01 g28144 ( .a(n31722), .o(n31935) );
ao12f01 g28145 ( .a(n31935), .b(n31726), .c(n31724), .o(n31936) );
no02f01 g28146 ( .a(n31936), .b(n31934), .o(n31937) );
na03f01 g28147 ( .a(n31937), .b(n31931), .c(n31749), .o(n31938) );
na02f01 g28148 ( .a(n31938), .b(n31730), .o(n31939) );
no02f01 g28149 ( .a(n31680), .b(n31352), .o(n31940) );
in01f01 g28150 ( .a(n31649), .o(n31941) );
na02f01 g28151 ( .a(n31941), .b(n31643), .o(n31942) );
ao12f01 g28152 ( .a(n31351), .b(n31679), .c(n31942), .o(n31943) );
no02f01 g28153 ( .a(n31943), .b(n31940), .o(n31944) );
no02f01 g28154 ( .a(n30385), .b(n30371), .o(n31945) );
no02f01 g28155 ( .a(n31945), .b(n31689), .o(n31946) );
na02f01 g28156 ( .a(n31945), .b(n31689), .o(n31947) );
in01f01 g28157 ( .a(n31947), .o(n31948) );
no02f01 g28158 ( .a(n31948), .b(n31946), .o(n31949) );
in01f01 g28159 ( .a(n31949), .o(n31950) );
no02f01 g28160 ( .a(n31950), .b(n31944), .o(n31951) );
in01f01 g28161 ( .a(n31951), .o(n31952) );
no03f01 g28162 ( .a(n31696), .b(n31685), .c(n31682), .o(n31953) );
na02f01 g28163 ( .a(n31950), .b(n31944), .o(n31954) );
in01f01 g28164 ( .a(n31954), .o(n31955) );
no02f01 g28165 ( .a(n31955), .b(n31953), .o(n31956) );
in01f01 g28166 ( .a(n31956), .o(n31957) );
ao12f01 g28167 ( .a(n31957), .b(n31952), .c(n31939), .o(n31958) );
no02f01 g28168 ( .a(n31958), .b(n31698), .o(n31959) );
na02f01 g28169 ( .a(n31664), .b(n31059), .o(n31960) );
na02f01 g28170 ( .a(n31664), .b(n30477), .o(n31961) );
oa12f01 g28171 ( .a(n31664), .b(n31114), .c(n31130), .o(n31962) );
na03f01 g28172 ( .a(n31962), .b(n31961), .c(n31960), .o(n31963) );
in01f01 g28173 ( .a(n31963), .o(n31964) );
ao12f01 g28174 ( .a(n31673), .b(n31964), .c(n31959), .o(n31965) );
no02f01 g28175 ( .a(n31666), .b(n30507), .o(n31966) );
ao12f01 g28176 ( .a(n31666), .b(n30497), .c(n30486), .o(n31967) );
no02f01 g28177 ( .a(n31967), .b(n31966), .o(n31968) );
in01f01 g28178 ( .a(n31968), .o(n31969) );
no02f01 g28179 ( .a(n31969), .b(n31965), .o(n31970) );
no02f01 g28180 ( .a(n31664), .b(n30506), .o(n31971) );
no02f01 g28181 ( .a(n31971), .b(n31034), .o(n31972) );
in01f01 g28182 ( .a(n31972), .o(n31973) );
oa12f01 g28183 ( .a(n31666), .b(n31973), .c(n31970), .o(n31974) );
ao12f01 g28184 ( .a(n31664), .b(n31072), .c(n31070), .o(n31975) );
ao12f01 g28185 ( .a(n31975), .b(n31970), .c(n31034), .o(n31976) );
na02f01 g28186 ( .a(n31976), .b(n31974), .o(n31977) );
no02f01 g28187 ( .a(n31977), .b(n31669), .o(n31978) );
in01f01 g28188 ( .a(n31698), .o(n31979) );
in01f01 g28189 ( .a(n31730), .o(n31980) );
in01f01 g28190 ( .a(n31800), .o(n31981) );
oa12f01 g28191 ( .a(n31247), .b(n31819), .c(n31810), .o(n31982) );
na03f01 g28192 ( .a(n31817), .b(n31811), .c(n30940), .o(n31983) );
in01f01 g28193 ( .a(n31827), .o(n31984) );
na03f01 g28194 ( .a(n31984), .b(n31983), .c(n31982), .o(n31985) );
ao12f01 g28195 ( .a(n31984), .b(n31983), .c(n31982), .o(n31986) );
no03f01 g28196 ( .a(n31816), .b(n31616), .c(n31245), .o(n31987) );
ao12f01 g28197 ( .a(n30928), .b(n31772), .c(n31767), .o(n31988) );
oa12f01 g28198 ( .a(n31839), .b(n31988), .c(n31987), .o(n31989) );
in01f01 g28199 ( .a(n31845), .o(n31990) );
no02f01 g28200 ( .a(n31769), .b(n30873), .o(n31991) );
no02f01 g28201 ( .a(n31610), .b(n31226), .o(n31992) );
no03f01 g28202 ( .a(n31992), .b(n31991), .c(n31860), .o(n31993) );
ao12f01 g28203 ( .a(n31993), .b(n31858), .c(n31852), .o(n31994) );
na03f01 g28204 ( .a(n31769), .b(n31768), .c(n31233), .o(n31995) );
oa12f01 g28205 ( .a(n30899), .b(n31610), .c(n31609), .o(n31996) );
in01f01 g28206 ( .a(n31872), .o(n31997) );
ao12f01 g28207 ( .a(n31997), .b(n31996), .c(n31995), .o(n31998) );
no02f01 g28208 ( .a(n31998), .b(n31994), .o(n31999) );
in01f01 g28209 ( .a(n31881), .o(n32000) );
no03f01 g28210 ( .a(n32000), .b(n31874), .c(n31999), .o(n32001) );
oa12f01 g28211 ( .a(n32000), .b(n31874), .c(n31999), .o(n32002) );
oa12f01 g28212 ( .a(n32002), .b(n32001), .c(n31990), .o(n32003) );
no03f01 g28213 ( .a(n31839), .b(n31988), .c(n31987), .o(n32004) );
ao12f01 g28214 ( .a(n32004), .b(n32003), .c(n31989), .o(n32005) );
oa12f01 g28215 ( .a(n31985), .b(n32005), .c(n31986), .o(n32006) );
in01f01 g28216 ( .a(n31899), .o(n32007) );
na02f01 g28217 ( .a(n31905), .b(n31808), .o(n32008) );
ao12f01 g28218 ( .a(n32008), .b(n32007), .c(n32006), .o(n32009) );
ao12f01 g28219 ( .a(n31902), .b(n32007), .c(n32006), .o(n32010) );
oa22f01 g28220 ( .a(n32010), .b(n31808), .c(n32009), .d(n31981), .o(n32011) );
in01f01 g28221 ( .a(n31919), .o(n32012) );
in01f01 g28222 ( .a(n31920), .o(n32013) );
na03f01 g28223 ( .a(n31793), .b(n31783), .c(n31781), .o(n32014) );
na02f01 g28224 ( .a(n32014), .b(n32013), .o(n32015) );
ao12f01 g28225 ( .a(n32015), .b(n32012), .c(n32011), .o(n32016) );
no03f01 g28226 ( .a(n31927), .b(n32016), .c(n31794), .o(n32017) );
in01f01 g28227 ( .a(n31930), .o(n32018) );
no03f01 g28228 ( .a(n32018), .b(n32017), .c(n31763), .o(n32019) );
in01f01 g28229 ( .a(n31936), .o(n32020) );
na02f01 g28230 ( .a(n32020), .b(n31729), .o(n32021) );
no03f01 g28231 ( .a(n32021), .b(n32019), .c(n31748), .o(n32022) );
no02f01 g28232 ( .a(n32022), .b(n31980), .o(n32023) );
oa12f01 g28233 ( .a(n31956), .b(n31951), .c(n32023), .o(n32024) );
na02f01 g28234 ( .a(n32024), .b(n31979), .o(n32025) );
oa12f01 g28235 ( .a(n31672), .b(n31963), .c(n32025), .o(n32026) );
na02f01 g28236 ( .a(n31968), .b(n32026), .o(n32027) );
ao12f01 g28237 ( .a(n31664), .b(n31972), .c(n32027), .o(n32028) );
in01f01 g28238 ( .a(n31975), .o(n32029) );
oa12f01 g28239 ( .a(n32029), .b(n32027), .c(n30516), .o(n32030) );
no02f01 g28240 ( .a(n32030), .b(n32028), .o(n32031) );
no02f01 g28241 ( .a(n32031), .b(n31668), .o(n32032) );
no02f01 g28242 ( .a(n32032), .b(n31978), .o(n32033) );
no02f01 g28243 ( .a(n32033), .b(n31607), .o(n32034) );
na02f01 g28244 ( .a(n32031), .b(n31668), .o(n32035) );
na02f01 g28245 ( .a(n31977), .b(n31669), .o(n32036) );
na02f01 g28246 ( .a(n32036), .b(n32035), .o(n32037) );
no02f01 g28247 ( .a(n32037), .b(n31606), .o(n32038) );
no02f01 g28248 ( .a(n32038), .b(n32034), .o(n32039) );
in01f01 g28249 ( .a(n31962), .o(n32040) );
no03f01 g28250 ( .a(n32040), .b(n31958), .c(n31698), .o(n32041) );
no02f01 g28251 ( .a(n31664), .b(n31059), .o(n32042) );
in01f01 g28252 ( .a(n31960), .o(n32043) );
no02f01 g28253 ( .a(n32043), .b(n32042), .o(n32044) );
in01f01 g28254 ( .a(n32044), .o(n32045) );
no03f01 g28255 ( .a(n32045), .b(n32041), .c(n31670), .o(n32046) );
in01f01 g28256 ( .a(n31670), .o(n32047) );
na03f01 g28257 ( .a(n31962), .b(n32024), .c(n31979), .o(n32048) );
ao12f01 g28258 ( .a(n32044), .b(n32048), .c(n32047), .o(n32049) );
no02f01 g28259 ( .a(n32049), .b(n32046), .o(n32050) );
na04f01 g28260 ( .a(n31962), .b(n31960), .c(n32024), .d(n31979), .o(n32051) );
no02f01 g28261 ( .a(n32042), .b(n31670), .o(n32052) );
in01f01 g28262 ( .a(n31961), .o(n32053) );
no02f01 g28263 ( .a(n31664), .b(n30477), .o(n32054) );
no02f01 g28264 ( .a(n32054), .b(n32053), .o(n32055) );
na03f01 g28265 ( .a(n32055), .b(n32052), .c(n32051), .o(n32056) );
no04f01 g28266 ( .a(n32040), .b(n32043), .c(n31958), .d(n31698), .o(n32057) );
in01f01 g28267 ( .a(n32052), .o(n32058) );
in01f01 g28268 ( .a(n32055), .o(n32059) );
oa12f01 g28269 ( .a(n32059), .b(n32058), .c(n32057), .o(n32060) );
na02f01 g28270 ( .a(n32060), .b(n32056), .o(n32061) );
in01f01 g28271 ( .a(n32061), .o(n32062) );
ao12f01 g28272 ( .a(n31607), .b(n32062), .c(n32050), .o(n32063) );
no02f01 g28273 ( .a(n31664), .b(n31114), .o(n32064) );
in01f01 g28274 ( .a(n32064), .o(n32065) );
in01f01 g28275 ( .a(n31130), .o(n32066) );
no02f01 g28276 ( .a(n31666), .b(n32066), .o(n32067) );
no02f01 g28277 ( .a(n31664), .b(n31130), .o(n32068) );
no02f01 g28278 ( .a(n32068), .b(n32067), .o(n32069) );
in01f01 g28279 ( .a(n31114), .o(n32070) );
no02f01 g28280 ( .a(n31666), .b(n32070), .o(n32071) );
in01f01 g28281 ( .a(n32071), .o(n32072) );
na03f01 g28282 ( .a(n32072), .b(n32024), .c(n31979), .o(n32073) );
na03f01 g28283 ( .a(n32073), .b(n32069), .c(n32065), .o(n32074) );
in01f01 g28284 ( .a(n32069), .o(n32075) );
no03f01 g28285 ( .a(n32071), .b(n31958), .c(n31698), .o(n32076) );
oa12f01 g28286 ( .a(n32075), .b(n32076), .c(n32064), .o(n32077) );
na02f01 g28287 ( .a(n32077), .b(n32074), .o(n32078) );
no02f01 g28288 ( .a(n32071), .b(n32064), .o(n32079) );
in01f01 g28289 ( .a(n32079), .o(n32080) );
no02f01 g28290 ( .a(n32080), .b(n31959), .o(n32081) );
no02f01 g28291 ( .a(n32079), .b(n32025), .o(n32082) );
no02f01 g28292 ( .a(n32082), .b(n32081), .o(n32083) );
in01f01 g28293 ( .a(n32083), .o(n32084) );
no02f01 g28294 ( .a(n32084), .b(n32078), .o(n32085) );
no02f01 g28295 ( .a(n32085), .b(n31607), .o(n32086) );
no02f01 g28296 ( .a(n32086), .b(n32063), .o(n32087) );
no02f01 g28297 ( .a(n31664), .b(n31070), .o(n32088) );
no02f01 g28298 ( .a(n31666), .b(n30486), .o(n32089) );
no02f01 g28299 ( .a(n32089), .b(n32088), .o(n32090) );
na02f01 g28300 ( .a(n32090), .b(n31965), .o(n32091) );
in01f01 g28301 ( .a(n32090), .o(n32092) );
na02f01 g28302 ( .a(n32092), .b(n32026), .o(n32093) );
na02f01 g28303 ( .a(n32093), .b(n32091), .o(n32094) );
no02f01 g28304 ( .a(n31666), .b(n30497), .o(n32095) );
no02f01 g28305 ( .a(n31664), .b(n31072), .o(n32096) );
no02f01 g28306 ( .a(n32096), .b(n32095), .o(n32097) );
in01f01 g28307 ( .a(n32089), .o(n32098) );
ao12f01 g28308 ( .a(n32088), .b(n32098), .c(n32026), .o(n32099) );
na02f01 g28309 ( .a(n32099), .b(n32097), .o(n32100) );
in01f01 g28310 ( .a(n32097), .o(n32101) );
in01f01 g28311 ( .a(n32088), .o(n32102) );
oa12f01 g28312 ( .a(n32102), .b(n32089), .c(n31965), .o(n32103) );
na02f01 g28313 ( .a(n32103), .b(n32101), .o(n32104) );
na02f01 g28314 ( .a(n32104), .b(n32100), .o(n32105) );
oa12f01 g28315 ( .a(n31606), .b(n32105), .c(n32094), .o(n32106) );
na02f01 g28316 ( .a(n32106), .b(n32087), .o(n32107) );
no02f01 g28317 ( .a(n31967), .b(n31963), .o(n32108) );
na02f01 g28318 ( .a(n32108), .b(n31959), .o(n32109) );
no02f01 g28319 ( .a(n31975), .b(n31673), .o(n32110) );
na02f01 g28320 ( .a(n32110), .b(n32109), .o(n32111) );
no02f01 g28321 ( .a(n31971), .b(n31966), .o(n32112) );
in01f01 g28322 ( .a(n32112), .o(n32113) );
no02f01 g28323 ( .a(n32113), .b(n32111), .o(n32114) );
na02f01 g28324 ( .a(n32113), .b(n32111), .o(n32115) );
in01f01 g28325 ( .a(n32115), .o(n32116) );
no02f01 g28326 ( .a(n32116), .b(n32114), .o(n32117) );
no02f01 g28327 ( .a(n31664), .b(n30516), .o(n32118) );
no02f01 g28328 ( .a(n31666), .b(n31034), .o(n32119) );
no02f01 g28329 ( .a(n32119), .b(n32118), .o(n32120) );
in01f01 g28330 ( .a(n32120), .o(n32121) );
ao12f01 g28331 ( .a(n31673), .b(n32108), .c(n31959), .o(n32122) );
no02f01 g28332 ( .a(n31975), .b(n31971), .o(n32123) );
oa12f01 g28333 ( .a(n32123), .b(n32122), .c(n31966), .o(n32124) );
no02f01 g28334 ( .a(n32124), .b(n32121), .o(n32125) );
na02f01 g28335 ( .a(n32124), .b(n32121), .o(n32126) );
in01f01 g28336 ( .a(n32126), .o(n32127) );
no02f01 g28337 ( .a(n32127), .b(n32125), .o(n32128) );
ao12f01 g28338 ( .a(n31607), .b(n32128), .c(n32117), .o(n32129) );
no02f01 g28339 ( .a(n32129), .b(n32107), .o(n32130) );
ao12f01 g28340 ( .a(n31951), .b(n31954), .c(n32023), .o(n32131) );
no02f01 g28341 ( .a(n31953), .b(n31698), .o(n32132) );
in01f01 g28342 ( .a(n32132), .o(n32133) );
no02f01 g28343 ( .a(n32133), .b(n32131), .o(n32134) );
na02f01 g28344 ( .a(n32133), .b(n32131), .o(n32135) );
in01f01 g28345 ( .a(n32135), .o(n32136) );
no02f01 g28346 ( .a(n32136), .b(n32134), .o(n32137) );
in01f01 g28347 ( .a(n32137), .o(n32138) );
no02f01 g28348 ( .a(n32138), .b(n31606), .o(n32139) );
no02f01 g28349 ( .a(n31596), .b(n6075), .o(n32140) );
no02f01 g28350 ( .a(n31596), .b(n_22641), .o(n32141) );
no02f01 g28351 ( .a(n32141), .b(n32140), .o(n32142) );
in01f01 g28352 ( .a(n32142), .o(n32143) );
no02f01 g28353 ( .a(n31586), .b(n6075), .o(n32144) );
no03f01 g28354 ( .a(n32144), .b(n31570), .c(n31560), .o(n32145) );
no02f01 g28355 ( .a(n31586), .b(n_22641), .o(n32146) );
no02f01 g28356 ( .a(n32146), .b(n31575), .o(n32147) );
in01f01 g28357 ( .a(n32147), .o(n32148) );
no03f01 g28358 ( .a(n32148), .b(n32145), .c(n32143), .o(n32149) );
in01f01 g28359 ( .a(n32149), .o(n32150) );
oa12f01 g28360 ( .a(n32143), .b(n32148), .c(n32145), .o(n32151) );
na02f01 g28361 ( .a(n32151), .b(n32150), .o(n32152) );
no02f01 g28362 ( .a(n32019), .b(n31748), .o(n32153) );
no02f01 g28363 ( .a(n32153), .b(n31728), .o(n32154) );
no02f01 g28364 ( .a(n32154), .b(n31936), .o(n32155) );
in01f01 g28365 ( .a(n32155), .o(n32156) );
no02f01 g28366 ( .a(n31934), .b(n31714), .o(n32157) );
no02f01 g28367 ( .a(n32157), .b(n32156), .o(n32158) );
na02f01 g28368 ( .a(n32157), .b(n32156), .o(n32159) );
in01f01 g28369 ( .a(n32159), .o(n32160) );
no02f01 g28370 ( .a(n32160), .b(n32158), .o(n32161) );
na02f01 g28371 ( .a(n32161), .b(n32152), .o(n32162) );
no02f01 g28372 ( .a(n32161), .b(n32152), .o(n32163) );
no02f01 g28373 ( .a(n32146), .b(n32144), .o(n32164) );
no02f01 g28374 ( .a(n32164), .b(n31576), .o(n32165) );
na02f01 g28375 ( .a(n32164), .b(n31576), .o(n32166) );
in01f01 g28376 ( .a(n32166), .o(n32167) );
no02f01 g28377 ( .a(n31936), .b(n31728), .o(n32168) );
in01f01 g28378 ( .a(n32168), .o(n32169) );
no02f01 g28379 ( .a(n32169), .b(n32153), .o(n32170) );
no03f01 g28380 ( .a(n32168), .b(n32019), .c(n31748), .o(n32171) );
no02f01 g28381 ( .a(n32171), .b(n32170), .o(n32172) );
no03f01 g28382 ( .a(n32172), .b(n32167), .c(n32165), .o(n32173) );
oa12f01 g28383 ( .a(n32162), .b(n32173), .c(n32163), .o(n32174) );
no02f01 g28384 ( .a(n31557), .b(n_22641), .o(n32175) );
no02f01 g28385 ( .a(n32175), .b(n31572), .o(n32176) );
na02f01 g28386 ( .a(n32176), .b(n31560), .o(n32177) );
no02f01 g28387 ( .a(n31569), .b(n_22641), .o(n32178) );
no02f01 g28388 ( .a(n32178), .b(n31570), .o(n32179) );
in01f01 g28389 ( .a(n32179), .o(n32180) );
na02f01 g28390 ( .a(n32180), .b(n32177), .o(n32181) );
in01f01 g28391 ( .a(n32181), .o(n32182) );
no02f01 g28392 ( .a(n32180), .b(n32177), .o(n32183) );
no02f01 g28393 ( .a(n32183), .b(n32182), .o(n32184) );
no02f01 g28394 ( .a(n32017), .b(n31763), .o(n32185) );
no02f01 g28395 ( .a(n32018), .b(n31748), .o(n32186) );
no02f01 g28396 ( .a(n32186), .b(n32185), .o(n32187) );
na02f01 g28397 ( .a(n32186), .b(n32185), .o(n32188) );
in01f01 g28398 ( .a(n32188), .o(n32189) );
no02f01 g28399 ( .a(n32189), .b(n32187), .o(n32190) );
in01f01 g28400 ( .a(n32190), .o(n32191) );
no02f01 g28401 ( .a(n32191), .b(n32184), .o(n32192) );
in01f01 g28402 ( .a(n32192), .o(n32193) );
na02f01 g28403 ( .a(n31547), .b(n31534), .o(n32194) );
in01f01 g28404 ( .a(n31572), .o(n32195) );
no02f01 g28405 ( .a(n32175), .b(n31558), .o(n32196) );
ao12f01 g28406 ( .a(n32196), .b(n32195), .c(n32194), .o(n32197) );
na03f01 g28407 ( .a(n32196), .b(n32195), .c(n32194), .o(n32198) );
in01f01 g28408 ( .a(n32198), .o(n32199) );
no02f01 g28409 ( .a(n32016), .b(n31794), .o(n32200) );
in01f01 g28410 ( .a(n32200), .o(n32201) );
no02f01 g28411 ( .a(n31927), .b(n31763), .o(n32202) );
no02f01 g28412 ( .a(n32202), .b(n32201), .o(n32203) );
na02f01 g28413 ( .a(n32202), .b(n32201), .o(n32204) );
in01f01 g28414 ( .a(n32204), .o(n32205) );
no02f01 g28415 ( .a(n32205), .b(n32203), .o(n32206) );
no03f01 g28416 ( .a(n32206), .b(n32199), .c(n32197), .o(n32207) );
in01f01 g28417 ( .a(n32207), .o(n32208) );
no02f01 g28418 ( .a(n31532), .b(n_22641), .o(n32209) );
no02f01 g28419 ( .a(n31545), .b(n_22641), .o(n32210) );
no02f01 g28420 ( .a(n32210), .b(n31546), .o(n32211) );
in01f01 g28421 ( .a(n32211), .o(n32212) );
oa12f01 g28422 ( .a(n32212), .b(n32209), .c(n31534), .o(n32213) );
no03f01 g28423 ( .a(n32212), .b(n32209), .c(n31534), .o(n32214) );
in01f01 g28424 ( .a(n32214), .o(n32215) );
ao12f01 g28425 ( .a(n31920), .b(n32012), .c(n32011), .o(n32216) );
no02f01 g28426 ( .a(n31923), .b(n31794), .o(n32217) );
no02f01 g28427 ( .a(n32217), .b(n32216), .o(n32218) );
na02f01 g28428 ( .a(n32217), .b(n32216), .o(n32219) );
in01f01 g28429 ( .a(n32219), .o(n32220) );
no02f01 g28430 ( .a(n32220), .b(n32218), .o(n32221) );
in01f01 g28431 ( .a(n32221), .o(n32222) );
ao12f01 g28432 ( .a(n32222), .b(n32215), .c(n32213), .o(n32223) );
in01f01 g28433 ( .a(n32223), .o(n32224) );
no02f01 g28434 ( .a(n32209), .b(n31533), .o(n32225) );
na02f01 g28435 ( .a(n32225), .b(n31522), .o(n32226) );
in01f01 g28436 ( .a(n32226), .o(n32227) );
no02f01 g28437 ( .a(n32225), .b(n31522), .o(n32228) );
no02f01 g28438 ( .a(n31920), .b(n31919), .o(n32229) );
no02f01 g28439 ( .a(n32229), .b(n31907), .o(n32230) );
na02f01 g28440 ( .a(n32229), .b(n31907), .o(n32231) );
in01f01 g28441 ( .a(n32231), .o(n32232) );
no02f01 g28442 ( .a(n32232), .b(n32230), .o(n32233) );
no03f01 g28443 ( .a(n32233), .b(n32228), .c(n32227), .o(n32234) );
in01f01 g28444 ( .a(n32234), .o(n32235) );
ao12f01 g28445 ( .a(n_22641), .b(n31495), .c(n31493), .o(n32236) );
oa12f01 g28446 ( .a(n_22641), .b(n31400), .c(n31398), .o(n32237) );
no03f01 g28447 ( .a(n31461), .b(n31460), .c(n30886), .o(n32238) );
ao12f01 g28448 ( .a(n31406), .b(n31404), .c(n31403), .o(n32239) );
no02f01 g28449 ( .a(n32239), .b(n32238), .o(n32240) );
no03f01 g28450 ( .a(n31472), .b(n31467), .c(n31465), .o(n32241) );
ao12f01 g28451 ( .a(n31466), .b(n31469), .c(n31468), .o(n32242) );
no02f01 g28452 ( .a(n32242), .b(n32241), .o(n32243) );
ao12f01 g28453 ( .a(n6075), .b(n32243), .c(n32240), .o(n32244) );
in01f01 g28454 ( .a(n31479), .o(n32245) );
ao12f01 g28455 ( .a(n6075), .b(n31480), .c(n32245), .o(n32246) );
no02f01 g28456 ( .a(n32246), .b(n32244), .o(n32247) );
na02f01 g28457 ( .a(n32247), .b(n32237), .o(n32248) );
in01f01 g28458 ( .a(n31398), .o(n32249) );
oa12f01 g28459 ( .a(n31397), .b(n31239), .c(n30914), .o(n32250) );
na02f01 g28460 ( .a(n32250), .b(n32249), .o(n32251) );
in01f01 g28461 ( .a(n31485), .o(n32252) );
oa12f01 g28462 ( .a(n6075), .b(n32252), .c(n32251), .o(n32253) );
ao12f01 g28463 ( .a(n31496), .b(n32253), .c(n32248), .o(n32254) );
no02f01 g28464 ( .a(n31502), .b(n_22641), .o(n32255) );
no02f01 g28465 ( .a(n32255), .b(n31503), .o(n32256) );
in01f01 g28466 ( .a(n32256), .o(n32257) );
oa12f01 g28467 ( .a(n32257), .b(n32254), .c(n32236), .o(n32258) );
oa12f01 g28468 ( .a(n6075), .b(n31494), .c(n31514), .o(n32259) );
na02f01 g28469 ( .a(n32253), .b(n32248), .o(n32260) );
oa12f01 g28470 ( .a(n_22641), .b(n31494), .c(n31514), .o(n32261) );
na02f01 g28471 ( .a(n32261), .b(n32260), .o(n32262) );
na03f01 g28472 ( .a(n32256), .b(n32262), .c(n32259), .o(n32263) );
no02f01 g28473 ( .a(n31986), .b(n31828), .o(n32264) );
no02f01 g28474 ( .a(n32264), .b(n32005), .o(n32265) );
na02f01 g28475 ( .a(n32264), .b(n32005), .o(n32266) );
in01f01 g28476 ( .a(n32266), .o(n32267) );
no02f01 g28477 ( .a(n32267), .b(n32265), .o(n32268) );
in01f01 g28478 ( .a(n32268), .o(n32269) );
ao12f01 g28479 ( .a(n32269), .b(n32263), .c(n32258), .o(n32270) );
in01f01 g28480 ( .a(n32270), .o(n32271) );
ao22f01 g28481 ( .a(n32259), .b(n32261), .c(n32253), .d(n32248), .o(n32272) );
no04f01 g28482 ( .a(n32236), .b(n31496), .c(n31486), .d(n31484), .o(n32273) );
no02f01 g28483 ( .a(n32004), .b(n31841), .o(n32274) );
no02f01 g28484 ( .a(n32274), .b(n31884), .o(n32275) );
na02f01 g28485 ( .a(n32274), .b(n31884), .o(n32276) );
in01f01 g28486 ( .a(n32276), .o(n32277) );
no02f01 g28487 ( .a(n32277), .b(n32275), .o(n32278) );
no03f01 g28488 ( .a(n32278), .b(n32273), .c(n32272), .o(n32279) );
in01f01 g28489 ( .a(n32279), .o(n32280) );
oa12f01 g28490 ( .a(n6075), .b(n31481), .c(n31479), .o(n32281) );
oa12f01 g28491 ( .a(n6075), .b(n31400), .c(n31398), .o(n32282) );
ao22f01 g28492 ( .a(n32282), .b(n32237), .c(n32281), .d(n31483), .o(n32283) );
ao12f01 g28493 ( .a(n_22641), .b(n31480), .c(n32245), .o(n32284) );
no02f01 g28494 ( .a(n31401), .b(n_22641), .o(n32285) );
no04f01 g28495 ( .a(n32285), .b(n32284), .c(n32247), .d(n31402), .o(n32286) );
no02f01 g28496 ( .a(n32000), .b(n31845), .o(n32287) );
no02f01 g28497 ( .a(n31881), .b(n31990), .o(n32288) );
no02f01 g28498 ( .a(n32288), .b(n32287), .o(n32289) );
no02f01 g28499 ( .a(n32289), .b(n31875), .o(n32290) );
na02f01 g28500 ( .a(n32289), .b(n31875), .o(n32291) );
in01f01 g28501 ( .a(n32291), .o(n32292) );
no02f01 g28502 ( .a(n32292), .b(n32290), .o(n32293) );
oa12f01 g28503 ( .a(n32293), .b(n32286), .c(n32283), .o(n32294) );
oa12f01 g28504 ( .a(n31475), .b(n32284), .c(n32246), .o(n32295) );
na03f01 g28505 ( .a(n32281), .b(n31482), .c(n32244), .o(n32296) );
no02f01 g28506 ( .a(n31874), .b(n31998), .o(n32297) );
no02f01 g28507 ( .a(n32297), .b(n31994), .o(n32298) );
na02f01 g28508 ( .a(n32297), .b(n31994), .o(n32299) );
in01f01 g28509 ( .a(n32299), .o(n32300) );
no02f01 g28510 ( .a(n32300), .b(n32298), .o(n32301) );
in01f01 g28511 ( .a(n32301), .o(n32302) );
na03f01 g28512 ( .a(n32302), .b(n32296), .c(n32295), .o(n32303) );
no03f01 g28513 ( .a(n32243), .b(n31463), .c(n6075), .o(n32304) );
ao12f01 g28514 ( .a(n32240), .b(n31474), .c(n_22641), .o(n32305) );
in01f01 g28515 ( .a(n31858), .o(n32306) );
ao12f01 g28516 ( .a(n31852), .b(n31862), .c(n31861), .o(n32307) );
no02f01 g28517 ( .a(n31863), .b(n31851), .o(n32308) );
no02f01 g28518 ( .a(n32308), .b(n32307), .o(n32309) );
no02f01 g28519 ( .a(n32309), .b(n32306), .o(n32310) );
na02f01 g28520 ( .a(n32309), .b(n32306), .o(n32311) );
in01f01 g28521 ( .a(n32311), .o(n32312) );
no02f01 g28522 ( .a(n32312), .b(n32310), .o(n32313) );
oa12f01 g28523 ( .a(n32313), .b(n32305), .c(n32304), .o(n32314) );
na02f01 g28524 ( .a(n32243), .b(n6075), .o(n32315) );
na02f01 g28525 ( .a(n32243), .b(n_22641), .o(n32316) );
no02f01 g28526 ( .a(n31856), .b(n30884), .o(n32317) );
no02f01 g28527 ( .a(n31857), .b(n31222), .o(n32318) );
no02f01 g28528 ( .a(n32318), .b(n32317), .o(n32319) );
in01f01 g28529 ( .a(n32319), .o(n32320) );
na03f01 g28530 ( .a(n32320), .b(n32316), .c(n32315), .o(n32321) );
no03f01 g28531 ( .a(n32313), .b(n32305), .c(n32304), .o(n32322) );
ao12f01 g28532 ( .a(n32322), .b(n32321), .c(n32314), .o(n32323) );
ao12f01 g28533 ( .a(n32302), .b(n32296), .c(n32295), .o(n32324) );
oa12f01 g28534 ( .a(n32303), .b(n32324), .c(n32323), .o(n32325) );
no03f01 g28535 ( .a(n32293), .b(n32286), .c(n32283), .o(n32326) );
oa12f01 g28536 ( .a(n32294), .b(n32326), .c(n32325), .o(n32327) );
in01f01 g28537 ( .a(n32272), .o(n32328) );
na04f01 g28538 ( .a(n32259), .b(n32261), .c(n32253), .d(n32248), .o(n32329) );
in01f01 g28539 ( .a(n32278), .o(n32330) );
ao12f01 g28540 ( .a(n32330), .b(n32329), .c(n32328), .o(n32331) );
oa12f01 g28541 ( .a(n32280), .b(n32331), .c(n32327), .o(n32332) );
ao12f01 g28542 ( .a(n32256), .b(n32262), .c(n32259), .o(n32333) );
no03f01 g28543 ( .a(n32257), .b(n32254), .c(n32236), .o(n32334) );
no03f01 g28544 ( .a(n32268), .b(n32334), .c(n32333), .o(n32335) );
oa12f01 g28545 ( .a(n32271), .b(n32335), .c(n32332), .o(n32336) );
na02f01 g28546 ( .a(n31518), .b(n_22641), .o(n32337) );
na02f01 g28547 ( .a(n31518), .b(n6075), .o(n32338) );
na02f01 g28548 ( .a(n32338), .b(n32337), .o(n32339) );
no02f01 g28549 ( .a(n32262), .b(n31503), .o(n32340) );
no03f01 g28550 ( .a(n32340), .b(n32339), .c(n31516), .o(n32341) );
ao12f01 g28551 ( .a(n31392), .b(n31389), .c(n31241), .o(n32342) );
in01f01 g28552 ( .a(n31393), .o(n32343) );
no02f01 g28553 ( .a(n32343), .b(n32342), .o(n32344) );
no02f01 g28554 ( .a(n32344), .b(n_22641), .o(n32345) );
no02f01 g28555 ( .a(n32345), .b(n31394), .o(n32346) );
in01f01 g28556 ( .a(n31503), .o(n32347) );
na02f01 g28557 ( .a(n32254), .b(n32347), .o(n32348) );
ao12f01 g28558 ( .a(n32346), .b(n32348), .c(n31517), .o(n32349) );
no02f01 g28559 ( .a(n31902), .b(n31899), .o(n32350) );
no02f01 g28560 ( .a(n32350), .b(n31887), .o(n32351) );
na02f01 g28561 ( .a(n32350), .b(n31887), .o(n32352) );
in01f01 g28562 ( .a(n32352), .o(n32353) );
no02f01 g28563 ( .a(n32353), .b(n32351), .o(n32354) );
oa12f01 g28564 ( .a(n32354), .b(n32349), .c(n32341), .o(n32355) );
in01f01 g28565 ( .a(n32355), .o(n32356) );
no02f01 g28566 ( .a(n31511), .b(n_22641), .o(n32357) );
no02f01 g28567 ( .a(n32357), .b(n31512), .o(n32358) );
in01f01 g28568 ( .a(n32358), .o(n32359) );
na02f01 g28569 ( .a(n32338), .b(n31517), .o(n32360) );
no03f01 g28570 ( .a(n32360), .b(n32359), .c(n31504), .o(n32361) );
no02f01 g28571 ( .a(n31503), .b(n31496), .o(n32362) );
na03f01 g28572 ( .a(n32362), .b(n32260), .c(n32337), .o(n32363) );
no02f01 g28573 ( .a(n32345), .b(n31516), .o(n32364) );
ao12f01 g28574 ( .a(n32358), .b(n32364), .c(n32363), .o(n32365) );
ao12f01 g28575 ( .a(n31899), .b(n31905), .c(n31887), .o(n32366) );
in01f01 g28576 ( .a(n32366), .o(n32367) );
no02f01 g28577 ( .a(n31808), .b(n31981), .o(n32368) );
no02f01 g28578 ( .a(n31809), .b(n31800), .o(n32369) );
no02f01 g28579 ( .a(n32369), .b(n32368), .o(n32370) );
no02f01 g28580 ( .a(n32370), .b(n32367), .o(n32371) );
na02f01 g28581 ( .a(n32370), .b(n32367), .o(n32372) );
in01f01 g28582 ( .a(n32372), .o(n32373) );
no02f01 g28583 ( .a(n32373), .b(n32371), .o(n32374) );
no03f01 g28584 ( .a(n32374), .b(n32365), .c(n32361), .o(n32375) );
no03f01 g28585 ( .a(n32354), .b(n32349), .c(n32341), .o(n32376) );
no02f01 g28586 ( .a(n32376), .b(n32375), .o(n32377) );
oa12f01 g28587 ( .a(n32377), .b(n32356), .c(n32336), .o(n32378) );
na03f01 g28588 ( .a(n32364), .b(n32358), .c(n32363), .o(n32379) );
oa12f01 g28589 ( .a(n32359), .b(n32360), .c(n31504), .o(n32380) );
in01f01 g28590 ( .a(n32374), .o(n32381) );
ao12f01 g28591 ( .a(n32381), .b(n32380), .c(n32379), .o(n32382) );
in01f01 g28592 ( .a(n32382), .o(n32383) );
oa12f01 g28593 ( .a(n32233), .b(n32228), .c(n32227), .o(n32384) );
na03f01 g28594 ( .a(n32384), .b(n32383), .c(n32378), .o(n32385) );
na03f01 g28595 ( .a(n32222), .b(n32215), .c(n32213), .o(n32386) );
na03f01 g28596 ( .a(n32386), .b(n32385), .c(n32235), .o(n32387) );
oa12f01 g28597 ( .a(n32206), .b(n32199), .c(n32197), .o(n32388) );
na03f01 g28598 ( .a(n32388), .b(n32387), .c(n32224), .o(n32389) );
no03f01 g28599 ( .a(n32190), .b(n32183), .c(n32182), .o(n32390) );
in01f01 g28600 ( .a(n32390), .o(n32391) );
na03f01 g28601 ( .a(n32391), .b(n32389), .c(n32208), .o(n32392) );
in01f01 g28602 ( .a(n32151), .o(n32393) );
no02f01 g28603 ( .a(n32393), .b(n32149), .o(n32394) );
in01f01 g28604 ( .a(n32161), .o(n32395) );
no02f01 g28605 ( .a(n32395), .b(n32394), .o(n32396) );
in01f01 g28606 ( .a(n32165), .o(n32397) );
in01f01 g28607 ( .a(n32172), .o(n32398) );
ao12f01 g28608 ( .a(n32398), .b(n32166), .c(n32397), .o(n32399) );
no02f01 g28609 ( .a(n32399), .b(n32396), .o(n32400) );
na03f01 g28610 ( .a(n32400), .b(n32392), .c(n32193), .o(n32401) );
na02f01 g28611 ( .a(n32401), .b(n32174), .o(n32402) );
no02f01 g28612 ( .a(n31602), .b(n31601), .o(n32403) );
no02f01 g28613 ( .a(n31599), .b(n31598), .o(n32404) );
no02f01 g28614 ( .a(n32404), .b(n32403), .o(n32405) );
in01f01 g28615 ( .a(n32405), .o(n32406) );
na02f01 g28616 ( .a(n32404), .b(n32403), .o(n32407) );
no02f01 g28617 ( .a(n31955), .b(n31951), .o(n32408) );
in01f01 g28618 ( .a(n32408), .o(n32409) );
no02f01 g28619 ( .a(n32409), .b(n31939), .o(n32410) );
no02f01 g28620 ( .a(n32408), .b(n32023), .o(n32411) );
no02f01 g28621 ( .a(n32411), .b(n32410), .o(n32412) );
in01f01 g28622 ( .a(n32412), .o(n32413) );
ao12f01 g28623 ( .a(n32413), .b(n32407), .c(n32406), .o(n32414) );
in01f01 g28624 ( .a(n32414), .o(n32415) );
na03f01 g28625 ( .a(n32413), .b(n32407), .c(n32406), .o(n32416) );
oa12f01 g28626 ( .a(n32416), .b(n32137), .c(n31607), .o(n32417) );
ao12f01 g28627 ( .a(n32417), .b(n32415), .c(n32402), .o(n32418) );
ao12f01 g28628 ( .a(n31606), .b(n32084), .c(n32078), .o(n32419) );
no02f01 g28629 ( .a(n32061), .b(n31606), .o(n32420) );
na03f01 g28630 ( .a(n32044), .b(n32048), .c(n32047), .o(n32421) );
oa12f01 g28631 ( .a(n32045), .b(n32041), .c(n31670), .o(n32422) );
na02f01 g28632 ( .a(n32422), .b(n32421), .o(n32423) );
no02f01 g28633 ( .a(n32423), .b(n31606), .o(n32424) );
no02f01 g28634 ( .a(n32424), .b(n32420), .o(n32425) );
in01f01 g28635 ( .a(n32425), .o(n32426) );
no04f01 g28636 ( .a(n32426), .b(n32419), .c(n32418), .d(n32139), .o(n32427) );
no02f01 g28637 ( .a(n32094), .b(n31606), .o(n32428) );
no02f01 g28638 ( .a(n32105), .b(n31606), .o(n32429) );
no02f01 g28639 ( .a(n32429), .b(n32428), .o(n32430) );
in01f01 g28640 ( .a(n32114), .o(n32431) );
na02f01 g28641 ( .a(n32115), .b(n32431), .o(n32432) );
no02f01 g28642 ( .a(n32432), .b(n31606), .o(n32433) );
in01f01 g28643 ( .a(n32128), .o(n32434) );
no02f01 g28644 ( .a(n32434), .b(n31606), .o(n32435) );
no02f01 g28645 ( .a(n32435), .b(n32433), .o(n32436) );
na03f01 g28646 ( .a(n32436), .b(n32430), .c(n32427), .o(n32437) );
na03f01 g28647 ( .a(n32437), .b(n32130), .c(n32039), .o(n32438) );
in01f01 g28648 ( .a(n32039), .o(n32439) );
in01f01 g28649 ( .a(n32130), .o(n32440) );
in01f01 g28650 ( .a(n32139), .o(n32441) );
in01f01 g28651 ( .a(n32174), .o(n32442) );
oa22f01 g28652 ( .a(n32285), .b(n31402), .c(n32284), .d(n32247), .o(n32443) );
na04f01 g28653 ( .a(n32282), .b(n32281), .c(n31483), .d(n32237), .o(n32444) );
in01f01 g28654 ( .a(n32293), .o(n32445) );
ao12f01 g28655 ( .a(n32445), .b(n32444), .c(n32443), .o(n32446) );
ao12f01 g28656 ( .a(n32244), .b(n32281), .c(n31482), .o(n32447) );
no03f01 g28657 ( .a(n32284), .b(n32246), .c(n31475), .o(n32448) );
no03f01 g28658 ( .a(n32301), .b(n32448), .c(n32447), .o(n32449) );
na03f01 g28659 ( .a(n31474), .b(n32240), .c(n_22641), .o(n32450) );
oa12f01 g28660 ( .a(n31463), .b(n32243), .c(n6075), .o(n32451) );
in01f01 g28661 ( .a(n32313), .o(n32452) );
ao12f01 g28662 ( .a(n32452), .b(n32451), .c(n32450), .o(n32453) );
no02f01 g28663 ( .a(n31474), .b(n_22641), .o(n32454) );
no02f01 g28664 ( .a(n31474), .b(n6075), .o(n32455) );
no03f01 g28665 ( .a(n32319), .b(n32455), .c(n32454), .o(n32456) );
na03f01 g28666 ( .a(n32452), .b(n32451), .c(n32450), .o(n32457) );
oa12f01 g28667 ( .a(n32457), .b(n32456), .c(n32453), .o(n32458) );
oa12f01 g28668 ( .a(n32301), .b(n32448), .c(n32447), .o(n32459) );
ao12f01 g28669 ( .a(n32449), .b(n32459), .c(n32458), .o(n32460) );
na03f01 g28670 ( .a(n32445), .b(n32444), .c(n32443), .o(n32461) );
ao12f01 g28671 ( .a(n32446), .b(n32461), .c(n32460), .o(n32462) );
oa12f01 g28672 ( .a(n32278), .b(n32273), .c(n32272), .o(n32463) );
ao12f01 g28673 ( .a(n32279), .b(n32463), .c(n32462), .o(n32464) );
na03f01 g28674 ( .a(n32269), .b(n32263), .c(n32258), .o(n32465) );
ao12f01 g28675 ( .a(n32270), .b(n32465), .c(n32464), .o(n32466) );
na03f01 g28676 ( .a(n32381), .b(n32380), .c(n32379), .o(n32467) );
na03f01 g28677 ( .a(n32348), .b(n32346), .c(n31517), .o(n32468) );
oa12f01 g28678 ( .a(n32339), .b(n32340), .c(n31516), .o(n32469) );
in01f01 g28679 ( .a(n32354), .o(n32470) );
na03f01 g28680 ( .a(n32470), .b(n32469), .c(n32468), .o(n32471) );
na02f01 g28681 ( .a(n32471), .b(n32467), .o(n32472) );
ao12f01 g28682 ( .a(n32472), .b(n32355), .c(n32466), .o(n32473) );
in01f01 g28683 ( .a(n32228), .o(n32474) );
in01f01 g28684 ( .a(n32233), .o(n32475) );
ao12f01 g28685 ( .a(n32475), .b(n32474), .c(n32226), .o(n32476) );
no03f01 g28686 ( .a(n32476), .b(n32382), .c(n32473), .o(n32477) );
in01f01 g28687 ( .a(n32213), .o(n32478) );
no03f01 g28688 ( .a(n32221), .b(n32214), .c(n32478), .o(n32479) );
no03f01 g28689 ( .a(n32479), .b(n32477), .c(n32234), .o(n32480) );
in01f01 g28690 ( .a(n32197), .o(n32481) );
in01f01 g28691 ( .a(n32206), .o(n32482) );
ao12f01 g28692 ( .a(n32482), .b(n32198), .c(n32481), .o(n32483) );
no03f01 g28693 ( .a(n32483), .b(n32480), .c(n32223), .o(n32484) );
no03f01 g28694 ( .a(n32390), .b(n32484), .c(n32207), .o(n32485) );
oa12f01 g28695 ( .a(n32172), .b(n32167), .c(n32165), .o(n32486) );
na02f01 g28696 ( .a(n32486), .b(n32162), .o(n32487) );
no03f01 g28697 ( .a(n32487), .b(n32485), .c(n32192), .o(n32488) );
no02f01 g28698 ( .a(n32488), .b(n32442), .o(n32489) );
in01f01 g28699 ( .a(n32417), .o(n32490) );
oa12f01 g28700 ( .a(n32490), .b(n32414), .c(n32489), .o(n32491) );
in01f01 g28701 ( .a(n32419), .o(n32492) );
na04f01 g28702 ( .a(n32425), .b(n32492), .c(n32491), .d(n32441), .o(n32493) );
in01f01 g28703 ( .a(n32430), .o(n32494) );
in01f01 g28704 ( .a(n32436), .o(n32495) );
no03f01 g28705 ( .a(n32495), .b(n32494), .c(n32493), .o(n32496) );
oa12f01 g28706 ( .a(n32439), .b(n32496), .c(n32440), .o(n32497) );
na02f01 g28707 ( .a(n32497), .b(n32438), .o(n403) );
no02f01 g28708 ( .a(n8693), .b(n8661), .o(n32499) );
in01f01 g28709 ( .a(n32499), .o(n32500) );
in01f01 g28710 ( .a(n8675), .o(n32501) );
no02f01 g28711 ( .a(n8753), .b(n32501), .o(n32502) );
no02f01 g28712 ( .a(n8756), .b(n8713), .o(n32503) );
na03f01 g28713 ( .a(n32503), .b(n32502), .c(n32500), .o(n32504) );
in01f01 g28714 ( .a(n32502), .o(n32505) );
in01f01 g28715 ( .a(n32503), .o(n32506) );
oa12f01 g28716 ( .a(n32506), .b(n32505), .c(n32499), .o(n32507) );
na02f01 g28717 ( .a(n32507), .b(n32504), .o(n408) );
na02f01 g28718 ( .a(n26754), .b(n7712), .o(n32509) );
na02f01 g28719 ( .a(n26754), .b(n7682), .o(n32510) );
oa12f01 g28720 ( .a(n7682), .b(n26835), .c(n26833), .o(n32511) );
oa12f01 g28721 ( .a(n7682), .b(n26827), .c(n26824), .o(n32512) );
oa12f01 g28722 ( .a(n27071), .b(n26818), .c(n26817), .o(n32513) );
na03f01 g28723 ( .a(n27069), .b(n26703), .c(n26701), .o(n32514) );
ao12f01 g28724 ( .a(n7712), .b(n32514), .c(n32513), .o(n32515) );
oa12f01 g28725 ( .a(n27101), .b(n26814), .c(n26758), .o(n32516) );
na03f01 g28726 ( .a(n27099), .b(n26692), .c(n26521), .o(n32517) );
ao12f01 g28727 ( .a(n7712), .b(n32517), .c(n32516), .o(n32518) );
oa12f01 g28728 ( .a(n7682), .b(n27059), .c(n26859), .o(n32519) );
oa12f01 g28729 ( .a(n7682), .b(n27094), .c(n27092), .o(n32520) );
na02f01 g28730 ( .a(n32520), .b(n32519), .o(n32521) );
no02f01 g28731 ( .a(n32521), .b(n32518), .o(n32522) );
oa12f01 g28732 ( .a(n7682), .b(n27077), .c(n27075), .o(n32523) );
na02f01 g28733 ( .a(n32523), .b(n32522), .o(n32524) );
no02f01 g28734 ( .a(n32524), .b(n32515), .o(n32525) );
oa12f01 g28735 ( .a(n7712), .b(n26827), .c(n26824), .o(n32526) );
ao12f01 g28736 ( .a(n7682), .b(n32514), .c(n32513), .o(n32527) );
na03f01 g28737 ( .a(n27076), .b(n26696), .c(n26516), .o(n32528) );
oa12f01 g28738 ( .a(n27074), .b(n26815), .c(n26515), .o(n32529) );
ao12f01 g28739 ( .a(n7682), .b(n32529), .c(n32528), .o(n32530) );
no02f01 g28740 ( .a(n32530), .b(n32527), .o(n32531) );
na02f01 g28741 ( .a(n32531), .b(n32526), .o(n32532) );
ao12f01 g28742 ( .a(n32532), .b(n32525), .c(n32512), .o(n32533) );
oa12f01 g28743 ( .a(n7712), .b(n26835), .c(n26833), .o(n32534) );
na02f01 g28744 ( .a(n32534), .b(n32533), .o(n32535) );
ao12f01 g28745 ( .a(n7712), .b(n26843), .c(n26842), .o(n32536) );
in01f01 g28746 ( .a(n32536), .o(n32537) );
na03f01 g28747 ( .a(n32537), .b(n32535), .c(n32511), .o(n32538) );
ao12f01 g28748 ( .a(n7682), .b(n26843), .c(n26842), .o(n32539) );
in01f01 g28749 ( .a(n32539), .o(n32540) );
na04f01 g28750 ( .a(n32540), .b(n32538), .c(n32510), .d(n32509), .o(n32541) );
na02f01 g28751 ( .a(n32510), .b(n32509), .o(n32542) );
in01f01 g28752 ( .a(n32511), .o(n32543) );
na03f01 g28753 ( .a(n26826), .b(n26707), .c(n26706), .o(n32544) );
oa12f01 g28754 ( .a(n26823), .b(n26820), .c(n26819), .o(n32545) );
ao12f01 g28755 ( .a(n7712), .b(n32545), .c(n32544), .o(n32546) );
oa12f01 g28756 ( .a(n7682), .b(n27072), .c(n27070), .o(n32547) );
in01f01 g28757 ( .a(n32524), .o(n32548) );
na02f01 g28758 ( .a(n32548), .b(n32547), .o(n32549) );
ao12f01 g28759 ( .a(n7682), .b(n32545), .c(n32544), .o(n32550) );
oa12f01 g28760 ( .a(n7712), .b(n27072), .c(n27070), .o(n32551) );
oa12f01 g28761 ( .a(n7712), .b(n27077), .c(n27075), .o(n32552) );
na02f01 g28762 ( .a(n32552), .b(n32551), .o(n32553) );
no02f01 g28763 ( .a(n32553), .b(n32550), .o(n32554) );
oa12f01 g28764 ( .a(n32554), .b(n32549), .c(n32546), .o(n32555) );
in01f01 g28765 ( .a(n32534), .o(n32556) );
no02f01 g28766 ( .a(n32556), .b(n32555), .o(n32557) );
no03f01 g28767 ( .a(n32536), .b(n32557), .c(n32543), .o(n32558) );
oa12f01 g28768 ( .a(n32542), .b(n32539), .c(n32558), .o(n32559) );
no03f01 g28769 ( .a(n17769), .b(n17650), .c(n17540), .o(n32560) );
ao12f01 g28770 ( .a(n17768), .b(n17651), .c(n17740), .o(n32561) );
no02f01 g28771 ( .a(n32561), .b(n32560), .o(n32562) );
in01f01 g28772 ( .a(n32562), .o(n32563) );
na03f01 g28773 ( .a(n32563), .b(n32559), .c(n32541), .o(n32564) );
no03f01 g28774 ( .a(n32539), .b(n32558), .c(n32542), .o(n32565) );
ao22f01 g28775 ( .a(n32540), .b(n32538), .c(n32510), .d(n32509), .o(n32566) );
oa12f01 g28776 ( .a(n32562), .b(n32566), .c(n32565), .o(n32567) );
no02f01 g28777 ( .a(n32539), .b(n32536), .o(n32568) );
no03f01 g28778 ( .a(n32568), .b(n32557), .c(n32543), .o(n32569) );
in01f01 g28779 ( .a(n32568), .o(n32570) );
ao12f01 g28780 ( .a(n32570), .b(n32535), .c(n32511), .o(n32571) );
no02f01 g28781 ( .a(n17552), .b(n17743), .o(n32572) );
no02f01 g28782 ( .a(n32572), .b(n17649), .o(n32573) );
na02f01 g28783 ( .a(n32572), .b(n17649), .o(n32574) );
in01f01 g28784 ( .a(n32574), .o(n32575) );
no02f01 g28785 ( .a(n32575), .b(n32573), .o(n32576) );
no03f01 g28786 ( .a(n32576), .b(n32571), .c(n32569), .o(n32577) );
na03f01 g28787 ( .a(n32534), .b(n32533), .c(n32511), .o(n32578) );
oa12f01 g28788 ( .a(n32555), .b(n32556), .c(n32543), .o(n32579) );
no02f01 g28789 ( .a(n17562), .b(n17746), .o(n32580) );
no02f01 g28790 ( .a(n17563), .b(n17557), .o(n32581) );
no02f01 g28791 ( .a(n32581), .b(n32580), .o(n32582) );
in01f01 g28792 ( .a(n32582), .o(n32583) );
ao12f01 g28793 ( .a(n17642), .b(n17644), .c(n17628), .o(n32584) );
no02f01 g28794 ( .a(n32584), .b(n32583), .o(n32585) );
na02f01 g28795 ( .a(n32584), .b(n32583), .o(n32586) );
in01f01 g28796 ( .a(n32586), .o(n32587) );
no02f01 g28797 ( .a(n32587), .b(n32585), .o(n32588) );
in01f01 g28798 ( .a(n32588), .o(n32589) );
na03f01 g28799 ( .a(n32589), .b(n32579), .c(n32578), .o(n32590) );
ao22f01 g28800 ( .a(n32531), .b(n32549), .c(n32526), .d(n32512), .o(n32591) );
no04f01 g28801 ( .a(n32553), .b(n32550), .c(n32525), .d(n32546), .o(n32592) );
no02f01 g28802 ( .a(n17765), .b(n17642), .o(n32593) );
no02f01 g28803 ( .a(n32593), .b(n17628), .o(n32594) );
na02f01 g28804 ( .a(n32593), .b(n17628), .o(n32595) );
in01f01 g28805 ( .a(n32595), .o(n32596) );
no02f01 g28806 ( .a(n32596), .b(n32594), .o(n32597) );
no03f01 g28807 ( .a(n32597), .b(n32592), .c(n32591), .o(n32598) );
no02f01 g28808 ( .a(n17625), .b(n17750), .o(n32599) );
no02f01 g28809 ( .a(n32599), .b(n17624), .o(n32600) );
na02f01 g28810 ( .a(n32599), .b(n17624), .o(n32601) );
in01f01 g28811 ( .a(n32601), .o(n32602) );
no02f01 g28812 ( .a(n32602), .b(n32600), .o(n32603) );
in01f01 g28813 ( .a(n32522), .o(n32604) );
ao12f01 g28814 ( .a(n32604), .b(n32552), .c(n32523), .o(n32605) );
ao12f01 g28815 ( .a(n7712), .b(n32529), .c(n32528), .o(n32606) );
no03f01 g28816 ( .a(n32530), .b(n32606), .c(n32522), .o(n32607) );
no03f01 g28817 ( .a(n32607), .b(n32605), .c(n32603), .o(n32608) );
oa12f01 g28818 ( .a(n32603), .b(n32607), .c(n32605), .o(n32609) );
ao12f01 g28819 ( .a(n26857), .b(n26856), .c(n26809), .o(n32610) );
no03f01 g28820 ( .a(n26852), .b(n26851), .c(n26684), .o(n32611) );
no02f01 g28821 ( .a(n32611), .b(n32610), .o(n32612) );
ao12f01 g28822 ( .a(n7712), .b(n27063), .c(n32612), .o(n32613) );
oa12f01 g28823 ( .a(n27093), .b(n26813), .c(n26529), .o(n32614) );
na03f01 g28824 ( .a(n27091), .b(n26689), .c(n26530), .o(n32615) );
ao12f01 g28825 ( .a(n7712), .b(n32615), .c(n32614), .o(n32616) );
no02f01 g28826 ( .a(n32616), .b(n32613), .o(n32617) );
ao12f01 g28827 ( .a(n7682), .b(n32517), .c(n32516), .o(n32618) );
oa12f01 g28828 ( .a(n32617), .b(n32618), .c(n32518), .o(n32619) );
oa12f01 g28829 ( .a(n7682), .b(n27102), .c(n27100), .o(n32620) );
oa12f01 g28830 ( .a(n7712), .b(n27102), .c(n27100), .o(n32621) );
na03f01 g28831 ( .a(n32621), .b(n32521), .c(n32620), .o(n32622) );
no02f01 g28832 ( .a(n17623), .b(n17757), .o(n32623) );
no02f01 g28833 ( .a(n32623), .b(n17752), .o(n32624) );
na02f01 g28834 ( .a(n32623), .b(n17752), .o(n32625) );
in01f01 g28835 ( .a(n32625), .o(n32626) );
no02f01 g28836 ( .a(n32626), .b(n32624), .o(n32627) );
in01f01 g28837 ( .a(n32627), .o(n32628) );
na03f01 g28838 ( .a(n32628), .b(n32622), .c(n32619), .o(n32629) );
ao12f01 g28839 ( .a(n32628), .b(n32622), .c(n32619), .o(n32630) );
oa12f01 g28840 ( .a(n7712), .b(n27094), .c(n27092), .o(n32631) );
ao12f01 g28841 ( .a(n32613), .b(n32631), .c(n32520), .o(n32632) );
ao12f01 g28842 ( .a(n7682), .b(n32615), .c(n32614), .o(n32633) );
no03f01 g28843 ( .a(n32633), .b(n32616), .c(n32519), .o(n32634) );
no02f01 g28844 ( .a(n17597), .b(n17594), .o(n32635) );
no02f01 g28845 ( .a(n32635), .b(n17611), .o(n32636) );
na02f01 g28846 ( .a(n32635), .b(n17611), .o(n32637) );
in01f01 g28847 ( .a(n32637), .o(n32638) );
no02f01 g28848 ( .a(n32638), .b(n32636), .o(n32639) );
no03f01 g28849 ( .a(n32639), .b(n32634), .c(n32632), .o(n32640) );
oa12f01 g28850 ( .a(n32639), .b(n32634), .c(n32632), .o(n32641) );
in01f01 g28851 ( .a(n17605), .o(n32642) );
no02f01 g28852 ( .a(n17609), .b(n32642), .o(n32643) );
na02f01 g28853 ( .a(n17609), .b(n32642), .o(n32644) );
in01f01 g28854 ( .a(n32644), .o(n32645) );
no02f01 g28855 ( .a(n32645), .b(n32643), .o(n32646) );
no02f01 g28856 ( .a(n32646), .b(n17602), .o(n32647) );
na02f01 g28857 ( .a(n32646), .b(n17602), .o(n32648) );
in01f01 g28858 ( .a(n32648), .o(n32649) );
no02f01 g28859 ( .a(n32649), .b(n32647), .o(n32650) );
no02f01 g28860 ( .a(n17601), .b(n17268), .o(n32651) );
na02f01 g28861 ( .a(n17601), .b(n17268), .o(n32652) );
in01f01 g28862 ( .a(n32652), .o(n32653) );
no02f01 g28863 ( .a(n32653), .b(n32651), .o(n32654) );
no02f01 g28864 ( .a(n32654), .b(n27063), .o(n32655) );
no02f01 g28865 ( .a(n32655), .b(n32650), .o(n32656) );
in01f01 g28866 ( .a(n32656), .o(n32657) );
na02f01 g28867 ( .a(n32655), .b(n32650), .o(n32658) );
in01f01 g28868 ( .a(n32658), .o(n32659) );
oa12f01 g28869 ( .a(n26859), .b(n27063), .c(n7712), .o(n32660) );
na03f01 g28870 ( .a(n27059), .b(n32612), .c(n7682), .o(n32661) );
na02f01 g28871 ( .a(n32661), .b(n32660), .o(n32662) );
oa12f01 g28872 ( .a(n32657), .b(n32662), .c(n32659), .o(n32663) );
ao12f01 g28873 ( .a(n32640), .b(n32663), .c(n32641), .o(n32664) );
oa12f01 g28874 ( .a(n32629), .b(n32664), .c(n32630), .o(n32665) );
ao12f01 g28875 ( .a(n32608), .b(n32665), .c(n32609), .o(n32666) );
na02f01 g28876 ( .a(n32552), .b(n32524), .o(n32667) );
oa12f01 g28877 ( .a(n32667), .b(n32527), .c(n32515), .o(n32668) );
ao12f01 g28878 ( .a(n32530), .b(n32523), .c(n32522), .o(n32669) );
na03f01 g28879 ( .a(n32669), .b(n32551), .c(n32547), .o(n32670) );
no03f01 g28880 ( .a(n17762), .b(n17626), .c(n17575), .o(n32671) );
ao12f01 g28881 ( .a(n17761), .b(n17627), .c(n17574), .o(n32672) );
no02f01 g28882 ( .a(n32672), .b(n32671), .o(n32673) );
in01f01 g28883 ( .a(n32673), .o(n32674) );
na03f01 g28884 ( .a(n32674), .b(n32670), .c(n32668), .o(n32675) );
ao12f01 g28885 ( .a(n32674), .b(n32670), .c(n32668), .o(n32676) );
ao12f01 g28886 ( .a(n32676), .b(n32675), .c(n32666), .o(n32677) );
oa12f01 g28887 ( .a(n32597), .b(n32592), .c(n32591), .o(n32678) );
ao12f01 g28888 ( .a(n32598), .b(n32678), .c(n32677), .o(n32679) );
ao12f01 g28889 ( .a(n32589), .b(n32579), .c(n32578), .o(n32680) );
ao12f01 g28890 ( .a(n32680), .b(n32679), .c(n32590), .o(n32681) );
oa12f01 g28891 ( .a(n32576), .b(n32571), .c(n32569), .o(n32682) );
ao12f01 g28892 ( .a(n32577), .b(n32682), .c(n32681), .o(n32683) );
na03f01 g28893 ( .a(n32683), .b(n32567), .c(n32564), .o(n32684) );
in01f01 g28894 ( .a(n32564), .o(n32685) );
ao12f01 g28895 ( .a(n32563), .b(n32559), .c(n32541), .o(n32686) );
na03f01 g28896 ( .a(n32570), .b(n32535), .c(n32511), .o(n32687) );
oa12f01 g28897 ( .a(n32568), .b(n32557), .c(n32543), .o(n32688) );
in01f01 g28898 ( .a(n32576), .o(n32689) );
na03f01 g28899 ( .a(n32689), .b(n32688), .c(n32687), .o(n32690) );
no03f01 g28900 ( .a(n32556), .b(n32555), .c(n32543), .o(n32691) );
ao12f01 g28901 ( .a(n32533), .b(n32534), .c(n32511), .o(n32692) );
no03f01 g28902 ( .a(n32588), .b(n32692), .c(n32691), .o(n32693) );
in01f01 g28903 ( .a(n32598), .o(n32694) );
in01f01 g28904 ( .a(n32603), .o(n32695) );
oa12f01 g28905 ( .a(n32522), .b(n32530), .c(n32606), .o(n32696) );
na03f01 g28906 ( .a(n32552), .b(n32523), .c(n32604), .o(n32697) );
na03f01 g28907 ( .a(n32697), .b(n32696), .c(n32695), .o(n32698) );
ao12f01 g28908 ( .a(n32695), .b(n32697), .c(n32696), .o(n32699) );
ao12f01 g28909 ( .a(n32521), .b(n32621), .c(n32620), .o(n32700) );
no03f01 g28910 ( .a(n32618), .b(n32617), .c(n32518), .o(n32701) );
no03f01 g28911 ( .a(n32627), .b(n32701), .c(n32700), .o(n32702) );
oa12f01 g28912 ( .a(n32627), .b(n32701), .c(n32700), .o(n32703) );
oa12f01 g28913 ( .a(n32519), .b(n32633), .c(n32616), .o(n32704) );
na03f01 g28914 ( .a(n32631), .b(n32520), .c(n32613), .o(n32705) );
in01f01 g28915 ( .a(n32639), .o(n32706) );
na03f01 g28916 ( .a(n32706), .b(n32705), .c(n32704), .o(n32707) );
ao12f01 g28917 ( .a(n32706), .b(n32705), .c(n32704), .o(n32708) );
in01f01 g28918 ( .a(n32660), .o(n32709) );
no03f01 g28919 ( .a(n27063), .b(n26859), .c(n7712), .o(n32710) );
no02f01 g28920 ( .a(n32710), .b(n32709), .o(n32711) );
ao12f01 g28921 ( .a(n32656), .b(n32711), .c(n32658), .o(n32712) );
oa12f01 g28922 ( .a(n32707), .b(n32712), .c(n32708), .o(n32713) );
ao12f01 g28923 ( .a(n32702), .b(n32713), .c(n32703), .o(n32714) );
oa12f01 g28924 ( .a(n32698), .b(n32714), .c(n32699), .o(n32715) );
ao12f01 g28925 ( .a(n32669), .b(n32551), .c(n32547), .o(n32716) );
no03f01 g28926 ( .a(n32667), .b(n32527), .c(n32515), .o(n32717) );
no03f01 g28927 ( .a(n32673), .b(n32717), .c(n32716), .o(n32718) );
oa12f01 g28928 ( .a(n32673), .b(n32717), .c(n32716), .o(n32719) );
oa12f01 g28929 ( .a(n32719), .b(n32718), .c(n32715), .o(n32720) );
oa22f01 g28930 ( .a(n32553), .b(n32525), .c(n32550), .d(n32546), .o(n32721) );
na04f01 g28931 ( .a(n32531), .b(n32526), .c(n32549), .d(n32512), .o(n32722) );
in01f01 g28932 ( .a(n32597), .o(n32723) );
ao12f01 g28933 ( .a(n32723), .b(n32722), .c(n32721), .o(n32724) );
oa12f01 g28934 ( .a(n32694), .b(n32724), .c(n32720), .o(n32725) );
oa12f01 g28935 ( .a(n32588), .b(n32692), .c(n32691), .o(n32726) );
oa12f01 g28936 ( .a(n32726), .b(n32725), .c(n32693), .o(n32727) );
ao12f01 g28937 ( .a(n32689), .b(n32688), .c(n32687), .o(n32728) );
oa12f01 g28938 ( .a(n32690), .b(n32728), .c(n32727), .o(n32729) );
oa12f01 g28939 ( .a(n32729), .b(n32686), .c(n32685), .o(n32730) );
na02f01 g28940 ( .a(n32730), .b(n32684), .o(n413) );
na03f01 g28941 ( .a(state_cordic_1_), .b(mux_while_ln12_psv_q_8_), .c(rst), .o(n32732) );
na02f01 g28942 ( .a(n32732), .b(sin_out_5), .o(n32733) );
in01f01 g28943 ( .a(n32732), .o(n32734) );
in01f01 g28944 ( .a(delay_xor_ln21_unr28_stage10_stallmux_q_3_), .o(n32735) );
in01f01 g28945 ( .a(n_44610), .o(n32736) );
no02f01 g28946 ( .a(n32736), .b(delay_xor_ln21_unr28_stage10_stallmux_q_2_), .o(n32737) );
in01f01 g28947 ( .a(n32737), .o(n32738) );
no02f01 g28948 ( .a(n32736), .b(delay_xor_ln21_unr28_stage10_stallmux_q_1_), .o(n32739) );
no02f01 g28949 ( .a(n32736), .b(delay_xor_ln21_unr28_stage10_stallmux_q_0_), .o(n32740) );
no02f01 g28950 ( .a(n32740), .b(n32739), .o(n32741) );
na02f01 g28951 ( .a(n32741), .b(n32738), .o(n32742) );
in01f01 g28952 ( .a(n32742), .o(n32743) );
ao12f01 g28953 ( .a(n32735), .b(n32743), .c(n_44610), .o(n32744) );
in01f01 g28954 ( .a(n32744), .o(n32745) );
no02f01 g28955 ( .a(n32745), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_14_), .o(n32746) );
no02f01 g28956 ( .a(n_44610), .b(n32735), .o(n32747) );
no02f01 g28957 ( .a(n32736), .b(delay_xor_ln21_unr28_stage10_stallmux_q_3_), .o(n32748) );
no02f01 g28958 ( .a(n32748), .b(n32747), .o(n32749) );
in01f01 g28959 ( .a(n32749), .o(n32750) );
no02f01 g28960 ( .a(n32750), .b(n32743), .o(n32751) );
no02f01 g28961 ( .a(n32749), .b(n32742), .o(n32752) );
no02f01 g28962 ( .a(n32752), .b(n32751), .o(n32753) );
no02f01 g28963 ( .a(n32753), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_3_), .o(n32754) );
in01f01 g28964 ( .a(n32754), .o(n32755) );
na02f01 g28965 ( .a(n32736), .b(delay_xor_ln21_unr28_stage10_stallmux_q_2_), .o(n32756) );
na02f01 g28966 ( .a(n32756), .b(n32738), .o(n32757) );
no02f01 g28967 ( .a(n32757), .b(n32741), .o(n32758) );
in01f01 g28968 ( .a(n32741), .o(n32759) );
in01f01 g28969 ( .a(n32756), .o(n32760) );
no02f01 g28970 ( .a(n32760), .b(n32737), .o(n32761) );
no02f01 g28971 ( .a(n32761), .b(n32759), .o(n32762) );
no02f01 g28972 ( .a(n32762), .b(n32758), .o(n32763) );
na02f01 g28973 ( .a(n32763), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_2_), .o(n32764) );
in01f01 g28974 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_1_), .o(n32765) );
in01f01 g28975 ( .a(delay_xor_ln21_unr28_stage10_stallmux_q_1_), .o(n32766) );
na02f01 g28976 ( .a(n_44610), .b(n32766), .o(n32767) );
na02f01 g28977 ( .a(n32740), .b(n32767), .o(n32768) );
no02f01 g28978 ( .a(n_44610), .b(n32766), .o(n32769) );
no02f01 g28979 ( .a(n32769), .b(n32739), .o(n32770) );
oa12f01 g28980 ( .a(n32768), .b(n32770), .c(n32740), .o(n32771) );
no02f01 g28981 ( .a(n32771), .b(n32765), .o(n32772) );
na02f01 g28982 ( .a(n32771), .b(n32765), .o(n32773) );
no02f01 g28983 ( .a(n_44610), .b(delay_xor_ln21_unr28_stage10_stallmux_q_0_), .o(n32774) );
na02f01 g28984 ( .a(n_44610), .b(delay_xor_ln21_unr28_stage10_stallmux_q_0_), .o(n32775) );
in01f01 g28985 ( .a(n32775), .o(n32776) );
no02f01 g28986 ( .a(n32776), .b(n32774), .o(n32777) );
in01f01 g28987 ( .a(n32777), .o(n32778) );
no02f01 g28988 ( .a(n32778), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_0_), .o(n32779) );
in01f01 g28989 ( .a(n32779), .o(n32780) );
ao12f01 g28990 ( .a(n32772), .b(n32780), .c(n32773), .o(n32781) );
in01f01 g28991 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_2_), .o(n32782) );
oa12f01 g28992 ( .a(n32782), .b(n32762), .c(n32758), .o(n32783) );
in01f01 g28993 ( .a(n32783), .o(n32784) );
oa12f01 g28994 ( .a(n32764), .b(n32784), .c(n32781), .o(n32785) );
in01f01 g28995 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_3_), .o(n32786) );
no03f01 g28996 ( .a(n32752), .b(n32751), .c(n32786), .o(n32787) );
oa12f01 g28997 ( .a(n32755), .b(n32787), .c(n32785), .o(n32788) );
no02f01 g28998 ( .a(n32745), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_6_), .o(n32789) );
ao12f01 g28999 ( .a(n32745), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_5_), .c(delay_sub_ln21_0_unr27_stage10_stallmux_q_4_), .o(n32790) );
no02f01 g29000 ( .a(n32790), .b(n32789), .o(n32791) );
in01f01 g29001 ( .a(n32791), .o(n32792) );
no02f01 g29002 ( .a(n32792), .b(n32788), .o(n32793) );
no02f01 g29003 ( .a(n32745), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_7_), .o(n32794) );
in01f01 g29004 ( .a(n32794), .o(n32795) );
in01f01 g29005 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_6_), .o(n32796) );
no02f01 g29006 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_5_), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_4_), .o(n32797) );
ao12f01 g29007 ( .a(n32744), .b(n32797), .c(n32796), .o(n32798) );
in01f01 g29008 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_7_), .o(n32799) );
no02f01 g29009 ( .a(n32744), .b(n32799), .o(n32800) );
no02f01 g29010 ( .a(n32800), .b(n32798), .o(n32801) );
in01f01 g29011 ( .a(n32801), .o(n32802) );
ao12f01 g29012 ( .a(n32802), .b(n32795), .c(n32793), .o(n32803) );
ao12f01 g29013 ( .a(n32745), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_8_), .c(delay_sub_ln21_0_unr27_stage10_stallmux_q_9_), .o(n32804) );
no02f01 g29014 ( .a(n32745), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_10_), .o(n32805) );
no02f01 g29015 ( .a(n32745), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_11_), .o(n32806) );
no03f01 g29016 ( .a(n32806), .b(n32805), .c(n32804), .o(n32807) );
in01f01 g29017 ( .a(n32807), .o(n32808) );
no02f01 g29018 ( .a(n32745), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_12_), .o(n32809) );
no02f01 g29019 ( .a(n32745), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_13_), .o(n32810) );
no03f01 g29020 ( .a(n32810), .b(n32809), .c(n32808), .o(n32811) );
in01f01 g29021 ( .a(n32811), .o(n32812) );
no03f01 g29022 ( .a(n32812), .b(n32803), .c(n32746), .o(n32813) );
no02f01 g29023 ( .a(n32745), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_15_), .o(n32814) );
in01f01 g29024 ( .a(n32814), .o(n32815) );
in01f01 g29025 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_12_), .o(n32816) );
in01f01 g29026 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_13_), .o(n32817) );
ao12f01 g29027 ( .a(n32744), .b(n32817), .c(n32816), .o(n32818) );
in01f01 g29028 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_11_), .o(n32819) );
in01f01 g29029 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_10_), .o(n32820) );
ao12f01 g29030 ( .a(n32744), .b(n32820), .c(n32819), .o(n32821) );
in01f01 g29031 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_9_), .o(n32822) );
in01f01 g29032 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_8_), .o(n32823) );
ao12f01 g29033 ( .a(n32744), .b(n32823), .c(n32822), .o(n32824) );
no02f01 g29034 ( .a(n32824), .b(n32821), .o(n32825) );
in01f01 g29035 ( .a(n32825), .o(n32826) );
no02f01 g29036 ( .a(n32826), .b(n32818), .o(n32827) );
in01f01 g29037 ( .a(n32827), .o(n32828) );
in01f01 g29038 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_15_), .o(n32829) );
in01f01 g29039 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_14_), .o(n32830) );
ao12f01 g29040 ( .a(n32744), .b(n32830), .c(n32829), .o(n32831) );
no02f01 g29041 ( .a(n32831), .b(n32828), .o(n32832) );
in01f01 g29042 ( .a(n32832), .o(n32833) );
ao12f01 g29043 ( .a(n32833), .b(n32815), .c(n32813), .o(n32834) );
no02f01 g29044 ( .a(n32745), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_18_), .o(n32835) );
ao12f01 g29045 ( .a(n32745), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_17_), .c(delay_sub_ln21_0_unr27_stage10_stallmux_q_16_), .o(n32836) );
no02f01 g29046 ( .a(n32745), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_19_), .o(n32837) );
no03f01 g29047 ( .a(n32837), .b(n32836), .c(n32835), .o(n32838) );
in01f01 g29048 ( .a(n32838), .o(n32839) );
no02f01 g29049 ( .a(n32745), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_21_), .o(n32840) );
no02f01 g29050 ( .a(n32745), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_20_), .o(n32841) );
no02f01 g29051 ( .a(n32841), .b(n32840), .o(n32842) );
in01f01 g29052 ( .a(n32842), .o(n32843) );
no02f01 g29053 ( .a(n32745), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_23_), .o(n32844) );
no02f01 g29054 ( .a(n32745), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_22_), .o(n32845) );
no04f01 g29055 ( .a(n32845), .b(n32844), .c(n32843), .d(n32839), .o(n32846) );
in01f01 g29056 ( .a(n32846), .o(n32847) );
no02f01 g29057 ( .a(n32847), .b(n32834), .o(n32848) );
in01f01 g29058 ( .a(n32848), .o(n32849) );
no02f01 g29059 ( .a(n32745), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_25_), .o(n32850) );
no02f01 g29060 ( .a(n32745), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_24_), .o(n32851) );
no02f01 g29061 ( .a(n32851), .b(n32850), .o(n32852) );
in01f01 g29062 ( .a(n32852), .o(n32853) );
no02f01 g29063 ( .a(n32745), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_26_), .o(n32854) );
no02f01 g29064 ( .a(n32745), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_27_), .o(n32855) );
no03f01 g29065 ( .a(n32855), .b(n32854), .c(n32853), .o(n32856) );
in01f01 g29066 ( .a(n32856), .o(n32857) );
no02f01 g29067 ( .a(n32745), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_30_), .o(n32858) );
no02f01 g29068 ( .a(n32745), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_28_), .o(n32859) );
no02f01 g29069 ( .a(n32745), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_29_), .o(n32860) );
no02f01 g29070 ( .a(n32860), .b(n32859), .o(n32861) );
in01f01 g29071 ( .a(n32861), .o(n32862) );
no04f01 g29072 ( .a(n32862), .b(n32858), .c(n32857), .d(n32849), .o(n32863) );
in01f01 g29073 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_16_), .o(n32864) );
in01f01 g29074 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_17_), .o(n32865) );
ao12f01 g29075 ( .a(n32744), .b(n32865), .c(n32864), .o(n32866) );
in01f01 g29076 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_19_), .o(n32867) );
in01f01 g29077 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_18_), .o(n32868) );
ao12f01 g29078 ( .a(n32744), .b(n32868), .c(n32867), .o(n32869) );
no02f01 g29079 ( .a(n32869), .b(n32866), .o(n32870) );
in01f01 g29080 ( .a(n32870), .o(n32871) );
in01f01 g29081 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_21_), .o(n32872) );
in01f01 g29082 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_20_), .o(n32873) );
ao12f01 g29083 ( .a(n32744), .b(n32873), .c(n32872), .o(n32874) );
no02f01 g29084 ( .a(n32874), .b(n32871), .o(n32875) );
in01f01 g29085 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_25_), .o(n32876) );
in01f01 g29086 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_24_), .o(n32877) );
ao12f01 g29087 ( .a(n32744), .b(n32877), .c(n32876), .o(n32878) );
in01f01 g29088 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_26_), .o(n32879) );
in01f01 g29089 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_27_), .o(n32880) );
ao12f01 g29090 ( .a(n32744), .b(n32880), .c(n32879), .o(n32881) );
in01f01 g29091 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_22_), .o(n32882) );
in01f01 g29092 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_23_), .o(n32883) );
ao12f01 g29093 ( .a(n32744), .b(n32883), .c(n32882), .o(n32884) );
no03f01 g29094 ( .a(n32884), .b(n32881), .c(n32878), .o(n32885) );
na02f01 g29095 ( .a(n32885), .b(n32875), .o(n32886) );
in01f01 g29096 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_28_), .o(n32887) );
in01f01 g29097 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_29_), .o(n32888) );
ao12f01 g29098 ( .a(n32744), .b(n32888), .c(n32887), .o(n32889) );
no02f01 g29099 ( .a(n32889), .b(n32886), .o(n32890) );
in01f01 g29100 ( .a(n32890), .o(n32891) );
na02f01 g29101 ( .a(n32745), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_30_), .o(n32892) );
in01f01 g29102 ( .a(n32892), .o(n32893) );
no03f01 g29103 ( .a(n32893), .b(n32891), .c(n32863), .o(n32894) );
no02f01 g29104 ( .a(n32745), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_31_), .o(n32895) );
na02f01 g29105 ( .a(n32745), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_31_), .o(n32896) );
in01f01 g29106 ( .a(n32896), .o(n32897) );
no02f01 g29107 ( .a(n32897), .b(n32895), .o(n32898) );
no02f01 g29108 ( .a(n32898), .b(n32894), .o(n32899) );
na02f01 g29109 ( .a(n32898), .b(n32894), .o(n32900) );
in01f01 g29110 ( .a(n32900), .o(n32901) );
no02f01 g29111 ( .a(n32901), .b(n32899), .o(n32902) );
in01f01 g29112 ( .a(delay_sub_ln23_0_unr28_stage10_stallmux_q), .o(n32903) );
no02f01 g29113 ( .a(n32902), .b(n32903), .o(n32904) );
no02f01 g29114 ( .a(n32744), .b(n32888), .o(n32905) );
no02f01 g29115 ( .a(n32905), .b(n32860), .o(n32906) );
in01f01 g29116 ( .a(n32906), .o(n32907) );
no02f01 g29117 ( .a(n32857), .b(n32847), .o(n32908) );
in01f01 g29118 ( .a(n32908), .o(n32909) );
no02f01 g29119 ( .a(n32909), .b(n32834), .o(n32910) );
in01f01 g29120 ( .a(n32910), .o(n32911) );
no02f01 g29121 ( .a(n32744), .b(n32887), .o(n32912) );
no02f01 g29122 ( .a(n32912), .b(n32886), .o(n32913) );
oa12f01 g29123 ( .a(n32913), .b(n32911), .c(n32859), .o(n32914) );
no02f01 g29124 ( .a(n32914), .b(n32907), .o(n32915) );
na02f01 g29125 ( .a(n32914), .b(n32907), .o(n32916) );
in01f01 g29126 ( .a(n32916), .o(n32917) );
no02f01 g29127 ( .a(n32917), .b(n32915), .o(n32918) );
no02f01 g29128 ( .a(n32918), .b(n32903), .o(n32919) );
no02f01 g29129 ( .a(n32893), .b(n32858), .o(n32920) );
ao12f01 g29130 ( .a(n32891), .b(n32910), .c(n32861), .o(n32921) );
na02f01 g29131 ( .a(n32921), .b(n32920), .o(n32922) );
in01f01 g29132 ( .a(n32922), .o(n32923) );
no02f01 g29133 ( .a(n32921), .b(n32920), .o(n32924) );
no02f01 g29134 ( .a(n32924), .b(n32923), .o(n32925) );
no02f01 g29135 ( .a(n32925), .b(n32903), .o(n32926) );
no02f01 g29136 ( .a(n32926), .b(n32919), .o(n32927) );
ao12f01 g29137 ( .a(n32904), .b(n32927), .c(n32902), .o(n32928) );
in01f01 g29138 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_6_), .o(n32929) );
in01f01 g29139 ( .a(delay_xor_ln22_unr28_stage10_stallmux_q_1_), .o(n32930) );
na02f01 g29140 ( .a(n_44610), .b(n32930), .o(n32931) );
in01f01 g29141 ( .a(delay_xor_ln22_unr28_stage10_stallmux_q_2_), .o(n32932) );
in01f01 g29142 ( .a(delay_xor_ln22_unr28_stage10_stallmux_q_0_), .o(n32933) );
oa12f01 g29143 ( .a(n_44610), .b(n32933), .c(n32932), .o(n32934) );
na02f01 g29144 ( .a(n32934), .b(n32931), .o(n32935) );
oa12f01 g29145 ( .a(delay_xor_ln22_unr28_stage10_stallmux_q_3_), .b(n32935), .c(n32736), .o(n32936) );
no02f01 g29146 ( .a(n32936), .b(n32929), .o(n32937) );
in01f01 g29147 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_5_), .o(n32938) );
in01f01 g29148 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_4_), .o(n32939) );
ao12f01 g29149 ( .a(n32936), .b(n32939), .c(n32938), .o(n32940) );
no02f01 g29150 ( .a(n32940), .b(n32937), .o(n32941) );
in01f01 g29151 ( .a(n32941), .o(n32942) );
in01f01 g29152 ( .a(n32936), .o(n32943) );
no02f01 g29153 ( .a(n32943), .b(delay_add_ln22_unr27_stage10_stallmux_q_6_), .o(n32944) );
na02f01 g29154 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_4_), .b(delay_add_ln22_unr27_stage10_stallmux_q_5_), .o(n32945) );
na02f01 g29155 ( .a(n32945), .b(n32936), .o(n32946) );
in01f01 g29156 ( .a(n32946), .o(n32947) );
no02f01 g29157 ( .a(n32947), .b(n32944), .o(n32948) );
in01f01 g29158 ( .a(delay_xor_ln22_unr28_stage10_stallmux_q_3_), .o(n32949) );
no02f01 g29159 ( .a(n_44610), .b(n32949), .o(n32950) );
no02f01 g29160 ( .a(n32736), .b(delay_xor_ln22_unr28_stage10_stallmux_q_3_), .o(n32951) );
no02f01 g29161 ( .a(n32951), .b(n32950), .o(n32952) );
na02f01 g29162 ( .a(n32952), .b(n32935), .o(n32953) );
no02f01 g29163 ( .a(n32952), .b(n32935), .o(n32954) );
in01f01 g29164 ( .a(n32954), .o(n32955) );
na02f01 g29165 ( .a(n32955), .b(n32953), .o(n32956) );
no02f01 g29166 ( .a(n32956), .b(delay_add_ln22_unr27_stage10_stallmux_q_3_), .o(n32957) );
in01f01 g29167 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_2_), .o(n32958) );
no02f01 g29168 ( .a(n_44610), .b(n32932), .o(n32959) );
no02f01 g29169 ( .a(n32736), .b(delay_xor_ln22_unr28_stage10_stallmux_q_2_), .o(n32960) );
no02f01 g29170 ( .a(n32960), .b(n32959), .o(n32961) );
ao12f01 g29171 ( .a(n32736), .b(delay_xor_ln22_unr28_stage10_stallmux_q_0_), .c(delay_xor_ln22_unr28_stage10_stallmux_q_1_), .o(n32962) );
no02f01 g29172 ( .a(n32961), .b(n32962), .o(n32963) );
no02f01 g29173 ( .a(delay_xor_ln22_unr28_stage10_stallmux_q_0_), .b(n32736), .o(n32964) );
in01f01 g29174 ( .a(n32964), .o(n32965) );
na02f01 g29175 ( .a(n32965), .b(n32931), .o(n32966) );
ao12f01 g29176 ( .a(n32963), .b(n32966), .c(n32961), .o(n32967) );
no02f01 g29177 ( .a(n32967), .b(n32958), .o(n32968) );
no02f01 g29178 ( .a(n32736), .b(delay_xor_ln22_unr28_stage10_stallmux_q_1_), .o(n32969) );
no02f01 g29179 ( .a(n_44610), .b(n32930), .o(n32970) );
no02f01 g29180 ( .a(n32970), .b(n32969), .o(n32971) );
na02f01 g29181 ( .a(n32971), .b(n32964), .o(n32972) );
oa12f01 g29182 ( .a(n32965), .b(n32970), .c(n32969), .o(n32973) );
na02f01 g29183 ( .a(n32973), .b(n32972), .o(n32974) );
na02f01 g29184 ( .a(n32974), .b(delay_add_ln22_unr27_stage10_stallmux_q_1_), .o(n32975) );
no02f01 g29185 ( .a(n32974), .b(delay_add_ln22_unr27_stage10_stallmux_q_1_), .o(n32976) );
in01f01 g29186 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_0_), .o(n32977) );
no02f01 g29187 ( .a(delay_xor_ln22_unr28_stage10_stallmux_q_0_), .b(n_44610), .o(n32978) );
no02f01 g29188 ( .a(n32933), .b(n32736), .o(n32979) );
no02f01 g29189 ( .a(n32979), .b(n32978), .o(n32980) );
in01f01 g29190 ( .a(n32980), .o(n32981) );
no02f01 g29191 ( .a(n32981), .b(n32977), .o(n32982) );
in01f01 g29192 ( .a(n32982), .o(n32983) );
oa12f01 g29193 ( .a(n32975), .b(n32983), .c(n32976), .o(n32984) );
na02f01 g29194 ( .a(n32967), .b(n32958), .o(n32985) );
ao12f01 g29195 ( .a(n32968), .b(n32985), .c(n32984), .o(n32986) );
in01f01 g29196 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_3_), .o(n32987) );
ao12f01 g29197 ( .a(n32987), .b(n32955), .c(n32953), .o(n32988) );
in01f01 g29198 ( .a(n32988), .o(n32989) );
ao12f01 g29199 ( .a(n32957), .b(n32989), .c(n32986), .o(n32990) );
ao12f01 g29200 ( .a(n32942), .b(n32990), .c(n32948), .o(n32991) );
no02f01 g29201 ( .a(n32943), .b(delay_add_ln22_unr27_stage10_stallmux_q_7_), .o(n32992) );
na02f01 g29202 ( .a(n32943), .b(delay_add_ln22_unr27_stage10_stallmux_q_7_), .o(n32993) );
in01f01 g29203 ( .a(n32993), .o(n32994) );
no02f01 g29204 ( .a(n32994), .b(n32992), .o(n32995) );
no02f01 g29205 ( .a(n32995), .b(n32991), .o(n32996) );
na02f01 g29206 ( .a(n32995), .b(n32991), .o(n32997) );
in01f01 g29207 ( .a(n32997), .o(n32998) );
no02f01 g29208 ( .a(n32998), .b(n32996), .o(n32999) );
in01f01 g29209 ( .a(n32999), .o(n33000) );
no02f01 g29210 ( .a(n33000), .b(n32928), .o(n33001) );
in01f01 g29211 ( .a(n32986), .o(n33002) );
no02f01 g29212 ( .a(n32988), .b(n32957), .o(n33003) );
in01f01 g29213 ( .a(n33003), .o(n33004) );
no02f01 g29214 ( .a(n33004), .b(n33002), .o(n33005) );
no02f01 g29215 ( .a(n33003), .b(n32986), .o(n33006) );
no02f01 g29216 ( .a(n33006), .b(n33005), .o(n33007) );
in01f01 g29217 ( .a(n33007), .o(n33008) );
no02f01 g29218 ( .a(n33008), .b(n32928), .o(n33009) );
in01f01 g29219 ( .a(n33009), .o(n33010) );
in01f01 g29220 ( .a(n32902), .o(n33011) );
no02f01 g29221 ( .a(n32927), .b(n33011), .o(n33012) );
no03f01 g29222 ( .a(n32926), .b(n32919), .c(n32902), .o(n33013) );
no02f01 g29223 ( .a(n33013), .b(n33012), .o(n33014) );
in01f01 g29224 ( .a(n32984), .o(n33015) );
in01f01 g29225 ( .a(n32985), .o(n33016) );
no02f01 g29226 ( .a(n33016), .b(n32968), .o(n33017) );
no02f01 g29227 ( .a(n33017), .b(n33015), .o(n33018) );
na02f01 g29228 ( .a(n33017), .b(n33015), .o(n33019) );
in01f01 g29229 ( .a(n33019), .o(n33020) );
no02f01 g29230 ( .a(n33020), .b(n33018), .o(n33021) );
no02f01 g29231 ( .a(n33021), .b(n33014), .o(n33022) );
in01f01 g29232 ( .a(n33021), .o(n33023) );
no03f01 g29233 ( .a(n33023), .b(n33013), .c(n33012), .o(n33024) );
in01f01 g29234 ( .a(n33024), .o(n33025) );
in01f01 g29235 ( .a(n32915), .o(n33026) );
na02f01 g29236 ( .a(n32916), .b(n33026), .o(n33027) );
na02f01 g29237 ( .a(n33027), .b(delay_sub_ln23_0_unr28_stage10_stallmux_q), .o(n33028) );
in01f01 g29238 ( .a(n32925), .o(n33029) );
na02f01 g29239 ( .a(n33029), .b(n33028), .o(n33030) );
na02f01 g29240 ( .a(n32925), .b(n32919), .o(n33031) );
na02f01 g29241 ( .a(n33031), .b(n33030), .o(n33032) );
in01f01 g29242 ( .a(n32975), .o(n33033) );
no03f01 g29243 ( .a(n32982), .b(n32976), .c(n33033), .o(n33034) );
in01f01 g29244 ( .a(n32976), .o(n33035) );
ao12f01 g29245 ( .a(n32983), .b(n33035), .c(n32975), .o(n33036) );
no02f01 g29246 ( .a(n33036), .b(n33034), .o(n33037) );
in01f01 g29247 ( .a(n33037), .o(n33038) );
no02f01 g29248 ( .a(n33038), .b(n33032), .o(n33039) );
no02f01 g29249 ( .a(n32980), .b(n32977), .o(n33040) );
no02f01 g29250 ( .a(n32981), .b(delay_add_ln22_unr27_stage10_stallmux_q_0_), .o(n33041) );
no02f01 g29251 ( .a(n33041), .b(n33040), .o(n33042) );
no02f01 g29252 ( .a(n33042), .b(n32918), .o(n33043) );
in01f01 g29253 ( .a(n33043), .o(n33044) );
na02f01 g29254 ( .a(n33038), .b(n33032), .o(n33045) );
oa12f01 g29255 ( .a(n33045), .b(n33044), .c(n33039), .o(n33046) );
ao12f01 g29256 ( .a(n33022), .b(n33046), .c(n33025), .o(n33047) );
in01f01 g29257 ( .a(n32928), .o(n33048) );
no02f01 g29258 ( .a(n33007), .b(n33048), .o(n33049) );
in01f01 g29259 ( .a(n33049), .o(n33050) );
na02f01 g29260 ( .a(n33050), .b(n33047), .o(n33051) );
na02f01 g29261 ( .a(n33051), .b(n33010), .o(n33052) );
no02f01 g29262 ( .a(n32936), .b(n32939), .o(n33053) );
no02f01 g29263 ( .a(n32943), .b(delay_add_ln22_unr27_stage10_stallmux_q_4_), .o(n33054) );
in01f01 g29264 ( .a(n33054), .o(n33055) );
ao12f01 g29265 ( .a(n33053), .b(n33055), .c(n32990), .o(n33056) );
in01f01 g29266 ( .a(n33056), .o(n33057) );
no02f01 g29267 ( .a(n32936), .b(n32938), .o(n33058) );
no02f01 g29268 ( .a(n32943), .b(delay_add_ln22_unr27_stage10_stallmux_q_5_), .o(n33059) );
no02f01 g29269 ( .a(n33059), .b(n33058), .o(n33060) );
in01f01 g29270 ( .a(n33060), .o(n33061) );
no02f01 g29271 ( .a(n33061), .b(n33057), .o(n33062) );
no02f01 g29272 ( .a(n33060), .b(n33056), .o(n33063) );
no02f01 g29273 ( .a(n33063), .b(n33062), .o(n33064) );
in01f01 g29274 ( .a(n33064), .o(n33065) );
no02f01 g29275 ( .a(n33054), .b(n33053), .o(n33066) );
in01f01 g29276 ( .a(n33066), .o(n33067) );
no02f01 g29277 ( .a(n33067), .b(n32990), .o(n33068) );
in01f01 g29278 ( .a(n32990), .o(n33069) );
no02f01 g29279 ( .a(n33066), .b(n33069), .o(n33070) );
no02f01 g29280 ( .a(n33070), .b(n33068), .o(n33071) );
in01f01 g29281 ( .a(n33071), .o(n33072) );
ao12f01 g29282 ( .a(n32928), .b(n33072), .c(n33065), .o(n33073) );
ao12f01 g29283 ( .a(n32940), .b(n32990), .c(n32946), .o(n33074) );
no02f01 g29284 ( .a(n32944), .b(n32937), .o(n33075) );
no02f01 g29285 ( .a(n33075), .b(n33074), .o(n33076) );
na02f01 g29286 ( .a(n33075), .b(n33074), .o(n33077) );
in01f01 g29287 ( .a(n33077), .o(n33078) );
no02f01 g29288 ( .a(n33078), .b(n33076), .o(n33079) );
in01f01 g29289 ( .a(n33079), .o(n33080) );
no02f01 g29290 ( .a(n33080), .b(n32928), .o(n33081) );
no02f01 g29291 ( .a(n33081), .b(n33073), .o(n33082) );
in01f01 g29292 ( .a(n33082), .o(n33083) );
no02f01 g29293 ( .a(n33083), .b(n33052), .o(n33084) );
in01f01 g29294 ( .a(n33084), .o(n33085) );
ao12f01 g29295 ( .a(n33048), .b(n33079), .c(n32999), .o(n33086) );
ao12f01 g29296 ( .a(n33048), .b(n33071), .c(n33064), .o(n33087) );
no02f01 g29297 ( .a(n33087), .b(n33086), .o(n33088) );
ao12f01 g29298 ( .a(n33001), .b(n33088), .c(n33085), .o(n33089) );
no02f01 g29299 ( .a(n32943), .b(delay_add_ln22_unr27_stage10_stallmux_q_10_), .o(n33090) );
no03f01 g29300 ( .a(n32992), .b(n32947), .c(n32944), .o(n33091) );
no02f01 g29301 ( .a(n32994), .b(n32942), .o(n33092) );
in01f01 g29302 ( .a(n33092), .o(n33093) );
ao12f01 g29303 ( .a(n33093), .b(n33091), .c(n32990), .o(n33094) );
ao12f01 g29304 ( .a(n32943), .b(delay_add_ln22_unr27_stage10_stallmux_q_8_), .c(delay_add_ln22_unr27_stage10_stallmux_q_9_), .o(n33095) );
no03f01 g29305 ( .a(n33095), .b(n33094), .c(n33090), .o(n33096) );
in01f01 g29306 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_10_), .o(n33097) );
no02f01 g29307 ( .a(n32936), .b(n33097), .o(n33098) );
in01f01 g29308 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_9_), .o(n33099) );
in01f01 g29309 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_8_), .o(n33100) );
ao12f01 g29310 ( .a(n32936), .b(n33100), .c(n33099), .o(n33101) );
no03f01 g29311 ( .a(n33101), .b(n33098), .c(n33096), .o(n33102) );
no02f01 g29312 ( .a(n32943), .b(delay_add_ln22_unr27_stage10_stallmux_q_11_), .o(n33103) );
in01f01 g29313 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_11_), .o(n33104) );
no02f01 g29314 ( .a(n32936), .b(n33104), .o(n33105) );
no02f01 g29315 ( .a(n33105), .b(n33103), .o(n33106) );
no02f01 g29316 ( .a(n33106), .b(n33102), .o(n33107) );
na02f01 g29317 ( .a(n33106), .b(n33102), .o(n33108) );
in01f01 g29318 ( .a(n33108), .o(n33109) );
no02f01 g29319 ( .a(n33109), .b(n33107), .o(n33110) );
in01f01 g29320 ( .a(n33110), .o(n33111) );
no02f01 g29321 ( .a(n33111), .b(n32928), .o(n33112) );
no02f01 g29322 ( .a(n32936), .b(n33100), .o(n33113) );
no02f01 g29323 ( .a(n32943), .b(delay_add_ln22_unr27_stage10_stallmux_q_8_), .o(n33114) );
no02f01 g29324 ( .a(n33114), .b(n33094), .o(n33115) );
no02f01 g29325 ( .a(n33115), .b(n33113), .o(n33116) );
no02f01 g29326 ( .a(n32943), .b(delay_add_ln22_unr27_stage10_stallmux_q_9_), .o(n33117) );
no02f01 g29327 ( .a(n32936), .b(n33099), .o(n33118) );
no02f01 g29328 ( .a(n33118), .b(n33117), .o(n33119) );
no02f01 g29329 ( .a(n33119), .b(n33116), .o(n33120) );
na02f01 g29330 ( .a(n33119), .b(n33116), .o(n33121) );
in01f01 g29331 ( .a(n33121), .o(n33122) );
no02f01 g29332 ( .a(n33122), .b(n33120), .o(n33123) );
in01f01 g29333 ( .a(n33123), .o(n33124) );
in01f01 g29334 ( .a(n33094), .o(n33125) );
no02f01 g29335 ( .a(n33114), .b(n33113), .o(n33126) );
in01f01 g29336 ( .a(n33126), .o(n33127) );
no02f01 g29337 ( .a(n33127), .b(n33125), .o(n33128) );
no02f01 g29338 ( .a(n33126), .b(n33094), .o(n33129) );
no02f01 g29339 ( .a(n33129), .b(n33128), .o(n33130) );
in01f01 g29340 ( .a(n33130), .o(n33131) );
ao12f01 g29341 ( .a(n32928), .b(n33131), .c(n33124), .o(n33132) );
no02f01 g29342 ( .a(n33095), .b(n33094), .o(n33133) );
no02f01 g29343 ( .a(n33098), .b(n33090), .o(n33134) );
in01f01 g29344 ( .a(n33134), .o(n33135) );
no03f01 g29345 ( .a(n33135), .b(n33101), .c(n33133), .o(n33136) );
no02f01 g29346 ( .a(n33101), .b(n33133), .o(n33137) );
no02f01 g29347 ( .a(n33134), .b(n33137), .o(n33138) );
no02f01 g29348 ( .a(n33138), .b(n33136), .o(n33139) );
in01f01 g29349 ( .a(n33139), .o(n33140) );
no02f01 g29350 ( .a(n33140), .b(n32928), .o(n33141) );
no03f01 g29351 ( .a(n33141), .b(n33132), .c(n33112), .o(n33142) );
na02f01 g29352 ( .a(n33142), .b(n33089), .o(n33143) );
ao12f01 g29353 ( .a(n33048), .b(n33139), .c(n33110), .o(n33144) );
ao12f01 g29354 ( .a(n33048), .b(n33130), .c(n33123), .o(n33145) );
no02f01 g29355 ( .a(n33145), .b(n33144), .o(n33146) );
na02f01 g29356 ( .a(n33146), .b(n33143), .o(n33147) );
no03f01 g29357 ( .a(n33103), .b(n33095), .c(n33090), .o(n33148) );
in01f01 g29358 ( .a(n33148), .o(n33149) );
no02f01 g29359 ( .a(n33149), .b(n33094), .o(n33150) );
in01f01 g29360 ( .a(n33150), .o(n33151) );
no02f01 g29361 ( .a(n32943), .b(delay_add_ln22_unr27_stage10_stallmux_q_12_), .o(n33152) );
no02f01 g29362 ( .a(n33152), .b(n33151), .o(n33153) );
ao12f01 g29363 ( .a(n32936), .b(n33097), .c(n33104), .o(n33154) );
no02f01 g29364 ( .a(n33154), .b(n33101), .o(n33155) );
in01f01 g29365 ( .a(n33155), .o(n33156) );
in01f01 g29366 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_12_), .o(n33157) );
no02f01 g29367 ( .a(n32936), .b(n33157), .o(n33158) );
no03f01 g29368 ( .a(n33158), .b(n33156), .c(n33153), .o(n33159) );
in01f01 g29369 ( .a(n33159), .o(n33160) );
no02f01 g29370 ( .a(n32943), .b(delay_add_ln22_unr27_stage10_stallmux_q_13_), .o(n33161) );
in01f01 g29371 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_13_), .o(n33162) );
no02f01 g29372 ( .a(n32936), .b(n33162), .o(n33163) );
no02f01 g29373 ( .a(n33163), .b(n33161), .o(n33164) );
in01f01 g29374 ( .a(n33164), .o(n33165) );
no02f01 g29375 ( .a(n33165), .b(n33160), .o(n33166) );
no02f01 g29376 ( .a(n33164), .b(n33159), .o(n33167) );
no02f01 g29377 ( .a(n33167), .b(n33166), .o(n33168) );
in01f01 g29378 ( .a(n33168), .o(n33169) );
no02f01 g29379 ( .a(n33169), .b(n32928), .o(n33170) );
no02f01 g29380 ( .a(n33158), .b(n33152), .o(n33171) );
in01f01 g29381 ( .a(n33171), .o(n33172) );
no03f01 g29382 ( .a(n33172), .b(n33156), .c(n33150), .o(n33173) );
ao12f01 g29383 ( .a(n33171), .b(n33155), .c(n33151), .o(n33174) );
no02f01 g29384 ( .a(n33174), .b(n33173), .o(n33175) );
in01f01 g29385 ( .a(n33175), .o(n33176) );
no02f01 g29386 ( .a(n33176), .b(n32928), .o(n33177) );
no02f01 g29387 ( .a(n33177), .b(n33170), .o(n33178) );
in01f01 g29388 ( .a(n33178), .o(n33179) );
ao12f01 g29389 ( .a(n32936), .b(n33157), .c(n33162), .o(n33180) );
no02f01 g29390 ( .a(n33180), .b(n33156), .o(n33181) );
in01f01 g29391 ( .a(n33181), .o(n33182) );
no02f01 g29392 ( .a(n33161), .b(n33152), .o(n33183) );
in01f01 g29393 ( .a(n33183), .o(n33184) );
no02f01 g29394 ( .a(n33184), .b(n33151), .o(n33185) );
no02f01 g29395 ( .a(n33185), .b(n33182), .o(n33186) );
in01f01 g29396 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_14_), .o(n33187) );
no02f01 g29397 ( .a(n32936), .b(n33187), .o(n33188) );
no02f01 g29398 ( .a(n32943), .b(delay_add_ln22_unr27_stage10_stallmux_q_14_), .o(n33189) );
no02f01 g29399 ( .a(n33189), .b(n33188), .o(n33190) );
no02f01 g29400 ( .a(n33190), .b(n33186), .o(n33191) );
na02f01 g29401 ( .a(n33190), .b(n33186), .o(n33192) );
in01f01 g29402 ( .a(n33192), .o(n33193) );
no02f01 g29403 ( .a(n33193), .b(n33191), .o(n33194) );
in01f01 g29404 ( .a(n33194), .o(n33195) );
no02f01 g29405 ( .a(n33195), .b(n32928), .o(n33196) );
in01f01 g29406 ( .a(n33189), .o(n33197) );
na02f01 g29407 ( .a(n33197), .b(n33185), .o(n33198) );
in01f01 g29408 ( .a(n33198), .o(n33199) );
no03f01 g29409 ( .a(n33199), .b(n33188), .c(n33182), .o(n33200) );
in01f01 g29410 ( .a(n33200), .o(n33201) );
no02f01 g29411 ( .a(n32943), .b(delay_add_ln22_unr27_stage10_stallmux_q_15_), .o(n33202) );
in01f01 g29412 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_15_), .o(n33203) );
no02f01 g29413 ( .a(n32936), .b(n33203), .o(n33204) );
no02f01 g29414 ( .a(n33204), .b(n33202), .o(n33205) );
in01f01 g29415 ( .a(n33205), .o(n33206) );
no02f01 g29416 ( .a(n33206), .b(n33201), .o(n33207) );
no02f01 g29417 ( .a(n33205), .b(n33200), .o(n33208) );
no02f01 g29418 ( .a(n33208), .b(n33207), .o(n33209) );
in01f01 g29419 ( .a(n33209), .o(n33210) );
no02f01 g29420 ( .a(n33210), .b(n32928), .o(n33211) );
no03f01 g29421 ( .a(n33211), .b(n33196), .c(n33179), .o(n33212) );
ao12f01 g29422 ( .a(n33048), .b(n33175), .c(n33168), .o(n33213) );
ao12f01 g29423 ( .a(n33048), .b(n33209), .c(n33194), .o(n33214) );
no02f01 g29424 ( .a(n33214), .b(n33213), .o(n33215) );
in01f01 g29425 ( .a(n33215), .o(n33216) );
ao12f01 g29426 ( .a(n33216), .b(n33212), .c(n33147), .o(n33217) );
no03f01 g29427 ( .a(n33202), .b(n33189), .c(n33184), .o(n33218) );
ao12f01 g29428 ( .a(n32936), .b(n33203), .c(n33187), .o(n33219) );
no02f01 g29429 ( .a(n33219), .b(n33182), .o(n33220) );
in01f01 g29430 ( .a(n33220), .o(n33221) );
ao12f01 g29431 ( .a(n33221), .b(n33218), .c(n33150), .o(n33222) );
ao12f01 g29432 ( .a(n32943), .b(delay_add_ln22_unr27_stage10_stallmux_q_17_), .c(delay_add_ln22_unr27_stage10_stallmux_q_16_), .o(n33223) );
no02f01 g29433 ( .a(n33223), .b(n33222), .o(n33224) );
no02f01 g29434 ( .a(n32943), .b(delay_add_ln22_unr27_stage10_stallmux_q_19_), .o(n33225) );
no02f01 g29435 ( .a(n32943), .b(delay_add_ln22_unr27_stage10_stallmux_q_18_), .o(n33226) );
no02f01 g29436 ( .a(n33226), .b(n33225), .o(n33227) );
na02f01 g29437 ( .a(n33227), .b(n33224), .o(n33228) );
no02f01 g29438 ( .a(n32943), .b(delay_add_ln22_unr27_stage10_stallmux_q_20_), .o(n33229) );
in01f01 g29439 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_16_), .o(n33230) );
in01f01 g29440 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_17_), .o(n33231) );
ao12f01 g29441 ( .a(n32936), .b(n33231), .c(n33230), .o(n33232) );
in01f01 g29442 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_19_), .o(n33233) );
in01f01 g29443 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_18_), .o(n33234) );
ao12f01 g29444 ( .a(n32936), .b(n33234), .c(n33233), .o(n33235) );
no02f01 g29445 ( .a(n33235), .b(n33232), .o(n33236) );
in01f01 g29446 ( .a(n33236), .o(n33237) );
in01f01 g29447 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_20_), .o(n33238) );
no02f01 g29448 ( .a(n32936), .b(n33238), .o(n33239) );
no02f01 g29449 ( .a(n33239), .b(n33237), .o(n33240) );
oa12f01 g29450 ( .a(n33240), .b(n33229), .c(n33228), .o(n33241) );
no02f01 g29451 ( .a(n32943), .b(delay_add_ln22_unr27_stage10_stallmux_q_21_), .o(n33242) );
in01f01 g29452 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_21_), .o(n33243) );
no02f01 g29453 ( .a(n32936), .b(n33243), .o(n33244) );
no02f01 g29454 ( .a(n33244), .b(n33242), .o(n33245) );
in01f01 g29455 ( .a(n33245), .o(n33246) );
no02f01 g29456 ( .a(n33246), .b(n33241), .o(n33247) );
na02f01 g29457 ( .a(n33246), .b(n33241), .o(n33248) );
in01f01 g29458 ( .a(n33248), .o(n33249) );
no02f01 g29459 ( .a(n33249), .b(n33247), .o(n33250) );
in01f01 g29460 ( .a(n33250), .o(n33251) );
no02f01 g29461 ( .a(n33251), .b(n32928), .o(n33252) );
in01f01 g29462 ( .a(n33222), .o(n33253) );
no02f01 g29463 ( .a(n32936), .b(n33230), .o(n33254) );
no02f01 g29464 ( .a(n32943), .b(delay_add_ln22_unr27_stage10_stallmux_q_16_), .o(n33255) );
no02f01 g29465 ( .a(n33255), .b(n33254), .o(n33256) );
in01f01 g29466 ( .a(n33256), .o(n33257) );
no02f01 g29467 ( .a(n33257), .b(n33253), .o(n33258) );
no02f01 g29468 ( .a(n33256), .b(n33222), .o(n33259) );
no02f01 g29469 ( .a(n33259), .b(n33258), .o(n33260) );
in01f01 g29470 ( .a(n33260), .o(n33261) );
no02f01 g29471 ( .a(n33261), .b(n32928), .o(n33262) );
ao12f01 g29472 ( .a(n32936), .b(n33243), .c(n33238), .o(n33263) );
no02f01 g29473 ( .a(n33263), .b(n33237), .o(n33264) );
in01f01 g29474 ( .a(n33264), .o(n33265) );
no02f01 g29475 ( .a(n33242), .b(n33229), .o(n33266) );
in01f01 g29476 ( .a(n33266), .o(n33267) );
no02f01 g29477 ( .a(n33267), .b(n33228), .o(n33268) );
no02f01 g29478 ( .a(n33268), .b(n33265), .o(n33269) );
no02f01 g29479 ( .a(n32943), .b(delay_add_ln22_unr27_stage10_stallmux_q_22_), .o(n33270) );
in01f01 g29480 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_22_), .o(n33271) );
no02f01 g29481 ( .a(n32936), .b(n33271), .o(n33272) );
no02f01 g29482 ( .a(n33272), .b(n33270), .o(n33273) );
no02f01 g29483 ( .a(n33273), .b(n33269), .o(n33274) );
na02f01 g29484 ( .a(n33273), .b(n33269), .o(n33275) );
in01f01 g29485 ( .a(n33275), .o(n33276) );
no02f01 g29486 ( .a(n33276), .b(n33274), .o(n33277) );
in01f01 g29487 ( .a(n33277), .o(n33278) );
no02f01 g29488 ( .a(n33278), .b(n32928), .o(n33279) );
in01f01 g29489 ( .a(n33270), .o(n33280) );
na02f01 g29490 ( .a(n33280), .b(n33268), .o(n33281) );
in01f01 g29491 ( .a(n33281), .o(n33282) );
no03f01 g29492 ( .a(n33282), .b(n33272), .c(n33265), .o(n33283) );
in01f01 g29493 ( .a(n33283), .o(n33284) );
no02f01 g29494 ( .a(n32943), .b(delay_add_ln22_unr27_stage10_stallmux_q_23_), .o(n33285) );
in01f01 g29495 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_23_), .o(n33286) );
no02f01 g29496 ( .a(n32936), .b(n33286), .o(n33287) );
no02f01 g29497 ( .a(n33287), .b(n33285), .o(n33288) );
in01f01 g29498 ( .a(n33288), .o(n33289) );
no02f01 g29499 ( .a(n33289), .b(n33284), .o(n33290) );
no02f01 g29500 ( .a(n33288), .b(n33283), .o(n33291) );
no02f01 g29501 ( .a(n33291), .b(n33290), .o(n33292) );
in01f01 g29502 ( .a(n33292), .o(n33293) );
no02f01 g29503 ( .a(n33293), .b(n32928), .o(n33294) );
no04f01 g29504 ( .a(n33294), .b(n33279), .c(n33262), .d(n33252), .o(n33295) );
no02f01 g29505 ( .a(n32936), .b(n33234), .o(n33296) );
no03f01 g29506 ( .a(n33226), .b(n33223), .c(n33222), .o(n33297) );
no03f01 g29507 ( .a(n33297), .b(n33296), .c(n33232), .o(n33298) );
in01f01 g29508 ( .a(n33298), .o(n33299) );
no02f01 g29509 ( .a(n32936), .b(n33233), .o(n33300) );
no02f01 g29510 ( .a(n33300), .b(n33225), .o(n33301) );
in01f01 g29511 ( .a(n33301), .o(n33302) );
no02f01 g29512 ( .a(n33302), .b(n33299), .o(n33303) );
no02f01 g29513 ( .a(n33301), .b(n33298), .o(n33304) );
no02f01 g29514 ( .a(n33304), .b(n33303), .o(n33305) );
in01f01 g29515 ( .a(n33305), .o(n33306) );
no02f01 g29516 ( .a(n33306), .b(n32928), .o(n33307) );
in01f01 g29517 ( .a(n33255), .o(n33308) );
ao12f01 g29518 ( .a(n33254), .b(n33308), .c(n33253), .o(n33309) );
in01f01 g29519 ( .a(n33309), .o(n33310) );
no02f01 g29520 ( .a(n32936), .b(n33231), .o(n33311) );
no02f01 g29521 ( .a(n32943), .b(delay_add_ln22_unr27_stage10_stallmux_q_17_), .o(n33312) );
no02f01 g29522 ( .a(n33312), .b(n33311), .o(n33313) );
in01f01 g29523 ( .a(n33313), .o(n33314) );
no02f01 g29524 ( .a(n33314), .b(n33310), .o(n33315) );
no02f01 g29525 ( .a(n33313), .b(n33309), .o(n33316) );
no02f01 g29526 ( .a(n33316), .b(n33315), .o(n33317) );
in01f01 g29527 ( .a(n33317), .o(n33318) );
no02f01 g29528 ( .a(n33318), .b(n32928), .o(n33319) );
in01f01 g29529 ( .a(n33228), .o(n33320) );
no02f01 g29530 ( .a(n33237), .b(n33320), .o(n33321) );
no02f01 g29531 ( .a(n33239), .b(n33229), .o(n33322) );
no02f01 g29532 ( .a(n33322), .b(n33321), .o(n33323) );
na02f01 g29533 ( .a(n33322), .b(n33321), .o(n33324) );
in01f01 g29534 ( .a(n33324), .o(n33325) );
no02f01 g29535 ( .a(n33325), .b(n33323), .o(n33326) );
in01f01 g29536 ( .a(n33326), .o(n33327) );
no02f01 g29537 ( .a(n33327), .b(n32928), .o(n33328) );
no02f01 g29538 ( .a(n33232), .b(n33224), .o(n33329) );
no02f01 g29539 ( .a(n33296), .b(n33226), .o(n33330) );
no02f01 g29540 ( .a(n33330), .b(n33329), .o(n33331) );
na02f01 g29541 ( .a(n33330), .b(n33329), .o(n33332) );
in01f01 g29542 ( .a(n33332), .o(n33333) );
no02f01 g29543 ( .a(n33333), .b(n33331), .o(n33334) );
in01f01 g29544 ( .a(n33334), .o(n33335) );
no02f01 g29545 ( .a(n33335), .b(n32928), .o(n33336) );
no04f01 g29546 ( .a(n33336), .b(n33328), .c(n33319), .d(n33307), .o(n33337) );
na02f01 g29547 ( .a(n33337), .b(n33295), .o(n33338) );
no02f01 g29548 ( .a(n33338), .b(n33217), .o(n33339) );
ao12f01 g29549 ( .a(n33048), .b(n33317), .c(n33260), .o(n33340) );
ao12f01 g29550 ( .a(n33048), .b(n33334), .c(n33305), .o(n33341) );
ao12f01 g29551 ( .a(n33048), .b(n33292), .c(n33277), .o(n33342) );
ao12f01 g29552 ( .a(n33048), .b(n33326), .c(n33250), .o(n33343) );
no04f01 g29553 ( .a(n33343), .b(n33342), .c(n33341), .d(n33340), .o(n33344) );
in01f01 g29554 ( .a(n33344), .o(n33345) );
no02f01 g29555 ( .a(n33345), .b(n33339), .o(n33346) );
in01f01 g29556 ( .a(n33346), .o(n33347) );
no03f01 g29557 ( .a(n33285), .b(n33270), .c(n33267), .o(n33348) );
in01f01 g29558 ( .a(n33348), .o(n33349) );
no02f01 g29559 ( .a(n33349), .b(n33228), .o(n33350) );
ao12f01 g29560 ( .a(n32936), .b(n33286), .c(n33271), .o(n33351) );
no02f01 g29561 ( .a(n33351), .b(n33265), .o(n33352) );
in01f01 g29562 ( .a(n33352), .o(n33353) );
no02f01 g29563 ( .a(n32943), .b(delay_add_ln22_unr27_stage10_stallmux_q_24_), .o(n33354) );
in01f01 g29564 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_24_), .o(n33355) );
no02f01 g29565 ( .a(n32936), .b(n33355), .o(n33356) );
no02f01 g29566 ( .a(n33356), .b(n33354), .o(n33357) );
in01f01 g29567 ( .a(n33357), .o(n33358) );
no03f01 g29568 ( .a(n33358), .b(n33353), .c(n33350), .o(n33359) );
in01f01 g29569 ( .a(n33350), .o(n33360) );
ao12f01 g29570 ( .a(n33357), .b(n33352), .c(n33360), .o(n33361) );
no02f01 g29571 ( .a(n33361), .b(n33359), .o(n33362) );
in01f01 g29572 ( .a(n33362), .o(n33363) );
no02f01 g29573 ( .a(n33363), .b(n32928), .o(n33364) );
no02f01 g29574 ( .a(n33354), .b(n33360), .o(n33365) );
no03f01 g29575 ( .a(n33365), .b(n33356), .c(n33353), .o(n33366) );
in01f01 g29576 ( .a(n33366), .o(n33367) );
no02f01 g29577 ( .a(n32943), .b(delay_add_ln22_unr27_stage10_stallmux_q_25_), .o(n33368) );
in01f01 g29578 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_25_), .o(n33369) );
no02f01 g29579 ( .a(n32936), .b(n33369), .o(n33370) );
no02f01 g29580 ( .a(n33370), .b(n33368), .o(n33371) );
in01f01 g29581 ( .a(n33371), .o(n33372) );
no02f01 g29582 ( .a(n33372), .b(n33367), .o(n33373) );
no02f01 g29583 ( .a(n33371), .b(n33366), .o(n33374) );
no02f01 g29584 ( .a(n33374), .b(n33373), .o(n33375) );
in01f01 g29585 ( .a(n33375), .o(n33376) );
no02f01 g29586 ( .a(n33376), .b(n32928), .o(n33377) );
no02f01 g29587 ( .a(n33377), .b(n33364), .o(n33378) );
no02f01 g29588 ( .a(n33368), .b(n33354), .o(n33379) );
in01f01 g29589 ( .a(n33379), .o(n33380) );
no02f01 g29590 ( .a(n32943), .b(delay_add_ln22_unr27_stage10_stallmux_q_26_), .o(n33381) );
no03f01 g29591 ( .a(n33381), .b(n33380), .c(n33360), .o(n33382) );
ao12f01 g29592 ( .a(n32936), .b(n33355), .c(n33369), .o(n33383) );
no02f01 g29593 ( .a(n33383), .b(n33353), .o(n33384) );
in01f01 g29594 ( .a(n33384), .o(n33385) );
in01f01 g29595 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_26_), .o(n33386) );
no02f01 g29596 ( .a(n32936), .b(n33386), .o(n33387) );
no03f01 g29597 ( .a(n33387), .b(n33385), .c(n33382), .o(n33388) );
in01f01 g29598 ( .a(n33388), .o(n33389) );
no02f01 g29599 ( .a(n32943), .b(delay_add_ln22_unr27_stage10_stallmux_q_27_), .o(n33390) );
in01f01 g29600 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_27_), .o(n33391) );
no02f01 g29601 ( .a(n32936), .b(n33391), .o(n33392) );
no02f01 g29602 ( .a(n33392), .b(n33390), .o(n33393) );
in01f01 g29603 ( .a(n33393), .o(n33394) );
no02f01 g29604 ( .a(n33394), .b(n33389), .o(n33395) );
no02f01 g29605 ( .a(n33393), .b(n33388), .o(n33396) );
no02f01 g29606 ( .a(n33396), .b(n33395), .o(n33397) );
in01f01 g29607 ( .a(n33397), .o(n33398) );
no02f01 g29608 ( .a(n33398), .b(n32928), .o(n33399) );
no02f01 g29609 ( .a(n33380), .b(n33360), .o(n33400) );
no02f01 g29610 ( .a(n33387), .b(n33381), .o(n33401) );
in01f01 g29611 ( .a(n33401), .o(n33402) );
no03f01 g29612 ( .a(n33402), .b(n33385), .c(n33400), .o(n33403) );
no02f01 g29613 ( .a(n33385), .b(n33400), .o(n33404) );
no02f01 g29614 ( .a(n33401), .b(n33404), .o(n33405) );
no02f01 g29615 ( .a(n33405), .b(n33403), .o(n33406) );
in01f01 g29616 ( .a(n33406), .o(n33407) );
no02f01 g29617 ( .a(n33407), .b(n32928), .o(n33408) );
no02f01 g29618 ( .a(n33408), .b(n33399), .o(n33409) );
na02f01 g29619 ( .a(n33409), .b(n33378), .o(n33410) );
no03f01 g29620 ( .a(n33390), .b(n33381), .c(n33380), .o(n33411) );
na02f01 g29621 ( .a(n33411), .b(n33350), .o(n33412) );
no02f01 g29622 ( .a(n32943), .b(delay_add_ln22_unr27_stage10_stallmux_q_28_), .o(n33413) );
no02f01 g29623 ( .a(n32943), .b(delay_add_ln22_unr27_stage10_stallmux_q_29_), .o(n33414) );
no02f01 g29624 ( .a(n33414), .b(n33413), .o(n33415) );
in01f01 g29625 ( .a(n33415), .o(n33416) );
no02f01 g29626 ( .a(n33416), .b(n33412), .o(n33417) );
ao12f01 g29627 ( .a(n32936), .b(n33386), .c(n33391), .o(n33418) );
no02f01 g29628 ( .a(n33418), .b(n33385), .o(n33419) );
in01f01 g29629 ( .a(n33419), .o(n33420) );
in01f01 g29630 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_28_), .o(n33421) );
in01f01 g29631 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_29_), .o(n33422) );
ao12f01 g29632 ( .a(n32936), .b(n33422), .c(n33421), .o(n33423) );
no03f01 g29633 ( .a(n33423), .b(n33420), .c(n33417), .o(n33424) );
no02f01 g29634 ( .a(n32943), .b(delay_add_ln22_unr27_stage10_stallmux_q_30_), .o(n33425) );
in01f01 g29635 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_30_), .o(n33426) );
no02f01 g29636 ( .a(n32936), .b(n33426), .o(n33427) );
no02f01 g29637 ( .a(n33427), .b(n33425), .o(n33428) );
na02f01 g29638 ( .a(n33428), .b(n33424), .o(n33429) );
no02f01 g29639 ( .a(n33428), .b(n33424), .o(n33430) );
in01f01 g29640 ( .a(n33430), .o(n33431) );
na02f01 g29641 ( .a(n33431), .b(n33429), .o(n33432) );
no02f01 g29642 ( .a(n33432), .b(n32928), .o(n33433) );
in01f01 g29643 ( .a(n33412), .o(n33434) );
no02f01 g29644 ( .a(n32936), .b(n33421), .o(n33435) );
no02f01 g29645 ( .a(n33435), .b(n33413), .o(n33436) );
in01f01 g29646 ( .a(n33436), .o(n33437) );
no03f01 g29647 ( .a(n33437), .b(n33420), .c(n33434), .o(n33438) );
ao12f01 g29648 ( .a(n33436), .b(n33419), .c(n33412), .o(n33439) );
no02f01 g29649 ( .a(n33439), .b(n33438), .o(n33440) );
in01f01 g29650 ( .a(n33440), .o(n33441) );
no02f01 g29651 ( .a(n33441), .b(n32928), .o(n33442) );
no02f01 g29652 ( .a(n32936), .b(n33422), .o(n33443) );
no02f01 g29653 ( .a(n33443), .b(n33414), .o(n33444) );
in01f01 g29654 ( .a(n33444), .o(n33445) );
no02f01 g29655 ( .a(n33435), .b(n33420), .o(n33446) );
oa12f01 g29656 ( .a(n33446), .b(n33413), .c(n33412), .o(n33447) );
no02f01 g29657 ( .a(n33447), .b(n33445), .o(n33448) );
in01f01 g29658 ( .a(n33448), .o(n33449) );
na02f01 g29659 ( .a(n33447), .b(n33445), .o(n33450) );
na02f01 g29660 ( .a(n33450), .b(n33449), .o(n33451) );
no02f01 g29661 ( .a(n33451), .b(n32928), .o(n33452) );
no02f01 g29662 ( .a(n33452), .b(n33442), .o(n33453) );
in01f01 g29663 ( .a(n33453), .o(n33454) );
no03f01 g29664 ( .a(n33454), .b(n33433), .c(n33410), .o(n33455) );
na02f01 g29665 ( .a(n33455), .b(n33347), .o(n33456) );
ao12f01 g29666 ( .a(n33048), .b(n33406), .c(n33397), .o(n33457) );
ao12f01 g29667 ( .a(n33048), .b(n33375), .c(n33362), .o(n33458) );
no02f01 g29668 ( .a(n33458), .b(n33457), .o(n33459) );
in01f01 g29669 ( .a(n33459), .o(n33460) );
in01f01 g29670 ( .a(n33429), .o(n33461) );
no02f01 g29671 ( .a(n33430), .b(n33461), .o(n33462) );
in01f01 g29672 ( .a(n33450), .o(n33463) );
no02f01 g29673 ( .a(n33463), .b(n33448), .o(n33464) );
ao12f01 g29674 ( .a(n33048), .b(n33464), .c(n33440), .o(n33465) );
in01f01 g29675 ( .a(n33465), .o(n33466) );
ao12f01 g29676 ( .a(n33048), .b(n33466), .c(n33462), .o(n33467) );
no02f01 g29677 ( .a(n33467), .b(n33460), .o(n33468) );
no02f01 g29678 ( .a(n33425), .b(n33416), .o(n33469) );
na02f01 g29679 ( .a(n33469), .b(n33434), .o(n33470) );
oa12f01 g29680 ( .a(n32943), .b(n33423), .c(delay_add_ln22_unr27_stage10_stallmux_q_30_), .o(n33471) );
na02f01 g29681 ( .a(n33471), .b(n33419), .o(n33472) );
ao12f01 g29682 ( .a(n33472), .b(n33469), .c(n33434), .o(n33473) );
in01f01 g29683 ( .a(n33473), .o(n33474) );
in01f01 g29684 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_31_), .o(n33475) );
no02f01 g29685 ( .a(n32936), .b(n33475), .o(n33476) );
no02f01 g29686 ( .a(n32943), .b(delay_add_ln22_unr27_stage10_stallmux_q_31_), .o(n33477) );
no02f01 g29687 ( .a(n33477), .b(n33476), .o(n33478) );
in01f01 g29688 ( .a(n33478), .o(n33479) );
no02f01 g29689 ( .a(n33479), .b(n33472), .o(n33480) );
ao22f01 g29690 ( .a(n33480), .b(n33470), .c(n33479), .d(n33474), .o(n33481) );
in01f01 g29691 ( .a(n33481), .o(n33482) );
no02f01 g29692 ( .a(n33482), .b(n32928), .o(n33483) );
no02f01 g29693 ( .a(n33481), .b(n33048), .o(n33484) );
no02f01 g29694 ( .a(n33484), .b(n33483), .o(n33485) );
na03f01 g29695 ( .a(n33485), .b(n33468), .c(n33456), .o(n33486) );
in01f01 g29696 ( .a(n33486), .o(n33487) );
ao12f01 g29697 ( .a(n33485), .b(n33468), .c(n33456), .o(n33488) );
no02f01 g29698 ( .a(n33488), .b(n33487), .o(n33489) );
na02f01 g29699 ( .a(n33489), .b(delay_sub_ln23_0_unr29_stage10_stallmux_q), .o(n33490) );
in01f01 g29700 ( .a(delay_sub_ln23_0_unr29_stage10_stallmux_q), .o(n33491) );
in01f01 g29701 ( .a(n33488), .o(n33492) );
na02f01 g29702 ( .a(n33492), .b(n33486), .o(n33493) );
na02f01 g29703 ( .a(n33493), .b(n33491), .o(n33494) );
no02f01 g29704 ( .a(n33462), .b(n33048), .o(n33495) );
no02f01 g29705 ( .a(n33495), .b(n33433), .o(n33496) );
no03f01 g29706 ( .a(n33410), .b(n33338), .c(n33217), .o(n33497) );
no02f01 g29707 ( .a(n33460), .b(n33345), .o(n33498) );
in01f01 g29708 ( .a(n33498), .o(n33499) );
no02f01 g29709 ( .a(n33499), .b(n33497), .o(n33500) );
no02f01 g29710 ( .a(n33500), .b(n33454), .o(n33501) );
in01f01 g29711 ( .a(n33501), .o(n33502) );
ao12f01 g29712 ( .a(n33496), .b(n33502), .c(n33466), .o(n33503) );
na03f01 g29713 ( .a(n33502), .b(n33496), .c(n33466), .o(n33504) );
in01f01 g29714 ( .a(n33504), .o(n33505) );
no02f01 g29715 ( .a(n33505), .b(n33503), .o(n33506) );
ao22f01 g29716 ( .a(n33506), .b(delay_sub_ln23_0_unr29_stage10_stallmux_q), .c(n33494), .d(n33490), .o(n33507) );
in01f01 g29717 ( .a(n33507), .o(n33508) );
no02f01 g29718 ( .a(n33481), .b(n32903), .o(n33509) );
no02f01 g29719 ( .a(n33464), .b(n32903), .o(n33510) );
ao12f01 g29720 ( .a(n33510), .b(n33432), .c(delay_sub_ln23_0_unr28_stage10_stallmux_q), .o(n33511) );
ao12f01 g29721 ( .a(n33509), .b(n33511), .c(n33481), .o(n33512) );
in01f01 g29722 ( .a(n33512), .o(n33513) );
no03f01 g29723 ( .a(n32787), .b(n32785), .c(n32754), .o(n33514) );
in01f01 g29724 ( .a(n32764), .o(n33515) );
na02f01 g29725 ( .a(n32736), .b(delay_xor_ln21_unr28_stage10_stallmux_q_1_), .o(n33516) );
ao12f01 g29726 ( .a(n32740), .b(n33516), .c(n32767), .o(n33517) );
ao12f01 g29727 ( .a(n33517), .b(n32740), .c(n32767), .o(n33518) );
na02f01 g29728 ( .a(n33518), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_1_), .o(n33519) );
no02f01 g29729 ( .a(n33518), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_1_), .o(n33520) );
oa12f01 g29730 ( .a(n33519), .b(n32779), .c(n33520), .o(n33521) );
ao12f01 g29731 ( .a(n33515), .b(n32783), .c(n33521), .o(n33522) );
in01f01 g29732 ( .a(n32787), .o(n33523) );
ao12f01 g29733 ( .a(n33522), .b(n33523), .c(n32755), .o(n33524) );
no02f01 g29734 ( .a(n33524), .b(n33514), .o(n33525) );
in01f01 g29735 ( .a(n33525), .o(n33526) );
no02f01 g29736 ( .a(n33526), .b(n33513), .o(n33527) );
in01f01 g29737 ( .a(n33527), .o(n33528) );
na02f01 g29738 ( .a(n33511), .b(n33482), .o(n33529) );
na02f01 g29739 ( .a(n33451), .b(delay_sub_ln23_0_unr28_stage10_stallmux_q), .o(n33530) );
oa12f01 g29740 ( .a(n33530), .b(n33462), .c(n32903), .o(n33531) );
na02f01 g29741 ( .a(n33531), .b(n33481), .o(n33532) );
na02f01 g29742 ( .a(n33532), .b(n33529), .o(n33533) );
no03f01 g29743 ( .a(n32784), .b(n33521), .c(n33515), .o(n33534) );
ao12f01 g29744 ( .a(n32781), .b(n32783), .c(n32764), .o(n33535) );
no02f01 g29745 ( .a(n33535), .b(n33534), .o(n33536) );
no02f01 g29746 ( .a(n33536), .b(n33533), .o(n33537) );
na02f01 g29747 ( .a(n33510), .b(n33462), .o(n33538) );
na02f01 g29748 ( .a(n33530), .b(n33432), .o(n33539) );
no03f01 g29749 ( .a(n32780), .b(n33520), .c(n32772), .o(n33540) );
ao12f01 g29750 ( .a(n32779), .b(n32773), .c(n33519), .o(n33541) );
no02f01 g29751 ( .a(n33541), .b(n33540), .o(n33542) );
in01f01 g29752 ( .a(n33542), .o(n33543) );
ao12f01 g29753 ( .a(n33543), .b(n33539), .c(n33538), .o(n33544) );
no02f01 g29754 ( .a(n32777), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_0_), .o(n33545) );
in01f01 g29755 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_0_), .o(n33546) );
no02f01 g29756 ( .a(n32778), .b(n33546), .o(n33547) );
no02f01 g29757 ( .a(n33547), .b(n33545), .o(n33548) );
no02f01 g29758 ( .a(n33548), .b(n33464), .o(n33549) );
na02f01 g29759 ( .a(n33539), .b(n33538), .o(n33550) );
no02f01 g29760 ( .a(n33542), .b(n33550), .o(n33551) );
in01f01 g29761 ( .a(n33551), .o(n33552) );
oa12f01 g29762 ( .a(n33552), .b(n33549), .c(n33544), .o(n33553) );
in01f01 g29763 ( .a(n33536), .o(n33554) );
ao12f01 g29764 ( .a(n33554), .b(n33532), .c(n33529), .o(n33555) );
in01f01 g29765 ( .a(n33555), .o(n33556) );
ao12f01 g29766 ( .a(n33537), .b(n33556), .c(n33553), .o(n33557) );
no02f01 g29767 ( .a(n33525), .b(n33512), .o(n33558) );
in01f01 g29768 ( .a(n33558), .o(n33559) );
na02f01 g29769 ( .a(n33559), .b(n33557), .o(n33560) );
na02f01 g29770 ( .a(n33560), .b(n33528), .o(n33561) );
ao12f01 g29771 ( .a(n32754), .b(n33523), .c(n33522), .o(n33562) );
in01f01 g29772 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_4_), .o(n33563) );
no02f01 g29773 ( .a(n32744), .b(n33563), .o(n33564) );
no02f01 g29774 ( .a(n32745), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_4_), .o(n33565) );
in01f01 g29775 ( .a(n33565), .o(n33566) );
ao12f01 g29776 ( .a(n33564), .b(n33566), .c(n33562), .o(n33567) );
in01f01 g29777 ( .a(n33567), .o(n33568) );
no02f01 g29778 ( .a(n32745), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_5_), .o(n33569) );
in01f01 g29779 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_5_), .o(n33570) );
no02f01 g29780 ( .a(n32744), .b(n33570), .o(n33571) );
no02f01 g29781 ( .a(n33571), .b(n33569), .o(n33572) );
in01f01 g29782 ( .a(n33572), .o(n33573) );
no02f01 g29783 ( .a(n33573), .b(n33568), .o(n33574) );
no02f01 g29784 ( .a(n33572), .b(n33567), .o(n33575) );
no02f01 g29785 ( .a(n33575), .b(n33574), .o(n33576) );
in01f01 g29786 ( .a(n33576), .o(n33577) );
no02f01 g29787 ( .a(n33577), .b(n33513), .o(n33578) );
no02f01 g29788 ( .a(n33565), .b(n33564), .o(n33579) );
no02f01 g29789 ( .a(n33579), .b(n32788), .o(n33580) );
na02f01 g29790 ( .a(n33579), .b(n32788), .o(n33581) );
in01f01 g29791 ( .a(n33581), .o(n33582) );
no02f01 g29792 ( .a(n33582), .b(n33580), .o(n33583) );
in01f01 g29793 ( .a(n33583), .o(n33584) );
no02f01 g29794 ( .a(n33584), .b(n33513), .o(n33585) );
oa22f01 g29795 ( .a(n32797), .b(n32744), .c(n32790), .d(n32788), .o(n33586) );
in01f01 g29796 ( .a(n33586), .o(n33587) );
no02f01 g29797 ( .a(n32744), .b(n32796), .o(n33588) );
no02f01 g29798 ( .a(n33588), .b(n32789), .o(n33589) );
no02f01 g29799 ( .a(n33589), .b(n33587), .o(n33590) );
na02f01 g29800 ( .a(n33589), .b(n33587), .o(n33591) );
in01f01 g29801 ( .a(n33591), .o(n33592) );
no02f01 g29802 ( .a(n33592), .b(n33590), .o(n33593) );
in01f01 g29803 ( .a(n33593), .o(n33594) );
no02f01 g29804 ( .a(n33594), .b(n33513), .o(n33595) );
no03f01 g29805 ( .a(n33595), .b(n33585), .c(n33578), .o(n33596) );
no02f01 g29806 ( .a(n32798), .b(n32793), .o(n33597) );
no02f01 g29807 ( .a(n32800), .b(n32794), .o(n33598) );
no02f01 g29808 ( .a(n33598), .b(n33597), .o(n33599) );
na02f01 g29809 ( .a(n33598), .b(n33597), .o(n33600) );
in01f01 g29810 ( .a(n33600), .o(n33601) );
no02f01 g29811 ( .a(n33601), .b(n33599), .o(n33602) );
in01f01 g29812 ( .a(n33602), .o(n33603) );
no02f01 g29813 ( .a(n33603), .b(n33513), .o(n33604) );
in01f01 g29814 ( .a(n33604), .o(n33605) );
na02f01 g29815 ( .a(n33605), .b(n33596), .o(n33606) );
ao12f01 g29816 ( .a(n33512), .b(n33602), .c(n33593), .o(n33607) );
ao12f01 g29817 ( .a(n33512), .b(n33583), .c(n33576), .o(n33608) );
no02f01 g29818 ( .a(n33608), .b(n33607), .o(n33609) );
oa12f01 g29819 ( .a(n33609), .b(n33606), .c(n33561), .o(n33610) );
na02f01 g29820 ( .a(n32791), .b(n33562), .o(n33611) );
oa12f01 g29821 ( .a(n32801), .b(n32794), .c(n33611), .o(n33612) );
no02f01 g29822 ( .a(n32744), .b(n32823), .o(n33613) );
no02f01 g29823 ( .a(n32745), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_8_), .o(n33614) );
in01f01 g29824 ( .a(n33614), .o(n33615) );
ao12f01 g29825 ( .a(n33613), .b(n33615), .c(n33612), .o(n33616) );
no02f01 g29826 ( .a(n32745), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_9_), .o(n33617) );
no02f01 g29827 ( .a(n32744), .b(n32822), .o(n33618) );
no02f01 g29828 ( .a(n33618), .b(n33617), .o(n33619) );
no02f01 g29829 ( .a(n33619), .b(n33616), .o(n33620) );
na02f01 g29830 ( .a(n33619), .b(n33616), .o(n33621) );
in01f01 g29831 ( .a(n33621), .o(n33622) );
no02f01 g29832 ( .a(n33622), .b(n33620), .o(n33623) );
in01f01 g29833 ( .a(n33623), .o(n33624) );
no02f01 g29834 ( .a(n33624), .b(n33513), .o(n33625) );
no02f01 g29835 ( .a(n33614), .b(n33613), .o(n33626) );
in01f01 g29836 ( .a(n33626), .o(n33627) );
no02f01 g29837 ( .a(n33627), .b(n33612), .o(n33628) );
no02f01 g29838 ( .a(n33626), .b(n32803), .o(n33629) );
no02f01 g29839 ( .a(n33629), .b(n33628), .o(n33630) );
in01f01 g29840 ( .a(n33630), .o(n33631) );
no02f01 g29841 ( .a(n33631), .b(n33513), .o(n33632) );
no02f01 g29842 ( .a(n33632), .b(n33625), .o(n33633) );
in01f01 g29843 ( .a(n33633), .o(n33634) );
no02f01 g29844 ( .a(n32744), .b(n32820), .o(n33635) );
no03f01 g29845 ( .a(n32805), .b(n32804), .c(n32803), .o(n33636) );
no03f01 g29846 ( .a(n33636), .b(n32824), .c(n33635), .o(n33637) );
no02f01 g29847 ( .a(n32744), .b(n32819), .o(n33638) );
no02f01 g29848 ( .a(n33638), .b(n32806), .o(n33639) );
no02f01 g29849 ( .a(n33639), .b(n33637), .o(n33640) );
na02f01 g29850 ( .a(n33639), .b(n33637), .o(n33641) );
in01f01 g29851 ( .a(n33641), .o(n33642) );
no02f01 g29852 ( .a(n33642), .b(n33640), .o(n33643) );
in01f01 g29853 ( .a(n33643), .o(n33644) );
no02f01 g29854 ( .a(n33644), .b(n33513), .o(n33645) );
no02f01 g29855 ( .a(n32804), .b(n32803), .o(n33646) );
no02f01 g29856 ( .a(n33635), .b(n32805), .o(n33647) );
in01f01 g29857 ( .a(n33647), .o(n33648) );
no03f01 g29858 ( .a(n33648), .b(n33646), .c(n32824), .o(n33649) );
no02f01 g29859 ( .a(n33646), .b(n32824), .o(n33650) );
no02f01 g29860 ( .a(n33647), .b(n33650), .o(n33651) );
no02f01 g29861 ( .a(n33651), .b(n33649), .o(n33652) );
in01f01 g29862 ( .a(n33652), .o(n33653) );
no02f01 g29863 ( .a(n33653), .b(n33513), .o(n33654) );
no03f01 g29864 ( .a(n33654), .b(n33645), .c(n33634), .o(n33655) );
na02f01 g29865 ( .a(n33655), .b(n33610), .o(n33656) );
ao12f01 g29866 ( .a(n33512), .b(n33630), .c(n33623), .o(n33657) );
ao12f01 g29867 ( .a(n33512), .b(n33652), .c(n33643), .o(n33658) );
no02f01 g29868 ( .a(n33658), .b(n33657), .o(n33659) );
na02f01 g29869 ( .a(n33659), .b(n33656), .o(n33660) );
no02f01 g29870 ( .a(n32744), .b(n32816), .o(n33661) );
no03f01 g29871 ( .a(n32809), .b(n32808), .c(n32803), .o(n33662) );
no03f01 g29872 ( .a(n33662), .b(n32826), .c(n33661), .o(n33663) );
in01f01 g29873 ( .a(n33663), .o(n33664) );
no02f01 g29874 ( .a(n32744), .b(n32817), .o(n33665) );
no02f01 g29875 ( .a(n33665), .b(n32810), .o(n33666) );
in01f01 g29876 ( .a(n33666), .o(n33667) );
no02f01 g29877 ( .a(n33667), .b(n33664), .o(n33668) );
no02f01 g29878 ( .a(n33666), .b(n33663), .o(n33669) );
no02f01 g29879 ( .a(n33669), .b(n33668), .o(n33670) );
in01f01 g29880 ( .a(n33670), .o(n33671) );
no02f01 g29881 ( .a(n33671), .b(n33513), .o(n33672) );
no02f01 g29882 ( .a(n32808), .b(n32803), .o(n33673) );
no02f01 g29883 ( .a(n33661), .b(n32809), .o(n33674) );
in01f01 g29884 ( .a(n33674), .o(n33675) );
no03f01 g29885 ( .a(n33675), .b(n33673), .c(n32826), .o(n33676) );
no02f01 g29886 ( .a(n33673), .b(n32826), .o(n33677) );
no02f01 g29887 ( .a(n33674), .b(n33677), .o(n33678) );
no02f01 g29888 ( .a(n33678), .b(n33676), .o(n33679) );
in01f01 g29889 ( .a(n33679), .o(n33680) );
no02f01 g29890 ( .a(n33680), .b(n33513), .o(n33681) );
no02f01 g29891 ( .a(n33681), .b(n33672), .o(n33682) );
na02f01 g29892 ( .a(n33682), .b(n33660), .o(n33683) );
no02f01 g29893 ( .a(n32744), .b(n32830), .o(n33684) );
no03f01 g29894 ( .a(n33684), .b(n32828), .c(n32813), .o(n33685) );
no02f01 g29895 ( .a(n32744), .b(n32829), .o(n33686) );
no02f01 g29896 ( .a(n33686), .b(n32814), .o(n33687) );
no02f01 g29897 ( .a(n33687), .b(n33685), .o(n33688) );
na02f01 g29898 ( .a(n33687), .b(n33685), .o(n33689) );
in01f01 g29899 ( .a(n33689), .o(n33690) );
no02f01 g29900 ( .a(n33690), .b(n33688), .o(n33691) );
in01f01 g29901 ( .a(n33691), .o(n33692) );
no02f01 g29902 ( .a(n33692), .b(n33513), .o(n33693) );
ao12f01 g29903 ( .a(n32828), .b(n32811), .c(n33612), .o(n33694) );
no02f01 g29904 ( .a(n33684), .b(n32746), .o(n33695) );
no02f01 g29905 ( .a(n33695), .b(n33694), .o(n33696) );
na02f01 g29906 ( .a(n33695), .b(n33694), .o(n33697) );
in01f01 g29907 ( .a(n33697), .o(n33698) );
no02f01 g29908 ( .a(n33698), .b(n33696), .o(n33699) );
in01f01 g29909 ( .a(n33699), .o(n33700) );
no02f01 g29910 ( .a(n33700), .b(n33513), .o(n33701) );
no02f01 g29911 ( .a(n33701), .b(n33693), .o(n33702) );
in01f01 g29912 ( .a(n33702), .o(n33703) );
ao12f01 g29913 ( .a(n33512), .b(n33679), .c(n33670), .o(n33704) );
ao12f01 g29914 ( .a(n33512), .b(n33699), .c(n33691), .o(n33705) );
no02f01 g29915 ( .a(n33705), .b(n33704), .o(n33706) );
oa12f01 g29916 ( .a(n33706), .b(n33703), .c(n33683), .o(n33707) );
in01f01 g29917 ( .a(n33707), .o(n33708) );
in01f01 g29918 ( .a(n32834), .o(n33709) );
no02f01 g29919 ( .a(n32744), .b(n32864), .o(n33710) );
no02f01 g29920 ( .a(n32745), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_16_), .o(n33711) );
in01f01 g29921 ( .a(n33711), .o(n33712) );
ao12f01 g29922 ( .a(n33710), .b(n33712), .c(n33709), .o(n33713) );
in01f01 g29923 ( .a(n33713), .o(n33714) );
no02f01 g29924 ( .a(n32745), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_17_), .o(n33715) );
no02f01 g29925 ( .a(n32744), .b(n32865), .o(n33716) );
no02f01 g29926 ( .a(n33716), .b(n33715), .o(n33717) );
in01f01 g29927 ( .a(n33717), .o(n33718) );
no02f01 g29928 ( .a(n33718), .b(n33714), .o(n33719) );
no02f01 g29929 ( .a(n33717), .b(n33713), .o(n33720) );
no02f01 g29930 ( .a(n33720), .b(n33719), .o(n33721) );
in01f01 g29931 ( .a(n33721), .o(n33722) );
no02f01 g29932 ( .a(n33711), .b(n33710), .o(n33723) );
no02f01 g29933 ( .a(n33723), .b(n32834), .o(n33724) );
na02f01 g29934 ( .a(n33723), .b(n32834), .o(n33725) );
in01f01 g29935 ( .a(n33725), .o(n33726) );
no02f01 g29936 ( .a(n33726), .b(n33724), .o(n33727) );
in01f01 g29937 ( .a(n33727), .o(n33728) );
ao12f01 g29938 ( .a(n33513), .b(n33728), .c(n33722), .o(n33729) );
no02f01 g29939 ( .a(n32744), .b(n32868), .o(n33730) );
no03f01 g29940 ( .a(n32836), .b(n32835), .c(n32834), .o(n33731) );
no03f01 g29941 ( .a(n33731), .b(n33730), .c(n32866), .o(n33732) );
no02f01 g29942 ( .a(n32744), .b(n32867), .o(n33733) );
no02f01 g29943 ( .a(n33733), .b(n32837), .o(n33734) );
no02f01 g29944 ( .a(n33734), .b(n33732), .o(n33735) );
na02f01 g29945 ( .a(n33734), .b(n33732), .o(n33736) );
in01f01 g29946 ( .a(n33736), .o(n33737) );
no02f01 g29947 ( .a(n33737), .b(n33735), .o(n33738) );
in01f01 g29948 ( .a(n33738), .o(n33739) );
no02f01 g29949 ( .a(n33739), .b(n33513), .o(n33740) );
no02f01 g29950 ( .a(n32836), .b(n32834), .o(n33741) );
no02f01 g29951 ( .a(n33730), .b(n32835), .o(n33742) );
in01f01 g29952 ( .a(n33742), .o(n33743) );
no03f01 g29953 ( .a(n33743), .b(n33741), .c(n32866), .o(n33744) );
no02f01 g29954 ( .a(n33741), .b(n32866), .o(n33745) );
no02f01 g29955 ( .a(n33742), .b(n33745), .o(n33746) );
no02f01 g29956 ( .a(n33746), .b(n33744), .o(n33747) );
in01f01 g29957 ( .a(n33747), .o(n33748) );
no02f01 g29958 ( .a(n33748), .b(n33513), .o(n33749) );
no03f01 g29959 ( .a(n33749), .b(n33740), .c(n33729), .o(n33750) );
in01f01 g29960 ( .a(n33750), .o(n33751) );
no02f01 g29961 ( .a(n33751), .b(n33708), .o(n33752) );
in01f01 g29962 ( .a(n33752), .o(n33753) );
no02f01 g29963 ( .a(n32744), .b(n32873), .o(n33754) );
no02f01 g29964 ( .a(n32839), .b(n32834), .o(n33755) );
in01f01 g29965 ( .a(n33755), .o(n33756) );
no02f01 g29966 ( .a(n33756), .b(n32841), .o(n33757) );
no03f01 g29967 ( .a(n33757), .b(n33754), .c(n32871), .o(n33758) );
no02f01 g29968 ( .a(n32744), .b(n32872), .o(n33759) );
no02f01 g29969 ( .a(n33759), .b(n32840), .o(n33760) );
no02f01 g29970 ( .a(n33760), .b(n33758), .o(n33761) );
na02f01 g29971 ( .a(n33760), .b(n33758), .o(n33762) );
in01f01 g29972 ( .a(n33762), .o(n33763) );
no02f01 g29973 ( .a(n33763), .b(n33761), .o(n33764) );
in01f01 g29974 ( .a(n33764), .o(n33765) );
no02f01 g29975 ( .a(n33765), .b(n33513), .o(n33766) );
no02f01 g29976 ( .a(n33754), .b(n32841), .o(n33767) );
in01f01 g29977 ( .a(n33767), .o(n33768) );
no03f01 g29978 ( .a(n33768), .b(n33755), .c(n32871), .o(n33769) );
ao12f01 g29979 ( .a(n33767), .b(n33756), .c(n32870), .o(n33770) );
no02f01 g29980 ( .a(n33770), .b(n33769), .o(n33771) );
in01f01 g29981 ( .a(n33771), .o(n33772) );
no02f01 g29982 ( .a(n33772), .b(n33513), .o(n33773) );
in01f01 g29983 ( .a(n32875), .o(n33774) );
no02f01 g29984 ( .a(n33756), .b(n32843), .o(n33775) );
no02f01 g29985 ( .a(n32744), .b(n32882), .o(n33776) );
no02f01 g29986 ( .a(n33776), .b(n32845), .o(n33777) );
in01f01 g29987 ( .a(n33777), .o(n33778) );
no03f01 g29988 ( .a(n33778), .b(n33775), .c(n33774), .o(n33779) );
no02f01 g29989 ( .a(n33775), .b(n33774), .o(n33780) );
no02f01 g29990 ( .a(n33777), .b(n33780), .o(n33781) );
no02f01 g29991 ( .a(n33781), .b(n33779), .o(n33782) );
in01f01 g29992 ( .a(n33782), .o(n33783) );
no02f01 g29993 ( .a(n33783), .b(n33513), .o(n33784) );
no03f01 g29994 ( .a(n33756), .b(n32845), .c(n32843), .o(n33785) );
no03f01 g29995 ( .a(n33785), .b(n33776), .c(n33774), .o(n33786) );
no02f01 g29996 ( .a(n32744), .b(n32883), .o(n33787) );
no02f01 g29997 ( .a(n33787), .b(n32844), .o(n33788) );
no02f01 g29998 ( .a(n33788), .b(n33786), .o(n33789) );
na02f01 g29999 ( .a(n33788), .b(n33786), .o(n33790) );
in01f01 g30000 ( .a(n33790), .o(n33791) );
no02f01 g30001 ( .a(n33791), .b(n33789), .o(n33792) );
in01f01 g30002 ( .a(n33792), .o(n33793) );
no02f01 g30003 ( .a(n33793), .b(n33513), .o(n33794) );
no04f01 g30004 ( .a(n33794), .b(n33784), .c(n33773), .d(n33766), .o(n33795) );
in01f01 g30005 ( .a(n33795), .o(n33796) );
no02f01 g30006 ( .a(n33796), .b(n33753), .o(n33797) );
ao12f01 g30007 ( .a(n33512), .b(n33727), .c(n33721), .o(n33798) );
ao12f01 g30008 ( .a(n33512), .b(n33747), .c(n33738), .o(n33799) );
no02f01 g30009 ( .a(n33799), .b(n33798), .o(n33800) );
in01f01 g30010 ( .a(n33800), .o(n33801) );
ao12f01 g30011 ( .a(n33512), .b(n33771), .c(n33764), .o(n33802) );
ao12f01 g30012 ( .a(n33512), .b(n33792), .c(n33782), .o(n33803) );
no03f01 g30013 ( .a(n33803), .b(n33802), .c(n33801), .o(n33804) );
in01f01 g30014 ( .a(n33804), .o(n33805) );
no02f01 g30015 ( .a(n33805), .b(n33797), .o(n33806) );
no02f01 g30016 ( .a(n32884), .b(n33774), .o(n33807) );
in01f01 g30017 ( .a(n33807), .o(n33808) );
no02f01 g30018 ( .a(n32744), .b(n32877), .o(n33809) );
no02f01 g30019 ( .a(n33809), .b(n32851), .o(n33810) );
in01f01 g30020 ( .a(n33810), .o(n33811) );
no03f01 g30021 ( .a(n33811), .b(n33808), .c(n32848), .o(n33812) );
ao12f01 g30022 ( .a(n33810), .b(n33807), .c(n32849), .o(n33813) );
no02f01 g30023 ( .a(n33813), .b(n33812), .o(n33814) );
in01f01 g30024 ( .a(n33814), .o(n33815) );
no02f01 g30025 ( .a(n33815), .b(n33513), .o(n33816) );
no02f01 g30026 ( .a(n32851), .b(n32849), .o(n33817) );
no03f01 g30027 ( .a(n33817), .b(n33808), .c(n33809), .o(n33818) );
in01f01 g30028 ( .a(n33818), .o(n33819) );
no02f01 g30029 ( .a(n32744), .b(n32876), .o(n33820) );
no02f01 g30030 ( .a(n33820), .b(n32850), .o(n33821) );
in01f01 g30031 ( .a(n33821), .o(n33822) );
no02f01 g30032 ( .a(n33822), .b(n33819), .o(n33823) );
no02f01 g30033 ( .a(n33821), .b(n33818), .o(n33824) );
no02f01 g30034 ( .a(n33824), .b(n33823), .o(n33825) );
in01f01 g30035 ( .a(n33825), .o(n33826) );
no02f01 g30036 ( .a(n33826), .b(n33513), .o(n33827) );
no02f01 g30037 ( .a(n33827), .b(n33816), .o(n33828) );
in01f01 g30038 ( .a(n33828), .o(n33829) );
no02f01 g30039 ( .a(n33829), .b(n33806), .o(n33830) );
ao12f01 g30040 ( .a(n33512), .b(n33825), .c(n33814), .o(n33831) );
no02f01 g30041 ( .a(n33808), .b(n32878), .o(n33832) );
in01f01 g30042 ( .a(n33832), .o(n33833) );
ao12f01 g30043 ( .a(n33833), .b(n32852), .c(n32848), .o(n33834) );
no02f01 g30044 ( .a(n32744), .b(n32879), .o(n33835) );
no02f01 g30045 ( .a(n33835), .b(n32854), .o(n33836) );
no02f01 g30046 ( .a(n33836), .b(n33834), .o(n33837) );
na02f01 g30047 ( .a(n33836), .b(n33834), .o(n33838) );
in01f01 g30048 ( .a(n33838), .o(n33839) );
no02f01 g30049 ( .a(n33839), .b(n33837), .o(n33840) );
in01f01 g30050 ( .a(n33840), .o(n33841) );
no02f01 g30051 ( .a(n33841), .b(n33513), .o(n33842) );
no02f01 g30052 ( .a(n33840), .b(n33512), .o(n33843) );
no02f01 g30053 ( .a(n33843), .b(n33842), .o(n33844) );
in01f01 g30054 ( .a(n33844), .o(n33845) );
no03f01 g30055 ( .a(n33845), .b(n33831), .c(n33830), .o(n33846) );
no02f01 g30056 ( .a(n33831), .b(n33830), .o(n33847) );
no02f01 g30057 ( .a(n33844), .b(n33847), .o(n33848) );
no02f01 g30058 ( .a(n33848), .b(n33846), .o(n33849) );
in01f01 g30059 ( .a(n33849), .o(n33850) );
no02f01 g30060 ( .a(n33850), .b(n33508), .o(n33851) );
in01f01 g30061 ( .a(n33851), .o(n33852) );
in01f01 g30062 ( .a(n33830), .o(n33853) );
no02f01 g30063 ( .a(n33843), .b(n33831), .o(n33854) );
oa12f01 g30064 ( .a(n33854), .b(n33842), .c(n33853), .o(n33855) );
in01f01 g30065 ( .a(n33855), .o(n33856) );
no03f01 g30066 ( .a(n32854), .b(n32853), .c(n32849), .o(n33857) );
no02f01 g30067 ( .a(n33833), .b(n33835), .o(n33858) );
in01f01 g30068 ( .a(n33858), .o(n33859) );
no02f01 g30069 ( .a(n32744), .b(n32880), .o(n33860) );
no02f01 g30070 ( .a(n33860), .b(n32855), .o(n33861) );
in01f01 g30071 ( .a(n33861), .o(n33862) );
no03f01 g30072 ( .a(n33862), .b(n33859), .c(n33857), .o(n33863) );
no02f01 g30073 ( .a(n33859), .b(n33857), .o(n33864) );
no02f01 g30074 ( .a(n33861), .b(n33864), .o(n33865) );
no02f01 g30075 ( .a(n33865), .b(n33863), .o(n33866) );
in01f01 g30076 ( .a(n33866), .o(n33867) );
no02f01 g30077 ( .a(n33867), .b(n33513), .o(n33868) );
no02f01 g30078 ( .a(n33866), .b(n33512), .o(n33869) );
no02f01 g30079 ( .a(n33869), .b(n33868), .o(n33870) );
no02f01 g30080 ( .a(n33870), .b(n33856), .o(n33871) );
na02f01 g30081 ( .a(n33870), .b(n33856), .o(n33872) );
in01f01 g30082 ( .a(n33872), .o(n33873) );
no03f01 g30083 ( .a(n33873), .b(n33871), .c(n33508), .o(n33874) );
no02f01 g30084 ( .a(n33814), .b(n33512), .o(n33875) );
no02f01 g30085 ( .a(n33816), .b(n33806), .o(n33876) );
no02f01 g30086 ( .a(n33876), .b(n33875), .o(n33877) );
no02f01 g30087 ( .a(n33825), .b(n33512), .o(n33878) );
no02f01 g30088 ( .a(n33878), .b(n33827), .o(n33879) );
no02f01 g30089 ( .a(n33879), .b(n33877), .o(n33880) );
na02f01 g30090 ( .a(n33879), .b(n33877), .o(n33881) );
in01f01 g30091 ( .a(n33881), .o(n33882) );
no02f01 g30092 ( .a(n33882), .b(n33880), .o(n33883) );
in01f01 g30093 ( .a(n33883), .o(n33884) );
in01f01 g30094 ( .a(n33806), .o(n33885) );
no02f01 g30095 ( .a(n33875), .b(n33816), .o(n33886) );
in01f01 g30096 ( .a(n33886), .o(n33887) );
no02f01 g30097 ( .a(n33887), .b(n33885), .o(n33888) );
no02f01 g30098 ( .a(n33886), .b(n33806), .o(n33889) );
no02f01 g30099 ( .a(n33889), .b(n33888), .o(n33890) );
in01f01 g30100 ( .a(n33890), .o(n33891) );
ao12f01 g30101 ( .a(n33508), .b(n33891), .c(n33884), .o(n33892) );
no02f01 g30102 ( .a(n33892), .b(n33874), .o(n33893) );
na02f01 g30103 ( .a(n33893), .b(n33852), .o(n33894) );
no02f01 g30104 ( .a(n32912), .b(n32859), .o(n33895) );
in01f01 g30105 ( .a(n33895), .o(n33896) );
no03f01 g30106 ( .a(n33896), .b(n32910), .c(n32886), .o(n33897) );
no02f01 g30107 ( .a(n32910), .b(n32886), .o(n33898) );
no02f01 g30108 ( .a(n33895), .b(n33898), .o(n33899) );
no02f01 g30109 ( .a(n33899), .b(n33897), .o(n33900) );
in01f01 g30110 ( .a(n33900), .o(n33901) );
no02f01 g30111 ( .a(n33901), .b(n33513), .o(n33902) );
no02f01 g30112 ( .a(n33868), .b(n33842), .o(n33903) );
na02f01 g30113 ( .a(n33903), .b(n33828), .o(n33904) );
no04f01 g30114 ( .a(n33904), .b(n33796), .c(n33751), .d(n33708), .o(n33905) );
ao12f01 g30115 ( .a(n33512), .b(n33866), .c(n33840), .o(n33906) );
no02f01 g30116 ( .a(n33906), .b(n33831), .o(n33907) );
in01f01 g30117 ( .a(n33907), .o(n33908) );
no02f01 g30118 ( .a(n33908), .b(n33805), .o(n33909) );
in01f01 g30119 ( .a(n33909), .o(n33910) );
no02f01 g30120 ( .a(n33910), .b(n33905), .o(n33911) );
no02f01 g30121 ( .a(n33900), .b(n33512), .o(n33912) );
in01f01 g30122 ( .a(n33912), .o(n33913) );
ao12f01 g30123 ( .a(n33902), .b(n33913), .c(n33911), .o(n33914) );
in01f01 g30124 ( .a(n33914), .o(n33915) );
no02f01 g30125 ( .a(n33513), .b(n33027), .o(n33916) );
no02f01 g30126 ( .a(n33512), .b(n32918), .o(n33917) );
no02f01 g30127 ( .a(n33917), .b(n33916), .o(n33918) );
no02f01 g30128 ( .a(n33918), .b(n33915), .o(n33919) );
na02f01 g30129 ( .a(n33918), .b(n33915), .o(n33920) );
in01f01 g30130 ( .a(n33920), .o(n33921) );
no02f01 g30131 ( .a(n33921), .b(n33919), .o(n33922) );
in01f01 g30132 ( .a(n33922), .o(n33923) );
in01f01 g30133 ( .a(n33911), .o(n33924) );
no02f01 g30134 ( .a(n33912), .b(n33902), .o(n33925) );
in01f01 g30135 ( .a(n33925), .o(n33926) );
no02f01 g30136 ( .a(n33926), .b(n33924), .o(n33927) );
no02f01 g30137 ( .a(n33925), .b(n33911), .o(n33928) );
no02f01 g30138 ( .a(n33928), .b(n33927), .o(n33929) );
in01f01 g30139 ( .a(n33929), .o(n33930) );
ao12f01 g30140 ( .a(n33508), .b(n33930), .c(n33923), .o(n33931) );
ao12f01 g30141 ( .a(n33512), .b(n33900), .c(n32918), .o(n33932) );
no02f01 g30142 ( .a(n33916), .b(n33902), .o(n33933) );
in01f01 g30143 ( .a(n33933), .o(n33934) );
no02f01 g30144 ( .a(n33934), .b(n33911), .o(n33935) );
no02f01 g30145 ( .a(n33513), .b(n33029), .o(n33936) );
no02f01 g30146 ( .a(n33512), .b(n32925), .o(n33937) );
no02f01 g30147 ( .a(n33937), .b(n33936), .o(n33938) );
in01f01 g30148 ( .a(n33938), .o(n33939) );
no03f01 g30149 ( .a(n33939), .b(n33935), .c(n33932), .o(n33940) );
oa12f01 g30150 ( .a(n33939), .b(n33935), .c(n33932), .o(n33941) );
in01f01 g30151 ( .a(n33941), .o(n33942) );
no02f01 g30152 ( .a(n33942), .b(n33940), .o(n33943) );
in01f01 g30153 ( .a(n33943), .o(n33944) );
no02f01 g30154 ( .a(n33944), .b(n33508), .o(n33945) );
no03f01 g30155 ( .a(n33945), .b(n33931), .c(n33894), .o(n33946) );
no02f01 g30156 ( .a(n33773), .b(n33766), .o(n33947) );
no02f01 g30157 ( .a(n33801), .b(n33752), .o(n33948) );
in01f01 g30158 ( .a(n33948), .o(n33949) );
ao12f01 g30159 ( .a(n33802), .b(n33949), .c(n33947), .o(n33950) );
in01f01 g30160 ( .a(n33950), .o(n33951) );
no02f01 g30161 ( .a(n33782), .b(n33512), .o(n33952) );
no02f01 g30162 ( .a(n33952), .b(n33784), .o(n33953) );
in01f01 g30163 ( .a(n33953), .o(n33954) );
no02f01 g30164 ( .a(n33954), .b(n33951), .o(n33955) );
no02f01 g30165 ( .a(n33953), .b(n33950), .o(n33956) );
no02f01 g30166 ( .a(n33956), .b(n33955), .o(n33957) );
in01f01 g30167 ( .a(n33957), .o(n33958) );
no02f01 g30168 ( .a(n33958), .b(n33508), .o(n33959) );
in01f01 g30169 ( .a(n33952), .o(n33960) );
ao12f01 g30170 ( .a(n33784), .b(n33950), .c(n33960), .o(n33961) );
no02f01 g30171 ( .a(n33792), .b(n33512), .o(n33962) );
no02f01 g30172 ( .a(n33962), .b(n33794), .o(n33963) );
in01f01 g30173 ( .a(n33963), .o(n33964) );
no02f01 g30174 ( .a(n33964), .b(n33961), .o(n33965) );
na02f01 g30175 ( .a(n33964), .b(n33961), .o(n33966) );
in01f01 g30176 ( .a(n33966), .o(n33967) );
no03f01 g30177 ( .a(n33967), .b(n33965), .c(n33508), .o(n33968) );
no02f01 g30178 ( .a(n33771), .b(n33512), .o(n33969) );
no02f01 g30179 ( .a(n33969), .b(n33801), .o(n33970) );
oa12f01 g30180 ( .a(n33970), .b(n33773), .c(n33753), .o(n33971) );
in01f01 g30181 ( .a(n33971), .o(n33972) );
no02f01 g30182 ( .a(n33764), .b(n33512), .o(n33973) );
no02f01 g30183 ( .a(n33973), .b(n33766), .o(n33974) );
no02f01 g30184 ( .a(n33974), .b(n33972), .o(n33975) );
na02f01 g30185 ( .a(n33974), .b(n33972), .o(n33976) );
in01f01 g30186 ( .a(n33976), .o(n33977) );
no02f01 g30187 ( .a(n33977), .b(n33975), .o(n33978) );
in01f01 g30188 ( .a(n33978), .o(n33979) );
no02f01 g30189 ( .a(n33969), .b(n33773), .o(n33980) );
no02f01 g30190 ( .a(n33980), .b(n33948), .o(n33981) );
na02f01 g30191 ( .a(n33980), .b(n33948), .o(n33982) );
in01f01 g30192 ( .a(n33982), .o(n33983) );
no02f01 g30193 ( .a(n33983), .b(n33981), .o(n33984) );
in01f01 g30194 ( .a(n33984), .o(n33985) );
ao12f01 g30195 ( .a(n33508), .b(n33985), .c(n33979), .o(n33986) );
no03f01 g30196 ( .a(n33986), .b(n33968), .c(n33959), .o(n33987) );
in01f01 g30197 ( .a(n33632), .o(n33988) );
no02f01 g30198 ( .a(n33630), .b(n33512), .o(n33989) );
ao12f01 g30199 ( .a(n33989), .b(n33988), .c(n33610), .o(n33990) );
in01f01 g30200 ( .a(n33990), .o(n33991) );
no02f01 g30201 ( .a(n33623), .b(n33512), .o(n33992) );
no02f01 g30202 ( .a(n33992), .b(n33625), .o(n33993) );
in01f01 g30203 ( .a(n33993), .o(n33994) );
no02f01 g30204 ( .a(n33994), .b(n33991), .o(n33995) );
no02f01 g30205 ( .a(n33993), .b(n33990), .o(n33996) );
no02f01 g30206 ( .a(n33996), .b(n33995), .o(n33997) );
in01f01 g30207 ( .a(n33997), .o(n33998) );
in01f01 g30208 ( .a(n33610), .o(n33999) );
no02f01 g30209 ( .a(n33989), .b(n33632), .o(n34000) );
no02f01 g30210 ( .a(n34000), .b(n33999), .o(n34001) );
na02f01 g30211 ( .a(n34000), .b(n33999), .o(n34002) );
in01f01 g30212 ( .a(n34002), .o(n34003) );
no02f01 g30213 ( .a(n34003), .b(n34001), .o(n34004) );
in01f01 g30214 ( .a(n34004), .o(n34005) );
ao12f01 g30215 ( .a(n33508), .b(n34005), .c(n33998), .o(n34006) );
in01f01 g30216 ( .a(n33596), .o(n34007) );
no02f01 g30217 ( .a(n33593), .b(n33512), .o(n34008) );
no02f01 g30218 ( .a(n33608), .b(n34008), .o(n34009) );
oa12f01 g30219 ( .a(n34009), .b(n34007), .c(n33561), .o(n34010) );
no02f01 g30220 ( .a(n33602), .b(n33512), .o(n34011) );
no02f01 g30221 ( .a(n34011), .b(n33604), .o(n34012) );
in01f01 g30222 ( .a(n34012), .o(n34013) );
no02f01 g30223 ( .a(n34013), .b(n34010), .o(n34014) );
na02f01 g30224 ( .a(n34013), .b(n34010), .o(n34015) );
in01f01 g30225 ( .a(n34015), .o(n34016) );
no02f01 g30226 ( .a(n34016), .b(n34014), .o(n34017) );
in01f01 g30227 ( .a(n34017), .o(n34018) );
no02f01 g30228 ( .a(n34018), .b(n33508), .o(n34019) );
in01f01 g30229 ( .a(n33561), .o(n34020) );
in01f01 g30230 ( .a(n33585), .o(n34021) );
no02f01 g30231 ( .a(n33583), .b(n33512), .o(n34022) );
ao12f01 g30232 ( .a(n34022), .b(n34021), .c(n34020), .o(n34023) );
in01f01 g30233 ( .a(n34023), .o(n34024) );
no02f01 g30234 ( .a(n33576), .b(n33512), .o(n34025) );
no02f01 g30235 ( .a(n34025), .b(n33578), .o(n34026) );
in01f01 g30236 ( .a(n34026), .o(n34027) );
no02f01 g30237 ( .a(n34027), .b(n34024), .o(n34028) );
no02f01 g30238 ( .a(n34026), .b(n34023), .o(n34029) );
no02f01 g30239 ( .a(n34029), .b(n34028), .o(n34030) );
no02f01 g30240 ( .a(n34022), .b(n33585), .o(n34031) );
no02f01 g30241 ( .a(n34031), .b(n33561), .o(n34032) );
na02f01 g30242 ( .a(n34031), .b(n33561), .o(n34033) );
in01f01 g30243 ( .a(n34033), .o(n34034) );
no02f01 g30244 ( .a(n34034), .b(n34032), .o(n34035) );
ao12f01 g30245 ( .a(n33507), .b(n34035), .c(n34030), .o(n34036) );
no03f01 g30246 ( .a(n33506), .b(n33493), .c(n33491), .o(n34037) );
in01f01 g30247 ( .a(n34037), .o(n34038) );
oa12f01 g30248 ( .a(n33493), .b(n33506), .c(n33491), .o(n34039) );
in01f01 g30249 ( .a(n33549), .o(n34040) );
no03f01 g30250 ( .a(n33551), .b(n34040), .c(n33544), .o(n34041) );
no02f01 g30251 ( .a(n33551), .b(n33544), .o(n34042) );
no02f01 g30252 ( .a(n34042), .b(n33549), .o(n34043) );
no02f01 g30253 ( .a(n34043), .b(n34041), .o(n34044) );
in01f01 g30254 ( .a(n34044), .o(n34045) );
ao12f01 g30255 ( .a(n34045), .b(n34039), .c(n34038), .o(n34046) );
in01f01 g30256 ( .a(n33506), .o(n34047) );
no02f01 g30257 ( .a(n34047), .b(delay_sub_ln23_0_unr29_stage10_stallmux_q), .o(n34048) );
no02f01 g30258 ( .a(n34047), .b(n33491), .o(n34049) );
in01f01 g30259 ( .a(n33548), .o(n34050) );
no02f01 g30260 ( .a(n34050), .b(n33464), .o(n34051) );
no02f01 g30261 ( .a(n33548), .b(n33451), .o(n34052) );
no02f01 g30262 ( .a(n34052), .b(n34051), .o(n34053) );
no03f01 g30263 ( .a(n34053), .b(n34049), .c(n34048), .o(n34054) );
na03f01 g30264 ( .a(n34045), .b(n34039), .c(n34038), .o(n34055) );
oa12f01 g30265 ( .a(n34055), .b(n34054), .c(n34046), .o(n34056) );
no02f01 g30266 ( .a(n33555), .b(n33537), .o(n34057) );
in01f01 g30267 ( .a(n34057), .o(n34058) );
no02f01 g30268 ( .a(n34058), .b(n33553), .o(n34059) );
na02f01 g30269 ( .a(n34058), .b(n33553), .o(n34060) );
in01f01 g30270 ( .a(n34060), .o(n34061) );
no02f01 g30271 ( .a(n34061), .b(n34059), .o(n34062) );
na02f01 g30272 ( .a(n34062), .b(n33507), .o(n34063) );
na02f01 g30273 ( .a(n34063), .b(n34056), .o(n34064) );
in01f01 g30274 ( .a(n33557), .o(n34065) );
no02f01 g30275 ( .a(n33558), .b(n33527), .o(n34066) );
in01f01 g30276 ( .a(n34066), .o(n34067) );
no02f01 g30277 ( .a(n34067), .b(n34065), .o(n34068) );
no02f01 g30278 ( .a(n34066), .b(n33557), .o(n34069) );
no02f01 g30279 ( .a(n34069), .b(n34068), .o(n34070) );
no02f01 g30280 ( .a(n34070), .b(n34064), .o(n34071) );
in01f01 g30281 ( .a(n34070), .o(n34072) );
no02f01 g30282 ( .a(n34062), .b(n33507), .o(n34073) );
no02f01 g30283 ( .a(n34073), .b(n34072), .o(n34074) );
in01f01 g30284 ( .a(n34074), .o(n34075) );
ao12f01 g30285 ( .a(n34075), .b(n34063), .c(n34056), .o(n34076) );
no02f01 g30286 ( .a(n34076), .b(n33507), .o(n34077) );
no02f01 g30287 ( .a(n34077), .b(n34071), .o(n34078) );
in01f01 g30288 ( .a(n34035), .o(n34079) );
no02f01 g30289 ( .a(n34079), .b(n33508), .o(n34080) );
in01f01 g30290 ( .a(n34030), .o(n34081) );
no02f01 g30291 ( .a(n34081), .b(n33508), .o(n34082) );
no02f01 g30292 ( .a(n33585), .b(n33578), .o(n34083) );
ao12f01 g30293 ( .a(n33608), .b(n34083), .c(n34020), .o(n34084) );
no02f01 g30294 ( .a(n34008), .b(n33595), .o(n34085) );
no02f01 g30295 ( .a(n34085), .b(n34084), .o(n34086) );
na02f01 g30296 ( .a(n34085), .b(n34084), .o(n34087) );
in01f01 g30297 ( .a(n34087), .o(n34088) );
no02f01 g30298 ( .a(n34088), .b(n34086), .o(n34089) );
in01f01 g30299 ( .a(n34089), .o(n34090) );
no02f01 g30300 ( .a(n34090), .b(n33508), .o(n34091) );
no04f01 g30301 ( .a(n34091), .b(n34082), .c(n34080), .d(n34078), .o(n34092) );
ao12f01 g30302 ( .a(n33507), .b(n34089), .c(n34017), .o(n34093) );
no03f01 g30303 ( .a(n34093), .b(n34092), .c(n34036), .o(n34094) );
ao12f01 g30304 ( .a(n33657), .b(n33633), .c(n33610), .o(n34095) );
no02f01 g30305 ( .a(n33652), .b(n33512), .o(n34096) );
no02f01 g30306 ( .a(n34096), .b(n33654), .o(n34097) );
no02f01 g30307 ( .a(n34097), .b(n34095), .o(n34098) );
na02f01 g30308 ( .a(n34097), .b(n34095), .o(n34099) );
in01f01 g30309 ( .a(n34099), .o(n34100) );
no02f01 g30310 ( .a(n34100), .b(n34098), .o(n34101) );
in01f01 g30311 ( .a(n34101), .o(n34102) );
no02f01 g30312 ( .a(n34102), .b(n33508), .o(n34103) );
no04f01 g30313 ( .a(n34103), .b(n34094), .c(n34019), .d(n34006), .o(n34104) );
no03f01 g30314 ( .a(n33654), .b(n33634), .c(n33999), .o(n34105) );
no03f01 g30315 ( .a(n34105), .b(n34096), .c(n33657), .o(n34106) );
no02f01 g30316 ( .a(n33643), .b(n33512), .o(n34107) );
no02f01 g30317 ( .a(n34107), .b(n33645), .o(n34108) );
no02f01 g30318 ( .a(n34108), .b(n34106), .o(n34109) );
na02f01 g30319 ( .a(n34108), .b(n34106), .o(n34110) );
in01f01 g30320 ( .a(n34110), .o(n34111) );
no02f01 g30321 ( .a(n34111), .b(n34109), .o(n34112) );
in01f01 g30322 ( .a(n34112), .o(n34113) );
no02f01 g30323 ( .a(n34113), .b(n33508), .o(n34114) );
in01f01 g30324 ( .a(n34114), .o(n34115) );
ao12f01 g30325 ( .a(n33704), .b(n33682), .c(n33660), .o(n34116) );
no02f01 g30326 ( .a(n33699), .b(n33512), .o(n34117) );
no02f01 g30327 ( .a(n34117), .b(n33701), .o(n34118) );
no02f01 g30328 ( .a(n34118), .b(n34116), .o(n34119) );
na02f01 g30329 ( .a(n34118), .b(n34116), .o(n34120) );
in01f01 g30330 ( .a(n34120), .o(n34121) );
no02f01 g30331 ( .a(n34121), .b(n34119), .o(n34122) );
in01f01 g30332 ( .a(n34122), .o(n34123) );
no02f01 g30333 ( .a(n34123), .b(n33508), .o(n34124) );
in01f01 g30334 ( .a(n33659), .o(n34125) );
no02f01 g30335 ( .a(n33679), .b(n33512), .o(n34126) );
no02f01 g30336 ( .a(n33681), .b(n33656), .o(n34127) );
no03f01 g30337 ( .a(n34127), .b(n34126), .c(n34125), .o(n34128) );
no02f01 g30338 ( .a(n33670), .b(n33512), .o(n34129) );
no02f01 g30339 ( .a(n34129), .b(n33672), .o(n34130) );
no02f01 g30340 ( .a(n34130), .b(n34128), .o(n34131) );
na02f01 g30341 ( .a(n34130), .b(n34128), .o(n34132) );
in01f01 g30342 ( .a(n34132), .o(n34133) );
no02f01 g30343 ( .a(n34133), .b(n34131), .o(n34134) );
in01f01 g30344 ( .a(n33660), .o(n34135) );
no02f01 g30345 ( .a(n34126), .b(n33681), .o(n34136) );
no02f01 g30346 ( .a(n34136), .b(n34135), .o(n34137) );
na02f01 g30347 ( .a(n34136), .b(n34135), .o(n34138) );
in01f01 g30348 ( .a(n34138), .o(n34139) );
no02f01 g30349 ( .a(n34139), .b(n34137), .o(n34140) );
no02f01 g30350 ( .a(n34140), .b(n34134), .o(n34141) );
no02f01 g30351 ( .a(n34141), .b(n33508), .o(n34142) );
in01f01 g30352 ( .a(n34117), .o(n34143) );
ao12f01 g30353 ( .a(n33701), .b(n34116), .c(n34143), .o(n34144) );
in01f01 g30354 ( .a(n34144), .o(n34145) );
no02f01 g30355 ( .a(n33691), .b(n33512), .o(n34146) );
no02f01 g30356 ( .a(n34146), .b(n33693), .o(n34147) );
no02f01 g30357 ( .a(n34147), .b(n34145), .o(n34148) );
na02f01 g30358 ( .a(n34147), .b(n34145), .o(n34149) );
in01f01 g30359 ( .a(n34149), .o(n34150) );
no02f01 g30360 ( .a(n34150), .b(n34148), .o(n34151) );
in01f01 g30361 ( .a(n34151), .o(n34152) );
no02f01 g30362 ( .a(n34152), .b(n33508), .o(n34153) );
no03f01 g30363 ( .a(n34153), .b(n34142), .c(n34124), .o(n34154) );
na03f01 g30364 ( .a(n34154), .b(n34115), .c(n34104), .o(n34155) );
ao12f01 g30365 ( .a(n33507), .b(n34112), .c(n34101), .o(n34156) );
ao12f01 g30366 ( .a(n33507), .b(n34004), .c(n33997), .o(n34157) );
no02f01 g30367 ( .a(n34157), .b(n34156), .o(n34158) );
in01f01 g30368 ( .a(n34158), .o(n34159) );
ao12f01 g30369 ( .a(n33507), .b(n34140), .c(n34134), .o(n34160) );
ao12f01 g30370 ( .a(n33507), .b(n34151), .c(n34122), .o(n34161) );
no03f01 g30371 ( .a(n34161), .b(n34160), .c(n34159), .o(n34162) );
na02f01 g30372 ( .a(n34162), .b(n34155), .o(n34163) );
in01f01 g30373 ( .a(n33729), .o(n34164) );
ao12f01 g30374 ( .a(n33798), .b(n34164), .c(n33707), .o(n34165) );
no02f01 g30375 ( .a(n33747), .b(n33512), .o(n34166) );
no02f01 g30376 ( .a(n34166), .b(n33749), .o(n34167) );
no02f01 g30377 ( .a(n34167), .b(n34165), .o(n34168) );
na02f01 g30378 ( .a(n34167), .b(n34165), .o(n34169) );
in01f01 g30379 ( .a(n34169), .o(n34170) );
no02f01 g30380 ( .a(n34170), .b(n34168), .o(n34171) );
in01f01 g30381 ( .a(n34171), .o(n34172) );
no02f01 g30382 ( .a(n34172), .b(n33508), .o(n34173) );
no03f01 g30383 ( .a(n33749), .b(n33729), .c(n33708), .o(n34174) );
no02f01 g30384 ( .a(n34166), .b(n33798), .o(n34175) );
in01f01 g30385 ( .a(n34175), .o(n34176) );
no02f01 g30386 ( .a(n33738), .b(n33512), .o(n34177) );
no02f01 g30387 ( .a(n34177), .b(n33740), .o(n34178) );
in01f01 g30388 ( .a(n34178), .o(n34179) );
no03f01 g30389 ( .a(n34179), .b(n34176), .c(n34174), .o(n34180) );
no02f01 g30390 ( .a(n34176), .b(n34174), .o(n34181) );
no02f01 g30391 ( .a(n34178), .b(n34181), .o(n34182) );
no02f01 g30392 ( .a(n34182), .b(n34180), .o(n34183) );
in01f01 g30393 ( .a(n34183), .o(n34184) );
no02f01 g30394 ( .a(n34184), .b(n33508), .o(n34185) );
no02f01 g30395 ( .a(n33727), .b(n33512), .o(n34186) );
no02f01 g30396 ( .a(n33728), .b(n33513), .o(n34187) );
in01f01 g30397 ( .a(n34187), .o(n34188) );
ao12f01 g30398 ( .a(n34186), .b(n34188), .c(n33707), .o(n34189) );
in01f01 g30399 ( .a(n34189), .o(n34190) );
no02f01 g30400 ( .a(n33722), .b(n33513), .o(n34191) );
no02f01 g30401 ( .a(n33721), .b(n33512), .o(n34192) );
no02f01 g30402 ( .a(n34192), .b(n34191), .o(n34193) );
in01f01 g30403 ( .a(n34193), .o(n34194) );
no02f01 g30404 ( .a(n34194), .b(n34190), .o(n34195) );
no02f01 g30405 ( .a(n34193), .b(n34189), .o(n34196) );
no02f01 g30406 ( .a(n34196), .b(n34195), .o(n34197) );
no02f01 g30407 ( .a(n34187), .b(n34186), .o(n34198) );
no02f01 g30408 ( .a(n34198), .b(n33708), .o(n34199) );
na02f01 g30409 ( .a(n34198), .b(n33708), .o(n34200) );
in01f01 g30410 ( .a(n34200), .o(n34201) );
no02f01 g30411 ( .a(n34201), .b(n34199), .o(n34202) );
no02f01 g30412 ( .a(n34202), .b(n34197), .o(n34203) );
no02f01 g30413 ( .a(n34203), .b(n33508), .o(n34204) );
no03f01 g30414 ( .a(n34204), .b(n34185), .c(n34173), .o(n34205) );
na04f01 g30415 ( .a(n34205), .b(n34163), .c(n33987), .d(n33946), .o(n34206) );
in01f01 g30416 ( .a(n33946), .o(n34207) );
in01f01 g30417 ( .a(n33987), .o(n34208) );
ao12f01 g30418 ( .a(n33507), .b(n34202), .c(n34197), .o(n34209) );
ao12f01 g30419 ( .a(n33507), .b(n34183), .c(n34171), .o(n34210) );
no02f01 g30420 ( .a(n34210), .b(n34209), .o(n34211) );
ao12f01 g30421 ( .a(n33507), .b(n33984), .c(n33978), .o(n34212) );
no02f01 g30422 ( .a(n33967), .b(n33965), .o(n34213) );
ao12f01 g30423 ( .a(n33507), .b(n34213), .c(n33957), .o(n34214) );
no02f01 g30424 ( .a(n34214), .b(n34212), .o(n34215) );
oa12f01 g30425 ( .a(n34215), .b(n34211), .c(n34208), .o(n34216) );
in01f01 g30426 ( .a(n34216), .o(n34217) );
ao12f01 g30427 ( .a(n33507), .b(n33890), .c(n33883), .o(n34218) );
no02f01 g30428 ( .a(n33873), .b(n33871), .o(n34219) );
no02f01 g30429 ( .a(n33849), .b(n33507), .o(n34220) );
in01f01 g30430 ( .a(n34220), .o(n34221) );
ao12f01 g30431 ( .a(n33507), .b(n34221), .c(n34219), .o(n34222) );
ao12f01 g30432 ( .a(n33507), .b(n33929), .c(n33922), .o(n34223) );
in01f01 g30433 ( .a(n34223), .o(n34224) );
ao12f01 g30434 ( .a(n33507), .b(n34224), .c(n33943), .o(n34225) );
no03f01 g30435 ( .a(n34225), .b(n34222), .c(n34218), .o(n34226) );
oa12f01 g30436 ( .a(n34226), .b(n34217), .c(n34207), .o(n34227) );
in01f01 g30437 ( .a(n34227), .o(n34228) );
no03f01 g30438 ( .a(n33936), .b(n33934), .c(n33904), .o(n34229) );
in01f01 g30439 ( .a(n34229), .o(n34230) );
no02f01 g30440 ( .a(n34230), .b(n33806), .o(n34231) );
no02f01 g30441 ( .a(n33932), .b(n33029), .o(n34232) );
oa12f01 g30442 ( .a(n33907), .b(n34232), .c(n33512), .o(n34233) );
no02f01 g30443 ( .a(n33513), .b(n33011), .o(n34234) );
no02f01 g30444 ( .a(n33512), .b(n32902), .o(n34235) );
no02f01 g30445 ( .a(n34235), .b(n34234), .o(n34236) );
in01f01 g30446 ( .a(n34236), .o(n34237) );
no03f01 g30447 ( .a(n34237), .b(n34233), .c(n34231), .o(n34238) );
oa12f01 g30448 ( .a(n34237), .b(n34233), .c(n34231), .o(n34239) );
in01f01 g30449 ( .a(n34239), .o(n34240) );
no02f01 g30450 ( .a(n34240), .b(n34238), .o(n34241) );
no02f01 g30451 ( .a(n34241), .b(n33507), .o(n34242) );
in01f01 g30452 ( .a(n34238), .o(n34243) );
na02f01 g30453 ( .a(n34239), .b(n34243), .o(n34244) );
no02f01 g30454 ( .a(n34244), .b(n33508), .o(n34245) );
no02f01 g30455 ( .a(n34245), .b(n34242), .o(n34246) );
na03f01 g30456 ( .a(n34246), .b(n34228), .c(n34206), .o(n34247) );
in01f01 g30457 ( .a(n34006), .o(n34248) );
in01f01 g30458 ( .a(n34019), .o(n34249) );
in01f01 g30459 ( .a(n34036), .o(n34250) );
oa22f01 g30460 ( .a(n34076), .b(n33507), .c(n34070), .d(n34064), .o(n34251) );
in01f01 g30461 ( .a(n34080), .o(n34252) );
in01f01 g30462 ( .a(n34082), .o(n34253) );
in01f01 g30463 ( .a(n34091), .o(n34254) );
na04f01 g30464 ( .a(n34254), .b(n34253), .c(n34252), .d(n34251), .o(n34255) );
in01f01 g30465 ( .a(n34093), .o(n34256) );
na03f01 g30466 ( .a(n34256), .b(n34255), .c(n34250), .o(n34257) );
in01f01 g30467 ( .a(n34103), .o(n34258) );
na04f01 g30468 ( .a(n34258), .b(n34257), .c(n34249), .d(n34248), .o(n34259) );
no02f01 g30469 ( .a(n34114), .b(n34259), .o(n34260) );
in01f01 g30470 ( .a(n34162), .o(n34261) );
ao12f01 g30471 ( .a(n34261), .b(n34154), .c(n34260), .o(n34262) );
in01f01 g30472 ( .a(n34205), .o(n34263) );
no04f01 g30473 ( .a(n34263), .b(n34262), .c(n34208), .d(n34207), .o(n34264) );
in01f01 g30474 ( .a(n34246), .o(n34265) );
oa12f01 g30475 ( .a(n34265), .b(n34227), .c(n34264), .o(n34266) );
ao12f01 g30476 ( .a(delay_sub_ln23_0_unr30_stage10_stallmux_q), .b(n34266), .c(n34247), .o(n34267) );
na03f01 g30477 ( .a(n34241), .b(n33944), .c(delay_sub_ln23_0_unr29_stage10_stallmux_q), .o(n34268) );
oa12f01 g30478 ( .a(n34244), .b(n33943), .c(n33491), .o(n34269) );
in01f01 g30479 ( .a(n33045), .o(n34270) );
no03f01 g30480 ( .a(n34270), .b(n33043), .c(n33039), .o(n34271) );
no02f01 g30481 ( .a(n34270), .b(n33039), .o(n34272) );
no02f01 g30482 ( .a(n34272), .b(n33044), .o(n34273) );
no02f01 g30483 ( .a(n34273), .b(n34271), .o(n34274) );
na03f01 g30484 ( .a(n34274), .b(n34269), .c(n34268), .o(n34275) );
no02f01 g30485 ( .a(n33944), .b(delay_sub_ln23_0_unr29_stage10_stallmux_q), .o(n34276) );
no02f01 g30486 ( .a(n33944), .b(n33491), .o(n34277) );
no02f01 g30487 ( .a(n33042), .b(n33027), .o(n34278) );
na02f01 g30488 ( .a(n33042), .b(n33027), .o(n34279) );
in01f01 g30489 ( .a(n34279), .o(n34280) );
no02f01 g30490 ( .a(n34280), .b(n34278), .o(n34281) );
no03f01 g30491 ( .a(n34281), .b(n34277), .c(n34276), .o(n34282) );
ao12f01 g30492 ( .a(n34274), .b(n34269), .c(n34268), .o(n34283) );
ao12f01 g30493 ( .a(n34283), .b(n34282), .c(n34275), .o(n34284) );
no02f01 g30494 ( .a(n34241), .b(delay_sub_ln23_0_unr29_stage10_stallmux_q), .o(n34285) );
no02f01 g30495 ( .a(n34244), .b(n33491), .o(n34286) );
oa22f01 g30496 ( .a(n34286), .b(n34285), .c(n33944), .d(n33491), .o(n34287) );
no02f01 g30497 ( .a(n33024), .b(n33022), .o(n34288) );
in01f01 g30498 ( .a(n34288), .o(n34289) );
no02f01 g30499 ( .a(n34289), .b(n33046), .o(n34290) );
na02f01 g30500 ( .a(n34289), .b(n33046), .o(n34291) );
in01f01 g30501 ( .a(n34291), .o(n34292) );
no02f01 g30502 ( .a(n34292), .b(n34290), .o(n34293) );
na02f01 g30503 ( .a(n34293), .b(n34287), .o(n34294) );
in01f01 g30504 ( .a(n34294), .o(n34295) );
no02f01 g30505 ( .a(n34293), .b(n34287), .o(n34296) );
no02f01 g30506 ( .a(n34296), .b(n34295), .o(n34297) );
no02f01 g30507 ( .a(n34297), .b(n34284), .o(n34298) );
na02f01 g30508 ( .a(n34297), .b(n34284), .o(n34299) );
in01f01 g30509 ( .a(n34299), .o(n34300) );
no02f01 g30510 ( .a(n34300), .b(n34298), .o(n34301) );
in01f01 g30511 ( .a(n34301), .o(n34302) );
no02f01 g30512 ( .a(n34302), .b(n34267), .o(n34303) );
in01f01 g30513 ( .a(delay_sub_ln23_0_unr30_stage10_stallmux_q), .o(n34304) );
no03f01 g30514 ( .a(n34265), .b(n34227), .c(n34264), .o(n34305) );
ao12f01 g30515 ( .a(n34246), .b(n34228), .c(n34206), .o(n34306) );
oa12f01 g30516 ( .a(n34304), .b(n34306), .c(n34305), .o(n34307) );
no03f01 g30517 ( .a(n34244), .b(n33943), .c(n33491), .o(n34308) );
in01f01 g30518 ( .a(n34269), .o(n34309) );
in01f01 g30519 ( .a(n34274), .o(n34310) );
no03f01 g30520 ( .a(n34310), .b(n34309), .c(n34308), .o(n34311) );
no03f01 g30521 ( .a(n34283), .b(n34282), .c(n34311), .o(n34312) );
in01f01 g30522 ( .a(n34282), .o(n34313) );
oa12f01 g30523 ( .a(n34310), .b(n34309), .c(n34308), .o(n34314) );
ao12f01 g30524 ( .a(n34313), .b(n34314), .c(n34275), .o(n34315) );
no02f01 g30525 ( .a(n34315), .b(n34312), .o(n34316) );
no02f01 g30526 ( .a(n34316), .b(n34307), .o(n34317) );
no03f01 g30527 ( .a(n34306), .b(n34305), .c(delay_sub_ln23_0_unr30_stage10_stallmux_q), .o(n34318) );
no03f01 g30528 ( .a(n34306), .b(n34305), .c(n34304), .o(n34319) );
no02f01 g30529 ( .a(n34277), .b(n34276), .o(n34320) );
no02f01 g30530 ( .a(n34281), .b(n34320), .o(n34321) );
na02f01 g30531 ( .a(n34281), .b(n34320), .o(n34322) );
in01f01 g30532 ( .a(n34322), .o(n34323) );
no02f01 g30533 ( .a(n34323), .b(n34321), .o(n34324) );
no03f01 g30534 ( .a(n34324), .b(n34319), .c(n34318), .o(n34325) );
na02f01 g30535 ( .a(n34316), .b(n34307), .o(n34326) );
ao12f01 g30536 ( .a(n34317), .b(n34326), .c(n34325), .o(n34327) );
no02f01 g30537 ( .a(n34327), .b(n34303), .o(n34328) );
no02f01 g30538 ( .a(n34295), .b(n34284), .o(n34329) );
no02f01 g30539 ( .a(n33049), .b(n33009), .o(n34330) );
no02f01 g30540 ( .a(n34330), .b(n33047), .o(n34331) );
na02f01 g30541 ( .a(n34330), .b(n33047), .o(n34332) );
in01f01 g30542 ( .a(n34332), .o(n34333) );
no02f01 g30543 ( .a(n34333), .b(n34331), .o(n34334) );
no02f01 g30544 ( .a(n34334), .b(n34287), .o(n34335) );
in01f01 g30545 ( .a(n34287), .o(n34336) );
in01f01 g30546 ( .a(n34334), .o(n34337) );
no02f01 g30547 ( .a(n34337), .b(n34336), .o(n34338) );
no04f01 g30548 ( .a(n34338), .b(n34335), .c(n34329), .d(n34296), .o(n34339) );
no02f01 g30549 ( .a(n34329), .b(n34296), .o(n34340) );
no02f01 g30550 ( .a(n34338), .b(n34335), .o(n34341) );
no02f01 g30551 ( .a(n34341), .b(n34340), .o(n34342) );
no02f01 g30552 ( .a(n34342), .b(n34339), .o(n34343) );
in01f01 g30553 ( .a(n34343), .o(n34344) );
no02f01 g30554 ( .a(n34301), .b(n34307), .o(n34345) );
no02f01 g30555 ( .a(n34345), .b(n34344), .o(n34346) );
oa12f01 g30556 ( .a(n34346), .b(n34327), .c(n34303), .o(n34347) );
ao22f01 g30557 ( .a(n34347), .b(n34267), .c(n34344), .d(n34328), .o(n34348) );
oa12f01 g30558 ( .a(n34334), .b(n34293), .c(n34287), .o(n34349) );
in01f01 g30559 ( .a(n34349), .o(n34350) );
oa12f01 g30560 ( .a(n34350), .b(n34295), .c(n34284), .o(n34351) );
ao22f01 g30561 ( .a(n34351), .b(n34336), .c(n34337), .d(n34329), .o(n34352) );
no02f01 g30562 ( .a(n33071), .b(n33048), .o(n34353) );
no02f01 g30563 ( .a(n33072), .b(n32928), .o(n34354) );
no02f01 g30564 ( .a(n34354), .b(n34353), .o(n34355) );
in01f01 g30565 ( .a(n34355), .o(n34356) );
ao12f01 g30566 ( .a(n34356), .b(n33051), .c(n33010), .o(n34357) );
no02f01 g30567 ( .a(n34355), .b(n33052), .o(n34358) );
no02f01 g30568 ( .a(n34358), .b(n34357), .o(n34359) );
no02f01 g30569 ( .a(n34359), .b(n34287), .o(n34360) );
in01f01 g30570 ( .a(n34359), .o(n34361) );
no02f01 g30571 ( .a(n34361), .b(n34336), .o(n34362) );
no02f01 g30572 ( .a(n34362), .b(n34360), .o(n34363) );
no02f01 g30573 ( .a(n34363), .b(n34352), .o(n34364) );
na02f01 g30574 ( .a(n34363), .b(n34352), .o(n34365) );
in01f01 g30575 ( .a(n34365), .o(n34366) );
no02f01 g30576 ( .a(n34366), .b(n34364), .o(n34367) );
in01f01 g30577 ( .a(n34367), .o(n34368) );
no02f01 g30578 ( .a(n34368), .b(n34267), .o(n34369) );
no02f01 g30579 ( .a(n34369), .b(n34348), .o(n34370) );
no02f01 g30580 ( .a(n34367), .b(n34307), .o(n34371) );
no02f01 g30581 ( .a(n34362), .b(n34352), .o(n34372) );
no02f01 g30582 ( .a(n34372), .b(n34360), .o(n34373) );
no02f01 g30583 ( .a(n34354), .b(n33052), .o(n34374) );
no02f01 g30584 ( .a(n34374), .b(n34353), .o(n34375) );
no02f01 g30585 ( .a(n33065), .b(n32928), .o(n34376) );
no02f01 g30586 ( .a(n33064), .b(n33048), .o(n34377) );
no02f01 g30587 ( .a(n34377), .b(n34376), .o(n34378) );
no02f01 g30588 ( .a(n34378), .b(n34375), .o(n34379) );
na02f01 g30589 ( .a(n34378), .b(n34375), .o(n34380) );
in01f01 g30590 ( .a(n34380), .o(n34381) );
no02f01 g30591 ( .a(n34381), .b(n34379), .o(n34382) );
na02f01 g30592 ( .a(n34382), .b(n34287), .o(n34383) );
in01f01 g30593 ( .a(n34383), .o(n34384) );
no02f01 g30594 ( .a(n34382), .b(n34287), .o(n34385) );
no02f01 g30595 ( .a(n34385), .b(n34384), .o(n34386) );
no02f01 g30596 ( .a(n34386), .b(n34373), .o(n34387) );
na02f01 g30597 ( .a(n34386), .b(n34373), .o(n34388) );
in01f01 g30598 ( .a(n34388), .o(n34389) );
no02f01 g30599 ( .a(n34389), .b(n34387), .o(n34390) );
no02f01 g30600 ( .a(n34390), .b(n34307), .o(n34391) );
in01f01 g30601 ( .a(n34390), .o(n34392) );
no02f01 g30602 ( .a(n34392), .b(n34267), .o(n34393) );
no02f01 g30603 ( .a(n34393), .b(n34391), .o(n34394) );
in01f01 g30604 ( .a(n34394), .o(n34395) );
no03f01 g30605 ( .a(n34395), .b(n34371), .c(n34370), .o(n34396) );
no02f01 g30606 ( .a(n34371), .b(n34370), .o(n34397) );
no02f01 g30607 ( .a(n34394), .b(n34397), .o(n34398) );
oa12f01 g30608 ( .a(n32734), .b(n34398), .c(n34396), .o(n34399) );
na02f01 g30609 ( .a(n34399), .b(n32733), .o(n418) );
no03f01 g30610 ( .a(n32505), .b(n32499), .c(n8756), .o(n34401) );
no02f01 g30611 ( .a(n8706), .b(n5973), .o(n34402) );
no02f01 g30612 ( .a(n34402), .b(n8708), .o(n34403) );
oa12f01 g30613 ( .a(n34403), .b(n34401), .c(n8713), .o(n34404) );
no02f01 g30614 ( .a(n34401), .b(n8713), .o(n34405) );
in01f01 g30615 ( .a(n34403), .o(n34406) );
na02f01 g30616 ( .a(n34406), .b(n34405), .o(n34407) );
na02f01 g30617 ( .a(n34407), .b(n34404), .o(n422) );
no02f01 g30618 ( .a(n9646), .b(n9645), .o(n1526) );
in01f01 g30619 ( .a(n1526), .o(n427) );
in01f01 g30620 ( .a(n6050), .o(n34411) );
no02f01 g30621 ( .a(n5889), .b(n5873), .o(n34412) );
na02f01 g30622 ( .a(n5889), .b(n5873), .o(n34413) );
in01f01 g30623 ( .a(n34413), .o(n34414) );
no02f01 g30624 ( .a(n34414), .b(n34412), .o(n34415) );
na02f01 g30625 ( .a(n34415), .b(n34411), .o(n34416) );
in01f01 g30626 ( .a(n34415), .o(n34417) );
na02f01 g30627 ( .a(n34417), .b(n6050), .o(n34418) );
na02f01 g30628 ( .a(n34418), .b(n34416), .o(n432) );
in01f01 g30629 ( .a(n_27923), .o(n34420) );
no02f01 g30630 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_30_), .b(n34420), .o(n34421) );
ao12f01 g30631 ( .a(n34420), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_13_), .c(delay_sub_ln23_0_unr20_stage7_stallmux_q_12_), .o(n34422) );
no02f01 g30632 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_11_), .b(n34420), .o(n34423) );
no02f01 g30633 ( .a(n34420), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_10_), .o(n34424) );
no02f01 g30634 ( .a(n34424), .b(n34423), .o(n34425) );
no02f01 g30635 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_9_), .b(n34420), .o(n34426) );
in01f01 g30636 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_8_), .o(n34427) );
no02f01 g30637 ( .a(n34427), .b(delay_sub_ln23_unr21_stage7_stallmux_q_1_), .o(n34428) );
in01f01 g30638 ( .a(n34428), .o(n34429) );
na02f01 g30639 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_9_), .b(n34420), .o(n34430) );
ao12f01 g30640 ( .a(n34426), .b(n34430), .c(n34429), .o(n34431) );
in01f01 g30641 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_10_), .o(n34432) );
in01f01 g30642 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_11_), .o(n34433) );
ao12f01 g30643 ( .a(n_27923), .b(n34433), .c(n34432), .o(n34434) );
oa12f01 g30644 ( .a(n34425), .b(n34434), .c(n34431), .o(n34435) );
in01f01 g30645 ( .a(n34435), .o(n34436) );
in01f01 g30646 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_3_), .o(n34437) );
in01f01 g30647 ( .a(n_186), .o(n34438) );
in01f01 g30648 ( .a(delay_sub_ln23_unr21_stage7_stallmux_q_1_), .o(n34439) );
na02f01 g30649 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_1_), .b(n34439), .o(n34440) );
no02f01 g30650 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_1_), .b(n34439), .o(n34441) );
oa12f01 g30651 ( .a(n34440), .b(n34441), .c(n34438), .o(n34442) );
no02f01 g30652 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_2_), .b(n34439), .o(n34443) );
in01f01 g30653 ( .a(n34443), .o(n34444) );
na02f01 g30654 ( .a(n34444), .b(n34442), .o(n34445) );
in01f01 g30655 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_2_), .o(n34446) );
no02f01 g30656 ( .a(n34446), .b(delay_sub_ln23_unr21_stage7_stallmux_q_1_), .o(n34447) );
in01f01 g30657 ( .a(n34447), .o(n34448) );
na02f01 g30658 ( .a(n34445), .b(n34448), .o(n34449) );
no02f01 g30659 ( .a(n34449), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_3_), .o(n34450) );
oa22f01 g30660 ( .a(n34450), .b(delay_sub_ln23_unr21_stage7_stallmux_q_1_), .c(n34445), .d(n34437), .o(n34451) );
no02f01 g30661 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_4_), .b(n34439), .o(n34452) );
in01f01 g30662 ( .a(n34452), .o(n34453) );
na02f01 g30663 ( .a(n34453), .b(n34451), .o(n34454) );
no02f01 g30664 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_5_), .b(n34439), .o(n34455) );
no02f01 g30665 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_6_), .b(n34439), .o(n34456) );
no02f01 g30666 ( .a(n34456), .b(n34455), .o(n34457) );
in01f01 g30667 ( .a(n34457), .o(n34458) );
no02f01 g30668 ( .a(n34458), .b(n34454), .o(n34459) );
no02f01 g30669 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_7_), .b(n34439), .o(n34460) );
in01f01 g30670 ( .a(n34460), .o(n34461) );
in01f01 g30671 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_4_), .o(n34462) );
in01f01 g30672 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_5_), .o(n34463) );
ao12f01 g30673 ( .a(delay_sub_ln23_unr21_stage7_stallmux_q_1_), .b(n34463), .c(n34462), .o(n34464) );
in01f01 g30674 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_6_), .o(n34465) );
in01f01 g30675 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_7_), .o(n34466) );
ao12f01 g30676 ( .a(delay_sub_ln23_unr21_stage7_stallmux_q_1_), .b(n34466), .c(n34465), .o(n34467) );
no02f01 g30677 ( .a(n34467), .b(n34464), .o(n34468) );
in01f01 g30678 ( .a(n34468), .o(n34469) );
ao12f01 g30679 ( .a(n34469), .b(n34461), .c(n34459), .o(n34470) );
no02f01 g30680 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_8_), .b(n34439), .o(n34471) );
no03f01 g30681 ( .a(n34471), .b(n34470), .c(n34426), .o(n34472) );
ao12f01 g30682 ( .a(n34436), .b(n34472), .c(n34425), .o(n34473) );
no02f01 g30683 ( .a(n34473), .b(n34422), .o(n34474) );
no02f01 g30684 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_15_), .b(n34420), .o(n34475) );
no02f01 g30685 ( .a(n34420), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_14_), .o(n34476) );
no02f01 g30686 ( .a(n34476), .b(n34475), .o(n34477) );
in01f01 g30687 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_12_), .o(n34478) );
in01f01 g30688 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_13_), .o(n34479) );
ao12f01 g30689 ( .a(n_27923), .b(n34479), .c(n34478), .o(n34480) );
in01f01 g30690 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_14_), .o(n34481) );
in01f01 g30691 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_15_), .o(n34482) );
ao12f01 g30692 ( .a(n_27923), .b(n34482), .c(n34481), .o(n34483) );
no02f01 g30693 ( .a(n34483), .b(n34480), .o(n34484) );
in01f01 g30694 ( .a(n34484), .o(n34485) );
ao12f01 g30695 ( .a(n34485), .b(n34477), .c(n34474), .o(n34486) );
ao12f01 g30696 ( .a(n34420), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_17_), .c(delay_sub_ln23_0_unr20_stage7_stallmux_q_16_), .o(n34487) );
no02f01 g30697 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_19_), .b(n34420), .o(n34488) );
no02f01 g30698 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_18_), .b(n34420), .o(n34489) );
no03f01 g30699 ( .a(n34489), .b(n34488), .c(n34487), .o(n34490) );
in01f01 g30700 ( .a(n34490), .o(n34491) );
no02f01 g30701 ( .a(n34491), .b(n34486), .o(n34492) );
no02f01 g30702 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_21_), .b(n34420), .o(n34493) );
no02f01 g30703 ( .a(n34420), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_20_), .o(n34494) );
no02f01 g30704 ( .a(n34494), .b(n34493), .o(n34495) );
in01f01 g30705 ( .a(n34495), .o(n34496) );
no02f01 g30706 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_23_), .b(n34420), .o(n34497) );
no02f01 g30707 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_22_), .b(n34420), .o(n34498) );
no03f01 g30708 ( .a(n34498), .b(n34497), .c(n34496), .o(n34499) );
na02f01 g30709 ( .a(n34499), .b(n34492), .o(n34500) );
no02f01 g30710 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_25_), .b(n34420), .o(n34501) );
no02f01 g30711 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_24_), .b(n34420), .o(n34502) );
no02f01 g30712 ( .a(n34502), .b(n34501), .o(n34503) );
in01f01 g30713 ( .a(n34503), .o(n34504) );
no02f01 g30714 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_26_), .b(n34420), .o(n34505) );
no02f01 g30715 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_27_), .b(n34420), .o(n34506) );
no03f01 g30716 ( .a(n34506), .b(n34505), .c(n34504), .o(n34507) );
in01f01 g30717 ( .a(n34507), .o(n34508) );
no02f01 g30718 ( .a(n34508), .b(n34500), .o(n34509) );
no02f01 g30719 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_28_), .b(n34420), .o(n34510) );
no02f01 g30720 ( .a(n34420), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_29_), .o(n34511) );
no02f01 g30721 ( .a(n34511), .b(n34510), .o(n34512) );
na02f01 g30722 ( .a(n34512), .b(n34509), .o(n34513) );
in01f01 g30723 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_19_), .o(n34514) );
no02f01 g30724 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_17_), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_16_), .o(n34515) );
na02f01 g30725 ( .a(n34515), .b(n34514), .o(n34516) );
oa12f01 g30726 ( .a(n34420), .b(n34516), .c(delay_sub_ln23_0_unr20_stage7_stallmux_q_18_), .o(n34517) );
in01f01 g30727 ( .a(n34517), .o(n34518) );
in01f01 g30728 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_20_), .o(n34519) );
in01f01 g30729 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_21_), .o(n34520) );
ao12f01 g30730 ( .a(n_27923), .b(n34520), .c(n34519), .o(n34521) );
no02f01 g30731 ( .a(n34521), .b(n34518), .o(n34522) );
in01f01 g30732 ( .a(n34522), .o(n34523) );
in01f01 g30733 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_22_), .o(n34524) );
in01f01 g30734 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_23_), .o(n34525) );
ao12f01 g30735 ( .a(n_27923), .b(n34525), .c(n34524), .o(n34526) );
no02f01 g30736 ( .a(n34526), .b(n34523), .o(n34527) );
in01f01 g30737 ( .a(n34527), .o(n34528) );
in01f01 g30738 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_25_), .o(n34529) );
in01f01 g30739 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_24_), .o(n34530) );
ao12f01 g30740 ( .a(n_27923), .b(n34530), .c(n34529), .o(n34531) );
no02f01 g30741 ( .a(n34531), .b(n34528), .o(n34532) );
in01f01 g30742 ( .a(n34532), .o(n34533) );
in01f01 g30743 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_27_), .o(n34534) );
in01f01 g30744 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_26_), .o(n34535) );
ao12f01 g30745 ( .a(n_27923), .b(n34535), .c(n34534), .o(n34536) );
no02f01 g30746 ( .a(n34536), .b(n34533), .o(n34537) );
in01f01 g30747 ( .a(n34537), .o(n34538) );
in01f01 g30748 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_30_), .o(n34539) );
in01f01 g30749 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_29_), .o(n34540) );
in01f01 g30750 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_28_), .o(n34541) );
ao12f01 g30751 ( .a(n_27923), .b(n34541), .c(n34540), .o(n34542) );
in01f01 g30752 ( .a(n34542), .o(n34543) );
ao12f01 g30753 ( .a(n_27923), .b(n34543), .c(n34539), .o(n34544) );
no02f01 g30754 ( .a(n34544), .b(n34538), .o(n34545) );
oa12f01 g30755 ( .a(n34545), .b(n34513), .c(n34421), .o(n34546) );
in01f01 g30756 ( .a(n34440), .o(n34547) );
no03f01 g30757 ( .a(n34441), .b(n34547), .c(n_186), .o(n34548) );
in01f01 g30758 ( .a(n34441), .o(n34549) );
ao12f01 g30759 ( .a(n34438), .b(n34549), .c(n34440), .o(n34550) );
no02f01 g30760 ( .a(n34550), .b(n34548), .o(n34551) );
na02f01 g30761 ( .a(n34551), .b(n34546), .o(n34552) );
na02f01 g30762 ( .a(n34552), .b(n34438), .o(n34553) );
no02f01 g30763 ( .a(n34551), .b(n34546), .o(n34554) );
in01f01 g30764 ( .a(n34554), .o(n34555) );
na02f01 g30765 ( .a(n34555), .b(n34553), .o(n34556) );
in01f01 g30766 ( .a(n34546), .o(n5380) );
no02f01 g30767 ( .a(n34443), .b(n34447), .o(n34558) );
in01f01 g30768 ( .a(n34558), .o(n34559) );
no02f01 g30769 ( .a(n34559), .b(n34442), .o(n34560) );
in01f01 g30770 ( .a(n34442), .o(n34561) );
no02f01 g30771 ( .a(n34558), .b(n34561), .o(n34562) );
no02f01 g30772 ( .a(n34562), .b(n34560), .o(n34563) );
in01f01 g30773 ( .a(n34563), .o(n34564) );
no02f01 g30774 ( .a(n34564), .b(n5380), .o(n34565) );
in01f01 g30775 ( .a(n34565), .o(n34566) );
na02f01 g30776 ( .a(n34566), .b(n34556), .o(n34567) );
no02f01 g30777 ( .a(n34437), .b(delay_sub_ln23_unr21_stage7_stallmux_q_1_), .o(n34568) );
no02f01 g30778 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_3_), .b(n34439), .o(n34569) );
no02f01 g30779 ( .a(n34569), .b(n34568), .o(n34570) );
in01f01 g30780 ( .a(n34570), .o(n34571) );
no02f01 g30781 ( .a(n34571), .b(n34449), .o(n34572) );
ao12f01 g30782 ( .a(n34570), .b(n34445), .c(n34448), .o(n34573) );
no02f01 g30783 ( .a(n34573), .b(n34572), .o(n34574) );
in01f01 g30784 ( .a(n34574), .o(n34575) );
no02f01 g30785 ( .a(n34563), .b(n34546), .o(n34576) );
in01f01 g30786 ( .a(n34576), .o(n34577) );
na02f01 g30787 ( .a(n34577), .b(n34567), .o(n34578) );
no02f01 g30788 ( .a(n34578), .b(n34575), .o(n34579) );
oa22f01 g30789 ( .a(n34579), .b(n34546), .c(n34574), .d(n34567), .o(n34580) );
no02f01 g30790 ( .a(n34462), .b(delay_sub_ln23_unr21_stage7_stallmux_q_1_), .o(n34581) );
no02f01 g30791 ( .a(n34581), .b(n34452), .o(n34582) );
in01f01 g30792 ( .a(n34582), .o(n34583) );
no02f01 g30793 ( .a(n34583), .b(n34451), .o(n34584) );
in01f01 g30794 ( .a(n34451), .o(n34585) );
no02f01 g30795 ( .a(n34582), .b(n34585), .o(n34586) );
no02f01 g30796 ( .a(n34586), .b(n34584), .o(n34587) );
in01f01 g30797 ( .a(n34587), .o(n34588) );
no02f01 g30798 ( .a(n34588), .b(n5380), .o(n34589) );
in01f01 g30799 ( .a(n34589), .o(n34590) );
na02f01 g30800 ( .a(n34590), .b(n34580), .o(n34591) );
ao12f01 g30801 ( .a(n34581), .b(n34453), .c(n34451), .o(n34592) );
no02f01 g30802 ( .a(n34463), .b(delay_sub_ln23_unr21_stage7_stallmux_q_1_), .o(n34593) );
no02f01 g30803 ( .a(n34593), .b(n34455), .o(n34594) );
no02f01 g30804 ( .a(n34594), .b(n34592), .o(n34595) );
na02f01 g30805 ( .a(n34594), .b(n34592), .o(n34596) );
in01f01 g30806 ( .a(n34596), .o(n34597) );
no02f01 g30807 ( .a(n34597), .b(n34595), .o(n34598) );
in01f01 g30808 ( .a(n34598), .o(n34599) );
no02f01 g30809 ( .a(n34599), .b(n5380), .o(n34600) );
in01f01 g30810 ( .a(n34464), .o(n34601) );
oa12f01 g30811 ( .a(n34601), .b(n34455), .c(n34454), .o(n34602) );
no02f01 g30812 ( .a(n34465), .b(delay_sub_ln23_unr21_stage7_stallmux_q_1_), .o(n34603) );
no02f01 g30813 ( .a(n34603), .b(n34456), .o(n34604) );
in01f01 g30814 ( .a(n34604), .o(n34605) );
no02f01 g30815 ( .a(n34605), .b(n34602), .o(n34606) );
na02f01 g30816 ( .a(n34605), .b(n34602), .o(n34607) );
in01f01 g30817 ( .a(n34607), .o(n34608) );
no02f01 g30818 ( .a(n34608), .b(n34606), .o(n34609) );
in01f01 g30819 ( .a(n34609), .o(n34610) );
no02f01 g30820 ( .a(n34610), .b(n5380), .o(n34611) );
no02f01 g30821 ( .a(n34611), .b(n34600), .o(n34612) );
in01f01 g30822 ( .a(n34612), .o(n34613) );
no02f01 g30823 ( .a(n34613), .b(n34591), .o(n34614) );
no03f01 g30824 ( .a(n34603), .b(n34464), .c(n34459), .o(n34615) );
in01f01 g30825 ( .a(n34615), .o(n34616) );
no02f01 g30826 ( .a(n34466), .b(delay_sub_ln23_unr21_stage7_stallmux_q_1_), .o(n34617) );
no02f01 g30827 ( .a(n34617), .b(n34460), .o(n34618) );
in01f01 g30828 ( .a(n34618), .o(n34619) );
no02f01 g30829 ( .a(n34619), .b(n34616), .o(n34620) );
no02f01 g30830 ( .a(n34618), .b(n34615), .o(n34621) );
no02f01 g30831 ( .a(n34621), .b(n34620), .o(n34622) );
in01f01 g30832 ( .a(n34622), .o(n34623) );
no02f01 g30833 ( .a(n34623), .b(n5380), .o(n34624) );
in01f01 g30834 ( .a(n34624), .o(n34625) );
na02f01 g30835 ( .a(n34625), .b(n34614), .o(n34626) );
ao12f01 g30836 ( .a(n34546), .b(n34598), .c(n34587), .o(n34627) );
ao12f01 g30837 ( .a(n34546), .b(n34622), .c(n34609), .o(n34628) );
no02f01 g30838 ( .a(n34628), .b(n34627), .o(n34629) );
na02f01 g30839 ( .a(n34629), .b(n34626), .o(n34630) );
no02f01 g30840 ( .a(n34471), .b(n34470), .o(n34631) );
no02f01 g30841 ( .a(n34631), .b(n34428), .o(n34632) );
in01f01 g30842 ( .a(n34426), .o(n34633) );
na02f01 g30843 ( .a(n34430), .b(n34633), .o(n34634) );
in01f01 g30844 ( .a(n34634), .o(n34635) );
no02f01 g30845 ( .a(n34635), .b(n34632), .o(n34636) );
na02f01 g30846 ( .a(n34635), .b(n34632), .o(n34637) );
in01f01 g30847 ( .a(n34637), .o(n34638) );
no02f01 g30848 ( .a(n34638), .b(n34636), .o(n34639) );
in01f01 g30849 ( .a(n34639), .o(n34640) );
no02f01 g30850 ( .a(n34640), .b(n34546), .o(n34641) );
in01f01 g30851 ( .a(n34470), .o(n34642) );
no02f01 g30852 ( .a(n34471), .b(n34428), .o(n34643) );
in01f01 g30853 ( .a(n34643), .o(n34644) );
no02f01 g30854 ( .a(n34644), .b(n34642), .o(n34645) );
no02f01 g30855 ( .a(n34643), .b(n34470), .o(n34646) );
no02f01 g30856 ( .a(n34646), .b(n34645), .o(n34647) );
in01f01 g30857 ( .a(n34647), .o(n34648) );
no02f01 g30858 ( .a(n34648), .b(n34546), .o(n34649) );
no02f01 g30859 ( .a(n34649), .b(n34641), .o(n34650) );
in01f01 g30860 ( .a(n34650), .o(n34651) );
in01f01 g30861 ( .a(n34424), .o(n34652) );
no02f01 g30862 ( .a(n_27923), .b(n34432), .o(n34653) );
no02f01 g30863 ( .a(n34472), .b(n34431), .o(n34654) );
in01f01 g30864 ( .a(n34654), .o(n34655) );
ao12f01 g30865 ( .a(n34653), .b(n34655), .c(n34652), .o(n34656) );
in01f01 g30866 ( .a(n34656), .o(n34657) );
no02f01 g30867 ( .a(n34433), .b(n_27923), .o(n34658) );
no02f01 g30868 ( .a(n34658), .b(n34423), .o(n34659) );
in01f01 g30869 ( .a(n34659), .o(n34660) );
no02f01 g30870 ( .a(n34660), .b(n34657), .o(n34661) );
no02f01 g30871 ( .a(n34659), .b(n34656), .o(n34662) );
no02f01 g30872 ( .a(n34662), .b(n34661), .o(n34663) );
in01f01 g30873 ( .a(n34663), .o(n34664) );
no02f01 g30874 ( .a(n34664), .b(n34546), .o(n34665) );
no02f01 g30875 ( .a(n34653), .b(n34424), .o(n34666) );
no02f01 g30876 ( .a(n34666), .b(n34654), .o(n34667) );
na02f01 g30877 ( .a(n34666), .b(n34654), .o(n34668) );
in01f01 g30878 ( .a(n34668), .o(n34669) );
no02f01 g30879 ( .a(n34669), .b(n34667), .o(n34670) );
in01f01 g30880 ( .a(n34670), .o(n34671) );
no02f01 g30881 ( .a(n34671), .b(n34546), .o(n34672) );
no03f01 g30882 ( .a(n34672), .b(n34665), .c(n34651), .o(n34673) );
na02f01 g30883 ( .a(n34673), .b(n34630), .o(n34674) );
no02f01 g30884 ( .a(n34478), .b(n_27923), .o(n34675) );
no02f01 g30885 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_12_), .b(n34420), .o(n34676) );
no02f01 g30886 ( .a(n34676), .b(n34473), .o(n34677) );
no02f01 g30887 ( .a(n34677), .b(n34675), .o(n34678) );
no02f01 g30888 ( .a(n34479), .b(n_27923), .o(n34679) );
no02f01 g30889 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_13_), .b(n34420), .o(n34680) );
no02f01 g30890 ( .a(n34680), .b(n34679), .o(n34681) );
no02f01 g30891 ( .a(n34681), .b(n34678), .o(n34682) );
na02f01 g30892 ( .a(n34681), .b(n34678), .o(n34683) );
in01f01 g30893 ( .a(n34683), .o(n34684) );
no02f01 g30894 ( .a(n34684), .b(n34682), .o(n34685) );
in01f01 g30895 ( .a(n34685), .o(n34686) );
no02f01 g30896 ( .a(n34686), .b(n34546), .o(n34687) );
no02f01 g30897 ( .a(n34676), .b(n34675), .o(n34688) );
no02f01 g30898 ( .a(n34688), .b(n34473), .o(n34689) );
na02f01 g30899 ( .a(n34688), .b(n34473), .o(n34690) );
in01f01 g30900 ( .a(n34690), .o(n34691) );
no02f01 g30901 ( .a(n34691), .b(n34689), .o(n34692) );
in01f01 g30902 ( .a(n34692), .o(n34693) );
no02f01 g30903 ( .a(n34693), .b(n34546), .o(n34694) );
no02f01 g30904 ( .a(n34694), .b(n34687), .o(n34695) );
in01f01 g30905 ( .a(n34695), .o(n34696) );
no02f01 g30906 ( .a(n34480), .b(n34474), .o(n34697) );
in01f01 g30907 ( .a(n34697), .o(n34698) );
no02f01 g30908 ( .a(n_27923), .b(n34481), .o(n34699) );
no02f01 g30909 ( .a(n34699), .b(n34476), .o(n34700) );
in01f01 g30910 ( .a(n34700), .o(n34701) );
no02f01 g30911 ( .a(n34701), .b(n34698), .o(n34702) );
no02f01 g30912 ( .a(n34700), .b(n34697), .o(n34703) );
no02f01 g30913 ( .a(n34703), .b(n34702), .o(n34704) );
in01f01 g30914 ( .a(n34704), .o(n34705) );
no02f01 g30915 ( .a(n34705), .b(n34546), .o(n34706) );
in01f01 g30916 ( .a(n34476), .o(n34707) );
oa12f01 g30917 ( .a(n34707), .b(n34698), .c(n34699), .o(n34708) );
no02f01 g30918 ( .a(n34482), .b(n_27923), .o(n34709) );
no02f01 g30919 ( .a(n34709), .b(n34475), .o(n34710) );
no02f01 g30920 ( .a(n34710), .b(n34708), .o(n34711) );
na02f01 g30921 ( .a(n34710), .b(n34708), .o(n34712) );
in01f01 g30922 ( .a(n34712), .o(n34713) );
no02f01 g30923 ( .a(n34713), .b(n34711), .o(n34714) );
in01f01 g30924 ( .a(n34714), .o(n34715) );
no02f01 g30925 ( .a(n34715), .b(n34546), .o(n34716) );
no04f01 g30926 ( .a(n34716), .b(n34706), .c(n34696), .d(n34674), .o(n34717) );
ao12f01 g30927 ( .a(n5380), .b(n34647), .c(n34639), .o(n34718) );
ao12f01 g30928 ( .a(n5380), .b(n34670), .c(n34663), .o(n34719) );
no02f01 g30929 ( .a(n34719), .b(n34718), .o(n34720) );
in01f01 g30930 ( .a(n34720), .o(n34721) );
ao12f01 g30931 ( .a(n5380), .b(n34692), .c(n34685), .o(n34722) );
no02f01 g30932 ( .a(n34722), .b(n34721), .o(n34723) );
in01f01 g30933 ( .a(n34723), .o(n34724) );
ao12f01 g30934 ( .a(n5380), .b(n34714), .c(n34704), .o(n34725) );
no02f01 g30935 ( .a(n34725), .b(n34724), .o(n34726) );
in01f01 g30936 ( .a(n34726), .o(n34727) );
no02f01 g30937 ( .a(n34727), .b(n34717), .o(n34728) );
in01f01 g30938 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_16_), .o(n34729) );
no02f01 g30939 ( .a(n_27923), .b(n34729), .o(n34730) );
no02f01 g30940 ( .a(n34420), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_16_), .o(n34731) );
no02f01 g30941 ( .a(n34731), .b(n34486), .o(n34732) );
no02f01 g30942 ( .a(n34732), .b(n34730), .o(n34733) );
in01f01 g30943 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_17_), .o(n34734) );
no02f01 g30944 ( .a(n34734), .b(n_27923), .o(n34735) );
no02f01 g30945 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_17_), .b(n34420), .o(n34736) );
no02f01 g30946 ( .a(n34736), .b(n34735), .o(n34737) );
no02f01 g30947 ( .a(n34737), .b(n34733), .o(n34738) );
na02f01 g30948 ( .a(n34737), .b(n34733), .o(n34739) );
in01f01 g30949 ( .a(n34739), .o(n34740) );
no02f01 g30950 ( .a(n34740), .b(n34738), .o(n34741) );
in01f01 g30951 ( .a(n34741), .o(n34742) );
no02f01 g30952 ( .a(n34742), .b(n34546), .o(n34743) );
in01f01 g30953 ( .a(n34486), .o(n34744) );
no02f01 g30954 ( .a(n34731), .b(n34730), .o(n34745) );
in01f01 g30955 ( .a(n34745), .o(n34746) );
no02f01 g30956 ( .a(n34746), .b(n34744), .o(n34747) );
no02f01 g30957 ( .a(n34745), .b(n34486), .o(n34748) );
no02f01 g30958 ( .a(n34748), .b(n34747), .o(n34749) );
in01f01 g30959 ( .a(n34749), .o(n34750) );
no02f01 g30960 ( .a(n34750), .b(n34546), .o(n34751) );
no02f01 g30961 ( .a(n34751), .b(n34743), .o(n34752) );
in01f01 g30962 ( .a(n34752), .o(n34753) );
no02f01 g30963 ( .a(n34487), .b(n34486), .o(n34754) );
no02f01 g30964 ( .a(n34515), .b(n_27923), .o(n34755) );
no02f01 g30965 ( .a(n34755), .b(n34754), .o(n34756) );
in01f01 g30966 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_18_), .o(n34757) );
no02f01 g30967 ( .a(n34757), .b(n_27923), .o(n34758) );
no02f01 g30968 ( .a(n34758), .b(n34489), .o(n34759) );
no02f01 g30969 ( .a(n34759), .b(n34756), .o(n34760) );
na02f01 g30970 ( .a(n34759), .b(n34756), .o(n34761) );
in01f01 g30971 ( .a(n34761), .o(n34762) );
no02f01 g30972 ( .a(n34762), .b(n34760), .o(n34763) );
in01f01 g30973 ( .a(n34763), .o(n34764) );
no02f01 g30974 ( .a(n34764), .b(n34546), .o(n34765) );
no03f01 g30975 ( .a(n34489), .b(n34487), .c(n34486), .o(n34766) );
no03f01 g30976 ( .a(n34766), .b(n34755), .c(n34758), .o(n34767) );
in01f01 g30977 ( .a(n34767), .o(n34768) );
no02f01 g30978 ( .a(n34514), .b(n_27923), .o(n34769) );
no02f01 g30979 ( .a(n34769), .b(n34488), .o(n34770) );
in01f01 g30980 ( .a(n34770), .o(n34771) );
no02f01 g30981 ( .a(n34771), .b(n34768), .o(n34772) );
no02f01 g30982 ( .a(n34770), .b(n34767), .o(n34773) );
no02f01 g30983 ( .a(n34773), .b(n34772), .o(n34774) );
in01f01 g30984 ( .a(n34774), .o(n34775) );
no02f01 g30985 ( .a(n34775), .b(n34546), .o(n34776) );
no03f01 g30986 ( .a(n34776), .b(n34765), .c(n34753), .o(n34777) );
in01f01 g30987 ( .a(n34777), .o(n34778) );
no02f01 g30988 ( .a(n34778), .b(n34728), .o(n34779) );
ao12f01 g30989 ( .a(n34523), .b(n34495), .c(n34492), .o(n34780) );
no02f01 g30990 ( .a(n34524), .b(n_27923), .o(n34781) );
no02f01 g30991 ( .a(n34781), .b(n34498), .o(n34782) );
no02f01 g30992 ( .a(n34782), .b(n34780), .o(n34783) );
na02f01 g30993 ( .a(n34782), .b(n34780), .o(n34784) );
in01f01 g30994 ( .a(n34784), .o(n34785) );
no03f01 g30995 ( .a(n34785), .b(n34783), .c(n34546), .o(n34786) );
in01f01 g30996 ( .a(n34492), .o(n34787) );
no03f01 g30997 ( .a(n34498), .b(n34496), .c(n34787), .o(n34788) );
no03f01 g30998 ( .a(n34788), .b(n34781), .c(n34523), .o(n34789) );
in01f01 g30999 ( .a(n34789), .o(n34790) );
no02f01 g31000 ( .a(n34525), .b(n_27923), .o(n34791) );
no02f01 g31001 ( .a(n34791), .b(n34497), .o(n34792) );
in01f01 g31002 ( .a(n34792), .o(n34793) );
no02f01 g31003 ( .a(n34793), .b(n34790), .o(n34794) );
no02f01 g31004 ( .a(n34792), .b(n34789), .o(n34795) );
no03f01 g31005 ( .a(n34795), .b(n34794), .c(n34546), .o(n34796) );
no02f01 g31006 ( .a(n_27923), .b(n34519), .o(n34797) );
no02f01 g31007 ( .a(n34797), .b(n34518), .o(n34798) );
oa12f01 g31008 ( .a(n34798), .b(n34494), .c(n34787), .o(n34799) );
in01f01 g31009 ( .a(n34799), .o(n34800) );
no02f01 g31010 ( .a(n34520), .b(n_27923), .o(n34801) );
no02f01 g31011 ( .a(n34801), .b(n34493), .o(n34802) );
no02f01 g31012 ( .a(n34802), .b(n34800), .o(n34803) );
na02f01 g31013 ( .a(n34802), .b(n34800), .o(n34804) );
in01f01 g31014 ( .a(n34804), .o(n34805) );
no03f01 g31015 ( .a(n34805), .b(n34803), .c(n34546), .o(n34806) );
no02f01 g31016 ( .a(n34797), .b(n34494), .o(n34807) );
in01f01 g31017 ( .a(n34807), .o(n34808) );
no03f01 g31018 ( .a(n34808), .b(n34518), .c(n34492), .o(n34809) );
ao12f01 g31019 ( .a(n34807), .b(n34517), .c(n34787), .o(n34810) );
no02f01 g31020 ( .a(n34810), .b(n34809), .o(n34811) );
in01f01 g31021 ( .a(n34811), .o(n34812) );
no02f01 g31022 ( .a(n34812), .b(n34546), .o(n34813) );
no04f01 g31023 ( .a(n34813), .b(n34806), .c(n34796), .d(n34786), .o(n34814) );
in01f01 g31024 ( .a(n34500), .o(n34815) );
no02f01 g31025 ( .a(n34530), .b(n_27923), .o(n34816) );
no02f01 g31026 ( .a(n34816), .b(n34502), .o(n34817) );
in01f01 g31027 ( .a(n34817), .o(n34818) );
no03f01 g31028 ( .a(n34818), .b(n34528), .c(n34815), .o(n34819) );
ao12f01 g31029 ( .a(n34817), .b(n34527), .c(n34500), .o(n34820) );
no02f01 g31030 ( .a(n34820), .b(n34819), .o(n34821) );
in01f01 g31031 ( .a(n34821), .o(n34822) );
no02f01 g31032 ( .a(n34822), .b(n34546), .o(n34823) );
in01f01 g31033 ( .a(n34823), .o(n34824) );
no02f01 g31034 ( .a(n34535), .b(n_27923), .o(n34825) );
no03f01 g31035 ( .a(n34505), .b(n34504), .c(n34500), .o(n34826) );
no03f01 g31036 ( .a(n34826), .b(n34825), .c(n34533), .o(n34827) );
no02f01 g31037 ( .a(n34534), .b(n_27923), .o(n34828) );
no02f01 g31038 ( .a(n34828), .b(n34506), .o(n34829) );
no02f01 g31039 ( .a(n34829), .b(n34827), .o(n34830) );
na02f01 g31040 ( .a(n34829), .b(n34827), .o(n34831) );
in01f01 g31041 ( .a(n34831), .o(n34832) );
no03f01 g31042 ( .a(n34832), .b(n34830), .c(n34546), .o(n34833) );
no02f01 g31043 ( .a(n34816), .b(n34528), .o(n34834) );
oa12f01 g31044 ( .a(n34834), .b(n34502), .c(n34500), .o(n34835) );
no02f01 g31045 ( .a(n34529), .b(n_27923), .o(n34836) );
no02f01 g31046 ( .a(n34836), .b(n34501), .o(n34837) );
in01f01 g31047 ( .a(n34837), .o(n34838) );
no02f01 g31048 ( .a(n34838), .b(n34835), .o(n34839) );
na02f01 g31049 ( .a(n34838), .b(n34835), .o(n34840) );
in01f01 g31050 ( .a(n34840), .o(n34841) );
no02f01 g31051 ( .a(n34841), .b(n34839), .o(n34842) );
in01f01 g31052 ( .a(n34842), .o(n34843) );
no02f01 g31053 ( .a(n34843), .b(n34546), .o(n34844) );
no02f01 g31054 ( .a(n34504), .b(n34500), .o(n34845) );
no02f01 g31055 ( .a(n34825), .b(n34505), .o(n34846) );
in01f01 g31056 ( .a(n34846), .o(n34847) );
no03f01 g31057 ( .a(n34847), .b(n34845), .c(n34533), .o(n34848) );
no02f01 g31058 ( .a(n34845), .b(n34533), .o(n34849) );
no02f01 g31059 ( .a(n34846), .b(n34849), .o(n34850) );
no03f01 g31060 ( .a(n34850), .b(n34848), .c(n34546), .o(n34851) );
no03f01 g31061 ( .a(n34851), .b(n34844), .c(n34833), .o(n34852) );
na04f01 g31062 ( .a(n34852), .b(n34824), .c(n34814), .d(n34779), .o(n34853) );
no02f01 g31063 ( .a(n34541), .b(n_27923), .o(n34854) );
no03f01 g31064 ( .a(n34510), .b(n34508), .c(n34500), .o(n34855) );
no03f01 g31065 ( .a(n34855), .b(n34854), .c(n34538), .o(n34856) );
in01f01 g31066 ( .a(n34856), .o(n34857) );
no02f01 g31067 ( .a(n_27923), .b(n34540), .o(n34858) );
no02f01 g31068 ( .a(n34858), .b(n34511), .o(n34859) );
in01f01 g31069 ( .a(n34859), .o(n34860) );
no02f01 g31070 ( .a(n34860), .b(n34857), .o(n34861) );
no02f01 g31071 ( .a(n34859), .b(n34856), .o(n34862) );
no03f01 g31072 ( .a(n34862), .b(n34861), .c(n34546), .o(n34863) );
no02f01 g31073 ( .a(n34854), .b(n34510), .o(n34864) );
in01f01 g31074 ( .a(n34864), .o(n34865) );
no03f01 g31075 ( .a(n34865), .b(n34538), .c(n34509), .o(n34866) );
no02f01 g31076 ( .a(n34538), .b(n34509), .o(n34867) );
no02f01 g31077 ( .a(n34864), .b(n34867), .o(n34868) );
no03f01 g31078 ( .a(n34868), .b(n34866), .c(n34546), .o(n34869) );
no02f01 g31079 ( .a(n34869), .b(n34863), .o(n34870) );
in01f01 g31080 ( .a(n34870), .o(n34871) );
na03f01 g31081 ( .a(n34543), .b(n34537), .c(n34513), .o(n34872) );
no02f01 g31082 ( .a(n34539), .b(n_27923), .o(n34873) );
no02f01 g31083 ( .a(n34873), .b(n34421), .o(n34874) );
in01f01 g31084 ( .a(n34874), .o(n34875) );
no02f01 g31085 ( .a(n34875), .b(n34872), .o(n34876) );
na02f01 g31086 ( .a(n34875), .b(n34872), .o(n34877) );
in01f01 g31087 ( .a(n34877), .o(n34878) );
no03f01 g31088 ( .a(n34878), .b(n34876), .c(n34546), .o(n34879) );
no02f01 g31089 ( .a(n34879), .b(n34871), .o(n34880) );
in01f01 g31090 ( .a(n34880), .o(n34881) );
no03f01 g31091 ( .a(n34775), .b(n34750), .c(n34742), .o(n34882) );
ao12f01 g31092 ( .a(n5380), .b(n34882), .c(n34763), .o(n34883) );
no02f01 g31093 ( .a(n34805), .b(n34803), .o(n34884) );
ao12f01 g31094 ( .a(n5380), .b(n34811), .c(n34884), .o(n34885) );
no02f01 g31095 ( .a(n34885), .b(n34883), .o(n34886) );
in01f01 g31096 ( .a(n34886), .o(n34887) );
no02f01 g31097 ( .a(n34785), .b(n34783), .o(n34888) );
no02f01 g31098 ( .a(n34795), .b(n34794), .o(n34889) );
ao12f01 g31099 ( .a(n5380), .b(n34889), .c(n34888), .o(n34890) );
no02f01 g31100 ( .a(n34890), .b(n34887), .o(n34891) );
in01f01 g31101 ( .a(n34891), .o(n34892) );
ao12f01 g31102 ( .a(n5380), .b(n34842), .c(n34821), .o(n34893) );
no02f01 g31103 ( .a(n34893), .b(n34892), .o(n34894) );
in01f01 g31104 ( .a(n34894), .o(n34895) );
no02f01 g31105 ( .a(n34832), .b(n34830), .o(n34896) );
no02f01 g31106 ( .a(n34850), .b(n34848), .o(n34897) );
ao12f01 g31107 ( .a(n5380), .b(n34897), .c(n34896), .o(n34898) );
no02f01 g31108 ( .a(n34898), .b(n34895), .o(n34899) );
in01f01 g31109 ( .a(n34899), .o(n34900) );
no02f01 g31110 ( .a(n34878), .b(n34876), .o(n34901) );
no02f01 g31111 ( .a(n34862), .b(n34861), .o(n34902) );
no02f01 g31112 ( .a(n34868), .b(n34866), .o(n34903) );
ao12f01 g31113 ( .a(n5380), .b(n34903), .c(n34902), .o(n34904) );
in01f01 g31114 ( .a(n34904), .o(n34905) );
ao12f01 g31115 ( .a(n5380), .b(n34905), .c(n34901), .o(n34906) );
no02f01 g31116 ( .a(n34906), .b(n34900), .o(n34907) );
oa12f01 g31117 ( .a(n34907), .b(n34881), .c(n34853), .o(n34908) );
no02f01 g31118 ( .a(n34609), .b(n34546), .o(n34909) );
no02f01 g31119 ( .a(n34909), .b(n34627), .o(n34910) );
in01f01 g31120 ( .a(n34910), .o(n34911) );
no02f01 g31121 ( .a(n34622), .b(n34546), .o(n34912) );
no02f01 g31122 ( .a(n34912), .b(n34624), .o(n34913) );
in01f01 g31123 ( .a(n34913), .o(n34914) );
no03f01 g31124 ( .a(n34914), .b(n34911), .c(n34614), .o(n34915) );
no02f01 g31125 ( .a(n34911), .b(n34614), .o(n34916) );
no02f01 g31126 ( .a(n34913), .b(n34916), .o(n34917) );
no02f01 g31127 ( .a(n34917), .b(n34915), .o(n34918) );
in01f01 g31128 ( .a(n34918), .o(n34919) );
no02f01 g31129 ( .a(n34919), .b(n34908), .o(n34920) );
no02f01 g31130 ( .a(n34587), .b(n34546), .o(n34921) );
ao12f01 g31131 ( .a(n34921), .b(n34590), .c(n34580), .o(n34922) );
no02f01 g31132 ( .a(n34598), .b(n34546), .o(n34923) );
no02f01 g31133 ( .a(n34923), .b(n34600), .o(n34924) );
no02f01 g31134 ( .a(n34924), .b(n34922), .o(n34925) );
na02f01 g31135 ( .a(n34924), .b(n34922), .o(n34926) );
in01f01 g31136 ( .a(n34926), .o(n34927) );
no02f01 g31137 ( .a(n34927), .b(n34925), .o(n34928) );
in01f01 g31138 ( .a(n34580), .o(n34929) );
no02f01 g31139 ( .a(n34921), .b(n34589), .o(n34930) );
no02f01 g31140 ( .a(n34930), .b(n34929), .o(n34931) );
na02f01 g31141 ( .a(n34930), .b(n34929), .o(n34932) );
in01f01 g31142 ( .a(n34932), .o(n34933) );
no02f01 g31143 ( .a(n34933), .b(n34931), .o(n34934) );
ao12f01 g31144 ( .a(n34908), .b(n34934), .c(n34928), .o(n34935) );
in01f01 g31145 ( .a(n34908), .o(n5978) );
na02f01 g31146 ( .a(n34555), .b(n34552), .o(n34937) );
ao12f01 g31147 ( .a(n34438), .b(n34937), .c(n34908), .o(n34938) );
no02f01 g31148 ( .a(n34937), .b(n34438), .o(n34939) );
ao12f01 g31149 ( .a(n_186), .b(n34555), .c(n34552), .o(n34940) );
no02f01 g31150 ( .a(n34940), .b(n34939), .o(n34941) );
no02f01 g31151 ( .a(n34941), .b(n34908), .o(n34942) );
in01f01 g31152 ( .a(n34556), .o(n34943) );
no02f01 g31153 ( .a(n34576), .b(n34565), .o(n34944) );
no02f01 g31154 ( .a(n34944), .b(n34943), .o(n34945) );
na02f01 g31155 ( .a(n34944), .b(n34943), .o(n34946) );
in01f01 g31156 ( .a(n34946), .o(n34947) );
no02f01 g31157 ( .a(n34947), .b(n34945), .o(n34948) );
in01f01 g31158 ( .a(n34948), .o(n34949) );
oa22f01 g31159 ( .a(n34949), .b(n5978), .c(n34942), .d(n34938), .o(n34950) );
in01f01 g31160 ( .a(n34950), .o(n34951) );
no02f01 g31161 ( .a(n34574), .b(n34546), .o(n34952) );
no02f01 g31162 ( .a(n34575), .b(n5380), .o(n34953) );
no02f01 g31163 ( .a(n34953), .b(n34952), .o(n34954) );
in01f01 g31164 ( .a(n34954), .o(n34955) );
no02f01 g31165 ( .a(n34955), .b(n34578), .o(n34956) );
na02f01 g31166 ( .a(n34955), .b(n34578), .o(n34957) );
in01f01 g31167 ( .a(n34957), .o(n34958) );
no02f01 g31168 ( .a(n34958), .b(n34956), .o(n34959) );
in01f01 g31169 ( .a(n34959), .o(n34960) );
no02f01 g31170 ( .a(n34948), .b(n34908), .o(n34961) );
in01f01 g31171 ( .a(n34961), .o(n34962) );
na03f01 g31172 ( .a(n34959), .b(n34962), .c(n34950), .o(n34963) );
ao22f01 g31173 ( .a(n34963), .b(n5978), .c(n34960), .d(n34951), .o(n34964) );
in01f01 g31174 ( .a(n34934), .o(n34965) );
no02f01 g31175 ( .a(n34965), .b(n5978), .o(n34966) );
in01f01 g31176 ( .a(n34928), .o(n34967) );
no02f01 g31177 ( .a(n34967), .b(n5978), .o(n34968) );
no02f01 g31178 ( .a(n34600), .b(n34591), .o(n34969) );
no02f01 g31179 ( .a(n34909), .b(n34611), .o(n34970) );
in01f01 g31180 ( .a(n34970), .o(n34971) );
no03f01 g31181 ( .a(n34971), .b(n34969), .c(n34627), .o(n34972) );
no02f01 g31182 ( .a(n34969), .b(n34627), .o(n34973) );
no02f01 g31183 ( .a(n34970), .b(n34973), .o(n34974) );
no02f01 g31184 ( .a(n34974), .b(n34972), .o(n34975) );
in01f01 g31185 ( .a(n34975), .o(n34976) );
no02f01 g31186 ( .a(n34976), .b(n5978), .o(n34977) );
no04f01 g31187 ( .a(n34977), .b(n34968), .c(n34966), .d(n34964), .o(n34978) );
ao12f01 g31188 ( .a(n34918), .b(n34975), .c(n5978), .o(n34979) );
no03f01 g31189 ( .a(n34979), .b(n34978), .c(n34935), .o(n34980) );
no02f01 g31190 ( .a(n34647), .b(n5380), .o(n34981) );
no02f01 g31191 ( .a(n34981), .b(n34649), .o(n34982) );
in01f01 g31192 ( .a(n34982), .o(n34983) );
no02f01 g31193 ( .a(n34983), .b(n34630), .o(n34984) );
in01f01 g31194 ( .a(n34630), .o(n34985) );
no02f01 g31195 ( .a(n34982), .b(n34985), .o(n34986) );
no02f01 g31196 ( .a(n34986), .b(n34984), .o(n34987) );
in01f01 g31197 ( .a(n34987), .o(n34988) );
in01f01 g31198 ( .a(n34649), .o(n34989) );
ao12f01 g31199 ( .a(n34981), .b(n34989), .c(n34630), .o(n34990) );
in01f01 g31200 ( .a(n34990), .o(n34991) );
no02f01 g31201 ( .a(n34639), .b(n5380), .o(n34992) );
no02f01 g31202 ( .a(n34992), .b(n34641), .o(n34993) );
in01f01 g31203 ( .a(n34993), .o(n34994) );
no02f01 g31204 ( .a(n34994), .b(n34991), .o(n34995) );
no02f01 g31205 ( .a(n34993), .b(n34990), .o(n34996) );
no02f01 g31206 ( .a(n34996), .b(n34995), .o(n34997) );
in01f01 g31207 ( .a(n34997), .o(n34998) );
ao12f01 g31208 ( .a(n34908), .b(n34998), .c(n34988), .o(n34999) );
no02f01 g31209 ( .a(n34651), .b(n34985), .o(n35000) );
in01f01 g31210 ( .a(n35000), .o(n35001) );
no02f01 g31211 ( .a(n34670), .b(n5380), .o(n35002) );
no02f01 g31212 ( .a(n35002), .b(n34718), .o(n35003) );
oa12f01 g31213 ( .a(n35003), .b(n35001), .c(n34672), .o(n35004) );
in01f01 g31214 ( .a(n35004), .o(n35005) );
no02f01 g31215 ( .a(n34663), .b(n5380), .o(n35006) );
no02f01 g31216 ( .a(n35006), .b(n34665), .o(n35007) );
no02f01 g31217 ( .a(n35007), .b(n35005), .o(n35008) );
na02f01 g31218 ( .a(n35007), .b(n35005), .o(n35009) );
in01f01 g31219 ( .a(n35009), .o(n35010) );
no02f01 g31220 ( .a(n35010), .b(n35008), .o(n35011) );
in01f01 g31221 ( .a(n35011), .o(n35012) );
no02f01 g31222 ( .a(n35012), .b(n34908), .o(n35013) );
no02f01 g31223 ( .a(n35000), .b(n34718), .o(n35014) );
no02f01 g31224 ( .a(n35002), .b(n34672), .o(n35015) );
no02f01 g31225 ( .a(n35015), .b(n35014), .o(n35016) );
na02f01 g31226 ( .a(n35015), .b(n35014), .o(n35017) );
in01f01 g31227 ( .a(n35017), .o(n35018) );
no02f01 g31228 ( .a(n35018), .b(n35016), .o(n35019) );
in01f01 g31229 ( .a(n35019), .o(n35020) );
no02f01 g31230 ( .a(n35020), .b(n34908), .o(n35021) );
no02f01 g31231 ( .a(n35021), .b(n35013), .o(n35022) );
in01f01 g31232 ( .a(n35022), .o(n35023) );
no04f01 g31233 ( .a(n35023), .b(n34999), .c(n34980), .d(n34920), .o(n35024) );
ao12f01 g31234 ( .a(n5978), .b(n34997), .c(n34987), .o(n35025) );
ao12f01 g31235 ( .a(n5978), .b(n35019), .c(n35011), .o(n35026) );
no02f01 g31236 ( .a(n35026), .b(n35025), .o(n35027) );
in01f01 g31237 ( .a(n35027), .o(n35028) );
no02f01 g31238 ( .a(n34692), .b(n5380), .o(n35029) );
no02f01 g31239 ( .a(n35029), .b(n34721), .o(n35030) );
oa12f01 g31240 ( .a(n35030), .b(n34694), .c(n34674), .o(n35031) );
in01f01 g31241 ( .a(n35031), .o(n35032) );
no02f01 g31242 ( .a(n34685), .b(n5380), .o(n35033) );
no02f01 g31243 ( .a(n35033), .b(n34687), .o(n35034) );
no02f01 g31244 ( .a(n35034), .b(n35032), .o(n35035) );
na02f01 g31245 ( .a(n35034), .b(n35032), .o(n35036) );
in01f01 g31246 ( .a(n35036), .o(n35037) );
no02f01 g31247 ( .a(n35037), .b(n35035), .o(n35038) );
na02f01 g31248 ( .a(n34720), .b(n34674), .o(n35039) );
no02f01 g31249 ( .a(n35029), .b(n34694), .o(n35040) );
in01f01 g31250 ( .a(n35040), .o(n35041) );
no02f01 g31251 ( .a(n35041), .b(n35039), .o(n35042) );
na02f01 g31252 ( .a(n35041), .b(n35039), .o(n35043) );
in01f01 g31253 ( .a(n35043), .o(n35044) );
no02f01 g31254 ( .a(n35044), .b(n35042), .o(n35045) );
no02f01 g31255 ( .a(n35045), .b(n35038), .o(n35046) );
oa22f01 g31256 ( .a(n35046), .b(n34908), .c(n35028), .d(n35024), .o(n35047) );
no02f01 g31257 ( .a(n34696), .b(n34674), .o(n35048) );
in01f01 g31258 ( .a(n35048), .o(n35049) );
no02f01 g31259 ( .a(n34704), .b(n5380), .o(n35050) );
no02f01 g31260 ( .a(n35050), .b(n34724), .o(n35051) );
oa12f01 g31261 ( .a(n35051), .b(n34706), .c(n35049), .o(n35052) );
no02f01 g31262 ( .a(n34714), .b(n5380), .o(n35053) );
no02f01 g31263 ( .a(n35053), .b(n34716), .o(n35054) );
in01f01 g31264 ( .a(n35054), .o(n35055) );
no02f01 g31265 ( .a(n35055), .b(n35052), .o(n35056) );
na02f01 g31266 ( .a(n35055), .b(n35052), .o(n35057) );
in01f01 g31267 ( .a(n35057), .o(n35058) );
no02f01 g31268 ( .a(n35058), .b(n35056), .o(n35059) );
in01f01 g31269 ( .a(n35059), .o(n35060) );
no02f01 g31270 ( .a(n35060), .b(n34908), .o(n35061) );
no02f01 g31271 ( .a(n34724), .b(n35048), .o(n35062) );
no02f01 g31272 ( .a(n35050), .b(n34706), .o(n35063) );
no02f01 g31273 ( .a(n35063), .b(n35062), .o(n35064) );
na02f01 g31274 ( .a(n35063), .b(n35062), .o(n35065) );
in01f01 g31275 ( .a(n35065), .o(n35066) );
no02f01 g31276 ( .a(n35066), .b(n35064), .o(n35067) );
in01f01 g31277 ( .a(n35067), .o(n35068) );
no02f01 g31278 ( .a(n35068), .b(n34908), .o(n35069) );
no02f01 g31279 ( .a(n35069), .b(n35061), .o(n35070) );
in01f01 g31280 ( .a(n35070), .o(n35071) );
ao12f01 g31281 ( .a(n5978), .b(n35045), .c(n35038), .o(n35072) );
ao12f01 g31282 ( .a(n5978), .b(n35067), .c(n35059), .o(n35073) );
no02f01 g31283 ( .a(n35073), .b(n35072), .o(n35074) );
oa12f01 g31284 ( .a(n35074), .b(n35071), .c(n35047), .o(n35075) );
in01f01 g31285 ( .a(n34728), .o(n35076) );
in01f01 g31286 ( .a(n34751), .o(n35077) );
no02f01 g31287 ( .a(n34749), .b(n5380), .o(n35078) );
ao12f01 g31288 ( .a(n35078), .b(n35077), .c(n35076), .o(n35079) );
in01f01 g31289 ( .a(n35079), .o(n35080) );
no02f01 g31290 ( .a(n34741), .b(n5380), .o(n35081) );
no02f01 g31291 ( .a(n35081), .b(n34743), .o(n35082) );
in01f01 g31292 ( .a(n35082), .o(n35083) );
no02f01 g31293 ( .a(n35083), .b(n35080), .o(n35084) );
no02f01 g31294 ( .a(n35082), .b(n35079), .o(n35085) );
no02f01 g31295 ( .a(n35085), .b(n35084), .o(n35086) );
in01f01 g31296 ( .a(n35086), .o(n35087) );
no02f01 g31297 ( .a(n35078), .b(n34751), .o(n35088) );
no02f01 g31298 ( .a(n35088), .b(n34728), .o(n35089) );
na02f01 g31299 ( .a(n35088), .b(n34728), .o(n35090) );
in01f01 g31300 ( .a(n35090), .o(n35091) );
no02f01 g31301 ( .a(n35091), .b(n35089), .o(n35092) );
in01f01 g31302 ( .a(n35092), .o(n35093) );
ao12f01 g31303 ( .a(n34908), .b(n35093), .c(n35087), .o(n35094) );
in01f01 g31304 ( .a(n35094), .o(n35095) );
no02f01 g31305 ( .a(n34753), .b(n34728), .o(n35096) );
in01f01 g31306 ( .a(n35096), .o(n35097) );
no02f01 g31307 ( .a(n34763), .b(n5380), .o(n35098) );
ao12f01 g31308 ( .a(n5380), .b(n34749), .c(n34741), .o(n35099) );
no02f01 g31309 ( .a(n35099), .b(n35098), .o(n35100) );
oa12f01 g31310 ( .a(n35100), .b(n35097), .c(n34765), .o(n35101) );
no02f01 g31311 ( .a(n34774), .b(n5380), .o(n35102) );
no02f01 g31312 ( .a(n35102), .b(n34776), .o(n35103) );
in01f01 g31313 ( .a(n35103), .o(n35104) );
no02f01 g31314 ( .a(n35104), .b(n35101), .o(n35105) );
na02f01 g31315 ( .a(n35104), .b(n35101), .o(n35106) );
in01f01 g31316 ( .a(n35106), .o(n35107) );
no03f01 g31317 ( .a(n35107), .b(n35105), .c(n34908), .o(n35108) );
no02f01 g31318 ( .a(n35098), .b(n34765), .o(n35109) );
in01f01 g31319 ( .a(n35109), .o(n35110) );
no03f01 g31320 ( .a(n35110), .b(n35099), .c(n35096), .o(n35111) );
no02f01 g31321 ( .a(n35099), .b(n35096), .o(n35112) );
no02f01 g31322 ( .a(n35109), .b(n35112), .o(n35113) );
no03f01 g31323 ( .a(n35113), .b(n35111), .c(n34908), .o(n35114) );
no02f01 g31324 ( .a(n35114), .b(n35108), .o(n35115) );
no02f01 g31325 ( .a(n34811), .b(n5380), .o(n35116) );
no02f01 g31326 ( .a(n35116), .b(n34813), .o(n35117) );
in01f01 g31327 ( .a(n35117), .o(n35118) );
no03f01 g31328 ( .a(n35118), .b(n34883), .c(n34779), .o(n35119) );
no02f01 g31329 ( .a(n34883), .b(n34779), .o(n35120) );
no02f01 g31330 ( .a(n35117), .b(n35120), .o(n35121) );
no03f01 g31331 ( .a(n35121), .b(n35119), .c(n34908), .o(n35122) );
in01f01 g31332 ( .a(n34779), .o(n35123) );
no02f01 g31333 ( .a(n34813), .b(n35123), .o(n35124) );
in01f01 g31334 ( .a(n35124), .o(n35125) );
no02f01 g31335 ( .a(n35116), .b(n34883), .o(n35126) );
na02f01 g31336 ( .a(n35126), .b(n35125), .o(n35127) );
no02f01 g31337 ( .a(n34884), .b(n5380), .o(n35128) );
no02f01 g31338 ( .a(n35128), .b(n34806), .o(n35129) );
in01f01 g31339 ( .a(n35129), .o(n35130) );
no02f01 g31340 ( .a(n35130), .b(n35127), .o(n35131) );
na02f01 g31341 ( .a(n35130), .b(n35127), .o(n35132) );
in01f01 g31342 ( .a(n35132), .o(n35133) );
no03f01 g31343 ( .a(n35133), .b(n35131), .c(n34908), .o(n35134) );
no02f01 g31344 ( .a(n35134), .b(n35122), .o(n35135) );
in01f01 g31345 ( .a(n35135), .o(n35136) );
no03f01 g31346 ( .a(n35125), .b(n34806), .c(n34786), .o(n35137) );
no02f01 g31347 ( .a(n34888), .b(n5380), .o(n35138) );
no02f01 g31348 ( .a(n35138), .b(n34887), .o(n35139) );
in01f01 g31349 ( .a(n35139), .o(n35140) );
no02f01 g31350 ( .a(n34889), .b(n5380), .o(n35141) );
no02f01 g31351 ( .a(n35141), .b(n34796), .o(n35142) );
in01f01 g31352 ( .a(n35142), .o(n35143) );
no03f01 g31353 ( .a(n35143), .b(n35140), .c(n35137), .o(n35144) );
no02f01 g31354 ( .a(n35140), .b(n35137), .o(n35145) );
no02f01 g31355 ( .a(n35142), .b(n35145), .o(n35146) );
no03f01 g31356 ( .a(n35146), .b(n35144), .c(n34908), .o(n35147) );
oa12f01 g31357 ( .a(n34886), .b(n35125), .c(n34806), .o(n35148) );
no02f01 g31358 ( .a(n35138), .b(n34786), .o(n35149) );
in01f01 g31359 ( .a(n35149), .o(n35150) );
no02f01 g31360 ( .a(n35150), .b(n35148), .o(n35151) );
na02f01 g31361 ( .a(n35150), .b(n35148), .o(n35152) );
in01f01 g31362 ( .a(n35152), .o(n35153) );
no03f01 g31363 ( .a(n35153), .b(n35151), .c(n34908), .o(n35154) );
no03f01 g31364 ( .a(n35154), .b(n35147), .c(n35136), .o(n35155) );
na04f01 g31365 ( .a(n35155), .b(n35115), .c(n35095), .d(n35075), .o(n35156) );
ao12f01 g31366 ( .a(n5978), .b(n35092), .c(n35086), .o(n35157) );
no02f01 g31367 ( .a(n35107), .b(n35105), .o(n35158) );
no02f01 g31368 ( .a(n35113), .b(n35111), .o(n35159) );
ao12f01 g31369 ( .a(n5978), .b(n35159), .c(n35158), .o(n35160) );
no02f01 g31370 ( .a(n35160), .b(n35157), .o(n35161) );
in01f01 g31371 ( .a(n35161), .o(n35162) );
no02f01 g31372 ( .a(n35121), .b(n35119), .o(n35163) );
no02f01 g31373 ( .a(n35133), .b(n35131), .o(n35164) );
ao12f01 g31374 ( .a(n5978), .b(n35164), .c(n35163), .o(n35165) );
no02f01 g31375 ( .a(n35146), .b(n35144), .o(n35166) );
no02f01 g31376 ( .a(n35153), .b(n35151), .o(n35167) );
ao12f01 g31377 ( .a(n5978), .b(n35167), .c(n35166), .o(n35168) );
no03f01 g31378 ( .a(n35168), .b(n35165), .c(n35162), .o(n35169) );
no02f01 g31379 ( .a(n34897), .b(n5380), .o(n35170) );
in01f01 g31380 ( .a(n35170), .o(n35171) );
in01f01 g31381 ( .a(n34814), .o(n35172) );
no03f01 g31382 ( .a(n34823), .b(n35172), .c(n35123), .o(n35173) );
in01f01 g31383 ( .a(n34844), .o(n35174) );
ao12f01 g31384 ( .a(n34895), .b(n35174), .c(n35173), .o(n35175) );
ao12f01 g31385 ( .a(n34851), .b(n35175), .c(n35171), .o(n35176) );
in01f01 g31386 ( .a(n35176), .o(n35177) );
no02f01 g31387 ( .a(n34896), .b(n5380), .o(n35178) );
no02f01 g31388 ( .a(n35178), .b(n34833), .o(n35179) );
no02f01 g31389 ( .a(n35179), .b(n35177), .o(n35180) );
na02f01 g31390 ( .a(n35179), .b(n35177), .o(n35181) );
in01f01 g31391 ( .a(n35181), .o(n35182) );
no02f01 g31392 ( .a(n35182), .b(n35180), .o(n35183) );
in01f01 g31393 ( .a(n35183), .o(n35184) );
no02f01 g31394 ( .a(n35184), .b(n34908), .o(n35185) );
no02f01 g31395 ( .a(n34821), .b(n5380), .o(n35186) );
no02f01 g31396 ( .a(n35186), .b(n34892), .o(n35187) );
in01f01 g31397 ( .a(n35187), .o(n35188) );
no02f01 g31398 ( .a(n34842), .b(n5380), .o(n35189) );
no02f01 g31399 ( .a(n35189), .b(n34844), .o(n35190) );
in01f01 g31400 ( .a(n35190), .o(n35191) );
no03f01 g31401 ( .a(n35191), .b(n35188), .c(n35173), .o(n35192) );
no02f01 g31402 ( .a(n35188), .b(n35173), .o(n35193) );
no02f01 g31403 ( .a(n35190), .b(n35193), .o(n35194) );
no02f01 g31404 ( .a(n35194), .b(n35192), .o(n35195) );
in01f01 g31405 ( .a(n35195), .o(n35196) );
no02f01 g31406 ( .a(n35172), .b(n35123), .o(n35197) );
no02f01 g31407 ( .a(n35186), .b(n34823), .o(n35198) );
in01f01 g31408 ( .a(n35198), .o(n35199) );
no03f01 g31409 ( .a(n35199), .b(n34892), .c(n35197), .o(n35200) );
no02f01 g31410 ( .a(n34892), .b(n35197), .o(n35201) );
no02f01 g31411 ( .a(n35198), .b(n35201), .o(n35202) );
no02f01 g31412 ( .a(n35202), .b(n35200), .o(n35203) );
in01f01 g31413 ( .a(n35203), .o(n35204) );
ao12f01 g31414 ( .a(n34908), .b(n35204), .c(n35196), .o(n35205) );
in01f01 g31415 ( .a(n35175), .o(n35206) );
no02f01 g31416 ( .a(n35170), .b(n34851), .o(n35207) );
in01f01 g31417 ( .a(n35207), .o(n35208) );
no02f01 g31418 ( .a(n35208), .b(n35206), .o(n35209) );
no02f01 g31419 ( .a(n35207), .b(n35175), .o(n35210) );
no03f01 g31420 ( .a(n35210), .b(n35209), .c(n34908), .o(n35211) );
no03f01 g31421 ( .a(n35211), .b(n35205), .c(n35185), .o(n35212) );
in01f01 g31422 ( .a(n35212), .o(n35213) );
ao12f01 g31423 ( .a(n35213), .b(n35169), .c(n35156), .o(n35214) );
in01f01 g31424 ( .a(n34853), .o(n35215) );
no02f01 g31425 ( .a(n34900), .b(n35215), .o(n35216) );
no02f01 g31426 ( .a(n34903), .b(n5380), .o(n35217) );
in01f01 g31427 ( .a(n35217), .o(n35218) );
ao12f01 g31428 ( .a(n34869), .b(n35218), .c(n35216), .o(n35219) );
no02f01 g31429 ( .a(n34902), .b(n5380), .o(n35220) );
no02f01 g31430 ( .a(n35220), .b(n34863), .o(n35221) );
in01f01 g31431 ( .a(n35221), .o(n35222) );
no02f01 g31432 ( .a(n35222), .b(n35219), .o(n35223) );
na02f01 g31433 ( .a(n35222), .b(n35219), .o(n35224) );
in01f01 g31434 ( .a(n35224), .o(n35225) );
no02f01 g31435 ( .a(n35225), .b(n35223), .o(n35226) );
in01f01 g31436 ( .a(n35226), .o(n35227) );
no02f01 g31437 ( .a(n35217), .b(n34869), .o(n35228) );
no02f01 g31438 ( .a(n35228), .b(n35216), .o(n35229) );
na02f01 g31439 ( .a(n35228), .b(n35216), .o(n35230) );
in01f01 g31440 ( .a(n35230), .o(n35231) );
no02f01 g31441 ( .a(n35231), .b(n35229), .o(n35232) );
in01f01 g31442 ( .a(n35232), .o(n35233) );
ao12f01 g31443 ( .a(n34908), .b(n35233), .c(n35227), .o(n35234) );
no02f01 g31444 ( .a(n34904), .b(n34900), .o(n35235) );
oa12f01 g31445 ( .a(n35235), .b(n34871), .c(n34853), .o(n35236) );
in01f01 g31446 ( .a(n35236), .o(n35237) );
no02f01 g31447 ( .a(n34901), .b(n5380), .o(n35238) );
no02f01 g31448 ( .a(n35238), .b(n34879), .o(n35239) );
no02f01 g31449 ( .a(n35239), .b(n35237), .o(n35240) );
na02f01 g31450 ( .a(n35239), .b(n35237), .o(n35241) );
in01f01 g31451 ( .a(n35241), .o(n35242) );
no03f01 g31452 ( .a(n35242), .b(n35240), .c(n34908), .o(n35243) );
no02f01 g31453 ( .a(n35243), .b(n35234), .o(n35244) );
no02f01 g31454 ( .a(n35242), .b(n35240), .o(n35245) );
ao12f01 g31455 ( .a(n5978), .b(n35232), .c(n35226), .o(n35246) );
in01f01 g31456 ( .a(n35246), .o(n35247) );
ao12f01 g31457 ( .a(n5978), .b(n35247), .c(n35245), .o(n35248) );
ao12f01 g31458 ( .a(n5978), .b(n35203), .c(n35195), .o(n35249) );
in01f01 g31459 ( .a(n35249), .o(n35250) );
no02f01 g31460 ( .a(n35210), .b(n35209), .o(n35251) );
no02f01 g31461 ( .a(n35251), .b(n5978), .o(n35252) );
oa12f01 g31462 ( .a(n34908), .b(n35252), .c(n35184), .o(n35253) );
na02f01 g31463 ( .a(n35253), .b(n35250), .o(n35254) );
no02f01 g31464 ( .a(n35254), .b(n35248), .o(n35255) );
in01f01 g31465 ( .a(n35255), .o(n35256) );
ao12f01 g31466 ( .a(n35256), .b(n35244), .c(n35214), .o(n4176) );
in01f01 g31467 ( .a(n4176), .o(n35258) );
no02f01 g31468 ( .a(n34978), .b(n34935), .o(n35259) );
no02f01 g31469 ( .a(n34975), .b(n34908), .o(n35260) );
in01f01 g31470 ( .a(n35260), .o(n35261) );
na02f01 g31471 ( .a(n35261), .b(n35259), .o(n35262) );
in01f01 g31472 ( .a(n35262), .o(n35263) );
no02f01 g31473 ( .a(n34918), .b(n5978), .o(n35264) );
no02f01 g31474 ( .a(n35264), .b(n34920), .o(n35265) );
no02f01 g31475 ( .a(n35265), .b(n35263), .o(n35266) );
na02f01 g31476 ( .a(n35265), .b(n35263), .o(n35267) );
in01f01 g31477 ( .a(n35267), .o(n35268) );
no02f01 g31478 ( .a(n35268), .b(n35266), .o(n35269) );
in01f01 g31479 ( .a(n35269), .o(n35270) );
no02f01 g31480 ( .a(n35270), .b(n35258), .o(n35271) );
in01f01 g31481 ( .a(n34941), .o(n35272) );
no02f01 g31482 ( .a(n35272), .b(n5978), .o(n35273) );
no03f01 g31483 ( .a(n34942), .b(n35273), .c(n_186), .o(n35274) );
no02f01 g31484 ( .a(n34942), .b(n35273), .o(n35275) );
no02f01 g31485 ( .a(n35275), .b(n34438), .o(n35276) );
no02f01 g31486 ( .a(n35276), .b(n35274), .o(n35277) );
in01f01 g31487 ( .a(n35277), .o(n35278) );
na02f01 g31488 ( .a(n35278), .b(n4176), .o(n35279) );
oa12f01 g31489 ( .a(n34438), .b(n35275), .c(n4176), .o(n35280) );
no02f01 g31490 ( .a(n34949), .b(n5978), .o(n35281) );
no04f01 g31491 ( .a(n34961), .b(n35281), .c(n34942), .d(n34938), .o(n35282) );
no02f01 g31492 ( .a(n34942), .b(n34938), .o(n35283) );
no02f01 g31493 ( .a(n34961), .b(n35281), .o(n35284) );
no02f01 g31494 ( .a(n35284), .b(n35283), .o(n35285) );
no02f01 g31495 ( .a(n35285), .b(n35282), .o(n35286) );
in01f01 g31496 ( .a(n35286), .o(n35287) );
no02f01 g31497 ( .a(n35287), .b(n4176), .o(n35288) );
ao12f01 g31498 ( .a(n35288), .b(n35280), .c(n35279), .o(n35289) );
no02f01 g31499 ( .a(n34961), .b(n34951), .o(n35290) );
no02f01 g31500 ( .a(n34959), .b(n34908), .o(n35291) );
no02f01 g31501 ( .a(n34960), .b(n5978), .o(n35292) );
no02f01 g31502 ( .a(n35292), .b(n35291), .o(n35293) );
no02f01 g31503 ( .a(n35293), .b(n35290), .o(n35294) );
na02f01 g31504 ( .a(n35293), .b(n35290), .o(n35295) );
in01f01 g31505 ( .a(n35295), .o(n35296) );
no02f01 g31506 ( .a(n35296), .b(n35294), .o(n35297) );
in01f01 g31507 ( .a(n35297), .o(n35298) );
na02f01 g31508 ( .a(n35298), .b(n35289), .o(n35299) );
no02f01 g31509 ( .a(n35286), .b(n35258), .o(n35300) );
no03f01 g31510 ( .a(n35300), .b(n35298), .c(n35289), .o(n35301) );
oa12f01 g31511 ( .a(n35299), .b(n35301), .c(n35258), .o(n35302) );
in01f01 g31512 ( .a(n34964), .o(n35303) );
no02f01 g31513 ( .a(n34934), .b(n34908), .o(n35304) );
no02f01 g31514 ( .a(n35304), .b(n34966), .o(n35305) );
in01f01 g31515 ( .a(n35305), .o(n35306) );
no02f01 g31516 ( .a(n35306), .b(n35303), .o(n35307) );
no02f01 g31517 ( .a(n35305), .b(n34964), .o(n35308) );
no02f01 g31518 ( .a(n35308), .b(n35307), .o(n35309) );
in01f01 g31519 ( .a(n35309), .o(n35310) );
no02f01 g31520 ( .a(n35310), .b(n4176), .o(n35311) );
in01f01 g31521 ( .a(n35311), .o(n35312) );
no02f01 g31522 ( .a(n34966), .b(n34964), .o(n35313) );
no02f01 g31523 ( .a(n35304), .b(n35313), .o(n35314) );
no02f01 g31524 ( .a(n34928), .b(n34908), .o(n35315) );
no02f01 g31525 ( .a(n35315), .b(n34968), .o(n35316) );
no02f01 g31526 ( .a(n35316), .b(n35314), .o(n35317) );
na02f01 g31527 ( .a(n35316), .b(n35314), .o(n35318) );
in01f01 g31528 ( .a(n35318), .o(n35319) );
no02f01 g31529 ( .a(n35319), .b(n35317), .o(n35320) );
in01f01 g31530 ( .a(n35320), .o(n35321) );
no02f01 g31531 ( .a(n35321), .b(n4176), .o(n35322) );
in01f01 g31532 ( .a(n35322), .o(n35323) );
na03f01 g31533 ( .a(n35323), .b(n35312), .c(n35302), .o(n35324) );
ao12f01 g31534 ( .a(n35258), .b(n35320), .c(n35309), .o(n35325) );
in01f01 g31535 ( .a(n35325), .o(n35326) );
na02f01 g31536 ( .a(n35326), .b(n35324), .o(n35327) );
no03f01 g31537 ( .a(n34968), .b(n34966), .c(n34964), .o(n35328) );
no02f01 g31538 ( .a(n35260), .b(n34977), .o(n35329) );
in01f01 g31539 ( .a(n35329), .o(n35330) );
no03f01 g31540 ( .a(n35330), .b(n35328), .c(n34935), .o(n35331) );
no02f01 g31541 ( .a(n35328), .b(n34935), .o(n35332) );
no02f01 g31542 ( .a(n35329), .b(n35332), .o(n35333) );
no02f01 g31543 ( .a(n35333), .b(n35331), .o(n35334) );
in01f01 g31544 ( .a(n35334), .o(n35335) );
no02f01 g31545 ( .a(n35335), .b(n35258), .o(n35336) );
in01f01 g31546 ( .a(n35336), .o(n35337) );
ao12f01 g31547 ( .a(n4176), .b(n35334), .c(n35269), .o(n35338) );
ao12f01 g31548 ( .a(n35338), .b(n35337), .c(n35327), .o(n35339) );
no02f01 g31549 ( .a(n34980), .b(n34920), .o(n35340) );
in01f01 g31550 ( .a(n35340), .o(n35341) );
no02f01 g31551 ( .a(n34987), .b(n5978), .o(n35342) );
no02f01 g31552 ( .a(n34988), .b(n34908), .o(n35343) );
no02f01 g31553 ( .a(n35343), .b(n35342), .o(n35344) );
no02f01 g31554 ( .a(n35344), .b(n35341), .o(n35345) );
na02f01 g31555 ( .a(n35344), .b(n35341), .o(n35346) );
in01f01 g31556 ( .a(n35346), .o(n35347) );
no02f01 g31557 ( .a(n35347), .b(n35345), .o(n35348) );
in01f01 g31558 ( .a(n35348), .o(n35349) );
in01f01 g31559 ( .a(n35343), .o(n35350) );
ao12f01 g31560 ( .a(n35342), .b(n35350), .c(n35340), .o(n35351) );
no02f01 g31561 ( .a(n34998), .b(n34908), .o(n35352) );
no02f01 g31562 ( .a(n34997), .b(n5978), .o(n35353) );
no02f01 g31563 ( .a(n35353), .b(n35352), .o(n35354) );
no02f01 g31564 ( .a(n35354), .b(n35351), .o(n35355) );
na02f01 g31565 ( .a(n35354), .b(n35351), .o(n35356) );
in01f01 g31566 ( .a(n35356), .o(n35357) );
no02f01 g31567 ( .a(n35357), .b(n35355), .o(n35358) );
in01f01 g31568 ( .a(n35358), .o(n35359) );
ao12f01 g31569 ( .a(n35258), .b(n35359), .c(n35349), .o(n35360) );
no02f01 g31570 ( .a(n34999), .b(n35341), .o(n35361) );
no02f01 g31571 ( .a(n35019), .b(n5978), .o(n35362) );
no02f01 g31572 ( .a(n35362), .b(n35021), .o(n35363) );
in01f01 g31573 ( .a(n35363), .o(n35364) );
no03f01 g31574 ( .a(n35364), .b(n35025), .c(n35361), .o(n35365) );
no02f01 g31575 ( .a(n35025), .b(n35361), .o(n35366) );
no02f01 g31576 ( .a(n35363), .b(n35366), .o(n35367) );
no02f01 g31577 ( .a(n35367), .b(n35365), .o(n35368) );
in01f01 g31578 ( .a(n35368), .o(n35369) );
no02f01 g31579 ( .a(n35369), .b(n35258), .o(n35370) );
no03f01 g31580 ( .a(n35021), .b(n34999), .c(n35341), .o(n35371) );
no02f01 g31581 ( .a(n35362), .b(n35025), .o(n35372) );
in01f01 g31582 ( .a(n35372), .o(n35373) );
no02f01 g31583 ( .a(n35011), .b(n5978), .o(n35374) );
no02f01 g31584 ( .a(n35374), .b(n35013), .o(n35375) );
in01f01 g31585 ( .a(n35375), .o(n35376) );
no03f01 g31586 ( .a(n35376), .b(n35373), .c(n35371), .o(n35377) );
no02f01 g31587 ( .a(n35373), .b(n35371), .o(n35378) );
no02f01 g31588 ( .a(n35375), .b(n35378), .o(n35379) );
no02f01 g31589 ( .a(n35379), .b(n35377), .o(n35380) );
in01f01 g31590 ( .a(n35380), .o(n35381) );
no02f01 g31591 ( .a(n35381), .b(n35258), .o(n35382) );
no02f01 g31592 ( .a(n35382), .b(n35370), .o(n35383) );
in01f01 g31593 ( .a(n35383), .o(n35384) );
no04f01 g31594 ( .a(n35384), .b(n35360), .c(n35339), .d(n35271), .o(n35385) );
ao12f01 g31595 ( .a(n4176), .b(n35358), .c(n35348), .o(n35386) );
ao12f01 g31596 ( .a(n4176), .b(n35380), .c(n35368), .o(n35387) );
no02f01 g31597 ( .a(n35387), .b(n35386), .o(n35388) );
in01f01 g31598 ( .a(n35388), .o(n35389) );
no02f01 g31599 ( .a(n35028), .b(n35024), .o(n35390) );
in01f01 g31600 ( .a(n35390), .o(n35391) );
no02f01 g31601 ( .a(n35045), .b(n5978), .o(n35392) );
na02f01 g31602 ( .a(n35045), .b(n5978), .o(n35393) );
ao12f01 g31603 ( .a(n35392), .b(n35393), .c(n35391), .o(n35394) );
in01f01 g31604 ( .a(n35038), .o(n35395) );
no02f01 g31605 ( .a(n35395), .b(n34908), .o(n35396) );
no02f01 g31606 ( .a(n35038), .b(n5978), .o(n35397) );
no02f01 g31607 ( .a(n35397), .b(n35396), .o(n35398) );
no02f01 g31608 ( .a(n35398), .b(n35394), .o(n35399) );
na02f01 g31609 ( .a(n35398), .b(n35394), .o(n35400) );
in01f01 g31610 ( .a(n35400), .o(n35401) );
no02f01 g31611 ( .a(n35401), .b(n35399), .o(n35402) );
in01f01 g31612 ( .a(n35402), .o(n35403) );
no02f01 g31613 ( .a(n35403), .b(n35258), .o(n35404) );
in01f01 g31614 ( .a(n35393), .o(n35405) );
no02f01 g31615 ( .a(n35405), .b(n35392), .o(n35406) );
in01f01 g31616 ( .a(n35406), .o(n35407) );
no02f01 g31617 ( .a(n35407), .b(n35391), .o(n35408) );
no02f01 g31618 ( .a(n35406), .b(n35390), .o(n35409) );
no02f01 g31619 ( .a(n35409), .b(n35408), .o(n35410) );
in01f01 g31620 ( .a(n35410), .o(n35411) );
no02f01 g31621 ( .a(n35411), .b(n35258), .o(n35412) );
no02f01 g31622 ( .a(n35412), .b(n35404), .o(n35413) );
oa12f01 g31623 ( .a(n35413), .b(n35389), .c(n35385), .o(n35414) );
no02f01 g31624 ( .a(n35067), .b(n5978), .o(n35415) );
in01f01 g31625 ( .a(n35415), .o(n35416) );
in01f01 g31626 ( .a(n35047), .o(n35417) );
no02f01 g31627 ( .a(n35072), .b(n35417), .o(n35418) );
ao12f01 g31628 ( .a(n35069), .b(n35418), .c(n35416), .o(n35419) );
no02f01 g31629 ( .a(n35059), .b(n5978), .o(n35420) );
no02f01 g31630 ( .a(n35420), .b(n35061), .o(n35421) );
in01f01 g31631 ( .a(n35421), .o(n35422) );
no02f01 g31632 ( .a(n35422), .b(n35419), .o(n35423) );
na02f01 g31633 ( .a(n35422), .b(n35419), .o(n35424) );
in01f01 g31634 ( .a(n35424), .o(n35425) );
no02f01 g31635 ( .a(n35425), .b(n35423), .o(n35426) );
in01f01 g31636 ( .a(n35426), .o(n35427) );
no02f01 g31637 ( .a(n35427), .b(n35258), .o(n35428) );
no02f01 g31638 ( .a(n35415), .b(n35069), .o(n35429) );
in01f01 g31639 ( .a(n35429), .o(n35430) );
no03f01 g31640 ( .a(n35430), .b(n35072), .c(n35417), .o(n35431) );
no02f01 g31641 ( .a(n35429), .b(n35418), .o(n35432) );
no02f01 g31642 ( .a(n35432), .b(n35431), .o(n35433) );
in01f01 g31643 ( .a(n35433), .o(n35434) );
no02f01 g31644 ( .a(n35434), .b(n35258), .o(n35435) );
no02f01 g31645 ( .a(n35435), .b(n35428), .o(n35436) );
in01f01 g31646 ( .a(n35436), .o(n35437) );
ao12f01 g31647 ( .a(n4176), .b(n35433), .c(n35426), .o(n35438) );
ao12f01 g31648 ( .a(n4176), .b(n35410), .c(n35402), .o(n35439) );
no02f01 g31649 ( .a(n35439), .b(n35438), .o(n35440) );
oa12f01 g31650 ( .a(n35440), .b(n35437), .c(n35414), .o(n35441) );
no02f01 g31651 ( .a(n35092), .b(n5978), .o(n35442) );
no02f01 g31652 ( .a(n35093), .b(n34908), .o(n35443) );
in01f01 g31653 ( .a(n35443), .o(n35444) );
ao12f01 g31654 ( .a(n35442), .b(n35444), .c(n35075), .o(n35445) );
in01f01 g31655 ( .a(n35445), .o(n35446) );
no02f01 g31656 ( .a(n35087), .b(n34908), .o(n35447) );
no02f01 g31657 ( .a(n35086), .b(n5978), .o(n35448) );
no02f01 g31658 ( .a(n35448), .b(n35447), .o(n35449) );
in01f01 g31659 ( .a(n35449), .o(n35450) );
no02f01 g31660 ( .a(n35450), .b(n35446), .o(n35451) );
no02f01 g31661 ( .a(n35449), .b(n35445), .o(n35452) );
no02f01 g31662 ( .a(n35452), .b(n35451), .o(n35453) );
in01f01 g31663 ( .a(n35453), .o(n35454) );
no02f01 g31664 ( .a(n35454), .b(n35258), .o(n35455) );
in01f01 g31665 ( .a(n35075), .o(n35456) );
no02f01 g31666 ( .a(n35443), .b(n35442), .o(n35457) );
no02f01 g31667 ( .a(n35457), .b(n35456), .o(n35458) );
na02f01 g31668 ( .a(n35457), .b(n35456), .o(n35459) );
in01f01 g31669 ( .a(n35459), .o(n35460) );
no02f01 g31670 ( .a(n35460), .b(n35458), .o(n35461) );
in01f01 g31671 ( .a(n35461), .o(n35462) );
no02f01 g31672 ( .a(n35462), .b(n35258), .o(n35463) );
no02f01 g31673 ( .a(n35463), .b(n35455), .o(n35464) );
in01f01 g31674 ( .a(n35464), .o(n35465) );
no02f01 g31675 ( .a(n35094), .b(n35456), .o(n35466) );
in01f01 g31676 ( .a(n35466), .o(n35467) );
no02f01 g31677 ( .a(n35159), .b(n5978), .o(n35468) );
no02f01 g31678 ( .a(n35468), .b(n35157), .o(n35469) );
oa12f01 g31679 ( .a(n35469), .b(n35114), .c(n35467), .o(n35470) );
no02f01 g31680 ( .a(n35158), .b(n5978), .o(n35471) );
no02f01 g31681 ( .a(n35471), .b(n35108), .o(n35472) );
in01f01 g31682 ( .a(n35472), .o(n35473) );
no02f01 g31683 ( .a(n35473), .b(n35470), .o(n35474) );
na02f01 g31684 ( .a(n35473), .b(n35470), .o(n35475) );
in01f01 g31685 ( .a(n35475), .o(n35476) );
no03f01 g31686 ( .a(n35476), .b(n35474), .c(n35258), .o(n35477) );
no02f01 g31687 ( .a(n35468), .b(n35114), .o(n35478) );
in01f01 g31688 ( .a(n35478), .o(n35479) );
no03f01 g31689 ( .a(n35479), .b(n35157), .c(n35466), .o(n35480) );
no02f01 g31690 ( .a(n35157), .b(n35466), .o(n35481) );
no02f01 g31691 ( .a(n35478), .b(n35481), .o(n35482) );
no02f01 g31692 ( .a(n35482), .b(n35480), .o(n35483) );
in01f01 g31693 ( .a(n35483), .o(n35484) );
no02f01 g31694 ( .a(n35484), .b(n35258), .o(n35485) );
no03f01 g31695 ( .a(n35485), .b(n35477), .c(n35465), .o(n35486) );
in01f01 g31696 ( .a(n35115), .o(n35487) );
no02f01 g31697 ( .a(n35487), .b(n35467), .o(n35488) );
in01f01 g31698 ( .a(n35488), .o(n35489) );
no02f01 g31699 ( .a(n35163), .b(n5978), .o(n35490) );
no02f01 g31700 ( .a(n35490), .b(n35162), .o(n35491) );
oa12f01 g31701 ( .a(n35491), .b(n35122), .c(n35489), .o(n35492) );
no02f01 g31702 ( .a(n35164), .b(n5978), .o(n35493) );
no02f01 g31703 ( .a(n35493), .b(n35134), .o(n35494) );
in01f01 g31704 ( .a(n35494), .o(n35495) );
no02f01 g31705 ( .a(n35495), .b(n35492), .o(n35496) );
na02f01 g31706 ( .a(n35495), .b(n35492), .o(n35497) );
in01f01 g31707 ( .a(n35497), .o(n35498) );
no03f01 g31708 ( .a(n35498), .b(n35496), .c(n35258), .o(n35499) );
no02f01 g31709 ( .a(n35162), .b(n35488), .o(n35500) );
no02f01 g31710 ( .a(n35490), .b(n35122), .o(n35501) );
no02f01 g31711 ( .a(n35501), .b(n35500), .o(n35502) );
na02f01 g31712 ( .a(n35501), .b(n35500), .o(n35503) );
in01f01 g31713 ( .a(n35503), .o(n35504) );
no02f01 g31714 ( .a(n35504), .b(n35502), .o(n35505) );
in01f01 g31715 ( .a(n35505), .o(n35506) );
no02f01 g31716 ( .a(n35506), .b(n35258), .o(n35507) );
no02f01 g31717 ( .a(n35507), .b(n35499), .o(n35508) );
in01f01 g31718 ( .a(n35508), .o(n35509) );
ao12f01 g31719 ( .a(n35162), .b(n35135), .c(n35488), .o(n35510) );
no02f01 g31720 ( .a(n35167), .b(n5978), .o(n35511) );
no02f01 g31721 ( .a(n35511), .b(n35165), .o(n35512) );
oa12f01 g31722 ( .a(n35512), .b(n35510), .c(n35154), .o(n35513) );
no02f01 g31723 ( .a(n35166), .b(n5978), .o(n35514) );
no02f01 g31724 ( .a(n35514), .b(n35147), .o(n35515) );
in01f01 g31725 ( .a(n35515), .o(n35516) );
no02f01 g31726 ( .a(n35516), .b(n35513), .o(n35517) );
na02f01 g31727 ( .a(n35516), .b(n35513), .o(n35518) );
in01f01 g31728 ( .a(n35518), .o(n35519) );
no03f01 g31729 ( .a(n35519), .b(n35517), .c(n35258), .o(n35520) );
in01f01 g31730 ( .a(n35510), .o(n35521) );
no02f01 g31731 ( .a(n35511), .b(n35154), .o(n35522) );
in01f01 g31732 ( .a(n35522), .o(n35523) );
no03f01 g31733 ( .a(n35523), .b(n35521), .c(n35165), .o(n35524) );
in01f01 g31734 ( .a(n35165), .o(n35525) );
ao12f01 g31735 ( .a(n35522), .b(n35510), .c(n35525), .o(n35526) );
no02f01 g31736 ( .a(n35526), .b(n35524), .o(n35527) );
in01f01 g31737 ( .a(n35527), .o(n35528) );
no02f01 g31738 ( .a(n35528), .b(n35258), .o(n35529) );
no03f01 g31739 ( .a(n35529), .b(n35520), .c(n35509), .o(n35530) );
na03f01 g31740 ( .a(n35530), .b(n35486), .c(n35441), .o(n35531) );
in01f01 g31741 ( .a(n35530), .o(n35532) );
no02f01 g31742 ( .a(n35476), .b(n35474), .o(n35533) );
ao12f01 g31743 ( .a(n4176), .b(n35483), .c(n35533), .o(n35534) );
ao12f01 g31744 ( .a(n4176), .b(n35461), .c(n35453), .o(n35535) );
no02f01 g31745 ( .a(n35535), .b(n35534), .o(n35536) );
no02f01 g31746 ( .a(n35498), .b(n35496), .o(n35537) );
ao12f01 g31747 ( .a(n4176), .b(n35505), .c(n35537), .o(n35538) );
no02f01 g31748 ( .a(n35519), .b(n35517), .o(n35539) );
ao12f01 g31749 ( .a(n4176), .b(n35527), .c(n35539), .o(n35540) );
no02f01 g31750 ( .a(n35540), .b(n35538), .o(n35541) );
oa12f01 g31751 ( .a(n35541), .b(n35536), .c(n35532), .o(n35542) );
in01f01 g31752 ( .a(n35542), .o(n35543) );
na02f01 g31753 ( .a(n35543), .b(n35531), .o(n35544) );
in01f01 g31754 ( .a(n35544), .o(n35545) );
in01f01 g31755 ( .a(n35156), .o(n35546) );
in01f01 g31756 ( .a(n35169), .o(n35547) );
no02f01 g31757 ( .a(n35547), .b(n35546), .o(n35548) );
no02f01 g31758 ( .a(n35203), .b(n5978), .o(n35549) );
no02f01 g31759 ( .a(n35204), .b(n34908), .o(n35550) );
no02f01 g31760 ( .a(n35550), .b(n35549), .o(n35551) );
no02f01 g31761 ( .a(n35551), .b(n35548), .o(n35552) );
na02f01 g31762 ( .a(n35551), .b(n35548), .o(n35553) );
in01f01 g31763 ( .a(n35553), .o(n35554) );
no02f01 g31764 ( .a(n35554), .b(n35552), .o(n35555) );
in01f01 g31765 ( .a(n35555), .o(n35556) );
no02f01 g31766 ( .a(n35556), .b(n35258), .o(n35557) );
no02f01 g31767 ( .a(n35555), .b(n4176), .o(n35558) );
no02f01 g31768 ( .a(n35558), .b(n35557), .o(n35559) );
na02f01 g31769 ( .a(n35559), .b(n35545), .o(n35560) );
in01f01 g31770 ( .a(n35559), .o(n35561) );
na02f01 g31771 ( .a(n35561), .b(n35544), .o(n35562) );
na02f01 g31772 ( .a(n35562), .b(n35560), .o(n437) );
no02f01 g31773 ( .a(n9634), .b(n9268), .o(n35564) );
in01f01 g31774 ( .a(n35564), .o(n35565) );
na02f01 g31775 ( .a(n35565), .b(n9431), .o(n35566) );
na02f01 g31776 ( .a(n35564), .b(n9633), .o(n35567) );
na02f01 g31777 ( .a(n35567), .b(n35566), .o(n442) );
no02f01 g31778 ( .a(n11817), .b(n11535), .o(n35569) );
no02f01 g31779 ( .a(n11841), .b(n11828), .o(n35570) );
in01f01 g31780 ( .a(n35570), .o(n35571) );
na02f01 g31781 ( .a(n35571), .b(n35569), .o(n35572) );
oa12f01 g31782 ( .a(n35570), .b(n11817), .c(n11535), .o(n35573) );
na02f01 g31783 ( .a(n35573), .b(n35572), .o(n447) );
no02f01 g31784 ( .a(n9621), .b(n9620), .o(n35575) );
in01f01 g31785 ( .a(n35575), .o(n35576) );
in01f01 g31786 ( .a(n9381), .o(n35577) );
ao12f01 g31787 ( .a(n9398), .b(n35577), .c(n35576), .o(n35578) );
in01f01 g31788 ( .a(n35578), .o(n35579) );
no02f01 g31789 ( .a(n9399), .b(n9394), .o(n35580) );
in01f01 g31790 ( .a(n35580), .o(n35581) );
na02f01 g31791 ( .a(n35581), .b(n35579), .o(n35582) );
na02f01 g31792 ( .a(n35580), .b(n35578), .o(n35583) );
na02f01 g31793 ( .a(n35583), .b(n35582), .o(n457) );
na03f01 g31794 ( .a(n32712), .b(n32641), .c(n32707), .o(n35585) );
oa12f01 g31795 ( .a(n32663), .b(n32708), .c(n32640), .o(n35586) );
na02f01 g31796 ( .a(n35586), .b(n35585), .o(n462) );
no02f01 g31797 ( .a(n9453), .b(n9225), .o(n35588) );
no02f01 g31798 ( .a(n9454), .b(n9224), .o(n35589) );
no02f01 g31799 ( .a(n35589), .b(n35588), .o(n35590) );
na02f01 g31800 ( .a(n35590), .b(n9636), .o(n35591) );
in01f01 g31801 ( .a(n35590), .o(n35592) );
na02f01 g31802 ( .a(n35592), .b(n9436), .o(n35593) );
na02f01 g31803 ( .a(n35593), .b(n35591), .o(n467) );
na02f01 g31804 ( .a(n32732), .b(cos_out_4), .o(n35595) );
no02f01 g31805 ( .a(n34336), .b(n33493), .o(n35596) );
no02f01 g31806 ( .a(n34287), .b(n33489), .o(n35597) );
no02f01 g31807 ( .a(n35597), .b(n35596), .o(n35598) );
no02f01 g31808 ( .a(n33130), .b(n33048), .o(n35599) );
no02f01 g31809 ( .a(n33131), .b(n32928), .o(n35600) );
in01f01 g31810 ( .a(n35600), .o(n35601) );
ao12f01 g31811 ( .a(n35599), .b(n35601), .c(n33089), .o(n35602) );
no02f01 g31812 ( .a(n33124), .b(n32928), .o(n35603) );
no02f01 g31813 ( .a(n33123), .b(n33048), .o(n35604) );
no02f01 g31814 ( .a(n35604), .b(n35603), .o(n35605) );
no02f01 g31815 ( .a(n35605), .b(n35602), .o(n35606) );
na02f01 g31816 ( .a(n35605), .b(n35602), .o(n35607) );
in01f01 g31817 ( .a(n35607), .o(n35608) );
no02f01 g31818 ( .a(n35608), .b(n35606), .o(n35609) );
in01f01 g31819 ( .a(n35609), .o(n35610) );
no02f01 g31820 ( .a(n35600), .b(n35599), .o(n35611) );
in01f01 g31821 ( .a(n35611), .o(n35612) );
no02f01 g31822 ( .a(n35612), .b(n33089), .o(n35613) );
in01f01 g31823 ( .a(n33089), .o(n35614) );
no02f01 g31824 ( .a(n35611), .b(n35614), .o(n35615) );
no02f01 g31825 ( .a(n35615), .b(n35613), .o(n35616) );
in01f01 g31826 ( .a(n35616), .o(n35617) );
ao12f01 g31827 ( .a(n34336), .b(n35617), .c(n35610), .o(n35618) );
no02f01 g31828 ( .a(n33079), .b(n33048), .o(n35619) );
no02f01 g31829 ( .a(n33087), .b(n35619), .o(n35620) );
na02f01 g31830 ( .a(n35620), .b(n33085), .o(n35621) );
no02f01 g31831 ( .a(n32999), .b(n33048), .o(n35622) );
no02f01 g31832 ( .a(n35622), .b(n33001), .o(n35623) );
in01f01 g31833 ( .a(n35623), .o(n35624) );
no02f01 g31834 ( .a(n35624), .b(n35621), .o(n35625) );
na02f01 g31835 ( .a(n35624), .b(n35621), .o(n35626) );
in01f01 g31836 ( .a(n35626), .o(n35627) );
no02f01 g31837 ( .a(n35627), .b(n35625), .o(n35628) );
in01f01 g31838 ( .a(n35628), .o(n35629) );
no02f01 g31839 ( .a(n35629), .b(n34336), .o(n35630) );
no02f01 g31840 ( .a(n33073), .b(n33052), .o(n35631) );
no02f01 g31841 ( .a(n35619), .b(n33081), .o(n35632) );
in01f01 g31842 ( .a(n35632), .o(n35633) );
no03f01 g31843 ( .a(n35633), .b(n35631), .c(n33087), .o(n35634) );
no02f01 g31844 ( .a(n35631), .b(n33087), .o(n35635) );
no02f01 g31845 ( .a(n35632), .b(n35635), .o(n35636) );
no02f01 g31846 ( .a(n35636), .b(n35634), .o(n35637) );
na02f01 g31847 ( .a(n35637), .b(n34287), .o(n35638) );
na02f01 g31848 ( .a(n35638), .b(n34383), .o(n35639) );
in01f01 g31849 ( .a(n35639), .o(n35640) );
na02f01 g31850 ( .a(n34382), .b(n34359), .o(n35641) );
na02f01 g31851 ( .a(n35641), .b(n34336), .o(n35642) );
in01f01 g31852 ( .a(n35642), .o(n35643) );
ao12f01 g31853 ( .a(n34287), .b(n35637), .c(n35628), .o(n35644) );
no02f01 g31854 ( .a(n35644), .b(n35643), .o(n35645) );
in01f01 g31855 ( .a(n35645), .o(n35646) );
ao12f01 g31856 ( .a(n35646), .b(n35640), .c(n34372), .o(n35647) );
no02f01 g31857 ( .a(n33132), .b(n35614), .o(n35648) );
in01f01 g31858 ( .a(n35648), .o(n35649) );
no02f01 g31859 ( .a(n33139), .b(n33048), .o(n35650) );
no02f01 g31860 ( .a(n33145), .b(n35650), .o(n35651) );
oa12f01 g31861 ( .a(n35651), .b(n35649), .c(n33141), .o(n35652) );
in01f01 g31862 ( .a(n35652), .o(n35653) );
no02f01 g31863 ( .a(n33110), .b(n33048), .o(n35654) );
no02f01 g31864 ( .a(n35654), .b(n33112), .o(n35655) );
no02f01 g31865 ( .a(n35655), .b(n35653), .o(n35656) );
na02f01 g31866 ( .a(n35655), .b(n35653), .o(n35657) );
in01f01 g31867 ( .a(n35657), .o(n35658) );
no02f01 g31868 ( .a(n35658), .b(n35656), .o(n35659) );
in01f01 g31869 ( .a(n35659), .o(n35660) );
no02f01 g31870 ( .a(n35660), .b(n34336), .o(n35661) );
no02f01 g31871 ( .a(n35648), .b(n33145), .o(n35662) );
no02f01 g31872 ( .a(n35650), .b(n33141), .o(n35663) );
no02f01 g31873 ( .a(n35663), .b(n35662), .o(n35664) );
na02f01 g31874 ( .a(n35663), .b(n35662), .o(n35665) );
in01f01 g31875 ( .a(n35665), .o(n35666) );
no02f01 g31876 ( .a(n35666), .b(n35664), .o(n35667) );
in01f01 g31877 ( .a(n35667), .o(n35668) );
no02f01 g31878 ( .a(n35668), .b(n34336), .o(n35669) );
no02f01 g31879 ( .a(n35669), .b(n35661), .o(n35670) );
in01f01 g31880 ( .a(n35670), .o(n35671) );
no04f01 g31881 ( .a(n35671), .b(n35647), .c(n35630), .d(n35618), .o(n35672) );
ao12f01 g31882 ( .a(n34287), .b(n35616), .c(n35609), .o(n35673) );
ao12f01 g31883 ( .a(n34287), .b(n35667), .c(n35659), .o(n35674) );
no02f01 g31884 ( .a(n35674), .b(n35673), .o(n35675) );
in01f01 g31885 ( .a(n35675), .o(n35676) );
no03f01 g31886 ( .a(n33213), .b(n33145), .c(n33144), .o(n35677) );
oa12f01 g31887 ( .a(n35677), .b(n33179), .c(n33143), .o(n35678) );
no02f01 g31888 ( .a(n33194), .b(n33048), .o(n35679) );
no02f01 g31889 ( .a(n35679), .b(n33196), .o(n35680) );
in01f01 g31890 ( .a(n35680), .o(n35681) );
no02f01 g31891 ( .a(n35681), .b(n35678), .o(n35682) );
in01f01 g31892 ( .a(n35678), .o(n35683) );
no02f01 g31893 ( .a(n35680), .b(n35683), .o(n35684) );
no02f01 g31894 ( .a(n35684), .b(n35682), .o(n35685) );
in01f01 g31895 ( .a(n35685), .o(n35686) );
no02f01 g31896 ( .a(n35686), .b(n34336), .o(n35687) );
in01f01 g31897 ( .a(n33177), .o(n35688) );
no02f01 g31898 ( .a(n33175), .b(n33048), .o(n35689) );
ao12f01 g31899 ( .a(n35689), .b(n35688), .c(n33147), .o(n35690) );
no02f01 g31900 ( .a(n33168), .b(n33048), .o(n35691) );
no02f01 g31901 ( .a(n35691), .b(n33170), .o(n35692) );
no02f01 g31902 ( .a(n35692), .b(n35690), .o(n35693) );
na02f01 g31903 ( .a(n35692), .b(n35690), .o(n35694) );
in01f01 g31904 ( .a(n35694), .o(n35695) );
no02f01 g31905 ( .a(n35695), .b(n35693), .o(n35696) );
no02f01 g31906 ( .a(n35689), .b(n33177), .o(n35697) );
in01f01 g31907 ( .a(n35697), .o(n35698) );
no02f01 g31908 ( .a(n35698), .b(n33147), .o(n35699) );
na02f01 g31909 ( .a(n35698), .b(n33147), .o(n35700) );
in01f01 g31910 ( .a(n35700), .o(n35701) );
no02f01 g31911 ( .a(n35701), .b(n35699), .o(n35702) );
no02f01 g31912 ( .a(n35702), .b(n35696), .o(n35703) );
no02f01 g31913 ( .a(n35703), .b(n34336), .o(n35704) );
no02f01 g31914 ( .a(n35678), .b(n35679), .o(n35705) );
no02f01 g31915 ( .a(n35705), .b(n33196), .o(n35706) );
in01f01 g31916 ( .a(n35706), .o(n35707) );
no02f01 g31917 ( .a(n33209), .b(n33048), .o(n35708) );
no02f01 g31918 ( .a(n35708), .b(n33211), .o(n35709) );
no02f01 g31919 ( .a(n35709), .b(n35707), .o(n35710) );
na02f01 g31920 ( .a(n35709), .b(n35707), .o(n35711) );
in01f01 g31921 ( .a(n35711), .o(n35712) );
no02f01 g31922 ( .a(n35712), .b(n35710), .o(n35713) );
in01f01 g31923 ( .a(n35713), .o(n35714) );
no02f01 g31924 ( .a(n35714), .b(n34336), .o(n35715) );
no03f01 g31925 ( .a(n35715), .b(n35704), .c(n35687), .o(n35716) );
oa12f01 g31926 ( .a(n35716), .b(n35676), .c(n35672), .o(n35717) );
ao12f01 g31927 ( .a(n34287), .b(n35702), .c(n35696), .o(n35718) );
ao12f01 g31928 ( .a(n34287), .b(n35713), .c(n35685), .o(n35719) );
no02f01 g31929 ( .a(n35719), .b(n35718), .o(n35720) );
no02f01 g31930 ( .a(n33262), .b(n33217), .o(n35721) );
in01f01 g31931 ( .a(n35721), .o(n35722) );
no02f01 g31932 ( .a(n35722), .b(n33319), .o(n35723) );
no02f01 g31933 ( .a(n33334), .b(n33048), .o(n35724) );
no02f01 g31934 ( .a(n35724), .b(n33336), .o(n35725) );
in01f01 g31935 ( .a(n35725), .o(n35726) );
no03f01 g31936 ( .a(n35726), .b(n35723), .c(n33340), .o(n35727) );
no02f01 g31937 ( .a(n35723), .b(n33340), .o(n35728) );
no02f01 g31938 ( .a(n35725), .b(n35728), .o(n35729) );
no02f01 g31939 ( .a(n35729), .b(n35727), .o(n35730) );
in01f01 g31940 ( .a(n35730), .o(n35731) );
no02f01 g31941 ( .a(n35731), .b(n34336), .o(n35732) );
in01f01 g31942 ( .a(n35732), .o(n35733) );
no03f01 g31943 ( .a(n35722), .b(n33336), .c(n33319), .o(n35734) );
in01f01 g31944 ( .a(n35734), .o(n35735) );
no02f01 g31945 ( .a(n35724), .b(n33340), .o(n35736) );
na02f01 g31946 ( .a(n35736), .b(n35735), .o(n35737) );
no02f01 g31947 ( .a(n33305), .b(n33048), .o(n35738) );
no02f01 g31948 ( .a(n35738), .b(n33307), .o(n35739) );
in01f01 g31949 ( .a(n35739), .o(n35740) );
no02f01 g31950 ( .a(n35740), .b(n35737), .o(n35741) );
na02f01 g31951 ( .a(n35740), .b(n35737), .o(n35742) );
in01f01 g31952 ( .a(n35742), .o(n35743) );
no02f01 g31953 ( .a(n35743), .b(n35741), .o(n35744) );
in01f01 g31954 ( .a(n35744), .o(n35745) );
no02f01 g31955 ( .a(n35745), .b(n34336), .o(n35746) );
no02f01 g31956 ( .a(n33260), .b(n33048), .o(n35747) );
no02f01 g31957 ( .a(n35747), .b(n35721), .o(n35748) );
no02f01 g31958 ( .a(n33317), .b(n33048), .o(n35749) );
no02f01 g31959 ( .a(n35749), .b(n33319), .o(n35750) );
no02f01 g31960 ( .a(n35750), .b(n35748), .o(n35751) );
na02f01 g31961 ( .a(n35750), .b(n35748), .o(n35752) );
in01f01 g31962 ( .a(n35752), .o(n35753) );
no02f01 g31963 ( .a(n35753), .b(n35751), .o(n35754) );
in01f01 g31964 ( .a(n35754), .o(n35755) );
in01f01 g31965 ( .a(n33217), .o(n35756) );
no02f01 g31966 ( .a(n35747), .b(n33262), .o(n35757) );
in01f01 g31967 ( .a(n35757), .o(n35758) );
no02f01 g31968 ( .a(n35758), .b(n35756), .o(n35759) );
no02f01 g31969 ( .a(n35757), .b(n33217), .o(n35760) );
no02f01 g31970 ( .a(n35760), .b(n35759), .o(n35761) );
in01f01 g31971 ( .a(n35761), .o(n35762) );
ao12f01 g31972 ( .a(n34336), .b(n35762), .c(n35755), .o(n35763) );
no02f01 g31973 ( .a(n35763), .b(n35746), .o(n35764) );
na02f01 g31974 ( .a(n35764), .b(n35733), .o(n35765) );
no02f01 g31975 ( .a(n33341), .b(n33340), .o(n35766) );
oa12f01 g31976 ( .a(n35766), .b(n35735), .c(n33307), .o(n35767) );
in01f01 g31977 ( .a(n35767), .o(n35768) );
no03f01 g31978 ( .a(n35768), .b(n33328), .c(n33252), .o(n35769) );
no02f01 g31979 ( .a(n33277), .b(n33048), .o(n35770) );
no02f01 g31980 ( .a(n35770), .b(n33279), .o(n35771) );
in01f01 g31981 ( .a(n35771), .o(n35772) );
no03f01 g31982 ( .a(n35772), .b(n35769), .c(n33343), .o(n35773) );
no02f01 g31983 ( .a(n35769), .b(n33343), .o(n35774) );
no02f01 g31984 ( .a(n35771), .b(n35774), .o(n35775) );
no02f01 g31985 ( .a(n35775), .b(n35773), .o(n35776) );
in01f01 g31986 ( .a(n35776), .o(n35777) );
no02f01 g31987 ( .a(n35777), .b(n34336), .o(n35778) );
in01f01 g31988 ( .a(n35770), .o(n35779) );
ao12f01 g31989 ( .a(n33279), .b(n35774), .c(n35779), .o(n35780) );
in01f01 g31990 ( .a(n35780), .o(n35781) );
no02f01 g31991 ( .a(n33292), .b(n33048), .o(n35782) );
no02f01 g31992 ( .a(n35782), .b(n33294), .o(n35783) );
no02f01 g31993 ( .a(n35783), .b(n35781), .o(n35784) );
na02f01 g31994 ( .a(n35783), .b(n35781), .o(n35785) );
in01f01 g31995 ( .a(n35785), .o(n35786) );
no03f01 g31996 ( .a(n35786), .b(n35784), .c(n34336), .o(n35787) );
in01f01 g31997 ( .a(n33328), .o(n35788) );
no02f01 g31998 ( .a(n33326), .b(n33048), .o(n35789) );
ao12f01 g31999 ( .a(n35789), .b(n35767), .c(n35788), .o(n35790) );
in01f01 g32000 ( .a(n35790), .o(n35791) );
no02f01 g32001 ( .a(n33250), .b(n33048), .o(n35792) );
no02f01 g32002 ( .a(n35792), .b(n33252), .o(n35793) );
in01f01 g32003 ( .a(n35793), .o(n35794) );
no02f01 g32004 ( .a(n35794), .b(n35791), .o(n35795) );
no02f01 g32005 ( .a(n35793), .b(n35790), .o(n35796) );
no02f01 g32006 ( .a(n35796), .b(n35795), .o(n35797) );
no02f01 g32007 ( .a(n35789), .b(n33328), .o(n35798) );
no02f01 g32008 ( .a(n35798), .b(n35768), .o(n35799) );
na02f01 g32009 ( .a(n35798), .b(n35768), .o(n35800) );
in01f01 g32010 ( .a(n35800), .o(n35801) );
no02f01 g32011 ( .a(n35801), .b(n35799), .o(n35802) );
no02f01 g32012 ( .a(n35802), .b(n35797), .o(n35803) );
no02f01 g32013 ( .a(n35803), .b(n34336), .o(n35804) );
no04f01 g32014 ( .a(n35804), .b(n35787), .c(n35778), .d(n35765), .o(n35805) );
in01f01 g32015 ( .a(n35805), .o(n35806) );
ao12f01 g32016 ( .a(n35806), .b(n35720), .c(n35717), .o(n35807) );
ao12f01 g32017 ( .a(n34287), .b(n35761), .c(n35754), .o(n35808) );
ao12f01 g32018 ( .a(n34287), .b(n35744), .c(n35730), .o(n35809) );
no02f01 g32019 ( .a(n35809), .b(n35808), .o(n35810) );
no02f01 g32020 ( .a(n35797), .b(n34287), .o(n35811) );
no02f01 g32021 ( .a(n35802), .b(n34287), .o(n35812) );
no02f01 g32022 ( .a(n35812), .b(n35811), .o(n35813) );
na02f01 g32023 ( .a(n35813), .b(n35810), .o(n35814) );
no02f01 g32024 ( .a(n35786), .b(n35784), .o(n35815) );
ao12f01 g32025 ( .a(n34287), .b(n35815), .c(n35776), .o(n35816) );
no02f01 g32026 ( .a(n35816), .b(n35814), .o(n35817) );
in01f01 g32027 ( .a(n35817), .o(n35818) );
ao12f01 g32028 ( .a(n33458), .b(n33378), .c(n33347), .o(n35819) );
in01f01 g32029 ( .a(n35819), .o(n35820) );
no02f01 g32030 ( .a(n33406), .b(n33048), .o(n35821) );
no02f01 g32031 ( .a(n35821), .b(n33408), .o(n35822) );
in01f01 g32032 ( .a(n35822), .o(n35823) );
no02f01 g32033 ( .a(n35823), .b(n35820), .o(n35824) );
no02f01 g32034 ( .a(n35822), .b(n35819), .o(n35825) );
no02f01 g32035 ( .a(n35825), .b(n35824), .o(n35826) );
in01f01 g32036 ( .a(n35826), .o(n35827) );
no02f01 g32037 ( .a(n35827), .b(n34336), .o(n35828) );
in01f01 g32038 ( .a(n35828), .o(n35829) );
in01f01 g32039 ( .a(n33364), .o(n35830) );
no02f01 g32040 ( .a(n33362), .b(n33048), .o(n35831) );
ao12f01 g32041 ( .a(n35831), .b(n35830), .c(n33347), .o(n35832) );
in01f01 g32042 ( .a(n35832), .o(n35833) );
no02f01 g32043 ( .a(n33375), .b(n33048), .o(n35834) );
no02f01 g32044 ( .a(n35834), .b(n33377), .o(n35835) );
in01f01 g32045 ( .a(n35835), .o(n35836) );
no02f01 g32046 ( .a(n35836), .b(n35833), .o(n35837) );
no02f01 g32047 ( .a(n35835), .b(n35832), .o(n35838) );
no02f01 g32048 ( .a(n35838), .b(n35837), .o(n35839) );
in01f01 g32049 ( .a(n35839), .o(n35840) );
no02f01 g32050 ( .a(n35831), .b(n33364), .o(n35841) );
no02f01 g32051 ( .a(n35841), .b(n33346), .o(n35842) );
na02f01 g32052 ( .a(n35841), .b(n33346), .o(n35843) );
in01f01 g32053 ( .a(n35843), .o(n35844) );
no02f01 g32054 ( .a(n35844), .b(n35842), .o(n35845) );
in01f01 g32055 ( .a(n35845), .o(n35846) );
ao12f01 g32056 ( .a(n34336), .b(n35846), .c(n35840), .o(n35847) );
in01f01 g32057 ( .a(n35821), .o(n35848) );
ao12f01 g32058 ( .a(n33408), .b(n35819), .c(n35848), .o(n35849) );
no02f01 g32059 ( .a(n33397), .b(n33048), .o(n35850) );
no02f01 g32060 ( .a(n35850), .b(n33399), .o(n35851) );
in01f01 g32061 ( .a(n35851), .o(n35852) );
no02f01 g32062 ( .a(n35852), .b(n35849), .o(n35853) );
na02f01 g32063 ( .a(n35852), .b(n35849), .o(n35854) );
in01f01 g32064 ( .a(n35854), .o(n35855) );
no02f01 g32065 ( .a(n35855), .b(n35853), .o(n35856) );
in01f01 g32066 ( .a(n35856), .o(n35857) );
no02f01 g32067 ( .a(n35857), .b(n34336), .o(n35858) );
no02f01 g32068 ( .a(n35858), .b(n35847), .o(n35859) );
na02f01 g32069 ( .a(n35859), .b(n35829), .o(n35860) );
no02f01 g32070 ( .a(n33440), .b(n33048), .o(n35861) );
in01f01 g32071 ( .a(n35861), .o(n35862) );
ao12f01 g32072 ( .a(n33442), .b(n33500), .c(n35862), .o(n35863) );
in01f01 g32073 ( .a(n35863), .o(n35864) );
no02f01 g32074 ( .a(n33464), .b(n33048), .o(n35865) );
no02f01 g32075 ( .a(n35865), .b(n33452), .o(n35866) );
no02f01 g32076 ( .a(n35866), .b(n35864), .o(n35867) );
na02f01 g32077 ( .a(n35866), .b(n35864), .o(n35868) );
in01f01 g32078 ( .a(n35868), .o(n35869) );
no02f01 g32079 ( .a(n35869), .b(n35867), .o(n35870) );
in01f01 g32080 ( .a(n35870), .o(n35871) );
no02f01 g32081 ( .a(n35861), .b(n33442), .o(n35872) );
in01f01 g32082 ( .a(n35872), .o(n35873) );
no03f01 g32083 ( .a(n35873), .b(n33499), .c(n33497), .o(n35874) );
no02f01 g32084 ( .a(n35872), .b(n33500), .o(n35875) );
no02f01 g32085 ( .a(n35875), .b(n35874), .o(n35876) );
in01f01 g32086 ( .a(n35876), .o(n35877) );
ao12f01 g32087 ( .a(n34336), .b(n35877), .c(n35871), .o(n35878) );
no02f01 g32088 ( .a(n34336), .b(n34047), .o(n35879) );
no03f01 g32089 ( .a(n35879), .b(n35878), .c(n35860), .o(n35880) );
oa12f01 g32090 ( .a(n35880), .b(n35818), .c(n35807), .o(n35881) );
no02f01 g32091 ( .a(n35877), .b(n35871), .o(n35882) );
ao12f01 g32092 ( .a(n34287), .b(n35882), .c(n33506), .o(n35883) );
no02f01 g32093 ( .a(n35826), .b(n34287), .o(n35884) );
in01f01 g32094 ( .a(n35884), .o(n35885) );
ao12f01 g32095 ( .a(n34287), .b(n35845), .c(n35839), .o(n35886) );
no02f01 g32096 ( .a(n35856), .b(n34287), .o(n35887) );
no02f01 g32097 ( .a(n35887), .b(n35886), .o(n35888) );
na02f01 g32098 ( .a(n35888), .b(n35885), .o(n35889) );
no02f01 g32099 ( .a(n35889), .b(n35883), .o(n35890) );
na03f01 g32100 ( .a(n35890), .b(n35881), .c(n35598), .o(n35891) );
in01f01 g32101 ( .a(n35598), .o(n35892) );
in01f01 g32102 ( .a(n35618), .o(n35893) );
in01f01 g32103 ( .a(n35630), .o(n35894) );
oa12f01 g32104 ( .a(n34314), .b(n34313), .c(n34311), .o(n35895) );
ao12f01 g32105 ( .a(n34349), .b(n34294), .c(n35895), .o(n35896) );
na02f01 g32106 ( .a(n34337), .b(n34329), .o(n35897) );
oa12f01 g32107 ( .a(n35897), .b(n35896), .c(n34287), .o(n35898) );
in01f01 g32108 ( .a(n34362), .o(n35899) );
na03f01 g32109 ( .a(n35640), .b(n35899), .c(n35898), .o(n35900) );
na02f01 g32110 ( .a(n35645), .b(n35900), .o(n35901) );
na04f01 g32111 ( .a(n35670), .b(n35901), .c(n35894), .d(n35893), .o(n35902) );
in01f01 g32112 ( .a(n35716), .o(n35903) );
ao12f01 g32113 ( .a(n35903), .b(n35675), .c(n35902), .o(n35904) );
in01f01 g32114 ( .a(n35720), .o(n35905) );
oa12f01 g32115 ( .a(n35805), .b(n35905), .c(n35904), .o(n35906) );
in01f01 g32116 ( .a(n35880), .o(n35907) );
ao12f01 g32117 ( .a(n35907), .b(n35817), .c(n35906), .o(n35908) );
in01f01 g32118 ( .a(n35890), .o(n35909) );
oa12f01 g32119 ( .a(n35892), .b(n35909), .c(n35908), .o(n35910) );
na02f01 g32120 ( .a(n35910), .b(n35891), .o(n35911) );
na02f01 g32121 ( .a(n35911), .b(n34304), .o(n35912) );
in01f01 g32122 ( .a(n34055), .o(n35913) );
no02f01 g32123 ( .a(n35913), .b(n34046), .o(n35914) );
no02f01 g32124 ( .a(n35914), .b(n34054), .o(n35915) );
na02f01 g32125 ( .a(n35914), .b(n34054), .o(n35916) );
in01f01 g32126 ( .a(n35916), .o(n35917) );
no02f01 g32127 ( .a(n35917), .b(n35915), .o(n35918) );
in01f01 g32128 ( .a(n35918), .o(n35919) );
na02f01 g32129 ( .a(n35919), .b(n35912), .o(n35920) );
no03f01 g32130 ( .a(n35909), .b(n35908), .c(n35892), .o(n35921) );
ao12f01 g32131 ( .a(n35598), .b(n35890), .c(n35881), .o(n35922) );
no03f01 g32132 ( .a(n35922), .b(n35921), .c(delay_sub_ln23_0_unr30_stage10_stallmux_q), .o(n35923) );
no03f01 g32133 ( .a(n35922), .b(n35921), .c(n34304), .o(n35924) );
no02f01 g32134 ( .a(n34049), .b(n34048), .o(n35925) );
no02f01 g32135 ( .a(n34053), .b(n35925), .o(n35926) );
na02f01 g32136 ( .a(n34053), .b(n35925), .o(n35927) );
in01f01 g32137 ( .a(n35927), .o(n35928) );
no02f01 g32138 ( .a(n35928), .b(n35926), .o(n35929) );
no03f01 g32139 ( .a(n35929), .b(n35924), .c(n35923), .o(n35930) );
no02f01 g32140 ( .a(n35922), .b(n35921), .o(n35931) );
no03f01 g32141 ( .a(n35919), .b(n35931), .c(delay_sub_ln23_0_unr30_stage10_stallmux_q), .o(n35932) );
oa12f01 g32142 ( .a(n35920), .b(n35932), .c(n35930), .o(n35933) );
in01f01 g32143 ( .a(n34063), .o(n35934) );
no03f01 g32144 ( .a(n34073), .b(n35934), .c(n34056), .o(n35935) );
no02f01 g32145 ( .a(n34054), .b(n34046), .o(n35936) );
no02f01 g32146 ( .a(n35913), .b(n35936), .o(n35937) );
no02f01 g32147 ( .a(n34073), .b(n35934), .o(n35938) );
no02f01 g32148 ( .a(n35938), .b(n35937), .o(n35939) );
no02f01 g32149 ( .a(n35939), .b(n35935), .o(n35940) );
in01f01 g32150 ( .a(n35940), .o(n35941) );
no02f01 g32151 ( .a(n35941), .b(n35912), .o(n35942) );
in01f01 g32152 ( .a(n35942), .o(n35943) );
no02f01 g32153 ( .a(n35931), .b(delay_sub_ln23_0_unr30_stage10_stallmux_q), .o(n35944) );
ao12f01 g32154 ( .a(n34073), .b(n34063), .c(n34056), .o(n35945) );
no02f01 g32155 ( .a(n34072), .b(n33508), .o(n35946) );
no02f01 g32156 ( .a(n34070), .b(n33507), .o(n35947) );
no02f01 g32157 ( .a(n35947), .b(n35946), .o(n35948) );
no02f01 g32158 ( .a(n35948), .b(n35945), .o(n35949) );
na02f01 g32159 ( .a(n35948), .b(n35945), .o(n35950) );
in01f01 g32160 ( .a(n35950), .o(n35951) );
no02f01 g32161 ( .a(n35951), .b(n35949), .o(n35952) );
na02f01 g32162 ( .a(n35952), .b(n35944), .o(n35953) );
na03f01 g32163 ( .a(n35953), .b(n35943), .c(n35933), .o(n35954) );
ao12f01 g32164 ( .a(n35944), .b(n35952), .c(n35940), .o(n35955) );
in01f01 g32165 ( .a(n35955), .o(n35956) );
na02f01 g32166 ( .a(n35956), .b(n35954), .o(n35957) );
no02f01 g32167 ( .a(n34035), .b(n33507), .o(n35958) );
no02f01 g32168 ( .a(n35958), .b(n34080), .o(n35959) );
in01f01 g32169 ( .a(n35959), .o(n35960) );
no02f01 g32170 ( .a(n35960), .b(n34251), .o(n35961) );
no02f01 g32171 ( .a(n35959), .b(n34078), .o(n35962) );
no02f01 g32172 ( .a(n35962), .b(n35961), .o(n35963) );
in01f01 g32173 ( .a(n35963), .o(n35964) );
no02f01 g32174 ( .a(n35964), .b(n35912), .o(n35965) );
no02f01 g32175 ( .a(n35963), .b(n35944), .o(n35966) );
no02f01 g32176 ( .a(n35966), .b(n35965), .o(n35967) );
in01f01 g32177 ( .a(n35967), .o(n35968) );
no02f01 g32178 ( .a(n35968), .b(n35957), .o(n35969) );
no02f01 g32179 ( .a(n35918), .b(n35944), .o(n35970) );
na03f01 g32180 ( .a(n35910), .b(n35891), .c(n34304), .o(n35971) );
na03f01 g32181 ( .a(n35910), .b(n35891), .c(delay_sub_ln23_0_unr30_stage10_stallmux_q), .o(n35972) );
in01f01 g32182 ( .a(n35929), .o(n35973) );
na03f01 g32183 ( .a(n35973), .b(n35972), .c(n35971), .o(n35974) );
in01f01 g32184 ( .a(n35932), .o(n35975) );
ao12f01 g32185 ( .a(n35970), .b(n35975), .c(n35974), .o(n35976) );
no02f01 g32186 ( .a(n35942), .b(n35976), .o(n35977) );
ao12f01 g32187 ( .a(n35955), .b(n35953), .c(n35977), .o(n35978) );
no02f01 g32188 ( .a(n35967), .b(n35978), .o(n35979) );
oa12f01 g32189 ( .a(n32734), .b(n35979), .c(n35969), .o(n35980) );
na02f01 g32190 ( .a(n35980), .b(n35595), .o(n472) );
in01f01 g32191 ( .a(n7413), .o(n35982) );
no02f01 g32192 ( .a(n7205), .b(n4338), .o(n35983) );
no02f01 g32193 ( .a(n7205), .b(n4370), .o(n35984) );
no02f01 g32194 ( .a(n35984), .b(n7418), .o(n35985) );
in01f01 g32195 ( .a(n35985), .o(n35986) );
no04f01 g32196 ( .a(n35986), .b(n35983), .c(n35982), .d(n7381), .o(n35987) );
ao12f01 g32197 ( .a(n7164), .b(n4263), .c(n4258), .o(n35988) );
oa12f01 g32198 ( .a(n7205), .b(n35988), .c(n4338), .o(n35989) );
na02f01 g32199 ( .a(n35989), .b(n7415), .o(n35990) );
no02f01 g32200 ( .a(n7205), .b(n4379_1), .o(n35991) );
no02f01 g32201 ( .a(n7164), .b(n4248), .o(n35992) );
no02f01 g32202 ( .a(n35992), .b(n35991), .o(n35993) );
in01f01 g32203 ( .a(n35993), .o(n35994) );
no03f01 g32204 ( .a(n35994), .b(n35990), .c(n35987), .o(n35995) );
no02f01 g32205 ( .a(n35990), .b(n35987), .o(n35996) );
no02f01 g32206 ( .a(n35993), .b(n35996), .o(n35997) );
no02f01 g32207 ( .a(n35997), .b(n35995), .o(n35998) );
no02f01 g32208 ( .a(n35998), .b(n3789), .o(n35999) );
in01f01 g32209 ( .a(n7425), .o(n36000) );
na03f01 g32210 ( .a(n36000), .b(n7455), .c(n7452), .o(n36001) );
no02f01 g32211 ( .a(n7164), .b(n4258), .o(n36002) );
no02f01 g32212 ( .a(n36002), .b(n35984), .o(n36003) );
in01f01 g32213 ( .a(n36003), .o(n36004) );
in01f01 g32214 ( .a(n7419), .o(n36005) );
ao12f01 g32215 ( .a(n7418), .b(n36005), .c(n7417), .o(n36006) );
no02f01 g32216 ( .a(n36006), .b(n36004), .o(n36007) );
na02f01 g32217 ( .a(n36006), .b(n36004), .o(n36008) );
in01f01 g32218 ( .a(n36008), .o(n36009) );
no02f01 g32219 ( .a(n36009), .b(n36007), .o(n36010) );
no02f01 g32220 ( .a(n36010), .b(n3789), .o(n36011) );
no02f01 g32221 ( .a(n36011), .b(n36001), .o(n36012) );
no02f01 g32222 ( .a(n36010), .b(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n36013) );
in01f01 g32223 ( .a(n36013), .o(n36014) );
no02f01 g32224 ( .a(n7164), .b(n4337), .o(n36015) );
no02f01 g32225 ( .a(n36015), .b(n35983), .o(n36016) );
in01f01 g32226 ( .a(n36016), .o(n36017) );
in01f01 g32227 ( .a(n35988), .o(n36018) );
oa12f01 g32228 ( .a(n36018), .b(n35986), .c(n7417), .o(n36019) );
no02f01 g32229 ( .a(n36019), .b(n36017), .o(n36020) );
na02f01 g32230 ( .a(n36019), .b(n36017), .o(n36021) );
in01f01 g32231 ( .a(n36021), .o(n36022) );
no02f01 g32232 ( .a(n36022), .b(n36020), .o(n36023) );
no02f01 g32233 ( .a(n36023), .b(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n36024) );
in01f01 g32234 ( .a(n36020), .o(n36025) );
na02f01 g32235 ( .a(n36021), .b(n36025), .o(n36026) );
no02f01 g32236 ( .a(n36026), .b(n3789), .o(n36027) );
no02f01 g32237 ( .a(n36027), .b(n36024), .o(n36028) );
na02f01 g32238 ( .a(n36028), .b(n36014), .o(n36029) );
oa12f01 g32239 ( .a(n3789), .b(n36029), .c(n36012), .o(n36030) );
na02f01 g32240 ( .a(n36026), .b(n3789), .o(n36031) );
na02f01 g32241 ( .a(n36023), .b(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n36032) );
na02f01 g32242 ( .a(n36032), .b(n36031), .o(n36033) );
ao12f01 g32243 ( .a(delay_sub_ln23_0_unr22_stage8_stallmux_q), .b(n7424), .c(n7409), .o(n36034) );
ao12f01 g32244 ( .a(n36034), .b(n36033), .c(n36012), .o(n36035) );
no02f01 g32245 ( .a(n35998), .b(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n36036) );
ao12f01 g32246 ( .a(n36036), .b(n36035), .c(n36030), .o(n36037) );
no02f01 g32247 ( .a(n36037), .b(n35999), .o(n36038) );
no02f01 g32248 ( .a(n4518_1), .b(n4389_1), .o(n36039) );
no02f01 g32249 ( .a(n4532), .b(n4344_1), .o(n36040) );
in01f01 g32250 ( .a(n4536), .o(n36041) );
ao12f01 g32251 ( .a(n36040), .b(n36041), .c(n36039), .o(n36042) );
no02f01 g32252 ( .a(n4525), .b(n4344_1), .o(n36043) );
no02f01 g32253 ( .a(n36043), .b(n4537), .o(n36044) );
no02f01 g32254 ( .a(n36044), .b(n36042), .o(n36045) );
na02f01 g32255 ( .a(n36044), .b(n36042), .o(n36046) );
in01f01 g32256 ( .a(n36046), .o(n36047) );
no02f01 g32257 ( .a(n36047), .b(n36045), .o(n36048) );
in01f01 g32258 ( .a(n36048), .o(n36049) );
no02f01 g32259 ( .a(n4536), .b(n36040), .o(n36050) );
in01f01 g32260 ( .a(n36050), .o(n36051) );
no02f01 g32261 ( .a(n36051), .b(n36039), .o(n36052) );
na02f01 g32262 ( .a(n36051), .b(n36039), .o(n36053) );
in01f01 g32263 ( .a(n36053), .o(n36054) );
no02f01 g32264 ( .a(n36054), .b(n36052), .o(n36055) );
in01f01 g32265 ( .a(n36055), .o(n36056) );
ao12f01 g32266 ( .a(n36038), .b(n36056), .c(n36049), .o(n36057) );
no03f01 g32267 ( .a(n7425), .b(n7410), .c(n7399), .o(n36058) );
in01f01 g32268 ( .a(n36011), .o(n36059) );
na02f01 g32269 ( .a(n36059), .b(n36058), .o(n36060) );
no02f01 g32270 ( .a(n36034), .b(n36013), .o(n36061) );
no02f01 g32271 ( .a(n36023), .b(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n36062) );
no02f01 g32272 ( .a(n36023), .b(n3789), .o(n36063) );
no02f01 g32273 ( .a(n36063), .b(n36062), .o(n36064) );
ao12f01 g32274 ( .a(n36064), .b(n36061), .c(n36060), .o(n36065) );
in01f01 g32275 ( .a(n36061), .o(n36066) );
in01f01 g32276 ( .a(n36064), .o(n36067) );
no03f01 g32277 ( .a(n36067), .b(n36066), .c(n36012), .o(n36068) );
no02f01 g32278 ( .a(n4512), .b(n4420), .o(n36069) );
no02f01 g32279 ( .a(n4677_1), .b(n4407), .o(n36070) );
no02f01 g32280 ( .a(n36070), .b(n36069), .o(n36071) );
na02f01 g32281 ( .a(n36070), .b(n36069), .o(n36072) );
in01f01 g32282 ( .a(n36072), .o(n36073) );
no02f01 g32283 ( .a(n36073), .b(n36071), .o(n36074) );
in01f01 g32284 ( .a(n36074), .o(n36075) );
no03f01 g32285 ( .a(n36075), .b(n36068), .c(n36065), .o(n36076) );
oa12f01 g32286 ( .a(n7523), .b(n7547), .c(n7438), .o(n36077) );
no02f01 g32287 ( .a(n36013), .b(n36011), .o(n36078) );
in01f01 g32288 ( .a(n36078), .o(n36079) );
oa12f01 g32289 ( .a(n36079), .b(n36034), .c(n36058), .o(n36080) );
in01f01 g32290 ( .a(n36034), .o(n36081) );
na03f01 g32291 ( .a(n36078), .b(n36081), .c(n36001), .o(n36082) );
na02f01 g32292 ( .a(n36082), .b(n36080), .o(n36083) );
no04f01 g32293 ( .a(n4511), .b(n4674), .c(n4429_1), .d(n4420), .o(n36084) );
ao22f01 g32294 ( .a(n4675), .b(n4652_1), .c(n4507), .d(n4430), .o(n36085) );
no02f01 g32295 ( .a(n36085), .b(n36084), .o(n36086) );
in01f01 g32296 ( .a(n36086), .o(n36087) );
no02f01 g32297 ( .a(n36087), .b(n36083), .o(n36088) );
in01f01 g32298 ( .a(n36088), .o(n36089) );
oa12f01 g32299 ( .a(n36075), .b(n36068), .c(n36065), .o(n36090) );
ao12f01 g32300 ( .a(n36086), .b(n36082), .c(n36080), .o(n36091) );
in01f01 g32301 ( .a(n36091), .o(n36092) );
na02f01 g32302 ( .a(n36092), .b(n36090), .o(n36093) );
ao12f01 g32303 ( .a(n36093), .b(n36089), .c(n36077), .o(n36094) );
no02f01 g32304 ( .a(n36036), .b(n35999), .o(n36095) );
na03f01 g32305 ( .a(n36095), .b(n36035), .c(n36030), .o(n36096) );
no02f01 g32306 ( .a(n36033), .b(n36013), .o(n36097) );
ao12f01 g32307 ( .a(delay_sub_ln23_0_unr22_stage8_stallmux_q), .b(n36097), .c(n36060), .o(n36098) );
oa12f01 g32308 ( .a(n36081), .b(n36028), .c(n36060), .o(n36099) );
in01f01 g32309 ( .a(n36095), .o(n36100) );
oa12f01 g32310 ( .a(n36100), .b(n36099), .c(n36098), .o(n36101) );
na02f01 g32311 ( .a(n36101), .b(n36096), .o(n36102) );
no04f01 g32312 ( .a(n4515), .b(n4678), .c(n4407), .d(n4398), .o(n36103) );
ao22f01 g32313 ( .a(n4679), .b(n4651), .c(n4513_1), .d(n4408), .o(n36104) );
no02f01 g32314 ( .a(n36104), .b(n36103), .o(n36105) );
in01f01 g32315 ( .a(n36105), .o(n36106) );
no02f01 g32316 ( .a(n36106), .b(n36102), .o(n36107) );
no02f01 g32317 ( .a(n4516), .b(n4398), .o(n36108) );
no02f01 g32318 ( .a(n4517), .b(n4389_1), .o(n36109) );
no02f01 g32319 ( .a(n36109), .b(n36108), .o(n36110) );
na02f01 g32320 ( .a(n36109), .b(n36108), .o(n36111) );
in01f01 g32321 ( .a(n36111), .o(n36112) );
no02f01 g32322 ( .a(n36112), .b(n36110), .o(n36113) );
in01f01 g32323 ( .a(n36113), .o(n36114) );
no02f01 g32324 ( .a(n36114), .b(n36038), .o(n36115) );
no04f01 g32325 ( .a(n36115), .b(n36107), .c(n36094), .d(n36076), .o(n36116) );
na02f01 g32326 ( .a(n36106), .b(n36102), .o(n36117) );
na02f01 g32327 ( .a(n36114), .b(n36038), .o(n36118) );
ao12f01 g32328 ( .a(n36115), .b(n36118), .c(n36117), .o(n36119) );
in01f01 g32329 ( .a(n35999), .o(n36120) );
no02f01 g32330 ( .a(n36099), .b(n36098), .o(n36121) );
oa12f01 g32331 ( .a(n36120), .b(n36036), .c(n36121), .o(n36122) );
ao12f01 g32332 ( .a(n36122), .b(n36055), .c(n36048), .o(n36123) );
no03f01 g32333 ( .a(n36123), .b(n36119), .c(n36116), .o(n36124) );
no02f01 g32334 ( .a(n4685), .b(n4684), .o(n36125) );
no02f01 g32335 ( .a(n4545), .b(n4344_1), .o(n36126) );
no02f01 g32336 ( .a(n36126), .b(n4547), .o(n36127) );
in01f01 g32337 ( .a(n36127), .o(n36128) );
no02f01 g32338 ( .a(n36128), .b(n36125), .o(n36129) );
in01f01 g32339 ( .a(n36125), .o(n36130) );
no02f01 g32340 ( .a(n36127), .b(n36130), .o(n36131) );
no02f01 g32341 ( .a(n36131), .b(n36129), .o(n36132) );
in01f01 g32342 ( .a(n36132), .o(n36133) );
ao12f01 g32343 ( .a(n36126), .b(n4548_1), .c(n36125), .o(n36134) );
no02f01 g32344 ( .a(n4568_1), .b(n4344_1), .o(n36135) );
no02f01 g32345 ( .a(n36135), .b(n4570), .o(n36136) );
no02f01 g32346 ( .a(n36136), .b(n36134), .o(n36137) );
na02f01 g32347 ( .a(n36136), .b(n36134), .o(n36138) );
in01f01 g32348 ( .a(n36138), .o(n36139) );
no02f01 g32349 ( .a(n36139), .b(n36137), .o(n36140) );
in01f01 g32350 ( .a(n36140), .o(n36141) );
ao12f01 g32351 ( .a(n36038), .b(n36141), .c(n36133), .o(n36142) );
no02f01 g32352 ( .a(n4556), .b(n4344_1), .o(n36143) );
in01f01 g32353 ( .a(n36143), .o(n36144) );
no03f01 g32354 ( .a(n4570), .b(n4547), .c(n36130), .o(n36145) );
no02f01 g32355 ( .a(n36145), .b(n4585), .o(n36146) );
ao12f01 g32356 ( .a(n4558_1), .b(n36146), .c(n36144), .o(n36147) );
no02f01 g32357 ( .a(n4579), .b(n4344_1), .o(n36148) );
no02f01 g32358 ( .a(n36148), .b(n4581), .o(n36149) );
in01f01 g32359 ( .a(n36149), .o(n36150) );
no02f01 g32360 ( .a(n36150), .b(n36147), .o(n36151) );
na02f01 g32361 ( .a(n36150), .b(n36147), .o(n36152) );
in01f01 g32362 ( .a(n36152), .o(n36153) );
no02f01 g32363 ( .a(n36153), .b(n36151), .o(n36154) );
na02f01 g32364 ( .a(n36154), .b(n36122), .o(n36155) );
in01f01 g32365 ( .a(n36155), .o(n36156) );
no02f01 g32366 ( .a(n36143), .b(n4558_1), .o(n36157) );
in01f01 g32367 ( .a(n36157), .o(n36158) );
no03f01 g32368 ( .a(n36158), .b(n36145), .c(n4585), .o(n36159) );
no02f01 g32369 ( .a(n36157), .b(n36146), .o(n36160) );
no02f01 g32370 ( .a(n36160), .b(n36159), .o(n36161) );
na02f01 g32371 ( .a(n36161), .b(n36122), .o(n36162) );
in01f01 g32372 ( .a(n36162), .o(n36163) );
no02f01 g32373 ( .a(n36163), .b(n36156), .o(n36164) );
in01f01 g32374 ( .a(n36164), .o(n36165) );
no04f01 g32375 ( .a(n36165), .b(n36142), .c(n36124), .d(n36057), .o(n36166) );
ao12f01 g32376 ( .a(n36122), .b(n36140), .c(n36132), .o(n36167) );
ao12f01 g32377 ( .a(n36122), .b(n36161), .c(n36154), .o(n36168) );
no02f01 g32378 ( .a(n36168), .b(n36167), .o(n36169) );
in01f01 g32379 ( .a(n36169), .o(n36170) );
no02f01 g32380 ( .a(n36170), .b(n36166), .o(n36171) );
in01f01 g32381 ( .a(n4609), .o(n36172) );
no02f01 g32382 ( .a(n4607), .b(n4344_1), .o(n36173) );
ao12f01 g32383 ( .a(n36173), .b(n36172), .c(n4587), .o(n36174) );
in01f01 g32384 ( .a(n36174), .o(n36175) );
no02f01 g32385 ( .a(n4600), .b(n4344_1), .o(n36176) );
no02f01 g32386 ( .a(n36176), .b(n4602), .o(n36177) );
in01f01 g32387 ( .a(n36177), .o(n36178) );
no02f01 g32388 ( .a(n36178), .b(n36175), .o(n36179) );
no02f01 g32389 ( .a(n36177), .b(n36174), .o(n36180) );
no02f01 g32390 ( .a(n36180), .b(n36179), .o(n36181) );
no02f01 g32391 ( .a(n36173), .b(n4609), .o(n36182) );
no02f01 g32392 ( .a(n36182), .b(n4689), .o(n36183) );
na02f01 g32393 ( .a(n36182), .b(n4689), .o(n36184) );
in01f01 g32394 ( .a(n36184), .o(n36185) );
no02f01 g32395 ( .a(n36185), .b(n36183), .o(n36186) );
no02f01 g32396 ( .a(n36186), .b(n36181), .o(n36187) );
no02f01 g32397 ( .a(n36187), .b(n36038), .o(n36188) );
no02f01 g32398 ( .a(n36188), .b(n36171), .o(n36189) );
no02f01 g32399 ( .a(n4627), .b(n4344_1), .o(n36190) );
no02f01 g32400 ( .a(n36190), .b(n4629), .o(n36191) );
in01f01 g32401 ( .a(n36191), .o(n36192) );
no03f01 g32402 ( .a(n36192), .b(n4633_1), .c(n4697_1), .o(n36193) );
in01f01 g32403 ( .a(n4633_1), .o(n36194) );
ao12f01 g32404 ( .a(n36191), .b(n36194), .c(n4723), .o(n36195) );
no02f01 g32405 ( .a(n36195), .b(n36193), .o(n36196) );
na02f01 g32406 ( .a(n36196), .b(n36122), .o(n36197) );
ao12f01 g32407 ( .a(n36122), .b(n36186), .c(n36181), .o(n36198) );
in01f01 g32408 ( .a(n36198), .o(n36199) );
in01f01 g32409 ( .a(n36196), .o(n36200) );
na02f01 g32410 ( .a(n36200), .b(n36038), .o(n36201) );
na02f01 g32411 ( .a(n36201), .b(n36199), .o(n36202) );
ao12f01 g32412 ( .a(n36202), .b(n36197), .c(n36189), .o(n36203) );
no02f01 g32413 ( .a(n4633_1), .b(n36190), .o(n36204) );
oa12f01 g32414 ( .a(n36204), .b(n4629), .c(n4723), .o(n36205) );
no02f01 g32415 ( .a(n4619), .b(n4344_1), .o(n36206) );
no02f01 g32416 ( .a(n36206), .b(n4621), .o(n36207) );
in01f01 g32417 ( .a(n36207), .o(n36208) );
no02f01 g32418 ( .a(n36208), .b(n36205), .o(n36209) );
na02f01 g32419 ( .a(n36208), .b(n36205), .o(n36210) );
in01f01 g32420 ( .a(n36210), .o(n36211) );
no02f01 g32421 ( .a(n36211), .b(n36209), .o(n36212) );
no02f01 g32422 ( .a(n36212), .b(n36122), .o(n36213) );
in01f01 g32423 ( .a(n36212), .o(n36214) );
no02f01 g32424 ( .a(n36214), .b(n36038), .o(n36215) );
no02f01 g32425 ( .a(n36215), .b(n36213), .o(n36216) );
na02f01 g32426 ( .a(n36216), .b(n36203), .o(n36217) );
in01f01 g32427 ( .a(n36203), .o(n36218) );
in01f01 g32428 ( .a(n36216), .o(n36219) );
na02f01 g32429 ( .a(n36219), .b(n36218), .o(n36220) );
na02f01 g32430 ( .a(n36220), .b(n36217), .o(n476) );
na02f01 g32431 ( .a(n32732), .b(cos_out_17), .o(n36222) );
no02f01 g32432 ( .a(n34202), .b(n33507), .o(n36223) );
na02f01 g32433 ( .a(n34202), .b(n33507), .o(n36224) );
in01f01 g32434 ( .a(n36224), .o(n36225) );
no02f01 g32435 ( .a(n36225), .b(n36223), .o(n36226) );
no02f01 g32436 ( .a(n36226), .b(n34262), .o(n36227) );
na02f01 g32437 ( .a(n36226), .b(n34262), .o(n36228) );
in01f01 g32438 ( .a(n36228), .o(n36229) );
no02f01 g32439 ( .a(n36229), .b(n36227), .o(n36230) );
no02f01 g32440 ( .a(n36230), .b(n35944), .o(n36231) );
no02f01 g32441 ( .a(n34080), .b(n34078), .o(n36232) );
no02f01 g32442 ( .a(n34030), .b(n33507), .o(n36233) );
no02f01 g32443 ( .a(n36233), .b(n34082), .o(n36234) );
in01f01 g32444 ( .a(n36234), .o(n36235) );
no03f01 g32445 ( .a(n36235), .b(n35958), .c(n36232), .o(n36236) );
no02f01 g32446 ( .a(n35958), .b(n36232), .o(n36237) );
no02f01 g32447 ( .a(n36234), .b(n36237), .o(n36238) );
no02f01 g32448 ( .a(n36238), .b(n36236), .o(n36239) );
in01f01 g32449 ( .a(n36239), .o(n36240) );
no02f01 g32450 ( .a(n36240), .b(n35912), .o(n36241) );
ao12f01 g32451 ( .a(n34036), .b(n34253), .c(n36232), .o(n36242) );
no02f01 g32452 ( .a(n34089), .b(n33507), .o(n36243) );
no02f01 g32453 ( .a(n36243), .b(n34091), .o(n36244) );
no02f01 g32454 ( .a(n36244), .b(n36242), .o(n36245) );
na02f01 g32455 ( .a(n36244), .b(n36242), .o(n36246) );
in01f01 g32456 ( .a(n36246), .o(n36247) );
no02f01 g32457 ( .a(n36247), .b(n36245), .o(n36248) );
in01f01 g32458 ( .a(n36248), .o(n36249) );
no02f01 g32459 ( .a(n36249), .b(n35912), .o(n36250) );
no02f01 g32460 ( .a(n36250), .b(n36241), .o(n36251) );
in01f01 g32461 ( .a(n36251), .o(n36252) );
no03f01 g32462 ( .a(n36252), .b(n35965), .c(n35978), .o(n36253) );
no03f01 g32463 ( .a(n36243), .b(n34092), .c(n34036), .o(n36254) );
in01f01 g32464 ( .a(n36254), .o(n36255) );
no02f01 g32465 ( .a(n34017), .b(n33507), .o(n36256) );
no02f01 g32466 ( .a(n36256), .b(n34019), .o(n36257) );
in01f01 g32467 ( .a(n36257), .o(n36258) );
no02f01 g32468 ( .a(n36258), .b(n36255), .o(n36259) );
no02f01 g32469 ( .a(n36257), .b(n36254), .o(n36260) );
no02f01 g32470 ( .a(n36260), .b(n36259), .o(n36261) );
in01f01 g32471 ( .a(n36261), .o(n36262) );
no02f01 g32472 ( .a(n36262), .b(n35912), .o(n36263) );
in01f01 g32473 ( .a(n36263), .o(n36264) );
ao12f01 g32474 ( .a(n35944), .b(n36261), .c(n36248), .o(n36265) );
ao12f01 g32475 ( .a(n35944), .b(n36239), .c(n35963), .o(n36266) );
no02f01 g32476 ( .a(n36266), .b(n36265), .o(n36267) );
in01f01 g32477 ( .a(n36267), .o(n36268) );
ao12f01 g32478 ( .a(n36268), .b(n36264), .c(n36253), .o(n36269) );
no02f01 g32479 ( .a(n34094), .b(n34019), .o(n36270) );
no02f01 g32480 ( .a(n34004), .b(n33507), .o(n36271) );
no02f01 g32481 ( .a(n34005), .b(n33508), .o(n36272) );
no02f01 g32482 ( .a(n36272), .b(n36271), .o(n36273) );
in01f01 g32483 ( .a(n36273), .o(n36274) );
no02f01 g32484 ( .a(n36274), .b(n36270), .o(n36275) );
no03f01 g32485 ( .a(n36273), .b(n34094), .c(n34019), .o(n36276) );
no02f01 g32486 ( .a(n36276), .b(n36275), .o(n36277) );
in01f01 g32487 ( .a(n36277), .o(n36278) );
no02f01 g32488 ( .a(n36278), .b(n35912), .o(n36279) );
in01f01 g32489 ( .a(n36272), .o(n36280) );
ao12f01 g32490 ( .a(n36271), .b(n36280), .c(n36270), .o(n36281) );
no02f01 g32491 ( .a(n33998), .b(n33508), .o(n36282) );
no02f01 g32492 ( .a(n33997), .b(n33507), .o(n36283) );
no02f01 g32493 ( .a(n36283), .b(n36282), .o(n36284) );
no02f01 g32494 ( .a(n36284), .b(n36281), .o(n36285) );
na02f01 g32495 ( .a(n36284), .b(n36281), .o(n36286) );
in01f01 g32496 ( .a(n36286), .o(n36287) );
no02f01 g32497 ( .a(n36287), .b(n36285), .o(n36288) );
in01f01 g32498 ( .a(n36288), .o(n36289) );
no02f01 g32499 ( .a(n36289), .b(n35912), .o(n36290) );
no02f01 g32500 ( .a(n36290), .b(n36279), .o(n36291) );
in01f01 g32501 ( .a(n36291), .o(n36292) );
no02f01 g32502 ( .a(n34101), .b(n33507), .o(n36293) );
no02f01 g32503 ( .a(n34157), .b(n36293), .o(n36294) );
na02f01 g32504 ( .a(n36294), .b(n34259), .o(n36295) );
in01f01 g32505 ( .a(n36295), .o(n36296) );
no02f01 g32506 ( .a(n34112), .b(n33507), .o(n36297) );
no02f01 g32507 ( .a(n36297), .b(n34114), .o(n36298) );
no02f01 g32508 ( .a(n36298), .b(n36296), .o(n36299) );
na02f01 g32509 ( .a(n36298), .b(n36296), .o(n36300) );
in01f01 g32510 ( .a(n36300), .o(n36301) );
no02f01 g32511 ( .a(n36301), .b(n36299), .o(n36302) );
in01f01 g32512 ( .a(n36302), .o(n36303) );
no02f01 g32513 ( .a(n36303), .b(n35912), .o(n36304) );
ao12f01 g32514 ( .a(n34157), .b(n36270), .c(n34248), .o(n36305) );
in01f01 g32515 ( .a(n36305), .o(n36306) );
no02f01 g32516 ( .a(n36293), .b(n34103), .o(n36307) );
in01f01 g32517 ( .a(n36307), .o(n36308) );
no02f01 g32518 ( .a(n36308), .b(n36306), .o(n36309) );
no02f01 g32519 ( .a(n36307), .b(n36305), .o(n36310) );
no02f01 g32520 ( .a(n36310), .b(n36309), .o(n36311) );
in01f01 g32521 ( .a(n36311), .o(n36312) );
no02f01 g32522 ( .a(n36312), .b(n35912), .o(n36313) );
no03f01 g32523 ( .a(n36313), .b(n36304), .c(n36292), .o(n36314) );
in01f01 g32524 ( .a(n36314), .o(n36315) );
no02f01 g32525 ( .a(n34140), .b(n33507), .o(n36316) );
no02f01 g32526 ( .a(n34159), .b(n34260), .o(n36317) );
in01f01 g32527 ( .a(n36317), .o(n36318) );
na02f01 g32528 ( .a(n34140), .b(n33507), .o(n36319) );
ao12f01 g32529 ( .a(n36316), .b(n36319), .c(n36318), .o(n36320) );
in01f01 g32530 ( .a(n36320), .o(n36321) );
in01f01 g32531 ( .a(n34134), .o(n36322) );
no02f01 g32532 ( .a(n36322), .b(n33508), .o(n36323) );
no02f01 g32533 ( .a(n34134), .b(n33507), .o(n36324) );
no02f01 g32534 ( .a(n36324), .b(n36323), .o(n36325) );
in01f01 g32535 ( .a(n36325), .o(n36326) );
no02f01 g32536 ( .a(n36326), .b(n36321), .o(n36327) );
no02f01 g32537 ( .a(n36325), .b(n36320), .o(n36328) );
no02f01 g32538 ( .a(n36328), .b(n36327), .o(n36329) );
in01f01 g32539 ( .a(n36329), .o(n36330) );
no02f01 g32540 ( .a(n36330), .b(n35912), .o(n36331) );
in01f01 g32541 ( .a(n36319), .o(n36332) );
no02f01 g32542 ( .a(n36332), .b(n36316), .o(n36333) );
no02f01 g32543 ( .a(n36333), .b(n36317), .o(n36334) );
na02f01 g32544 ( .a(n36333), .b(n36317), .o(n36335) );
in01f01 g32545 ( .a(n36335), .o(n36336) );
no02f01 g32546 ( .a(n36336), .b(n36334), .o(n36337) );
in01f01 g32547 ( .a(n36337), .o(n36338) );
no02f01 g32548 ( .a(n36338), .b(n35912), .o(n36339) );
no02f01 g32549 ( .a(n36339), .b(n36331), .o(n36340) );
in01f01 g32550 ( .a(n36340), .o(n36341) );
no02f01 g32551 ( .a(n34122), .b(n33507), .o(n36342) );
in01f01 g32552 ( .a(n36342), .o(n36343) );
no02f01 g32553 ( .a(n36317), .b(n34142), .o(n36344) );
no02f01 g32554 ( .a(n36344), .b(n34160), .o(n36345) );
ao12f01 g32555 ( .a(n34124), .b(n36345), .c(n36343), .o(n36346) );
in01f01 g32556 ( .a(n36346), .o(n36347) );
no02f01 g32557 ( .a(n34151), .b(n33507), .o(n36348) );
no02f01 g32558 ( .a(n36348), .b(n34153), .o(n36349) );
no02f01 g32559 ( .a(n36349), .b(n36347), .o(n36350) );
na02f01 g32560 ( .a(n36349), .b(n36347), .o(n36351) );
in01f01 g32561 ( .a(n36351), .o(n36352) );
no02f01 g32562 ( .a(n36352), .b(n36350), .o(n36353) );
in01f01 g32563 ( .a(n36353), .o(n36354) );
no02f01 g32564 ( .a(n36354), .b(n35912), .o(n36355) );
no02f01 g32565 ( .a(n36342), .b(n34124), .o(n36356) );
in01f01 g32566 ( .a(n36356), .o(n36357) );
no03f01 g32567 ( .a(n36357), .b(n36344), .c(n34160), .o(n36358) );
no02f01 g32568 ( .a(n36356), .b(n36345), .o(n36359) );
no02f01 g32569 ( .a(n36359), .b(n36358), .o(n36360) );
in01f01 g32570 ( .a(n36360), .o(n36361) );
no02f01 g32571 ( .a(n36361), .b(n35912), .o(n36362) );
no03f01 g32572 ( .a(n36362), .b(n36355), .c(n36341), .o(n36363) );
in01f01 g32573 ( .a(n36363), .o(n36364) );
no03f01 g32574 ( .a(n36364), .b(n36315), .c(n36269), .o(n36365) );
ao12f01 g32575 ( .a(n35944), .b(n36311), .c(n36302), .o(n36366) );
ao12f01 g32576 ( .a(n35944), .b(n36288), .c(n36277), .o(n36367) );
no02f01 g32577 ( .a(n36367), .b(n36366), .o(n36368) );
in01f01 g32578 ( .a(n36368), .o(n36369) );
ao12f01 g32579 ( .a(n35944), .b(n36337), .c(n36329), .o(n36370) );
ao12f01 g32580 ( .a(n35944), .b(n36360), .c(n36353), .o(n36371) );
no03f01 g32581 ( .a(n36371), .b(n36370), .c(n36369), .o(n36372) );
in01f01 g32582 ( .a(n36372), .o(n36373) );
no02f01 g32583 ( .a(n36373), .b(n36365), .o(n36374) );
in01f01 g32584 ( .a(n36230), .o(n36375) );
no02f01 g32585 ( .a(n36375), .b(n35912), .o(n36376) );
no02f01 g32586 ( .a(n36376), .b(n36374), .o(n36377) );
ao12f01 g32587 ( .a(n36223), .b(n36224), .c(n34163), .o(n36378) );
in01f01 g32588 ( .a(n36378), .o(n36379) );
in01f01 g32589 ( .a(n34197), .o(n36380) );
no02f01 g32590 ( .a(n36380), .b(n33508), .o(n36381) );
no02f01 g32591 ( .a(n34197), .b(n33507), .o(n36382) );
no02f01 g32592 ( .a(n36382), .b(n36381), .o(n36383) );
in01f01 g32593 ( .a(n36383), .o(n36384) );
no02f01 g32594 ( .a(n36384), .b(n36379), .o(n36385) );
no02f01 g32595 ( .a(n36383), .b(n36378), .o(n36386) );
no02f01 g32596 ( .a(n36386), .b(n36385), .o(n36387) );
in01f01 g32597 ( .a(n36387), .o(n36388) );
no02f01 g32598 ( .a(n36388), .b(n35912), .o(n36389) );
no02f01 g32599 ( .a(n36387), .b(n35944), .o(n36390) );
no02f01 g32600 ( .a(n36390), .b(n36389), .o(n36391) );
in01f01 g32601 ( .a(n36391), .o(n36392) );
no03f01 g32602 ( .a(n36392), .b(n36377), .c(n36231), .o(n36393) );
no02f01 g32603 ( .a(n36377), .b(n36231), .o(n36394) );
no02f01 g32604 ( .a(n36391), .b(n36394), .o(n36395) );
oa12f01 g32605 ( .a(n32734), .b(n36395), .c(n36393), .o(n36396) );
na02f01 g32606 ( .a(n36396), .b(n36222), .o(n481) );
no02f01 g32607 ( .a(n9591), .b(n9231), .o(n36398) );
no02f01 g32608 ( .a(n36398), .b(n9241), .o(n36399) );
in01f01 g32609 ( .a(n36399), .o(n5638) );
no02f01 g32610 ( .a(n4201), .b(n936), .o(n36401) );
no02f01 g32611 ( .a(n36401), .b(n5638), .o(n36402) );
in01f01 g32612 ( .a(n36401), .o(n36403) );
no02f01 g32613 ( .a(n36403), .b(n36399), .o(n36404) );
no02f01 g32614 ( .a(n36404), .b(n36402), .o(n485) );
no02f01 g32615 ( .a(n22028), .b(n21661), .o(n36406) );
no02f01 g32616 ( .a(n22034), .b(n21662), .o(n36407) );
no02f01 g32617 ( .a(n36407), .b(n36406), .o(n36408) );
no02f01 g32618 ( .a(n22046), .b(n21665), .o(n36409) );
in01f01 g32619 ( .a(n36409), .o(n36410) );
oa12f01 g32620 ( .a(n22028), .b(n22031), .c(n21666), .o(n36411) );
na03f01 g32621 ( .a(n36411), .b(n36410), .c(n36408), .o(n36412) );
in01f01 g32622 ( .a(n36408), .o(n36413) );
no02f01 g32623 ( .a(n22031), .b(n21666), .o(n36414) );
no02f01 g32624 ( .a(n36414), .b(n22034), .o(n36415) );
oa12f01 g32625 ( .a(n36413), .b(n36415), .c(n36409), .o(n36416) );
ao12f01 g32626 ( .a(n11514), .b(n36416), .c(n36412), .o(n36417) );
no03f01 g32627 ( .a(n36415), .b(n36409), .c(n36413), .o(n36418) );
ao12f01 g32628 ( .a(n36408), .b(n36411), .c(n36410), .o(n36419) );
oa12f01 g32629 ( .a(n11514), .b(n36419), .c(n36418), .o(n36420) );
oa12f01 g32630 ( .a(n11514), .b(n22452), .c(n22048), .o(n36421) );
no02f01 g32631 ( .a(n22433), .b(n22014), .o(n36422) );
ao12f01 g32632 ( .a(n22429), .b(n22044), .c(n22008), .o(n36423) );
oa12f01 g32633 ( .a(n11514), .b(n36423), .c(n36422), .o(n36424) );
na03f01 g32634 ( .a(n36424), .b(n25594), .c(n25582), .o(n36425) );
no03f01 g32635 ( .a(n25612), .b(n25595), .c(n25592), .o(n36426) );
na02f01 g32636 ( .a(n36426), .b(n36425), .o(n36427) );
oa12f01 g32637 ( .a(n11515), .b(n22052), .c(n22051), .o(n36428) );
oa12f01 g32638 ( .a(n11515), .b(n22445), .c(n22443), .o(n36429) );
na02f01 g32639 ( .a(n36429), .b(n36428), .o(n36430) );
ao12f01 g32640 ( .a(n36430), .b(n36427), .c(n36421), .o(n36431) );
oa12f01 g32641 ( .a(n36420), .b(n36431), .c(n36417), .o(n36432) );
no02f01 g32642 ( .a(n36432), .b(n21954), .o(n36433) );
oa12f01 g32643 ( .a(n11515), .b(n36419), .c(n36418), .o(n36434) );
ao12f01 g32644 ( .a(n11515), .b(n36416), .c(n36412), .o(n36435) );
ao12f01 g32645 ( .a(n11515), .b(n22446), .c(n22053), .o(n36436) );
oa12f01 g32646 ( .a(n25594), .b(n25590), .c(n11515), .o(n36437) );
no02f01 g32647 ( .a(n36437), .b(n25611), .o(n36438) );
oa12f01 g32648 ( .a(n11515), .b(n36423), .c(n36422), .o(n36439) );
ao12f01 g32649 ( .a(n25595), .b(n22401), .c(n11515), .o(n36440) );
na02f01 g32650 ( .a(n36440), .b(n36439), .o(n36441) );
no02f01 g32651 ( .a(n36441), .b(n36438), .o(n36442) );
ao12f01 g32652 ( .a(n11514), .b(n22047), .c(n22039), .o(n36443) );
ao12f01 g32653 ( .a(n11514), .b(n22451), .c(n22450), .o(n36444) );
no02f01 g32654 ( .a(n36444), .b(n36443), .o(n36445) );
oa12f01 g32655 ( .a(n36445), .b(n36442), .c(n36436), .o(n36446) );
ao12f01 g32656 ( .a(n36435), .b(n36446), .c(n36434), .o(n36447) );
no02f01 g32657 ( .a(n36447), .b(n21962), .o(n36448) );
no02f01 g32658 ( .a(n36448), .b(n36433), .o(n36449) );
in01f01 g32659 ( .a(n21914), .o(n36450) );
na02f01 g32660 ( .a(n25596), .b(n25593), .o(n36451) );
na02f01 g32661 ( .a(n25586), .b(n25584), .o(n36452) );
na02f01 g32662 ( .a(n36452), .b(n36451), .o(n36453) );
no02f01 g32663 ( .a(n36453), .b(n36450), .o(n36454) );
no02f01 g32664 ( .a(n25620), .b(n36454), .o(n36455) );
in01f01 g32665 ( .a(n21922), .o(n36456) );
na02f01 g32666 ( .a(n25617), .b(n25615), .o(n36457) );
na02f01 g32667 ( .a(n36457), .b(n36456), .o(n36458) );
na02f01 g32668 ( .a(n25607), .b(n25599), .o(n36459) );
na03f01 g32669 ( .a(n36459), .b(n36458), .c(n25601), .o(n36460) );
ao22f01 g32670 ( .a(n36460), .b(n25619), .c(n36455), .d(n25605), .o(n36461) );
no02f01 g32671 ( .a(n22446), .b(n11515), .o(n36462) );
ao12f01 g32672 ( .a(n11515), .b(n22047), .c(n22039), .o(n36463) );
no02f01 g32673 ( .a(n36443), .b(n36463), .o(n36464) );
no03f01 g32674 ( .a(n36444), .b(n36441), .c(n36438), .o(n36465) );
no03f01 g32675 ( .a(n36465), .b(n36464), .c(n36462), .o(n36466) );
na02f01 g32676 ( .a(n22452), .b(n11514), .o(n36467) );
oa12f01 g32677 ( .a(n11514), .b(n22052), .c(n22051), .o(n36468) );
na02f01 g32678 ( .a(n36428), .b(n36468), .o(n36469) );
na03f01 g32679 ( .a(n36429), .b(n36426), .c(n36425), .o(n36470) );
ao12f01 g32680 ( .a(n36469), .b(n36470), .c(n36467), .o(n36471) );
no03f01 g32681 ( .a(n36471), .b(n36466), .c(n21939), .o(n36472) );
na03f01 g32682 ( .a(n36470), .b(n36469), .c(n36467), .o(n36473) );
oa12f01 g32683 ( .a(n36464), .b(n36465), .c(n36462), .o(n36474) );
na03f01 g32684 ( .a(n36474), .b(n36473), .c(n21968), .o(n36475) );
na02f01 g32685 ( .a(n36429), .b(n36467), .o(n36476) );
na02f01 g32686 ( .a(n36476), .b(n36427), .o(n36477) );
no02f01 g32687 ( .a(n36444), .b(n36462), .o(n36478) );
na02f01 g32688 ( .a(n36478), .b(n36442), .o(n36479) );
na03f01 g32689 ( .a(n36479), .b(n36477), .c(n21846), .o(n36480) );
na02f01 g32690 ( .a(n36480), .b(n36475), .o(n36481) );
ao12f01 g32691 ( .a(n21968), .b(n36474), .c(n36473), .o(n36482) );
ao12f01 g32692 ( .a(n21846), .b(n36479), .c(n36477), .o(n36483) );
no02f01 g32693 ( .a(n36483), .b(n36482), .o(n36484) );
oa22f01 g32694 ( .a(n36484), .b(n36472), .c(n36481), .d(n36461), .o(n36485) );
oa12f01 g32695 ( .a(n36421), .b(n36430), .c(n36427), .o(n36486) );
na03f01 g32696 ( .a(n36486), .b(n36420), .c(n36434), .o(n36487) );
ao12f01 g32697 ( .a(n36436), .b(n36445), .c(n36442), .o(n36488) );
oa12f01 g32698 ( .a(n36488), .b(n36435), .c(n36417), .o(n36489) );
ao12f01 g32699 ( .a(n21965), .b(n36489), .c(n36487), .o(n36490) );
no02f01 g32700 ( .a(n36490), .b(n36485), .o(n36491) );
no03f01 g32701 ( .a(n36488), .b(n36435), .c(n36417), .o(n36492) );
ao12f01 g32702 ( .a(n36486), .b(n36420), .c(n36434), .o(n36493) );
no03f01 g32703 ( .a(n36493), .b(n36492), .c(n22098), .o(n36494) );
oa12f01 g32704 ( .a(n36449), .b(n36494), .c(n36491), .o(n36495) );
in01f01 g32705 ( .a(n36449), .o(n36496) );
na03f01 g32706 ( .a(n25619), .b(n25605), .c(n25599), .o(n36497) );
oa12f01 g32707 ( .a(n25603), .b(n14332), .c(n13891), .o(n36498) );
no02f01 g32708 ( .a(n36498), .b(n36454), .o(n36499) );
no03f01 g32709 ( .a(n36499), .b(n25618), .c(n25600), .o(n36500) );
oa12f01 g32710 ( .a(n36497), .b(n36500), .c(n25620), .o(n36501) );
no02f01 g32711 ( .a(n36478), .b(n36442), .o(n36502) );
no02f01 g32712 ( .a(n36476), .b(n36427), .o(n36503) );
no03f01 g32713 ( .a(n36503), .b(n36502), .c(n21932), .o(n36504) );
no02f01 g32714 ( .a(n36504), .b(n36472), .o(n36505) );
oa12f01 g32715 ( .a(n21939), .b(n36471), .c(n36466), .o(n36506) );
oa12f01 g32716 ( .a(n21932), .b(n36503), .c(n36502), .o(n36507) );
na02f01 g32717 ( .a(n36507), .b(n36506), .o(n36508) );
ao22f01 g32718 ( .a(n36508), .b(n36475), .c(n36505), .d(n36501), .o(n36509) );
oa12f01 g32719 ( .a(n22098), .b(n36493), .c(n36492), .o(n36510) );
na02f01 g32720 ( .a(n36510), .b(n36509), .o(n36511) );
na03f01 g32721 ( .a(n36489), .b(n36487), .c(n21965), .o(n36512) );
na03f01 g32722 ( .a(n36512), .b(n36511), .c(n36496), .o(n36513) );
na02f01 g32723 ( .a(n36513), .b(n36495), .o(n490) );
no02f01 g32724 ( .a(n29937), .b(n24563), .o(n36515) );
no02f01 g32725 ( .a(n29938), .b(n25005), .o(n36516) );
no02f01 g32726 ( .a(n36516), .b(n36515), .o(n36517) );
no02f01 g32727 ( .a(n29937), .b(n24543), .o(n36518) );
in01f01 g32728 ( .a(n36518), .o(n36519) );
no02f01 g32729 ( .a(n30132), .b(n29943), .o(n36520) );
no02f01 g32730 ( .a(n29938), .b(n24538), .o(n36521) );
in01f01 g32731 ( .a(n36521), .o(n36522) );
na02f01 g32732 ( .a(n36522), .b(n36520), .o(n36523) );
na03f01 g32733 ( .a(n36523), .b(n36519), .c(n36517), .o(n36524) );
ao12f01 g32734 ( .a(n36517), .b(n36523), .c(n36519), .o(n36525) );
in01f01 g32735 ( .a(n36525), .o(n36526) );
na02f01 g32736 ( .a(n36526), .b(n36524), .o(n495) );
no02f01 g32737 ( .a(n9743), .b(n5001), .o(n36528) );
no02f01 g32738 ( .a(n36528), .b(n9745), .o(n36529) );
na02f01 g32739 ( .a(n36529), .b(n9724), .o(n36530) );
no03f01 g32740 ( .a(n6935), .b(n6933), .c(n6924), .o(n36531) );
oa22f01 g32741 ( .a(n36531), .b(n6934), .c(n6932), .d(n6923), .o(n36532) );
in01f01 g32742 ( .a(n6948), .o(n36533) );
in01f01 g32743 ( .a(n6983), .o(n36534) );
na04f01 g32744 ( .a(n36534), .b(n6970), .c(n36533), .d(n36532), .o(n36535) );
ao12f01 g32745 ( .a(n9673), .b(n6987), .c(n36535), .o(n36536) );
oa22f01 g32746 ( .a(n9695), .b(n6934), .c(n9678), .d(n36536), .o(n36537) );
in01f01 g32747 ( .a(n9719), .o(n36538) );
oa12f01 g32748 ( .a(n9722), .b(n36538), .c(n36537), .o(n36539) );
in01f01 g32749 ( .a(n36529), .o(n36540) );
na02f01 g32750 ( .a(n36540), .b(n36539), .o(n36541) );
na02f01 g32751 ( .a(n36541), .b(n36530), .o(n500) );
na02f01 g32752 ( .a(n32732), .b(sin_out_9), .o(n36543) );
no02f01 g32753 ( .a(n35647), .b(n35630), .o(n36544) );
in01f01 g32754 ( .a(n36544), .o(n36545) );
no02f01 g32755 ( .a(n35616), .b(n34287), .o(n36546) );
no02f01 g32756 ( .a(n35617), .b(n34336), .o(n36547) );
no02f01 g32757 ( .a(n36547), .b(n36546), .o(n36548) );
no02f01 g32758 ( .a(n36548), .b(n36545), .o(n36549) );
na02f01 g32759 ( .a(n36548), .b(n36545), .o(n36550) );
in01f01 g32760 ( .a(n36550), .o(n36551) );
no02f01 g32761 ( .a(n36551), .b(n36549), .o(n36552) );
no02f01 g32762 ( .a(n36552), .b(n34307), .o(n36553) );
in01f01 g32763 ( .a(n34303), .o(n36554) );
in01f01 g32764 ( .a(n34316), .o(n36555) );
na02f01 g32765 ( .a(n36555), .b(n34267), .o(n36556) );
na03f01 g32766 ( .a(n34266), .b(n34247), .c(n34304), .o(n36557) );
na03f01 g32767 ( .a(n34266), .b(n34247), .c(delay_sub_ln23_0_unr30_stage10_stallmux_q), .o(n36558) );
in01f01 g32768 ( .a(n34324), .o(n36559) );
na03f01 g32769 ( .a(n36559), .b(n36558), .c(n36557), .o(n36560) );
no02f01 g32770 ( .a(n36555), .b(n34267), .o(n36561) );
oa12f01 g32771 ( .a(n36556), .b(n36561), .c(n36560), .o(n36562) );
na02f01 g32772 ( .a(n36562), .b(n36554), .o(n36563) );
in01f01 g32773 ( .a(n34346), .o(n36564) );
ao12f01 g32774 ( .a(n36564), .b(n36562), .c(n36554), .o(n36565) );
oa22f01 g32775 ( .a(n36565), .b(n34307), .c(n34343), .d(n36563), .o(n36566) );
in01f01 g32776 ( .a(n34369), .o(n36567) );
in01f01 g32777 ( .a(n34393), .o(n36568) );
na02f01 g32778 ( .a(n34383), .b(n34372), .o(n36569) );
na02f01 g32779 ( .a(n36569), .b(n35642), .o(n36570) );
no02f01 g32780 ( .a(n35637), .b(n34287), .o(n36571) );
in01f01 g32781 ( .a(n36571), .o(n36572) );
na02f01 g32782 ( .a(n36572), .b(n35638), .o(n36573) );
no02f01 g32783 ( .a(n36573), .b(n36570), .o(n36574) );
na02f01 g32784 ( .a(n36573), .b(n36570), .o(n36575) );
in01f01 g32785 ( .a(n36575), .o(n36576) );
no02f01 g32786 ( .a(n36576), .b(n36574), .o(n36577) );
in01f01 g32787 ( .a(n36577), .o(n36578) );
no02f01 g32788 ( .a(n36578), .b(n34267), .o(n36579) );
in01f01 g32789 ( .a(n36579), .o(n36580) );
na04f01 g32790 ( .a(n36580), .b(n36568), .c(n36567), .d(n36566), .o(n36581) );
na03f01 g32791 ( .a(n36572), .b(n35642), .c(n35900), .o(n36582) );
in01f01 g32792 ( .a(n36582), .o(n36583) );
no02f01 g32793 ( .a(n35628), .b(n34287), .o(n36584) );
no02f01 g32794 ( .a(n36584), .b(n35630), .o(n36585) );
no02f01 g32795 ( .a(n36585), .b(n36583), .o(n36586) );
na02f01 g32796 ( .a(n36585), .b(n36583), .o(n36587) );
in01f01 g32797 ( .a(n36587), .o(n36588) );
no02f01 g32798 ( .a(n36588), .b(n36586), .o(n36589) );
in01f01 g32799 ( .a(n36589), .o(n36590) );
no02f01 g32800 ( .a(n36590), .b(n34267), .o(n36591) );
ao12f01 g32801 ( .a(n34307), .b(n36589), .c(n36577), .o(n36592) );
ao12f01 g32802 ( .a(n34307), .b(n34390), .c(n34367), .o(n36593) );
no02f01 g32803 ( .a(n36593), .b(n36592), .o(n36594) );
oa12f01 g32804 ( .a(n36594), .b(n36591), .c(n36581), .o(n36595) );
in01f01 g32805 ( .a(n36552), .o(n36596) );
no02f01 g32806 ( .a(n36596), .b(n34267), .o(n36597) );
in01f01 g32807 ( .a(n36597), .o(n36598) );
ao12f01 g32808 ( .a(n36553), .b(n36598), .c(n36595), .o(n36599) );
in01f01 g32809 ( .a(n36599), .o(n36600) );
in01f01 g32810 ( .a(n36547), .o(n36601) );
ao12f01 g32811 ( .a(n36546), .b(n36601), .c(n36544), .o(n36602) );
in01f01 g32812 ( .a(n36602), .o(n36603) );
no02f01 g32813 ( .a(n35609), .b(n34287), .o(n36604) );
no02f01 g32814 ( .a(n35610), .b(n34336), .o(n36605) );
no02f01 g32815 ( .a(n36605), .b(n36604), .o(n36606) );
in01f01 g32816 ( .a(n36606), .o(n36607) );
no02f01 g32817 ( .a(n36607), .b(n36603), .o(n36608) );
no02f01 g32818 ( .a(n36606), .b(n36602), .o(n36609) );
no02f01 g32819 ( .a(n36609), .b(n36608), .o(n36610) );
no02f01 g32820 ( .a(n36610), .b(n34307), .o(n36611) );
in01f01 g32821 ( .a(n36610), .o(n36612) );
no02f01 g32822 ( .a(n36612), .b(n34267), .o(n36613) );
no02f01 g32823 ( .a(n36613), .b(n36611), .o(n36614) );
in01f01 g32824 ( .a(n36614), .o(n36615) );
no02f01 g32825 ( .a(n36615), .b(n36600), .o(n36616) );
no02f01 g32826 ( .a(n36614), .b(n36599), .o(n36617) );
oa12f01 g32827 ( .a(n32734), .b(n36617), .c(n36616), .o(n36618) );
na02f01 g32828 ( .a(n36618), .b(n36543), .o(n505) );
in01f01 g32829 ( .a(n25355), .o(n36620) );
in01f01 g32830 ( .a(n25377), .o(n36621) );
no02f01 g32831 ( .a(n25369), .b(n24980), .o(n36622) );
no02f01 g32832 ( .a(n25367), .b(n25366), .o(n36623) );
no02f01 g32833 ( .a(n36623), .b(n36622), .o(n36624) );
in01f01 g32834 ( .a(n25376), .o(n36625) );
in01f01 g32835 ( .a(n25378), .o(n36626) );
na03f01 g32836 ( .a(n24979), .b(n24975), .c(n25365), .o(n36627) );
na02f01 g32837 ( .a(n36627), .b(n36626), .o(n36628) );
in01f01 g32838 ( .a(n25391), .o(n36629) );
in01f01 g32839 ( .a(n25402), .o(n36630) );
oa12f01 g32840 ( .a(n24476), .b(n25410), .c(n25409), .o(n36631) );
na03f01 g32841 ( .a(n25404), .b(n25403), .c(n24449), .o(n36632) );
in01f01 g32842 ( .a(n25414), .o(n36633) );
ao12f01 g32843 ( .a(n36633), .b(n36632), .c(n36631), .o(n36634) );
no02f01 g32844 ( .a(n25448), .b(n25445), .o(n36635) );
ao12f01 g32845 ( .a(n36635), .b(n25458), .c(n25449), .o(n36636) );
in01f01 g32846 ( .a(n25461), .o(n36637) );
oa12f01 g32847 ( .a(n36637), .b(n36636), .c(n36634), .o(n36638) );
ao12f01 g32848 ( .a(n24477), .b(n24491), .c(n25394), .o(n36639) );
in01f01 g32849 ( .a(n25395), .o(n36640) );
oa12f01 g32850 ( .a(n25400), .b(n36640), .c(n36639), .o(n36641) );
ao12f01 g32851 ( .a(n36630), .b(n36641), .c(n36638), .o(n36642) );
oa12f01 g32852 ( .a(n25381), .b(n24970), .c(n25384), .o(n36643) );
in01f01 g32853 ( .a(n25385), .o(n36644) );
in01f01 g32854 ( .a(n25390), .o(n36645) );
ao12f01 g32855 ( .a(n36645), .b(n36644), .c(n36643), .o(n36646) );
oa12f01 g32856 ( .a(n36629), .b(n36646), .c(n36642), .o(n36647) );
no03f01 g32857 ( .a(n24494), .b(n24973), .c(n24432), .o(n36648) );
no02f01 g32858 ( .a(n25467), .b(n24493), .o(n36649) );
oa12f01 g32859 ( .a(n25472), .b(n36649), .c(n36648), .o(n36650) );
na02f01 g32860 ( .a(n36650), .b(n36647), .o(n36651) );
in01f01 g32861 ( .a(n25480), .o(n36652) );
ao12f01 g32862 ( .a(n36628), .b(n36652), .c(n36651), .o(n36653) );
ao12f01 g32863 ( .a(n25479), .b(n25476), .c(n36651), .o(n36654) );
oa22f01 g32864 ( .a(n36654), .b(n36653), .c(n36625), .d(n36624), .o(n36655) );
oa22f01 g32865 ( .a(n24520), .b(n24506), .c(n24519), .d(n24965), .o(n36656) );
na04f01 g32866 ( .a(n24991), .b(n24990), .c(n24985), .d(n24420), .o(n36657) );
in01f01 g32867 ( .a(n25362), .o(n36658) );
ao12f01 g32868 ( .a(n36658), .b(n36657), .c(n36656), .o(n36659) );
ao12f01 g32869 ( .a(n36659), .b(n36655), .c(n36621), .o(n36660) );
oa12f01 g32870 ( .a(n25354), .b(n25349), .c(n25347), .o(n36661) );
oa12f01 g32871 ( .a(n36661), .b(n36660), .c(n25363), .o(n36662) );
oa22f01 g32872 ( .a(n25336), .b(n24989), .c(n25335), .d(n25334), .o(n36663) );
in01f01 g32873 ( .a(n25337), .o(n36664) );
ao12f01 g32874 ( .a(n25341), .b(n36664), .c(n36663), .o(n36665) );
ao12f01 g32875 ( .a(n36665), .b(n36662), .c(n36620), .o(n36666) );
no02f01 g32876 ( .a(n36666), .b(n25343), .o(n36667) );
no02f01 g32877 ( .a(n25518), .b(n25504), .o(n36668) );
no02f01 g32878 ( .a(n36668), .b(n36667), .o(n36669) );
na02f01 g32879 ( .a(n36668), .b(n36667), .o(n36670) );
in01f01 g32880 ( .a(n36670), .o(n36671) );
no02f01 g32881 ( .a(n36671), .b(n36669), .o(n36672) );
na02f01 g32882 ( .a(n36672), .b(n6037), .o(n36673) );
in01f01 g32883 ( .a(n36672), .o(n4156) );
na02f01 g32884 ( .a(n4156), .b(n5873), .o(n36675) );
na02f01 g32885 ( .a(n36675), .b(n36673), .o(n509) );
in01f01 g32886 ( .a(n14160), .o(n36677) );
no02f01 g32887 ( .a(n14190), .b(n14174), .o(n36678) );
no02f01 g32888 ( .a(n36678), .b(n36677), .o(n36679) );
na02f01 g32889 ( .a(n36678), .b(n36677), .o(n36680) );
in01f01 g32890 ( .a(n36680), .o(n36681) );
no02f01 g32891 ( .a(n36681), .b(n36679), .o(n36682) );
na02f01 g32892 ( .a(n36682), .b(n2589), .o(n36683) );
in01f01 g32893 ( .a(n36682), .o(n4256) );
na02f01 g32894 ( .a(n4256), .b(n4116), .o(n36685) );
na02f01 g32895 ( .a(n36685), .b(n36683), .o(n514) );
in01f01 g32896 ( .a(n28064), .o(n36687) );
no02f01 g32897 ( .a(n29491), .b(n36687), .o(n36688) );
no02f01 g32898 ( .a(n29460), .b(n28064), .o(n36689) );
no02f01 g32899 ( .a(n36689), .b(n36688), .o(n36690) );
ao12f01 g32900 ( .a(n29460), .b(n28477), .c(n28026), .o(n36691) );
no02f01 g32901 ( .a(n28496), .b(n27983), .o(n36692) );
no02f01 g32902 ( .a(n36692), .b(n29491), .o(n36693) );
ao12f01 g32903 ( .a(n36693), .b(n29624), .c(n29632), .o(n36694) );
no02f01 g32904 ( .a(n29491), .b(n28018), .o(n36695) );
no02f01 g32905 ( .a(n29491), .b(n28003), .o(n36696) );
no02f01 g32906 ( .a(n36696), .b(n36695), .o(n36697) );
ao12f01 g32907 ( .a(n29460), .b(n28496), .c(n27983), .o(n36698) );
ao12f01 g32908 ( .a(n29460), .b(n28053), .c(n28513), .o(n36699) );
no02f01 g32909 ( .a(n36699), .b(n36698), .o(n36700) );
in01f01 g32910 ( .a(n36700), .o(n36701) );
ao12f01 g32911 ( .a(n36701), .b(n36697), .c(n36694), .o(n36702) );
no02f01 g32912 ( .a(n29491), .b(n28565), .o(n36703) );
no02f01 g32913 ( .a(n29491), .b(n28036), .o(n36704) );
no02f01 g32914 ( .a(n36704), .b(n36703), .o(n36705) );
in01f01 g32915 ( .a(n36705), .o(n36706) );
no02f01 g32916 ( .a(n36706), .b(n36702), .o(n36707) );
no02f01 g32917 ( .a(n29460), .b(n28461), .o(n36708) );
no03f01 g32918 ( .a(n36708), .b(n36707), .c(n36691), .o(n36709) );
no02f01 g32919 ( .a(n29491), .b(n28462), .o(n36710) );
oa12f01 g32920 ( .a(n36690), .b(n36710), .c(n36709), .o(n36711) );
in01f01 g32921 ( .a(n36690), .o(n36712) );
in01f01 g32922 ( .a(n36691), .o(n36713) );
oa22f01 g32923 ( .a(n36692), .b(n29491), .c(n29625), .d(n29622), .o(n36714) );
in01f01 g32924 ( .a(n36697), .o(n36715) );
oa12f01 g32925 ( .a(n36700), .b(n36715), .c(n36714), .o(n36716) );
na02f01 g32926 ( .a(n36705), .b(n36716), .o(n36717) );
in01f01 g32927 ( .a(n36708), .o(n36718) );
na03f01 g32928 ( .a(n36718), .b(n36717), .c(n36713), .o(n36719) );
in01f01 g32929 ( .a(n36710), .o(n36720) );
na03f01 g32930 ( .a(n36720), .b(n36719), .c(n36712), .o(n36721) );
na02f01 g32931 ( .a(n36721), .b(n36711), .o(n36722) );
no02f01 g32932 ( .a(n36722), .b(n29430), .o(n36723) );
ao12f01 g32933 ( .a(n36712), .b(n36720), .c(n36719), .o(n36724) );
no03f01 g32934 ( .a(n36710), .b(n36709), .c(n36690), .o(n36725) );
no02f01 g32935 ( .a(n36725), .b(n36724), .o(n36726) );
no02f01 g32936 ( .a(n36726), .b(n29639), .o(n36727) );
no02f01 g32937 ( .a(n36727), .b(n36723), .o(n36728) );
in01f01 g32938 ( .a(n36728), .o(n36729) );
na02f01 g32939 ( .a(n36717), .b(n36713), .o(n36730) );
no02f01 g32940 ( .a(n36710), .b(n36708), .o(n36731) );
in01f01 g32941 ( .a(n36731), .o(n36732) );
na02f01 g32942 ( .a(n36732), .b(n36730), .o(n36733) );
no02f01 g32943 ( .a(n36707), .b(n36691), .o(n36734) );
na02f01 g32944 ( .a(n36731), .b(n36734), .o(n36735) );
na02f01 g32945 ( .a(n36735), .b(n36733), .o(n36736) );
no02f01 g32946 ( .a(n36736), .b(n29430), .o(n36737) );
in01f01 g32947 ( .a(n36737), .o(n36738) );
no02f01 g32948 ( .a(n29663), .b(n29636), .o(n36739) );
in01f01 g32949 ( .a(n36739), .o(n36740) );
no02f01 g32950 ( .a(n29460), .b(n28053), .o(n36741) );
no02f01 g32951 ( .a(n36741), .b(n36695), .o(n36742) );
no02f01 g32952 ( .a(n29460), .b(n28513), .o(n36743) );
no03f01 g32953 ( .a(n36743), .b(n36698), .c(n36694), .o(n36744) );
no03f01 g32954 ( .a(n36744), .b(n36742), .c(n36696), .o(n36745) );
in01f01 g32955 ( .a(n36696), .o(n36746) );
in01f01 g32956 ( .a(n36742), .o(n36747) );
in01f01 g32957 ( .a(n36698), .o(n36748) );
in01f01 g32958 ( .a(n36743), .o(n36749) );
na03f01 g32959 ( .a(n36749), .b(n36748), .c(n36714), .o(n36750) );
ao12f01 g32960 ( .a(n36747), .b(n36750), .c(n36746), .o(n36751) );
no02f01 g32961 ( .a(n36751), .b(n36745), .o(n36752) );
na02f01 g32962 ( .a(n36752), .b(n29639), .o(n36753) );
in01f01 g32963 ( .a(n36753), .o(n36754) );
no02f01 g32964 ( .a(n36743), .b(n36696), .o(n36755) );
ao12f01 g32965 ( .a(n36755), .b(n36748), .c(n36714), .o(n36756) );
in01f01 g32966 ( .a(n36755), .o(n36757) );
no03f01 g32967 ( .a(n36757), .b(n36698), .c(n36694), .o(n36758) );
no02f01 g32968 ( .a(n36758), .b(n36756), .o(n36759) );
in01f01 g32969 ( .a(n36759), .o(n36760) );
no02f01 g32970 ( .a(n36760), .b(n29430), .o(n36761) );
no03f01 g32971 ( .a(n36761), .b(n36754), .c(n36740), .o(n36762) );
no02f01 g32972 ( .a(n29460), .b(n28477), .o(n36763) );
no02f01 g32973 ( .a(n36763), .b(n36704), .o(n36764) );
in01f01 g32974 ( .a(n36764), .o(n36765) );
no02f01 g32975 ( .a(n29460), .b(n28026), .o(n36766) );
no02f01 g32976 ( .a(n36703), .b(n36702), .o(n36767) );
no03f01 g32977 ( .a(n36767), .b(n36766), .c(n36765), .o(n36768) );
in01f01 g32978 ( .a(n36768), .o(n36769) );
oa12f01 g32979 ( .a(n36765), .b(n36767), .c(n36766), .o(n36770) );
na02f01 g32980 ( .a(n36770), .b(n36769), .o(n36771) );
no02f01 g32981 ( .a(n36766), .b(n36703), .o(n36772) );
no02f01 g32982 ( .a(n36772), .b(n36702), .o(n36773) );
in01f01 g32983 ( .a(n36773), .o(n36774) );
na02f01 g32984 ( .a(n36772), .b(n36702), .o(n36775) );
na02f01 g32985 ( .a(n36775), .b(n36774), .o(n36776) );
ao12f01 g32986 ( .a(n29430), .b(n36776), .c(n36771), .o(n36777) );
in01f01 g32987 ( .a(n36777), .o(n36778) );
na04f01 g32988 ( .a(n36778), .b(n36762), .c(n29614), .d(n29721), .o(n36779) );
oa12f01 g32989 ( .a(n29430), .b(n29662), .c(n29635), .o(n36780) );
na02f01 g32990 ( .a(n36780), .b(n29645), .o(n36781) );
ao12f01 g32991 ( .a(n29639), .b(n36759), .c(n36752), .o(n36782) );
no02f01 g32992 ( .a(n36782), .b(n36781), .o(n36783) );
oa12f01 g32993 ( .a(n29430), .b(n36776), .c(n36771), .o(n36784) );
na02f01 g32994 ( .a(n36784), .b(n36783), .o(n36785) );
in01f01 g32995 ( .a(n36785), .o(n36786) );
no02f01 g32996 ( .a(n36731), .b(n36734), .o(n36787) );
no02f01 g32997 ( .a(n36732), .b(n36730), .o(n36788) );
no02f01 g32998 ( .a(n36788), .b(n36787), .o(n36789) );
no02f01 g32999 ( .a(n36789), .b(n29639), .o(n36790) );
in01f01 g33000 ( .a(n36790), .o(n36791) );
na03f01 g33001 ( .a(n36791), .b(n36786), .c(n36779), .o(n36792) );
na03f01 g33002 ( .a(n36792), .b(n36738), .c(n36729), .o(n36793) );
in01f01 g33003 ( .a(n36762), .o(n36794) );
no04f01 g33004 ( .a(n36777), .b(n36794), .c(n29615), .d(n29578), .o(n36795) );
no03f01 g33005 ( .a(n36790), .b(n36785), .c(n36795), .o(n36796) );
oa12f01 g33006 ( .a(n36728), .b(n36796), .c(n36737), .o(n36797) );
na03f01 g33007 ( .a(n36797), .b(n36793), .c(n_27923), .o(n36798) );
no03f01 g33008 ( .a(n36796), .b(n36737), .c(n36728), .o(n36799) );
ao12f01 g33009 ( .a(n36729), .b(n36792), .c(n36738), .o(n36800) );
oa12f01 g33010 ( .a(n34420), .b(n36800), .c(n36799), .o(n36801) );
na02f01 g33011 ( .a(n36801), .b(n36798), .o(n519) );
no02f01 g33012 ( .a(n31664), .b(n30597), .o(n36803) );
no02f01 g33013 ( .a(n31666), .b(n30568), .o(n36804) );
no02f01 g33014 ( .a(n36804), .b(n36803), .o(n36805) );
in01f01 g33015 ( .a(n36805), .o(n36806) );
no02f01 g33016 ( .a(n31666), .b(n31011), .o(n36807) );
no02f01 g33017 ( .a(n36807), .b(n31667), .o(n36808) );
in01f01 g33018 ( .a(n36808), .o(n36809) );
no02f01 g33019 ( .a(n36809), .b(n32031), .o(n36810) );
no02f01 g33020 ( .a(n31666), .b(n30441), .o(n36811) );
no02f01 g33021 ( .a(n31666), .b(n30543), .o(n36812) );
no02f01 g33022 ( .a(n36812), .b(n36811), .o(n36813) );
in01f01 g33023 ( .a(n30441), .o(n36814) );
ao12f01 g33024 ( .a(n31664), .b(n30542), .c(n36814), .o(n36815) );
ao12f01 g33025 ( .a(n31664), .b(n30535), .c(n30525), .o(n36816) );
no02f01 g33026 ( .a(n36816), .b(n36815), .o(n36817) );
in01f01 g33027 ( .a(n36817), .o(n36818) );
ao12f01 g33028 ( .a(n36818), .b(n36813), .c(n36810), .o(n36819) );
no02f01 g33029 ( .a(n31666), .b(n30575), .o(n36820) );
no02f01 g33030 ( .a(n36820), .b(n36819), .o(n36821) );
no02f01 g33031 ( .a(n31664), .b(n30574), .o(n36822) );
no02f01 g33032 ( .a(n36822), .b(n36821), .o(n36823) );
in01f01 g33033 ( .a(n36823), .o(n36824) );
no02f01 g33034 ( .a(n36824), .b(n36806), .o(n36825) );
no02f01 g33035 ( .a(n36823), .b(n36805), .o(n36826) );
no02f01 g33036 ( .a(n36826), .b(n36825), .o(n36827) );
no02f01 g33037 ( .a(n36827), .b(n31607), .o(n36828) );
in01f01 g33038 ( .a(n36827), .o(n36829) );
no02f01 g33039 ( .a(n36829), .b(n31606), .o(n36830) );
no02f01 g33040 ( .a(n36830), .b(n36828), .o(n36831) );
in01f01 g33041 ( .a(n36831), .o(n36832) );
in01f01 g33042 ( .a(n36819), .o(n36833) );
no02f01 g33043 ( .a(n36822), .b(n36820), .o(n36834) );
in01f01 g33044 ( .a(n36834), .o(n36835) );
no02f01 g33045 ( .a(n36835), .b(n36833), .o(n36836) );
no02f01 g33046 ( .a(n36834), .b(n36819), .o(n36837) );
no02f01 g33047 ( .a(n36837), .b(n36836), .o(n36838) );
in01f01 g33048 ( .a(n36838), .o(n36839) );
no02f01 g33049 ( .a(n36839), .b(n31606), .o(n36840) );
in01f01 g33050 ( .a(n36840), .o(n36841) );
in01f01 g33051 ( .a(n36816), .o(n36842) );
oa12f01 g33052 ( .a(n36842), .b(n36809), .c(n32031), .o(n36843) );
no02f01 g33053 ( .a(n31664), .b(n30542), .o(n36844) );
no02f01 g33054 ( .a(n36844), .b(n36812), .o(n36845) );
in01f01 g33055 ( .a(n36845), .o(n36846) );
na02f01 g33056 ( .a(n36846), .b(n36843), .o(n36847) );
no02f01 g33057 ( .a(n36846), .b(n36843), .o(n36848) );
in01f01 g33058 ( .a(n36848), .o(n36849) );
na02f01 g33059 ( .a(n36849), .b(n36847), .o(n36850) );
no02f01 g33060 ( .a(n36850), .b(n31606), .o(n36851) );
in01f01 g33061 ( .a(n36851), .o(n36852) );
no02f01 g33062 ( .a(n31664), .b(n36814), .o(n36853) );
no02f01 g33063 ( .a(n36853), .b(n36811), .o(n36854) );
in01f01 g33064 ( .a(n36854), .o(n36855) );
no02f01 g33065 ( .a(n36843), .b(n36844), .o(n36856) );
no02f01 g33066 ( .a(n36856), .b(n36812), .o(n36857) );
no02f01 g33067 ( .a(n36857), .b(n36855), .o(n36858) );
in01f01 g33068 ( .a(n36858), .o(n36859) );
na02f01 g33069 ( .a(n36857), .b(n36855), .o(n36860) );
na02f01 g33070 ( .a(n36860), .b(n36859), .o(n36861) );
no02f01 g33071 ( .a(n36861), .b(n31606), .o(n36862) );
no02f01 g33072 ( .a(n31664), .b(n30535), .o(n36863) );
no02f01 g33073 ( .a(n36863), .b(n36807), .o(n36864) );
in01f01 g33074 ( .a(n31667), .o(n36865) );
ao12f01 g33075 ( .a(n31665), .b(n31977), .c(n36865), .o(n36866) );
na02f01 g33076 ( .a(n36866), .b(n36864), .o(n36867) );
in01f01 g33077 ( .a(n36864), .o(n36868) );
no02f01 g33078 ( .a(n32031), .b(n31667), .o(n36869) );
oa12f01 g33079 ( .a(n36868), .b(n36869), .c(n31665), .o(n36870) );
na02f01 g33080 ( .a(n36870), .b(n36867), .o(n36871) );
ao12f01 g33081 ( .a(n31606), .b(n36871), .c(n32037), .o(n36872) );
no02f01 g33082 ( .a(n36872), .b(n36862), .o(n36873) );
na02f01 g33083 ( .a(n36873), .b(n36852), .o(n36874) );
in01f01 g33084 ( .a(n36874), .o(n36875) );
na04f01 g33085 ( .a(n36875), .b(n32436), .c(n32430), .d(n32427), .o(n36876) );
in01f01 g33086 ( .a(n36871), .o(n36877) );
ao12f01 g33087 ( .a(n31607), .b(n36877), .c(n32033), .o(n36878) );
in01f01 g33088 ( .a(n36847), .o(n36879) );
no02f01 g33089 ( .a(n36848), .b(n36879), .o(n36880) );
in01f01 g33090 ( .a(n36860), .o(n36881) );
no02f01 g33091 ( .a(n36881), .b(n36858), .o(n36882) );
ao12f01 g33092 ( .a(n31607), .b(n36882), .c(n36880), .o(n36883) );
no02f01 g33093 ( .a(n36883), .b(n36878), .o(n36884) );
na02f01 g33094 ( .a(n36884), .b(n32130), .o(n36885) );
in01f01 g33095 ( .a(n36885), .o(n36886) );
no02f01 g33096 ( .a(n36838), .b(n31607), .o(n36887) );
in01f01 g33097 ( .a(n36887), .o(n36888) );
na03f01 g33098 ( .a(n36888), .b(n36886), .c(n36876), .o(n36889) );
na03f01 g33099 ( .a(n36889), .b(n36841), .c(n36832), .o(n36890) );
no04f01 g33100 ( .a(n36874), .b(n32495), .c(n32494), .d(n32493), .o(n36891) );
no03f01 g33101 ( .a(n36887), .b(n36885), .c(n36891), .o(n36892) );
oa12f01 g33102 ( .a(n36831), .b(n36892), .c(n36840), .o(n36893) );
na02f01 g33103 ( .a(n36893), .b(n36890), .o(n524) );
no03f01 g33104 ( .a(n4799), .b(n4775), .c(n4756_1), .o(n36895) );
in01f01 g33105 ( .a(n36895), .o(n36896) );
no02f01 g33106 ( .a(n7069), .b(n4340), .o(n36897) );
no02f01 g33107 ( .a(n7086), .b(n7077), .o(n36898) );
no02f01 g33108 ( .a(n36898), .b(n4340), .o(n36899) );
no04f01 g33109 ( .a(n36899), .b(n36897), .c(n36896), .d(n4727_1), .o(n36900) );
ao12f01 g33110 ( .a(n4344_1), .b(n4797), .c(n4773), .o(n36901) );
no02f01 g33111 ( .a(n36901), .b(n4757), .o(n36902) );
ao12f01 g33112 ( .a(n4344_1), .b(n7086), .c(n7077), .o(n36903) );
oa12f01 g33113 ( .a(n4340), .b(n36903), .c(n7069), .o(n36904) );
na02f01 g33114 ( .a(n36904), .b(n36902), .o(n36905) );
no02f01 g33115 ( .a(n7060), .b(n4344_1), .o(n36906) );
no02f01 g33116 ( .a(n7091), .b(n4340), .o(n36907) );
no02f01 g33117 ( .a(n36907), .b(n36906), .o(n36908) );
in01f01 g33118 ( .a(n36908), .o(n36909) );
no03f01 g33119 ( .a(n36909), .b(n36905), .c(n36900), .o(n36910) );
no02f01 g33120 ( .a(n36905), .b(n36900), .o(n36911) );
no02f01 g33121 ( .a(n36908), .b(n36911), .o(n36912) );
no02f01 g33122 ( .a(n36912), .b(n36910), .o(n36913) );
no02f01 g33123 ( .a(n36913), .b(n3789), .o(n36914) );
na02f01 g33124 ( .a(n36902), .b(n4701), .o(n36915) );
ao12f01 g33125 ( .a(n36915), .b(n36895), .c(n4725), .o(n36916) );
in01f01 g33126 ( .a(n36916), .o(n36917) );
no02f01 g33127 ( .a(n7077), .b(n4344_1), .o(n36918) );
no02f01 g33128 ( .a(n7078), .b(n4340), .o(n36919) );
no02f01 g33129 ( .a(n36919), .b(n36918), .o(n36920) );
in01f01 g33130 ( .a(n36920), .o(n36921) );
no02f01 g33131 ( .a(n36921), .b(n36917), .o(n36922) );
na02f01 g33132 ( .a(n36921), .b(n36917), .o(n36923) );
in01f01 g33133 ( .a(n36923), .o(n36924) );
no02f01 g33134 ( .a(n36924), .b(n36922), .o(n36925) );
no02f01 g33135 ( .a(n36925), .b(n3789), .o(n36926) );
no03f01 g33136 ( .a(n36926), .b(n4808), .c(n4787), .o(n36927) );
no02f01 g33137 ( .a(n7086), .b(n4344_1), .o(n36928) );
no02f01 g33138 ( .a(n7095), .b(n4340), .o(n36929) );
no02f01 g33139 ( .a(n36929), .b(n36928), .o(n36930) );
in01f01 g33140 ( .a(n36930), .o(n36931) );
in01f01 g33141 ( .a(n36918), .o(n36932) );
ao12f01 g33142 ( .a(n36919), .b(n36916), .c(n36932), .o(n36933) );
no02f01 g33143 ( .a(n36933), .b(n36931), .o(n36934) );
na02f01 g33144 ( .a(n36933), .b(n36931), .o(n36935) );
in01f01 g33145 ( .a(n36935), .o(n36936) );
no02f01 g33146 ( .a(n36936), .b(n36934), .o(n36937) );
no02f01 g33147 ( .a(n36937), .b(n3789), .o(n36938) );
in01f01 g33148 ( .a(n36938), .o(n36939) );
na02f01 g33149 ( .a(n36939), .b(n36927), .o(n36940) );
no02f01 g33150 ( .a(n36937), .b(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n36941) );
in01f01 g33151 ( .a(n36941), .o(n36942) );
no02f01 g33152 ( .a(n36916), .b(n36899), .o(n36943) );
no02f01 g33153 ( .a(n36943), .b(n36903), .o(n36944) );
no02f01 g33154 ( .a(n7068), .b(n4344_1), .o(n36945) );
no02f01 g33155 ( .a(n36945), .b(n36897), .o(n36946) );
na02f01 g33156 ( .a(n36946), .b(n36944), .o(n36947) );
in01f01 g33157 ( .a(n36947), .o(n36948) );
no02f01 g33158 ( .a(n36946), .b(n36944), .o(n36949) );
no02f01 g33159 ( .a(n36949), .b(n36948), .o(n36950) );
na02f01 g33160 ( .a(n36950), .b(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n36951) );
no02f01 g33161 ( .a(n36950), .b(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n36952) );
in01f01 g33162 ( .a(n36952), .o(n36953) );
na02f01 g33163 ( .a(n36953), .b(n36951), .o(n36954) );
in01f01 g33164 ( .a(n36954), .o(n36955) );
na03f01 g33165 ( .a(n36955), .b(n36942), .c(n36940), .o(n36956) );
ao12f01 g33166 ( .a(delay_sub_ln23_0_unr22_stage8_stallmux_q), .b(n36925), .c(n4807), .o(n36957) );
in01f01 g33167 ( .a(n36957), .o(n36958) );
oa12f01 g33168 ( .a(n36958), .b(n36955), .c(n36940), .o(n36959) );
ao12f01 g33169 ( .a(n36959), .b(n36956), .c(n3789), .o(n36960) );
no02f01 g33170 ( .a(n36913), .b(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n36961) );
no02f01 g33171 ( .a(n36961), .b(n36960), .o(n36962) );
no02f01 g33172 ( .a(n36962), .b(n36914), .o(n36963) );
no02f01 g33173 ( .a(n7241), .b(n7164), .o(n36964) );
no02f01 g33174 ( .a(n7242), .b(n7205), .o(n36965) );
no02f01 g33175 ( .a(n36965), .b(n36964), .o(n36966) );
no02f01 g33176 ( .a(n36966), .b(n7232), .o(n36967) );
na02f01 g33177 ( .a(n36966), .b(n7232), .o(n36968) );
in01f01 g33178 ( .a(n36968), .o(n36969) );
no02f01 g33179 ( .a(n36969), .b(n36967), .o(n36970) );
no02f01 g33180 ( .a(n36970), .b(n36963), .o(n36971) );
in01f01 g33181 ( .a(n36963), .o(n36972) );
no02f01 g33182 ( .a(n36957), .b(n36941), .o(n36973) );
na02f01 g33183 ( .a(n36973), .b(n36940), .o(n36974) );
no02f01 g33184 ( .a(n36950), .b(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n36975) );
no02f01 g33185 ( .a(n36950), .b(n3789), .o(n36976) );
no02f01 g33186 ( .a(n36976), .b(n36975), .o(n36977) );
in01f01 g33187 ( .a(n36977), .o(n36978) );
na02f01 g33188 ( .a(n36978), .b(n36974), .o(n36979) );
no02f01 g33189 ( .a(n36978), .b(n36974), .o(n36980) );
in01f01 g33190 ( .a(n36980), .o(n36981) );
na02f01 g33191 ( .a(n36981), .b(n36979), .o(n36982) );
no03f01 g33192 ( .a(n7355), .b(n7154), .c(n7126), .o(n36983) );
ao12f01 g33193 ( .a(n7354), .b(n7155), .c(n7342), .o(n36984) );
no02f01 g33194 ( .a(n36984), .b(n36983), .o(n36985) );
no02f01 g33195 ( .a(n36985), .b(n36982), .o(n36986) );
in01f01 g33196 ( .a(n36986), .o(n36987) );
no02f01 g33197 ( .a(n36957), .b(n36927), .o(n36988) );
no02f01 g33198 ( .a(n36941), .b(n36938), .o(n36989) );
na02f01 g33199 ( .a(n36989), .b(n36988), .o(n36990) );
no02f01 g33200 ( .a(n36989), .b(n36988), .o(n36991) );
in01f01 g33201 ( .a(n36991), .o(n36992) );
na02f01 g33202 ( .a(n36992), .b(n36990), .o(n36993) );
no03f01 g33203 ( .a(n7153), .b(n7352), .c(n7134), .o(n36994) );
ao12f01 g33204 ( .a(n7150), .b(n7353), .c(n7135), .o(n36995) );
no02f01 g33205 ( .a(n36995), .b(n36994), .o(n36996) );
no02f01 g33206 ( .a(n36996), .b(n36993), .o(n36997) );
no02f01 g33207 ( .a(n36925), .b(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n36998) );
no02f01 g33208 ( .a(n36998), .b(n36926), .o(n36999) );
in01f01 g33209 ( .a(n36999), .o(n37000) );
no02f01 g33210 ( .a(n4808), .b(n4787), .o(n37001) );
no03f01 g33211 ( .a(n37001), .b(n37000), .c(n4809), .o(n37002) );
in01f01 g33212 ( .a(n37002), .o(n37003) );
oa12f01 g33213 ( .a(n37000), .b(n37001), .c(n4809), .o(n37004) );
no03f01 g33214 ( .a(n7351), .b(n7148), .c(n7146), .o(n37005) );
ao12f01 g33215 ( .a(n7347), .b(n7149), .c(n7343), .o(n37006) );
no02f01 g33216 ( .a(n37006), .b(n37005), .o(n37007) );
in01f01 g33217 ( .a(n37007), .o(n37008) );
na03f01 g33218 ( .a(n37008), .b(n37004), .c(n37003), .o(n37009) );
ao12f01 g33219 ( .a(n4891), .b(n4971), .c(n4974), .o(n37010) );
ao12f01 g33220 ( .a(n37008), .b(n37004), .c(n37003), .o(n37011) );
oa12f01 g33221 ( .a(n37009), .b(n37011), .c(n37010), .o(n37012) );
na02f01 g33222 ( .a(n36996), .b(n36993), .o(n37013) );
ao12f01 g33223 ( .a(n36997), .b(n37013), .c(n37012), .o(n37014) );
in01f01 g33224 ( .a(n36985), .o(n37015) );
ao12f01 g33225 ( .a(n37015), .b(n36981), .c(n36979), .o(n37016) );
oa12f01 g33226 ( .a(n36987), .b(n37016), .c(n37014), .o(n37017) );
no02f01 g33227 ( .a(n36961), .b(n36914), .o(n37018) );
na02f01 g33228 ( .a(n37018), .b(n36960), .o(n37019) );
na02f01 g33229 ( .a(n36956), .b(n3789), .o(n37020) );
in01f01 g33230 ( .a(n36959), .o(n37021) );
na02f01 g33231 ( .a(n37021), .b(n37020), .o(n37022) );
in01f01 g33232 ( .a(n37018), .o(n37023) );
na02f01 g33233 ( .a(n37023), .b(n37022), .o(n37024) );
na02f01 g33234 ( .a(n37024), .b(n37019), .o(n37025) );
no02f01 g33235 ( .a(n7158), .b(n7115), .o(n37026) );
no02f01 g33236 ( .a(n37026), .b(n7156), .o(n37027) );
na02f01 g33237 ( .a(n37026), .b(n7156), .o(n37028) );
in01f01 g33238 ( .a(n37028), .o(n37029) );
no02f01 g33239 ( .a(n37029), .b(n37027), .o(n37030) );
na02f01 g33240 ( .a(n37030), .b(n37025), .o(n37031) );
no02f01 g33241 ( .a(n7160), .b(n7337), .o(n37032) );
no02f01 g33242 ( .a(n37032), .b(n7358), .o(n37033) );
na02f01 g33243 ( .a(n37032), .b(n7358), .o(n37034) );
in01f01 g33244 ( .a(n37034), .o(n37035) );
no02f01 g33245 ( .a(n37035), .b(n37033), .o(n37036) );
na02f01 g33246 ( .a(n37036), .b(n36963), .o(n37037) );
na03f01 g33247 ( .a(n37037), .b(n37031), .c(n37017), .o(n37038) );
no02f01 g33248 ( .a(n37030), .b(n37025), .o(n37039) );
no02f01 g33249 ( .a(n37036), .b(n36963), .o(n37040) );
oa12f01 g33250 ( .a(n37037), .b(n37040), .c(n37039), .o(n37041) );
na02f01 g33251 ( .a(n37041), .b(n37038), .o(n37042) );
no02f01 g33252 ( .a(n7179), .b(n7164), .o(n37043) );
in01f01 g33253 ( .a(n7183), .o(n37044) );
no03f01 g33254 ( .a(n37044), .b(n37043), .c(n7360), .o(n37045) );
no02f01 g33255 ( .a(n37044), .b(n37043), .o(n37046) );
no02f01 g33256 ( .a(n37046), .b(n7161), .o(n37047) );
no02f01 g33257 ( .a(n37047), .b(n37045), .o(n37048) );
no02f01 g33258 ( .a(n37048), .b(n36963), .o(n37049) );
ao12f01 g33259 ( .a(n37043), .b(n7183), .c(n7360), .o(n37050) );
in01f01 g33260 ( .a(n7182), .o(n37051) );
no02f01 g33261 ( .a(n7172), .b(n7164), .o(n37052) );
no02f01 g33262 ( .a(n37052), .b(n37051), .o(n37053) );
no02f01 g33263 ( .a(n37053), .b(n37050), .o(n37054) );
na02f01 g33264 ( .a(n37053), .b(n37050), .o(n37055) );
in01f01 g33265 ( .a(n37055), .o(n37056) );
no02f01 g33266 ( .a(n37056), .b(n37054), .o(n37057) );
in01f01 g33267 ( .a(n37057), .o(n37058) );
no02f01 g33268 ( .a(n37058), .b(n37049), .o(n37059) );
na03f01 g33269 ( .a(n37059), .b(n37041), .c(n37038), .o(n37060) );
no02f01 g33270 ( .a(n37057), .b(n37048), .o(n37061) );
ao22f01 g33271 ( .a(n37061), .b(n37042), .c(n37060), .d(n36972), .o(n37062) );
in01f01 g33272 ( .a(n7203), .o(n37063) );
no02f01 g33273 ( .a(n7202), .b(n7164), .o(n37064) );
no02f01 g33274 ( .a(n37064), .b(n37063), .o(n37065) );
in01f01 g33275 ( .a(n37065), .o(n37066) );
no02f01 g33276 ( .a(n37066), .b(n7185), .o(n37067) );
no02f01 g33277 ( .a(n37065), .b(n7362), .o(n37068) );
no02f01 g33278 ( .a(n37068), .b(n37067), .o(n37069) );
in01f01 g33279 ( .a(n37069), .o(n37070) );
oa12f01 g33280 ( .a(n7203), .b(n37064), .c(n7185), .o(n37071) );
in01f01 g33281 ( .a(n7196), .o(n37072) );
no02f01 g33282 ( .a(n7195), .b(n7164), .o(n37073) );
no02f01 g33283 ( .a(n37073), .b(n37072), .o(n37074) );
no02f01 g33284 ( .a(n37074), .b(n37071), .o(n37075) );
na02f01 g33285 ( .a(n37074), .b(n37071), .o(n37076) );
in01f01 g33286 ( .a(n37076), .o(n37077) );
no02f01 g33287 ( .a(n37077), .b(n37075), .o(n37078) );
in01f01 g33288 ( .a(n37078), .o(n37079) );
ao12f01 g33289 ( .a(n36972), .b(n37079), .c(n37070), .o(n37080) );
na02f01 g33290 ( .a(n7225), .b(n7205), .o(n37081) );
in01f01 g33291 ( .a(n7204), .o(n37082) );
ao12f01 g33292 ( .a(n7229), .b(n37082), .c(n7185), .o(n37083) );
ao12f01 g33293 ( .a(n7226), .b(n37083), .c(n37081), .o(n37084) );
no02f01 g33294 ( .a(n7215), .b(n7164), .o(n37085) );
no02f01 g33295 ( .a(n37085), .b(n7217), .o(n37086) );
in01f01 g33296 ( .a(n37086), .o(n37087) );
no02f01 g33297 ( .a(n37087), .b(n37084), .o(n37088) );
na02f01 g33298 ( .a(n37087), .b(n37084), .o(n37089) );
in01f01 g33299 ( .a(n37089), .o(n37090) );
no02f01 g33300 ( .a(n37090), .b(n37088), .o(n37091) );
in01f01 g33301 ( .a(n37091), .o(n37092) );
no02f01 g33302 ( .a(n37092), .b(n36972), .o(n37093) );
in01f01 g33303 ( .a(n7226), .o(n37094) );
na02f01 g33304 ( .a(n37081), .b(n37094), .o(n37095) );
in01f01 g33305 ( .a(n37095), .o(n37096) );
no02f01 g33306 ( .a(n37096), .b(n37083), .o(n37097) );
na02f01 g33307 ( .a(n37096), .b(n37083), .o(n37098) );
in01f01 g33308 ( .a(n37098), .o(n37099) );
no02f01 g33309 ( .a(n37099), .b(n37097), .o(n37100) );
in01f01 g33310 ( .a(n37100), .o(n37101) );
no02f01 g33311 ( .a(n37101), .b(n36972), .o(n37102) );
no03f01 g33312 ( .a(n37102), .b(n37093), .c(n37080), .o(n37103) );
in01f01 g33313 ( .a(n37103), .o(n37104) );
ao12f01 g33314 ( .a(n36963), .b(n37078), .c(n37069), .o(n37105) );
ao12f01 g33315 ( .a(n36963), .b(n37100), .c(n37091), .o(n37106) );
no02f01 g33316 ( .a(n37106), .b(n37105), .o(n37107) );
oa12f01 g33317 ( .a(n37107), .b(n37104), .c(n37062), .o(n37108) );
in01f01 g33318 ( .a(n36970), .o(n37109) );
no02f01 g33319 ( .a(n37109), .b(n36972), .o(n37110) );
in01f01 g33320 ( .a(n37110), .o(n37111) );
ao12f01 g33321 ( .a(n36971), .b(n37111), .c(n37108), .o(n37112) );
no02f01 g33322 ( .a(n36965), .b(n7232), .o(n37113) );
no02f01 g33323 ( .a(n7252), .b(n7205), .o(n37114) );
no02f01 g33324 ( .a(n7251), .b(n7164), .o(n37115) );
no02f01 g33325 ( .a(n37115), .b(n37114), .o(n37116) );
in01f01 g33326 ( .a(n37116), .o(n37117) );
no03f01 g33327 ( .a(n37117), .b(n37113), .c(n36964), .o(n37118) );
no02f01 g33328 ( .a(n37113), .b(n36964), .o(n37119) );
no02f01 g33329 ( .a(n37116), .b(n37119), .o(n37120) );
no02f01 g33330 ( .a(n37120), .b(n37118), .o(n37121) );
no02f01 g33331 ( .a(n37121), .b(n36963), .o(n37122) );
in01f01 g33332 ( .a(n37121), .o(n37123) );
no02f01 g33333 ( .a(n37123), .b(n36972), .o(n37124) );
no02f01 g33334 ( .a(n37124), .b(n37122), .o(n37125) );
na02f01 g33335 ( .a(n37125), .b(n37112), .o(n37126) );
in01f01 g33336 ( .a(n37112), .o(n37127) );
in01f01 g33337 ( .a(n37125), .o(n37128) );
na02f01 g33338 ( .a(n37128), .b(n37127), .o(n37129) );
na02f01 g33339 ( .a(n37129), .b(n37126), .o(n529) );
no02f01 g33340 ( .a(n25217), .b(n25023), .o(n37131) );
no02f01 g33341 ( .a(n25293), .b(n24613), .o(n37132) );
no02f01 g33342 ( .a(n37132), .b(n37131), .o(n37133) );
na02f01 g33343 ( .a(n25537), .b(n25286), .o(n37134) );
na03f01 g33344 ( .a(n37134), .b(n25201), .c(n25189), .o(n37135) );
na03f01 g33345 ( .a(n37135), .b(n37133), .c(n25297), .o(n37136) );
in01f01 g33346 ( .a(n37133), .o(n37137) );
in01f01 g33347 ( .a(n25322), .o(n37138) );
na03f01 g33348 ( .a(n25321), .b(n25309), .c(n25307), .o(n37139) );
na02f01 g33349 ( .a(n25531), .b(n37139), .o(n37140) );
oa12f01 g33350 ( .a(n37138), .b(n37140), .c(n25528), .o(n37141) );
in01f01 g33351 ( .a(n25535), .o(n37142) );
na02f01 g33352 ( .a(n25563), .b(n25231), .o(n37143) );
no04f01 g33353 ( .a(n37143), .b(n37142), .c(n37141), .d(n25261), .o(n37144) );
no02f01 g33354 ( .a(n37144), .b(n25569), .o(n37145) );
no03f01 g33355 ( .a(n37145), .b(n25561), .c(n25557), .o(n37146) );
oa12f01 g33356 ( .a(n37137), .b(n37146), .c(n25573), .o(n37147) );
na02f01 g33357 ( .a(n37147), .b(n37136), .o(n534) );
in01f01 g33358 ( .a(delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(n37149) );
no02f01 g33359 ( .a(n36972), .b(n36026), .o(n37150) );
no02f01 g33360 ( .a(n36963), .b(n36023), .o(n37151) );
no02f01 g33361 ( .a(n37151), .b(n37150), .o(n37152) );
in01f01 g33362 ( .a(n36990), .o(n37153) );
no02f01 g33363 ( .a(n36991), .b(n37153), .o(n37154) );
in01f01 g33364 ( .a(n36996), .o(n37155) );
na02f01 g33365 ( .a(n37155), .b(n37154), .o(n37156) );
in01f01 g33366 ( .a(n37009), .o(n37157) );
oa12f01 g33367 ( .a(n4973), .b(n4994), .c(n4895), .o(n37158) );
in01f01 g33368 ( .a(n37004), .o(n37159) );
oa12f01 g33369 ( .a(n37007), .b(n37159), .c(n37002), .o(n37160) );
ao12f01 g33370 ( .a(n37157), .b(n37160), .c(n37158), .o(n37161) );
no02f01 g33371 ( .a(n37155), .b(n37154), .o(n37162) );
oa12f01 g33372 ( .a(n37156), .b(n37162), .c(n37161), .o(n37163) );
in01f01 g33373 ( .a(n37016), .o(n37164) );
ao12f01 g33374 ( .a(n36986), .b(n37164), .c(n37163), .o(n37165) );
in01f01 g33375 ( .a(n37019), .o(n37166) );
no02f01 g33376 ( .a(n37018), .b(n36960), .o(n37167) );
no02f01 g33377 ( .a(n37167), .b(n37166), .o(n37168) );
in01f01 g33378 ( .a(n37030), .o(n37169) );
no02f01 g33379 ( .a(n37169), .b(n37168), .o(n37170) );
in01f01 g33380 ( .a(n37037), .o(n37171) );
no03f01 g33381 ( .a(n37171), .b(n37170), .c(n37165), .o(n37172) );
na02f01 g33382 ( .a(n37169), .b(n37168), .o(n37173) );
in01f01 g33383 ( .a(n37040), .o(n37174) );
ao12f01 g33384 ( .a(n37171), .b(n37174), .c(n37173), .o(n37175) );
no02f01 g33385 ( .a(n37175), .b(n37172), .o(n37176) );
in01f01 g33386 ( .a(n37059), .o(n37177) );
no03f01 g33387 ( .a(n37177), .b(n37175), .c(n37172), .o(n37178) );
in01f01 g33388 ( .a(n37061), .o(n37179) );
oa22f01 g33389 ( .a(n37179), .b(n37176), .c(n37178), .d(n36963), .o(n37180) );
in01f01 g33390 ( .a(n37107), .o(n37181) );
ao12f01 g33391 ( .a(n37181), .b(n37103), .c(n37180), .o(n37182) );
no02f01 g33392 ( .a(n37124), .b(n37110), .o(n37183) );
in01f01 g33393 ( .a(n37183), .o(n37184) );
no02f01 g33394 ( .a(n7253), .b(n7232), .o(n37185) );
no02f01 g33395 ( .a(n7271), .b(n7164), .o(n37186) );
no02f01 g33396 ( .a(n37186), .b(n7273), .o(n37187) );
in01f01 g33397 ( .a(n37187), .o(n37188) );
no03f01 g33398 ( .a(n37188), .b(n37185), .c(n7308), .o(n37189) );
no02f01 g33399 ( .a(n37185), .b(n7308), .o(n37190) );
no02f01 g33400 ( .a(n37187), .b(n37190), .o(n37191) );
no02f01 g33401 ( .a(n37191), .b(n37189), .o(n37192) );
in01f01 g33402 ( .a(n37192), .o(n37193) );
no02f01 g33403 ( .a(n37193), .b(n36972), .o(n37194) );
no03f01 g33404 ( .a(n7273), .b(n7253), .c(n7232), .o(n37195) );
no02f01 g33405 ( .a(n37186), .b(n7308), .o(n37196) );
in01f01 g33406 ( .a(n37196), .o(n37197) );
no02f01 g33407 ( .a(n7262), .b(n7164), .o(n37198) );
no02f01 g33408 ( .a(n37198), .b(n7264), .o(n37199) );
in01f01 g33409 ( .a(n37199), .o(n37200) );
no03f01 g33410 ( .a(n37200), .b(n37197), .c(n37195), .o(n37201) );
no02f01 g33411 ( .a(n37197), .b(n37195), .o(n37202) );
no02f01 g33412 ( .a(n37199), .b(n37202), .o(n37203) );
no02f01 g33413 ( .a(n37203), .b(n37201), .o(n37204) );
in01f01 g33414 ( .a(n37204), .o(n37205) );
no02f01 g33415 ( .a(n37205), .b(n36972), .o(n37206) );
no03f01 g33416 ( .a(n37206), .b(n37194), .c(n37184), .o(n37207) );
in01f01 g33417 ( .a(n37207), .o(n37208) );
no02f01 g33418 ( .a(n7294), .b(n7164), .o(n37209) );
no02f01 g33419 ( .a(n7275), .b(n7232), .o(n37210) );
no02f01 g33420 ( .a(n7311), .b(n37210), .o(n37211) );
no02f01 g33421 ( .a(n37211), .b(n7296), .o(n37212) );
no02f01 g33422 ( .a(n37212), .b(n37209), .o(n37213) );
no02f01 g33423 ( .a(n7285), .b(n7164), .o(n37214) );
no02f01 g33424 ( .a(n37214), .b(n7287), .o(n37215) );
no02f01 g33425 ( .a(n37215), .b(n37213), .o(n37216) );
na02f01 g33426 ( .a(n37215), .b(n37213), .o(n37217) );
in01f01 g33427 ( .a(n37217), .o(n37218) );
no02f01 g33428 ( .a(n37218), .b(n37216), .o(n37219) );
in01f01 g33429 ( .a(n37219), .o(n37220) );
no02f01 g33430 ( .a(n37220), .b(n36972), .o(n37221) );
no02f01 g33431 ( .a(n37209), .b(n7296), .o(n37222) );
no02f01 g33432 ( .a(n37222), .b(n37211), .o(n37223) );
na02f01 g33433 ( .a(n37222), .b(n37211), .o(n37224) );
in01f01 g33434 ( .a(n37224), .o(n37225) );
no02f01 g33435 ( .a(n37225), .b(n37223), .o(n37226) );
in01f01 g33436 ( .a(n37226), .o(n37227) );
no02f01 g33437 ( .a(n37227), .b(n36972), .o(n37228) );
no02f01 g33438 ( .a(n37228), .b(n37221), .o(n37229) );
in01f01 g33439 ( .a(n37229), .o(n37230) );
no02f01 g33440 ( .a(n36972), .b(n7444), .o(n37231) );
no02f01 g33441 ( .a(n7370), .b(n7369), .o(n37232) );
no02f01 g33442 ( .a(n7332), .b(n7300), .o(n37233) );
no02f01 g33443 ( .a(n37233), .b(n37232), .o(n37234) );
na02f01 g33444 ( .a(n37233), .b(n37232), .o(n37235) );
in01f01 g33445 ( .a(n37235), .o(n37236) );
no02f01 g33446 ( .a(n37236), .b(n37234), .o(n37237) );
in01f01 g33447 ( .a(n37237), .o(n37238) );
no02f01 g33448 ( .a(n37238), .b(n36972), .o(n37239) );
no02f01 g33449 ( .a(n37239), .b(n37231), .o(n37240) );
in01f01 g33450 ( .a(n37240), .o(n37241) );
no04f01 g33451 ( .a(n37241), .b(n37230), .c(n37208), .d(n37182), .o(n37242) );
no02f01 g33452 ( .a(n36972), .b(n7454), .o(n37243) );
no02f01 g33453 ( .a(n7448), .b(n7447), .o(n37244) );
in01f01 g33454 ( .a(n37244), .o(n37245) );
ao12f01 g33455 ( .a(n36972), .b(n37245), .c(n7445), .o(n37246) );
no02f01 g33456 ( .a(n36972), .b(n7397), .o(n37247) );
no03f01 g33457 ( .a(n37247), .b(n37246), .c(n37243), .o(n37248) );
na02f01 g33458 ( .a(n37248), .b(n37242), .o(n37249) );
ao12f01 g33459 ( .a(n36963), .b(n37121), .c(n36970), .o(n37250) );
ao12f01 g33460 ( .a(n36963), .b(n37204), .c(n37192), .o(n37251) );
no02f01 g33461 ( .a(n37251), .b(n37250), .o(n37252) );
in01f01 g33462 ( .a(n37252), .o(n37253) );
ao12f01 g33463 ( .a(n36963), .b(n37226), .c(n37219), .o(n37254) );
no02f01 g33464 ( .a(n37254), .b(n37253), .o(n37255) );
in01f01 g33465 ( .a(n37255), .o(n37256) );
ao12f01 g33466 ( .a(n36963), .b(n37237), .c(n7373), .o(n37257) );
no02f01 g33467 ( .a(n37257), .b(n37256), .o(n37258) );
in01f01 g33468 ( .a(n37258), .o(n37259) );
ao12f01 g33469 ( .a(n36963), .b(n37244), .c(n7383), .o(n37260) );
ao12f01 g33470 ( .a(n36963), .b(n7409), .c(n7326), .o(n37261) );
no02f01 g33471 ( .a(n37261), .b(n37260), .o(n37262) );
in01f01 g33472 ( .a(n37262), .o(n37263) );
no02f01 g33473 ( .a(n37263), .b(n37259), .o(n37264) );
na02f01 g33474 ( .a(n37264), .b(n37249), .o(n37265) );
in01f01 g33475 ( .a(n36010), .o(n37266) );
no02f01 g33476 ( .a(n36972), .b(n37266), .o(n37267) );
in01f01 g33477 ( .a(n7424), .o(n37268) );
no02f01 g33478 ( .a(n36972), .b(n37268), .o(n37269) );
no02f01 g33479 ( .a(n37269), .b(n37267), .o(n37270) );
na02f01 g33480 ( .a(n37270), .b(n37265), .o(n37271) );
ao12f01 g33481 ( .a(n36963), .b(n36010), .c(n7424), .o(n37272) );
in01f01 g33482 ( .a(n37272), .o(n37273) );
na03f01 g33483 ( .a(n37273), .b(n37271), .c(n37152), .o(n37274) );
in01f01 g33484 ( .a(n37152), .o(n37275) );
na02f01 g33485 ( .a(n37273), .b(n37271), .o(n37276) );
na02f01 g33486 ( .a(n37276), .b(n37275), .o(n37277) );
ao12f01 g33487 ( .a(n37149), .b(n37277), .c(n37274), .o(n37278) );
ao12f01 g33488 ( .a(delay_sub_ln23_0_unr23_stage8_stallmux_q), .b(n37277), .c(n37274), .o(n37279) );
no02f01 g33489 ( .a(n36963), .b(n7326), .o(n37280) );
no02f01 g33490 ( .a(n37280), .b(n37247), .o(n37281) );
in01f01 g33491 ( .a(n37281), .o(n37282) );
na04f01 g33492 ( .a(n37240), .b(n37229), .c(n37207), .d(n37108), .o(n37283) );
oa12f01 g33493 ( .a(n37258), .b(n37246), .c(n37283), .o(n37284) );
no03f01 g33494 ( .a(n37284), .b(n37282), .c(n37260), .o(n37285) );
in01f01 g33495 ( .a(n37260), .o(n37286) );
in01f01 g33496 ( .a(n37246), .o(n37287) );
ao12f01 g33497 ( .a(n37259), .b(n37287), .c(n37242), .o(n37288) );
ao12f01 g33498 ( .a(n37281), .b(n37288), .c(n37286), .o(n37289) );
oa12f01 g33499 ( .a(delay_sub_ln23_0_unr23_stage8_stallmux_q), .b(n37289), .c(n37285), .o(n37290) );
no02f01 g33500 ( .a(n36972), .b(n37245), .o(n37291) );
no02f01 g33501 ( .a(n36963), .b(n37244), .o(n37292) );
no02f01 g33502 ( .a(n37292), .b(n37291), .o(n37293) );
in01f01 g33503 ( .a(n37293), .o(n37294) );
no02f01 g33504 ( .a(n36972), .b(n7445), .o(n37295) );
no02f01 g33505 ( .a(n37295), .b(n37283), .o(n37296) );
no02f01 g33506 ( .a(n36963), .b(n7383), .o(n37297) );
no02f01 g33507 ( .a(n37297), .b(n37259), .o(n37298) );
in01f01 g33508 ( .a(n37298), .o(n37299) );
no03f01 g33509 ( .a(n37299), .b(n37296), .c(n37294), .o(n37300) );
in01f01 g33510 ( .a(n37295), .o(n37301) );
na02f01 g33511 ( .a(n37301), .b(n37242), .o(n37302) );
ao12f01 g33512 ( .a(n37293), .b(n37298), .c(n37302), .o(n37303) );
oa12f01 g33513 ( .a(delay_sub_ln23_0_unr23_stage8_stallmux_q), .b(n37303), .c(n37300), .o(n37304) );
no02f01 g33514 ( .a(n37295), .b(n37297), .o(n37305) );
no02f01 g33515 ( .a(n37259), .b(n37242), .o(n37306) );
na02f01 g33516 ( .a(n37306), .b(n37305), .o(n37307) );
in01f01 g33517 ( .a(n37305), .o(n37308) );
na02f01 g33518 ( .a(n37258), .b(n37283), .o(n37309) );
na02f01 g33519 ( .a(n37309), .b(n37308), .o(n37310) );
na02f01 g33520 ( .a(n37310), .b(n37307), .o(n5988) );
na02f01 g33521 ( .a(n5988), .b(delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(n37312) );
na03f01 g33522 ( .a(n37312), .b(n37304), .c(n37290), .o(n37313) );
in01f01 g33523 ( .a(n37247), .o(n37314) );
na02f01 g33524 ( .a(n37284), .b(n37314), .o(n37315) );
no02f01 g33525 ( .a(n37280), .b(n37260), .o(n37316) );
no02f01 g33526 ( .a(n36963), .b(n7409), .o(n37317) );
no02f01 g33527 ( .a(n37317), .b(n37243), .o(n37318) );
na03f01 g33528 ( .a(n37318), .b(n37316), .c(n37315), .o(n37319) );
no02f01 g33529 ( .a(n37288), .b(n37247), .o(n37320) );
in01f01 g33530 ( .a(n37316), .o(n37321) );
in01f01 g33531 ( .a(n37318), .o(n37322) );
oa12f01 g33532 ( .a(n37322), .b(n37321), .c(n37320), .o(n37323) );
ao12f01 g33533 ( .a(n37149), .b(n37323), .c(n37319), .o(n37324) );
in01f01 g33534 ( .a(n37248), .o(n37325) );
no02f01 g33535 ( .a(n37325), .b(n37283), .o(n37326) );
in01f01 g33536 ( .a(n37264), .o(n37327) );
no02f01 g33537 ( .a(n37327), .b(n37326), .o(n37328) );
no02f01 g33538 ( .a(n36963), .b(n7424), .o(n37329) );
no02f01 g33539 ( .a(n37329), .b(n37269), .o(n37330) );
na02f01 g33540 ( .a(n37330), .b(n37328), .o(n37331) );
in01f01 g33541 ( .a(n37330), .o(n37332) );
na02f01 g33542 ( .a(n37332), .b(n37265), .o(n37333) );
ao12f01 g33543 ( .a(n37149), .b(n37333), .c(n37331), .o(n37334) );
in01f01 g33544 ( .a(n37269), .o(n37335) );
in01f01 g33545 ( .a(n37329), .o(n37336) );
na03f01 g33546 ( .a(n37336), .b(n37264), .c(n37249), .o(n37337) );
no02f01 g33547 ( .a(n36963), .b(n36010), .o(n37338) );
no02f01 g33548 ( .a(n37338), .b(n37267), .o(n37339) );
in01f01 g33549 ( .a(n37339), .o(n37340) );
na03f01 g33550 ( .a(n37340), .b(n37337), .c(n37335), .o(n37341) );
no03f01 g33551 ( .a(n37329), .b(n37327), .c(n37326), .o(n37342) );
oa12f01 g33552 ( .a(n37339), .b(n37342), .c(n37269), .o(n37343) );
ao12f01 g33553 ( .a(n37149), .b(n37343), .c(n37341), .o(n37344) );
no04f01 g33554 ( .a(n37344), .b(n37334), .c(n37324), .d(n37313), .o(n37345) );
oa12f01 g33555 ( .a(n37345), .b(n37279), .c(n37278), .o(n37346) );
no02f01 g33556 ( .a(n37279), .b(n37278), .o(n37347) );
na03f01 g33557 ( .a(n37288), .b(n37281), .c(n37286), .o(n37348) );
oa12f01 g33558 ( .a(n37282), .b(n37284), .c(n37260), .o(n37349) );
ao12f01 g33559 ( .a(n37149), .b(n37349), .c(n37348), .o(n37350) );
na03f01 g33560 ( .a(n37298), .b(n37302), .c(n37293), .o(n37351) );
oa12f01 g33561 ( .a(n37294), .b(n37299), .c(n37296), .o(n37352) );
ao12f01 g33562 ( .a(n37149), .b(n37352), .c(n37351), .o(n37353) );
no02f01 g33563 ( .a(n37309), .b(n37308), .o(n37354) );
no02f01 g33564 ( .a(n37306), .b(n37305), .o(n37355) );
no02f01 g33565 ( .a(n37355), .b(n37354), .o(n37356) );
no02f01 g33566 ( .a(n37356), .b(n37149), .o(n37357) );
no03f01 g33567 ( .a(n37357), .b(n37353), .c(n37350), .o(n37358) );
no03f01 g33568 ( .a(n37322), .b(n37321), .c(n37320), .o(n37359) );
ao12f01 g33569 ( .a(n37318), .b(n37316), .c(n37315), .o(n37360) );
oa12f01 g33570 ( .a(delay_sub_ln23_0_unr23_stage8_stallmux_q), .b(n37360), .c(n37359), .o(n37361) );
in01f01 g33571 ( .a(n37334), .o(n37362) );
no03f01 g33572 ( .a(n37339), .b(n37342), .c(n37269), .o(n37363) );
ao12f01 g33573 ( .a(n37340), .b(n37337), .c(n37335), .o(n37364) );
oa12f01 g33574 ( .a(delay_sub_ln23_0_unr23_stage8_stallmux_q), .b(n37364), .c(n37363), .o(n37365) );
na04f01 g33575 ( .a(n37365), .b(n37362), .c(n37361), .d(n37358), .o(n37366) );
na02f01 g33576 ( .a(n37366), .b(n37347), .o(n37367) );
na02f01 g33577 ( .a(n37367), .b(n37346), .o(n539) );
no02f01 g33578 ( .a(n7011), .b(n6934), .o(n37369) );
no02f01 g33579 ( .a(n37369), .b(n7013), .o(n37370) );
in01f01 g33580 ( .a(n37370), .o(n37371) );
na02f01 g33581 ( .a(n37371), .b(n6990), .o(n37372) );
na02f01 g33582 ( .a(n37370), .b(n6989), .o(n37373) );
na02f01 g33583 ( .a(n37373), .b(n37372), .o(n544) );
in01f01 g33584 ( .a(n8421), .o(n37375) );
no02f01 g33585 ( .a(n37375), .b(cordic_combinational_sub_ln23_0_unr16_z_0_), .o(n37376) );
in01f01 g33586 ( .a(n8430), .o(n37377) );
oa22f01 g33587 ( .a(n37377), .b(n8429), .c(n37376), .d(n8420), .o(n37378) );
no02f01 g33588 ( .a(n37377), .b(n8429), .o(n37379) );
na02f01 g33589 ( .a(n37379), .b(n8422), .o(n37380) );
na02f01 g33590 ( .a(n37380), .b(n37378), .o(n549) );
in01f01 g33591 ( .a(n9233), .o(n37382) );
no03f01 g33592 ( .a(n9224), .b(n8899), .c(beta_31), .o(n37383) );
no02f01 g33593 ( .a(n9225), .b(n8899), .o(n37384) );
no02f01 g33594 ( .a(n9608), .b(n37384), .o(n37385) );
in01f01 g33595 ( .a(n37385), .o(n37386) );
no02f01 g33596 ( .a(n37386), .b(n37383), .o(n37387) );
ao12f01 g33597 ( .a(n9234), .b(n37387), .c(n37382), .o(n37388) );
no02f01 g33598 ( .a(n9594), .b(n8862), .o(n37389) );
no02f01 g33599 ( .a(n9595), .b(n8899), .o(n37390) );
no02f01 g33600 ( .a(n37390), .b(n37389), .o(n37391) );
in01f01 g33601 ( .a(n37391), .o(n3623) );
no02f01 g33602 ( .a(n3623), .b(n37388), .o(n37393) );
na02f01 g33603 ( .a(n3623), .b(n37388), .o(n37394) );
in01f01 g33604 ( .a(n37394), .o(n37395) );
no02f01 g33605 ( .a(n37395), .b(n37393), .o(n37396) );
in01f01 g33606 ( .a(n37396), .o(n554) );
no02f01 g33607 ( .a(n9595), .b(n4201), .o(n37398) );
no02f01 g33608 ( .a(n9594), .b(n9591), .o(n37399) );
no02f01 g33609 ( .a(n37399), .b(n37398), .o(n37400) );
in01f01 g33610 ( .a(n37400), .o(n559) );
no02f01 g33611 ( .a(n27136), .b(n26440), .o(n37402) );
in01f01 g33612 ( .a(n27133), .o(n37403) );
na02f01 g33613 ( .a(n27134), .b(n37403), .o(n37404) );
no02f01 g33614 ( .a(n37404), .b(n26441), .o(n37405) );
no02f01 g33615 ( .a(n37405), .b(n37402), .o(n37406) );
no02f01 g33616 ( .a(n27144), .b(n26440), .o(n37407) );
in01f01 g33617 ( .a(n37407), .o(n37408) );
na02f01 g33618 ( .a(n27124), .b(n27112), .o(n37409) );
na02f01 g33619 ( .a(n27140), .b(n26718), .o(n37410) );
in01f01 g33620 ( .a(n27143), .o(n37411) );
na02f01 g33621 ( .a(n37411), .b(n37410), .o(n37412) );
no02f01 g33622 ( .a(n37412), .b(n26441), .o(n37413) );
in01f01 g33623 ( .a(n37413), .o(n37414) );
na02f01 g33624 ( .a(n37414), .b(n37409), .o(n37415) );
na03f01 g33625 ( .a(n37415), .b(n37408), .c(n37406), .o(n37416) );
in01f01 g33626 ( .a(n37406), .o(n37417) );
no02f01 g33627 ( .a(n27248), .b(n27239), .o(n37418) );
oa12f01 g33628 ( .a(n37408), .b(n37413), .c(n37418), .o(n37419) );
na02f01 g33629 ( .a(n37419), .b(n37417), .o(n37420) );
na03f01 g33630 ( .a(n37420), .b(n37416), .c(n1821), .o(n37421) );
na02f01 g33631 ( .a(n37420), .b(n37416), .o(n2781) );
na02f01 g33632 ( .a(n2781), .b(n8066), .o(n37423) );
na02f01 g33633 ( .a(n37423), .b(n37421), .o(n564) );
in01f01 g33634 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_27_), .o(n37425) );
no02f01 g33635 ( .a(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .b(n37425), .o(n37426) );
in01f01 g33636 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_14_), .o(n37427) );
in01f01 g33637 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_5_), .o(n37428) );
in01f01 g33638 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_2_), .o(n37429) );
in01f01 g33639 ( .a(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .o(n37430) );
in01f01 g33640 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_0_), .o(n37431) );
no02f01 g33641 ( .a(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .b(n37431), .o(n37432) );
no02f01 g33642 ( .a(n37430), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_0_), .o(n37433) );
in01f01 g33643 ( .a(n37433), .o(n37434) );
ao12f01 g33644 ( .a(n37432), .b(n37434), .c(delay_sub_ln23_0_unr26_stage9_stallmux_q_1_), .o(n37435) );
no02f01 g33645 ( .a(n37430), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_1_), .o(n37436) );
no02f01 g33646 ( .a(n37436), .b(n37435), .o(n37437) );
no02f01 g33647 ( .a(n37437), .b(n37430), .o(n37438) );
no02f01 g33648 ( .a(n37438), .b(n37429), .o(n37439) );
na02f01 g33649 ( .a(n37430), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_1_), .o(n37440) );
in01f01 g33650 ( .a(n37440), .o(n37441) );
no02f01 g33651 ( .a(n37441), .b(n37437), .o(n37442) );
no02f01 g33652 ( .a(n37442), .b(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .o(n37443) );
no02f01 g33653 ( .a(n37443), .b(n37439), .o(n37444) );
na03f01 g33654 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_5_), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_3_), .c(delay_sub_ln23_0_unr28_stage9_stallmux_q_4_), .o(n37445) );
ao12f01 g33655 ( .a(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .b(n37444), .c(n37428), .o(n37447) );
ao12f01 g33656 ( .a(n37444), .b(n37445), .c(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .o(n37448) );
oa12f01 g33657 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_6_), .b(n37448), .c(n37430), .o(n37449) );
in01f01 g33658 ( .a(n37449), .o(n37450) );
in01f01 g33659 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_4_), .o(n37451) );
in01f01 g33660 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_3_), .o(n37452) );
ao12f01 g33661 ( .a(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .b(n37452), .c(n37451), .o(n37453) );
no03f01 g33662 ( .a(n37453), .b(n37450), .c(n37447), .o(n37454) );
in01f01 g33663 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_8_), .o(n37455) );
in01f01 g33664 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_7_), .o(n37456) );
no02f01 g33665 ( .a(n37456), .b(n37455), .o(n37457) );
ao12f01 g33666 ( .a(n37430), .b(n37457), .c(delay_sub_ln23_0_unr28_stage9_stallmux_q_9_), .o(n37458) );
no02f01 g33667 ( .a(n37458), .b(n37454), .o(n37459) );
in01f01 g33668 ( .a(n37459), .o(n37460) );
no02f01 g33669 ( .a(n37430), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_10_), .o(n37461) );
no02f01 g33670 ( .a(n37461), .b(n37460), .o(n37462) );
in01f01 g33671 ( .a(n37462), .o(n37463) );
ao12f01 g33672 ( .a(n37430), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_11_), .c(delay_sub_ln23_0_unr28_stage9_stallmux_q_12_), .o(n37464) );
no02f01 g33673 ( .a(n37464), .b(n37463), .o(n37465) );
in01f01 g33674 ( .a(n37465), .o(n37466) );
no02f01 g33675 ( .a(n37430), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_13_), .o(n37467) );
no02f01 g33676 ( .a(n37467), .b(n37466), .o(n37468) );
na02f01 g33677 ( .a(n37430), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_13_), .o(n37469) );
in01f01 g33678 ( .a(n37469), .o(n37470) );
no02f01 g33679 ( .a(n37470), .b(n37468), .o(n37471) );
ao12f01 g33680 ( .a(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .b(n37471), .c(n37427), .o(n37472) );
ao12f01 g33681 ( .a(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .b(n37456), .c(n37455), .o(n37473) );
in01f01 g33682 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_10_), .o(n37474) );
in01f01 g33683 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_9_), .o(n37475) );
ao12f01 g33684 ( .a(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .b(n37475), .c(n37474), .o(n37476) );
no02f01 g33685 ( .a(n37476), .b(n37473), .o(n37477) );
in01f01 g33686 ( .a(n37477), .o(n37478) );
in01f01 g33687 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_12_), .o(n37479) );
in01f01 g33688 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_11_), .o(n37480) );
ao12f01 g33689 ( .a(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .b(n37480), .c(n37479), .o(n37481) );
no02f01 g33690 ( .a(n37481), .b(n37478), .o(n37482) );
in01f01 g33691 ( .a(n37482), .o(n37483) );
ao12f01 g33692 ( .a(n37483), .b(n37468), .c(delay_sub_ln23_0_unr28_stage9_stallmux_q_14_), .o(n37484) );
in01f01 g33693 ( .a(n37484), .o(n37485) );
no02f01 g33694 ( .a(n37485), .b(n37472), .o(n37486) );
in01f01 g33695 ( .a(n37486), .o(n37487) );
ao12f01 g33696 ( .a(n37430), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_15_), .c(delay_sub_ln23_0_unr28_stage9_stallmux_q_16_), .o(n37488) );
no02f01 g33697 ( .a(n37430), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_18_), .o(n37489) );
no02f01 g33698 ( .a(n37430), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_17_), .o(n37490) );
no03f01 g33699 ( .a(n37490), .b(n37489), .c(n37488), .o(n37491) );
na02f01 g33700 ( .a(n37491), .b(n37487), .o(n37492) );
ao12f01 g33701 ( .a(n37430), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_19_), .c(delay_sub_ln23_0_unr28_stage9_stallmux_q_20_), .o(n37493) );
no02f01 g33702 ( .a(n37493), .b(n37492), .o(n37494) );
in01f01 g33703 ( .a(n37494), .o(n37495) );
no02f01 g33704 ( .a(n37430), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_21_), .o(n37496) );
no02f01 g33705 ( .a(n37496), .b(n37495), .o(n37497) );
in01f01 g33706 ( .a(n37497), .o(n37498) );
no02f01 g33707 ( .a(n37430), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_22_), .o(n37499) );
no02f01 g33708 ( .a(n37499), .b(n37498), .o(n37500) );
in01f01 g33709 ( .a(n37500), .o(n37501) );
ao12f01 g33710 ( .a(n37430), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_24_), .c(delay_sub_ln23_0_unr28_stage9_stallmux_q_23_), .o(n37502) );
no02f01 g33711 ( .a(n37502), .b(n37501), .o(n37503) );
in01f01 g33712 ( .a(n37503), .o(n37504) );
no02f01 g33713 ( .a(n37430), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_25_), .o(n37505) );
no02f01 g33714 ( .a(n37505), .b(n37504), .o(n37506) );
in01f01 g33715 ( .a(n37506), .o(n37507) );
no02f01 g33716 ( .a(n37430), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_26_), .o(n37508) );
no02f01 g33717 ( .a(n37430), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_27_), .o(n37509) );
no03f01 g33718 ( .a(n37509), .b(n37508), .c(n37507), .o(n37510) );
no02f01 g33719 ( .a(n37510), .b(n37426), .o(n37511) );
in01f01 g33720 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_16_), .o(n37512) );
in01f01 g33721 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_15_), .o(n37513) );
ao12f01 g33722 ( .a(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .b(n37513), .c(n37512), .o(n37514) );
in01f01 g33723 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_17_), .o(n37515) );
in01f01 g33724 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_18_), .o(n37516) );
ao12f01 g33725 ( .a(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .b(n37516), .c(n37515), .o(n37517) );
no02f01 g33726 ( .a(n37517), .b(n37514), .o(n37518) );
in01f01 g33727 ( .a(n37518), .o(n37519) );
in01f01 g33728 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_20_), .o(n37520) );
in01f01 g33729 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_19_), .o(n37521) );
ao12f01 g33730 ( .a(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .b(n37521), .c(n37520), .o(n37522) );
no02f01 g33731 ( .a(n37522), .b(n37519), .o(n37523) );
in01f01 g33732 ( .a(n37523), .o(n37524) );
in01f01 g33733 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_22_), .o(n37525) );
in01f01 g33734 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_21_), .o(n37526) );
ao12f01 g33735 ( .a(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .b(n37526), .c(n37525), .o(n37527) );
no02f01 g33736 ( .a(n37527), .b(n37524), .o(n37528) );
in01f01 g33737 ( .a(n37528), .o(n37529) );
in01f01 g33738 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_23_), .o(n37530) );
in01f01 g33739 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_24_), .o(n37531) );
ao12f01 g33740 ( .a(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .b(n37531), .c(n37530), .o(n37532) );
no02f01 g33741 ( .a(n37532), .b(n37529), .o(n37533) );
in01f01 g33742 ( .a(n37533), .o(n37534) );
in01f01 g33743 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_26_), .o(n37535) );
in01f01 g33744 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_25_), .o(n37536) );
ao12f01 g33745 ( .a(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .b(n37536), .c(n37535), .o(n37537) );
no02f01 g33746 ( .a(n37537), .b(n37534), .o(n37538) );
no02f01 g33747 ( .a(n37430), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_28_), .o(n37539) );
in01f01 g33748 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_28_), .o(n37540) );
no02f01 g33749 ( .a(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .b(n37540), .o(n37541) );
no02f01 g33750 ( .a(n37541), .b(n37539), .o(n37542) );
ao12f01 g33751 ( .a(n37542), .b(n37538), .c(n37511), .o(n37543) );
in01f01 g33752 ( .a(n37538), .o(n37544) );
in01f01 g33753 ( .a(n37542), .o(n37545) );
no04f01 g33754 ( .a(n37545), .b(n37544), .c(n37510), .d(n37426), .o(n37546) );
no02f01 g33755 ( .a(n37546), .b(n37543), .o(n37547) );
no02f01 g33756 ( .a(n37508), .b(n37507), .o(n37548) );
in01f01 g33757 ( .a(n37548), .o(n37549) );
no02f01 g33758 ( .a(n37509), .b(n37426), .o(n37550) );
na03f01 g33759 ( .a(n37550), .b(n37538), .c(n37549), .o(n37551) );
in01f01 g33760 ( .a(n37550), .o(n37552) );
oa12f01 g33761 ( .a(n37552), .b(n37544), .c(n37548), .o(n37553) );
na02f01 g33762 ( .a(n37553), .b(n37551), .o(n37554) );
no02f01 g33763 ( .a(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .b(n37536), .o(n37555) );
no03f01 g33764 ( .a(n37555), .b(n37534), .c(n37506), .o(n37556) );
no02f01 g33765 ( .a(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .b(n37535), .o(n37557) );
no02f01 g33766 ( .a(n37557), .b(n37508), .o(n37558) );
na02f01 g33767 ( .a(n37558), .b(n37556), .o(n37559) );
in01f01 g33768 ( .a(n37556), .o(n37560) );
in01f01 g33769 ( .a(n37558), .o(n37561) );
na02f01 g33770 ( .a(n37561), .b(n37560), .o(n37562) );
na02f01 g33771 ( .a(n37562), .b(n37559), .o(n37563) );
no02f01 g33772 ( .a(n37555), .b(n37505), .o(n37564) );
na03f01 g33773 ( .a(n37564), .b(n37533), .c(n37504), .o(n37565) );
in01f01 g33774 ( .a(n37564), .o(n37566) );
oa12f01 g33775 ( .a(n37566), .b(n37534), .c(n37503), .o(n37567) );
na02f01 g33776 ( .a(n37567), .b(n37565), .o(n37568) );
no02f01 g33777 ( .a(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .b(n37526), .o(n37569) );
no02f01 g33778 ( .a(n37569), .b(n37496), .o(n37570) );
na03f01 g33779 ( .a(n37570), .b(n37518), .c(n37495), .o(n37571) );
in01f01 g33780 ( .a(n37570), .o(n37572) );
oa12f01 g33781 ( .a(n37572), .b(n37519), .c(n37494), .o(n37573) );
na02f01 g33782 ( .a(n37573), .b(n37571), .o(n37574) );
in01f01 g33783 ( .a(n37490), .o(n37575) );
no02f01 g33784 ( .a(n37488), .b(n37486), .o(n37576) );
in01f01 g33785 ( .a(n37514), .o(n37577) );
no02f01 g33786 ( .a(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .b(n37515), .o(n37578) );
in01f01 g33787 ( .a(n37578), .o(n37579) );
na02f01 g33788 ( .a(n37579), .b(n37577), .o(n37580) );
ao12f01 g33789 ( .a(n37580), .b(n37576), .c(n37575), .o(n37581) );
in01f01 g33790 ( .a(n37581), .o(n37582) );
no02f01 g33791 ( .a(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .b(n37516), .o(n37583) );
no02f01 g33792 ( .a(n37583), .b(n37489), .o(n37584) );
in01f01 g33793 ( .a(n37584), .o(n37585) );
na02f01 g33794 ( .a(n37585), .b(n37582), .o(n37586) );
na02f01 g33795 ( .a(n37584), .b(n37581), .o(n37587) );
na02f01 g33796 ( .a(n37587), .b(n37586), .o(n37588) );
no02f01 g33797 ( .a(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .b(n37513), .o(n37589) );
no02f01 g33798 ( .a(n37430), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_15_), .o(n37590) );
no02f01 g33799 ( .a(n37590), .b(n37486), .o(n37591) );
no02f01 g33800 ( .a(n37591), .b(n37589), .o(n37592) );
no02f01 g33801 ( .a(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .b(n37512), .o(n37593) );
no02f01 g33802 ( .a(n37430), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_16_), .o(n37594) );
no02f01 g33803 ( .a(n37594), .b(n37593), .o(n37595) );
no02f01 g33804 ( .a(n37595), .b(n37592), .o(n37596) );
na02f01 g33805 ( .a(n37595), .b(n37592), .o(n37597) );
in01f01 g33806 ( .a(n37597), .o(n37598) );
no02f01 g33807 ( .a(n37598), .b(n37596), .o(n37599) );
no02f01 g33808 ( .a(n37590), .b(n37589), .o(n37600) );
in01f01 g33809 ( .a(n37600), .o(n37601) );
no02f01 g33810 ( .a(n37601), .b(n37487), .o(n37602) );
no02f01 g33811 ( .a(n37600), .b(n37486), .o(n37603) );
no02f01 g33812 ( .a(n37603), .b(n37602), .o(n37604) );
na02f01 g33813 ( .a(n37482), .b(n37471), .o(n37605) );
in01f01 g33814 ( .a(n37605), .o(n37606) );
no02f01 g33815 ( .a(n37430), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_14_), .o(n37607) );
no02f01 g33816 ( .a(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .b(n37427), .o(n37608) );
no02f01 g33817 ( .a(n37608), .b(n37607), .o(n37609) );
no02f01 g33818 ( .a(n37609), .b(n37606), .o(n37610) );
na02f01 g33819 ( .a(n37609), .b(n37606), .o(n37611) );
in01f01 g33820 ( .a(n37611), .o(n37612) );
no02f01 g33821 ( .a(n37612), .b(n37610), .o(n37613) );
na03f01 g33822 ( .a(n37613), .b(n37604), .c(n37599), .o(n37614) );
no03f01 g33823 ( .a(n37569), .b(n37524), .c(n37497), .o(n37615) );
in01f01 g33824 ( .a(n37615), .o(n37616) );
no02f01 g33825 ( .a(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .b(n37525), .o(n37617) );
no02f01 g33826 ( .a(n37617), .b(n37499), .o(n37618) );
in01f01 g33827 ( .a(n37618), .o(n37619) );
no02f01 g33828 ( .a(n37619), .b(n37616), .o(n37620) );
no02f01 g33829 ( .a(n37618), .b(n37615), .o(n37621) );
no02f01 g33830 ( .a(n37621), .b(n37620), .o(n37622) );
no02f01 g33831 ( .a(n37578), .b(n37490), .o(n37623) );
in01f01 g33832 ( .a(n37623), .o(n37624) );
no03f01 g33833 ( .a(n37624), .b(n37576), .c(n37514), .o(n37625) );
no02f01 g33834 ( .a(n37576), .b(n37514), .o(n37626) );
no02f01 g33835 ( .a(n37623), .b(n37626), .o(n37627) );
no02f01 g33836 ( .a(n37627), .b(n37625), .o(n37628) );
na02f01 g33837 ( .a(n37518), .b(n37492), .o(n37629) );
no02f01 g33838 ( .a(n37430), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_20_), .o(n37630) );
no02f01 g33839 ( .a(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .b(n37520), .o(n37631) );
no02f01 g33840 ( .a(n37631), .b(n37630), .o(n37632) );
in01f01 g33841 ( .a(n37632), .o(n37633) );
no02f01 g33842 ( .a(n37633), .b(n37629), .o(n37634) );
in01f01 g33843 ( .a(n37629), .o(n37635) );
no02f01 g33844 ( .a(n37632), .b(n37635), .o(n37636) );
no02f01 g33845 ( .a(n37636), .b(n37634), .o(n37637) );
no02f01 g33846 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_19_), .b(n37430), .o(n37638) );
no02f01 g33847 ( .a(n37521), .b(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .o(n37639) );
no02f01 g33848 ( .a(n37639), .b(n37638), .o(n37640) );
no02f01 g33849 ( .a(n37640), .b(n37635), .o(n37641) );
in01f01 g33850 ( .a(n37640), .o(n37642) );
no02f01 g33851 ( .a(n37642), .b(n37629), .o(n37643) );
no02f01 g33852 ( .a(n37643), .b(n37641), .o(n37644) );
na04f01 g33853 ( .a(n37644), .b(n37637), .c(n37628), .d(n37622), .o(n37645) );
no04f01 g33854 ( .a(n37645), .b(n37614), .c(n37588), .d(n37574), .o(n37646) );
no02f01 g33855 ( .a(n37529), .b(n37500), .o(n37647) );
no02f01 g33856 ( .a(n37430), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_23_), .o(n37648) );
no02f01 g33857 ( .a(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .b(n37530), .o(n37649) );
no02f01 g33858 ( .a(n37649), .b(n37648), .o(n37650) );
no02f01 g33859 ( .a(n37650), .b(n37647), .o(n37651) );
in01f01 g33860 ( .a(n37647), .o(n37652) );
in01f01 g33861 ( .a(n37650), .o(n37653) );
no02f01 g33862 ( .a(n37653), .b(n37652), .o(n37654) );
no02f01 g33863 ( .a(n37654), .b(n37651), .o(n37655) );
no02f01 g33864 ( .a(n37430), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_24_), .o(n37656) );
no02f01 g33865 ( .a(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .b(n37531), .o(n37657) );
no02f01 g33866 ( .a(n37657), .b(n37656), .o(n37658) );
no02f01 g33867 ( .a(n37658), .b(n37647), .o(n37659) );
in01f01 g33868 ( .a(n37658), .o(n37660) );
no02f01 g33869 ( .a(n37660), .b(n37652), .o(n37661) );
no02f01 g33870 ( .a(n37661), .b(n37659), .o(n37662) );
na03f01 g33871 ( .a(n37662), .b(n37655), .c(n37646), .o(n37663) );
no04f01 g33872 ( .a(n37663), .b(n37568), .c(n37563), .d(n37554), .o(n37664) );
ao12f01 g33873 ( .a(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .b(n37511), .c(n37540), .o(n37665) );
ao12f01 g33874 ( .a(n37544), .b(n37510), .c(delay_sub_ln23_0_unr28_stage9_stallmux_q_28_), .o(n37666) );
in01f01 g33875 ( .a(n37666), .o(n37667) );
no02f01 g33876 ( .a(n37667), .b(n37665), .o(n2377) );
ao12f01 g33877 ( .a(n2377), .b(n37664), .c(n37547), .o(n37669) );
in01f01 g33878 ( .a(delay_sub_ln23_0_unr26_stage9_stallmux_q_1_), .o(n37670) );
in01f01 g33879 ( .a(n2377), .o(n37671) );
in01f01 g33880 ( .a(n37435), .o(n37672) );
no02f01 g33881 ( .a(n37441), .b(n37436), .o(n37673) );
in01f01 g33882 ( .a(n37673), .o(n37674) );
no02f01 g33883 ( .a(n37674), .b(n37672), .o(n37675) );
no02f01 g33884 ( .a(n37673), .b(n37435), .o(n37676) );
no02f01 g33885 ( .a(n37676), .b(n37675), .o(n37677) );
no02f01 g33886 ( .a(n37433), .b(n37432), .o(n37678) );
na03f01 g33887 ( .a(n37678), .b(delay_sub_ln23_0_unr26_stage9_stallmux_q_0_), .c(n37670), .o(n37679) );
no02f01 g33888 ( .a(n37679), .b(n37677), .o(n37680) );
oa22f01 g33889 ( .a(n37680), .b(n37671), .c(delay_sub_ln23_0_unr26_stage9_stallmux_q_0_), .d(n37670), .o(n37681) );
in01f01 g33890 ( .a(n37681), .o(n37682) );
in01f01 g33891 ( .a(n37444), .o(n37683) );
no02f01 g33892 ( .a(n37430), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_4_), .o(n37684) );
no02f01 g33893 ( .a(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .b(n37451), .o(n37685) );
no02f01 g33894 ( .a(n37685), .b(n37684), .o(n37686) );
in01f01 g33895 ( .a(n37686), .o(n37687) );
no02f01 g33896 ( .a(n37687), .b(n37683), .o(n37688) );
no02f01 g33897 ( .a(n37686), .b(n37444), .o(n37689) );
no02f01 g33898 ( .a(n37689), .b(n37688), .o(n37690) );
no02f01 g33899 ( .a(n37430), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_2_), .o(n37691) );
no02f01 g33900 ( .a(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .b(n37429), .o(n37692) );
no02f01 g33901 ( .a(n37692), .b(n37691), .o(n37693) );
in01f01 g33902 ( .a(n37693), .o(n37694) );
no03f01 g33903 ( .a(n37694), .b(n37441), .c(n37437), .o(n37695) );
no02f01 g33904 ( .a(n37693), .b(n37442), .o(n37696) );
no02f01 g33905 ( .a(n37696), .b(n37695), .o(n37697) );
no02f01 g33906 ( .a(n37697), .b(n37690), .o(n37698) );
no02f01 g33907 ( .a(n37428), .b(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .o(n37699) );
no02f01 g33908 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_5_), .b(n37430), .o(n37700) );
no02f01 g33909 ( .a(n37700), .b(n37699), .o(n37701) );
na02f01 g33910 ( .a(n37701), .b(n37444), .o(n37702) );
in01f01 g33911 ( .a(n37701), .o(n37703) );
na02f01 g33912 ( .a(n37703), .b(n37683), .o(n37704) );
na02f01 g33913 ( .a(n37704), .b(n37702), .o(n37705) );
no02f01 g33914 ( .a(n37430), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_3_), .o(n37706) );
no02f01 g33915 ( .a(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .b(n37452), .o(n37707) );
no02f01 g33916 ( .a(n37707), .b(n37706), .o(n37708) );
na02f01 g33917 ( .a(n37708), .b(n37444), .o(n37709) );
in01f01 g33918 ( .a(n37708), .o(n37710) );
na02f01 g33919 ( .a(n37710), .b(n37683), .o(n37711) );
na02f01 g33920 ( .a(n37711), .b(n37709), .o(n37712) );
na04f01 g33921 ( .a(n37712), .b(n37705), .c(n37698), .d(n37682), .o(n37713) );
in01f01 g33922 ( .a(n37678), .o(n37714) );
no02f01 g33923 ( .a(n37714), .b(delay_sub_ln23_0_unr26_stage9_stallmux_q_1_), .o(n37715) );
no02f01 g33924 ( .a(n37678), .b(n37670), .o(n37716) );
no02f01 g33925 ( .a(n37716), .b(n37715), .o(n37717) );
na04f01 g33926 ( .a(n37697), .b(n37690), .c(n37717), .d(n37677), .o(n37718) );
no04f01 g33927 ( .a(n37718), .b(n37712), .c(n37705), .d(n37682), .o(n37719) );
oa12f01 g33928 ( .a(n37713), .b(n37719), .c(n2377), .o(n37720) );
no02f01 g33929 ( .a(n37470), .b(n37467), .o(n37721) );
in01f01 g33930 ( .a(n37721), .o(n37722) );
no03f01 g33931 ( .a(n37722), .b(n37483), .c(n37465), .o(n37723) );
ao12f01 g33932 ( .a(n37721), .b(n37482), .c(n37466), .o(n37724) );
no02f01 g33933 ( .a(n37724), .b(n37723), .o(n37725) );
no02f01 g33934 ( .a(n37478), .b(n37462), .o(n37726) );
no02f01 g33935 ( .a(n37430), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_11_), .o(n37727) );
no02f01 g33936 ( .a(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .b(n37480), .o(n37728) );
no02f01 g33937 ( .a(n37728), .b(n37727), .o(n37729) );
no02f01 g33938 ( .a(n37729), .b(n37726), .o(n37730) );
in01f01 g33939 ( .a(n37726), .o(n37731) );
in01f01 g33940 ( .a(n37729), .o(n37732) );
no02f01 g33941 ( .a(n37732), .b(n37731), .o(n37733) );
no02f01 g33942 ( .a(n37733), .b(n37730), .o(n37734) );
no02f01 g33943 ( .a(n37430), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_12_), .o(n37735) );
no02f01 g33944 ( .a(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .b(n37479), .o(n37736) );
no02f01 g33945 ( .a(n37736), .b(n37735), .o(n37737) );
in01f01 g33946 ( .a(n37737), .o(n37738) );
no02f01 g33947 ( .a(n37738), .b(n37731), .o(n37739) );
no02f01 g33948 ( .a(n37737), .b(n37726), .o(n37740) );
no02f01 g33949 ( .a(n37740), .b(n37739), .o(n37741) );
no02f01 g33950 ( .a(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .b(n37475), .o(n37742) );
no03f01 g33951 ( .a(n37742), .b(n37473), .c(n37459), .o(n37743) );
no02f01 g33952 ( .a(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .b(n37474), .o(n37744) );
no02f01 g33953 ( .a(n37744), .b(n37461), .o(n37745) );
na02f01 g33954 ( .a(n37745), .b(n37743), .o(n37746) );
in01f01 g33955 ( .a(n37743), .o(n37747) );
in01f01 g33956 ( .a(n37745), .o(n37748) );
na02f01 g33957 ( .a(n37748), .b(n37747), .o(n37749) );
na02f01 g33958 ( .a(n37749), .b(n37746), .o(n37750) );
no03f01 g33959 ( .a(n37453), .b(n37699), .c(n37448), .o(n37751) );
no02f01 g33960 ( .a(n37430), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_6_), .o(n37752) );
na02f01 g33961 ( .a(n37430), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_6_), .o(n37753) );
in01f01 g33962 ( .a(n37753), .o(n37754) );
no02f01 g33963 ( .a(n37754), .b(n37752), .o(n37755) );
no02f01 g33964 ( .a(n37755), .b(n37751), .o(n37756) );
na02f01 g33965 ( .a(n37755), .b(n37751), .o(n37757) );
in01f01 g33966 ( .a(n37757), .o(n37758) );
no02f01 g33967 ( .a(n37758), .b(n37756), .o(n37759) );
no02f01 g33968 ( .a(n37430), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_9_), .o(n37760) );
no02f01 g33969 ( .a(n37742), .b(n37760), .o(n37761) );
no02f01 g33970 ( .a(n37761), .b(n37454), .o(n37762) );
na02f01 g33971 ( .a(n37761), .b(n37454), .o(n37763) );
in01f01 g33972 ( .a(n37763), .o(n37764) );
no02f01 g33973 ( .a(n37764), .b(n37762), .o(n37765) );
no02f01 g33974 ( .a(n37430), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_8_), .o(n37766) );
no02f01 g33975 ( .a(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .b(n37455), .o(n37767) );
no02f01 g33976 ( .a(n37767), .b(n37766), .o(n37768) );
no02f01 g33977 ( .a(n37768), .b(n37454), .o(n37769) );
in01f01 g33978 ( .a(n37454), .o(n37770) );
in01f01 g33979 ( .a(n37768), .o(n37771) );
no02f01 g33980 ( .a(n37771), .b(n37770), .o(n37772) );
no02f01 g33981 ( .a(n37772), .b(n37769), .o(n37773) );
no02f01 g33982 ( .a(n37430), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_7_), .o(n37774) );
no02f01 g33983 ( .a(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .b(n37456), .o(n37775) );
no02f01 g33984 ( .a(n37775), .b(n37774), .o(n37776) );
no02f01 g33985 ( .a(n37776), .b(n37454), .o(n37777) );
in01f01 g33986 ( .a(n37776), .o(n37778) );
no02f01 g33987 ( .a(n37778), .b(n37770), .o(n37779) );
no02f01 g33988 ( .a(n37779), .b(n37777), .o(n37780) );
no04f01 g33989 ( .a(n37780), .b(n37773), .c(n37765), .d(n37759), .o(n37781) );
na02f01 g33990 ( .a(n37781), .b(n37750), .o(n37782) );
no04f01 g33991 ( .a(n37782), .b(n37741), .c(n37734), .d(n37725), .o(n37783) );
na02f01 g33992 ( .a(n37783), .b(n37720), .o(n37784) );
na04f01 g33993 ( .a(n37780), .b(n37773), .c(n37765), .d(n37759), .o(n37785) );
no02f01 g33994 ( .a(n37785), .b(n37750), .o(n37786) );
na04f01 g33995 ( .a(n37786), .b(n37741), .c(n37734), .d(n37725), .o(n37787) );
oa12f01 g33996 ( .a(n37671), .b(n37787), .c(n37720), .o(n37788) );
no03f01 g33997 ( .a(n37644), .b(n37637), .c(n37628), .o(n37789) );
no03f01 g33998 ( .a(n37613), .b(n37604), .c(n37599), .o(n37790) );
na04f01 g33999 ( .a(n37790), .b(n37789), .c(n37588), .d(n37574), .o(n37791) );
ao22f01 g34000 ( .a(n37791), .b(n2377), .c(n37788), .d(n37784), .o(n37792) );
no03f01 g34001 ( .a(n37662), .b(n37655), .c(n37622), .o(n37793) );
na04f01 g34002 ( .a(n37793), .b(n37568), .c(n37563), .d(n37554), .o(n37794) );
oa12f01 g34003 ( .a(n2377), .b(n37794), .c(n37547), .o(n37795) );
oa12f01 g34004 ( .a(n37795), .b(n37792), .c(n37669), .o(n569) );
in01f01 g34005 ( .a(n8518), .o(n37797) );
in01f01 g34006 ( .a(n8484), .o(n37798) );
in01f01 g34007 ( .a(n8485), .o(n37799) );
no02f01 g34008 ( .a(n37799), .b(n37798), .o(n37800) );
in01f01 g34009 ( .a(n37800), .o(n37801) );
no02f01 g34010 ( .a(n8508), .b(n37801), .o(n37802) );
ao12f01 g34011 ( .a(n8471), .b(n8533), .c(n8516), .o(n37803) );
ao12f01 g34012 ( .a(n37803), .b(n37802), .c(n37797), .o(n37804) );
in01f01 g34013 ( .a(n37804), .o(n37805) );
no02f01 g34014 ( .a(n8528), .b(n8471), .o(n37806) );
no02f01 g34015 ( .a(n37806), .b(n8530), .o(n37807) );
in01f01 g34016 ( .a(n37807), .o(n37808) );
na02f01 g34017 ( .a(n37808), .b(n37805), .o(n37809) );
na02f01 g34018 ( .a(n37807), .b(n37804), .o(n37810) );
na02f01 g34019 ( .a(n37810), .b(n37809), .o(n574) );
ao12f01 g34020 ( .a(n32538), .b(n26754), .c(n7682), .o(n37812) );
na02f01 g34021 ( .a(n37412), .b(n7682), .o(n37813) );
oa12f01 g34022 ( .a(n7682), .b(n27135), .c(n27133), .o(n37814) );
na03f01 g34023 ( .a(n37814), .b(n37813), .c(n37812), .o(n37815) );
oa12f01 g34024 ( .a(n7712), .b(n26844), .c(n26754), .o(n37816) );
na02f01 g34025 ( .a(n37412), .b(n7712), .o(n37817) );
na02f01 g34026 ( .a(n37817), .b(n37816), .o(n37818) );
ao12f01 g34027 ( .a(n37818), .b(n37404), .c(n7712), .o(n37819) );
na02f01 g34028 ( .a(n37819), .b(n37815), .o(n37820) );
in01f01 g34029 ( .a(n27158), .o(n37821) );
ao12f01 g34030 ( .a(n7712), .b(n27159), .c(n37821), .o(n37822) );
no02f01 g34031 ( .a(n27169), .b(n7712), .o(n37823) );
no02f01 g34032 ( .a(n37823), .b(n37822), .o(n37824) );
na02f01 g34033 ( .a(n37824), .b(n37820), .o(n37825) );
no02f01 g34034 ( .a(n27189), .b(n7712), .o(n37826) );
oa12f01 g34035 ( .a(n7712), .b(n27160), .c(n27158), .o(n37827) );
na02f01 g34036 ( .a(n27153), .b(n7712), .o(n37828) );
na02f01 g34037 ( .a(n37828), .b(n37827), .o(n37829) );
oa12f01 g34038 ( .a(n7712), .b(n27188), .c(n27186), .o(n37830) );
in01f01 g34039 ( .a(n37830), .o(n37831) );
in01f01 g34040 ( .a(n27180), .o(n37832) );
ao12f01 g34041 ( .a(n7682), .b(n27181), .c(n37832), .o(n37833) );
no03f01 g34042 ( .a(n37833), .b(n37831), .c(n37829), .o(n37834) );
oa12f01 g34043 ( .a(n37834), .b(n37826), .c(n37825), .o(n37835) );
no02f01 g34044 ( .a(n27183), .b(n7712), .o(n37836) );
in01f01 g34045 ( .a(n37836), .o(n37837) );
no02f01 g34046 ( .a(n26738), .b(n7712), .o(n37838) );
in01f01 g34047 ( .a(n37838), .o(n37839) );
no02f01 g34048 ( .a(n26504), .b(n25954), .o(n37840) );
in01f01 g34049 ( .a(n25954), .o(n37841) );
no02f01 g34050 ( .a(n26502), .b(n37841), .o(n37842) );
no02f01 g34051 ( .a(n37842), .b(n37840), .o(n37843) );
in01f01 g34052 ( .a(n37843), .o(n37844) );
in01f01 g34053 ( .a(n26503), .o(n37845) );
in01f01 g34054 ( .a(n26732), .o(n37846) );
na03f01 g34055 ( .a(n37846), .b(n27173), .c(n37845), .o(n37847) );
in01f01 g34056 ( .a(n26729), .o(n37848) );
no02f01 g34057 ( .a(n26508), .b(n26442), .o(n37849) );
no02f01 g34058 ( .a(n37849), .b(n26504), .o(n37850) );
no02f01 g34059 ( .a(n37850), .b(n37848), .o(n37851) );
oa12f01 g34060 ( .a(n37851), .b(n37847), .c(n26726), .o(n37852) );
na02f01 g34061 ( .a(n37852), .b(n37844), .o(n37853) );
in01f01 g34062 ( .a(n37853), .o(n37854) );
no02f01 g34063 ( .a(n37852), .b(n37844), .o(n37855) );
no02f01 g34064 ( .a(n37855), .b(n37854), .o(n37856) );
in01f01 g34065 ( .a(n37856), .o(n37857) );
na02f01 g34066 ( .a(n37857), .b(n7682), .o(n37858) );
na04f01 g34067 ( .a(n37858), .b(n37839), .c(n37837), .d(n37835), .o(n37859) );
no02f01 g34068 ( .a(n26738), .b(n7682), .o(n37860) );
no02f01 g34069 ( .a(n37856), .b(n7682), .o(n37861) );
no02f01 g34070 ( .a(n37861), .b(n37860), .o(n37862) );
in01f01 g34071 ( .a(n37858), .o(n37863) );
no02f01 g34072 ( .a(n37861), .b(n37863), .o(n37864) );
na03f01 g34073 ( .a(n37864), .b(n37862), .c(n37859), .o(n37865) );
na02f01 g34074 ( .a(n37837), .b(n37835), .o(n37866) );
na02f01 g34075 ( .a(n37858), .b(n37839), .o(n37867) );
oa12f01 g34076 ( .a(n37862), .b(n37867), .c(n37866), .o(n37868) );
in01f01 g34077 ( .a(n37864), .o(n37869) );
na02f01 g34078 ( .a(n37869), .b(n37868), .o(n37870) );
na02f01 g34079 ( .a(n37870), .b(n37865), .o(n37871) );
ao12f01 g34080 ( .a(n37871), .b(n26327), .c(n26874), .o(n37872) );
no02f01 g34081 ( .a(n26287), .b(n26279), .o(n37873) );
no02f01 g34082 ( .a(n26293), .b(n26290), .o(n37874) );
no02f01 g34083 ( .a(n37874), .b(n37873), .o(n37875) );
in01f01 g34084 ( .a(n37875), .o(n37876) );
na02f01 g34085 ( .a(n37876), .b(n37871), .o(n37877) );
no02f01 g34086 ( .a(n17825), .b(n17824), .o(n37878) );
in01f01 g34087 ( .a(n37878), .o(n37879) );
in01f01 g34088 ( .a(n37860), .o(n37880) );
na03f01 g34089 ( .a(n37839), .b(n37837), .c(n37835), .o(n37881) );
na03f01 g34090 ( .a(n37881), .b(n37864), .c(n37880), .o(n37882) );
na02f01 g34091 ( .a(n32558), .b(n32510), .o(n37883) );
no02f01 g34092 ( .a(n27144), .b(n7712), .o(n37884) );
ao12f01 g34093 ( .a(n7712), .b(n27134), .c(n37403), .o(n37885) );
no03f01 g34094 ( .a(n37885), .b(n37884), .c(n37883), .o(n37886) );
in01f01 g34095 ( .a(n37816), .o(n37887) );
no02f01 g34096 ( .a(n27144), .b(n7682), .o(n37888) );
no02f01 g34097 ( .a(n37888), .b(n37887), .o(n37889) );
oa12f01 g34098 ( .a(n37889), .b(n27136), .c(n7682), .o(n37890) );
no02f01 g34099 ( .a(n37890), .b(n37886), .o(n37891) );
no03f01 g34100 ( .a(n37823), .b(n37822), .c(n37891), .o(n37892) );
in01f01 g34101 ( .a(n37826), .o(n37893) );
ao12f01 g34102 ( .a(n7682), .b(n27159), .c(n37821), .o(n37894) );
no02f01 g34103 ( .a(n27169), .b(n7682), .o(n37895) );
no02f01 g34104 ( .a(n37895), .b(n37894), .o(n37896) );
oa12f01 g34105 ( .a(n7712), .b(n27182), .c(n27180), .o(n37897) );
na03f01 g34106 ( .a(n37897), .b(n37830), .c(n37896), .o(n37898) );
ao12f01 g34107 ( .a(n37898), .b(n37893), .c(n37892), .o(n37899) );
no03f01 g34108 ( .a(n37838), .b(n37836), .c(n37899), .o(n37900) );
oa12f01 g34109 ( .a(n37869), .b(n37900), .c(n37860), .o(n37901) );
ao12f01 g34110 ( .a(n37879), .b(n37901), .c(n37882), .o(n37902) );
na03f01 g34111 ( .a(n37901), .b(n37882), .c(n37879), .o(n37903) );
no02f01 g34112 ( .a(n17836), .b(n17835), .o(n37904) );
in01f01 g34113 ( .a(n37904), .o(n37905) );
no02f01 g34114 ( .a(n37836), .b(n37899), .o(n37906) );
no02f01 g34115 ( .a(n37860), .b(n37838), .o(n37907) );
in01f01 g34116 ( .a(n37907), .o(n37908) );
no02f01 g34117 ( .a(n37908), .b(n37906), .o(n37909) );
no02f01 g34118 ( .a(n37907), .b(n37866), .o(n37910) );
no02f01 g34119 ( .a(n37910), .b(n37909), .o(n37911) );
na02f01 g34120 ( .a(n37911), .b(n37905), .o(n37912) );
ao12f01 g34121 ( .a(n37902), .b(n37912), .c(n37903), .o(n37913) );
ao12f01 g34122 ( .a(n37871), .b(n37874), .c(n37873), .o(n37914) );
oa12f01 g34123 ( .a(n37877), .b(n37914), .c(n37913), .o(n37915) );
no03f01 g34124 ( .a(n37900), .b(n37869), .c(n37860), .o(n37916) );
ao12f01 g34125 ( .a(n37864), .b(n37881), .c(n37880), .o(n37917) );
oa12f01 g34126 ( .a(n37878), .b(n37917), .c(n37916), .o(n37918) );
no03f01 g34127 ( .a(n37831), .b(n37829), .c(n37892), .o(n37919) );
no02f01 g34128 ( .a(n37836), .b(n37833), .o(n37920) );
oa12f01 g34129 ( .a(n37920), .b(n37919), .c(n37826), .o(n37921) );
na03f01 g34130 ( .a(n37830), .b(n37896), .c(n37825), .o(n37922) );
in01f01 g34131 ( .a(n37920), .o(n37923) );
na03f01 g34132 ( .a(n37923), .b(n37922), .c(n37893), .o(n37924) );
ao12f01 g34133 ( .a(n17830), .b(n37924), .c(n37921), .o(n37925) );
no02f01 g34134 ( .a(n37894), .b(n37822), .o(n37926) );
no03f01 g34135 ( .a(n37895), .b(n37890), .c(n37886), .o(n37927) );
oa12f01 g34136 ( .a(n37926), .b(n37927), .c(n37823), .o(n37928) );
na02f01 g34137 ( .a(n27153), .b(n7682), .o(n37929) );
oa12f01 g34138 ( .a(n7682), .b(n27160), .c(n27158), .o(n37930) );
na02f01 g34139 ( .a(n37827), .b(n37930), .o(n37931) );
na03f01 g34140 ( .a(n37828), .b(n37819), .c(n37815), .o(n37932) );
na03f01 g34141 ( .a(n37932), .b(n37931), .c(n37929), .o(n37933) );
no02f01 g34142 ( .a(n17691), .b(n17784), .o(n37934) );
in01f01 g34143 ( .a(n37934), .o(n37935) );
ao12f01 g34144 ( .a(n17674), .b(n17676), .c(n17804), .o(n37936) );
no02f01 g34145 ( .a(n37936), .b(n37935), .o(n37937) );
na02f01 g34146 ( .a(n37936), .b(n37935), .o(n37938) );
in01f01 g34147 ( .a(n37938), .o(n37939) );
no02f01 g34148 ( .a(n37939), .b(n37937), .o(n37940) );
in01f01 g34149 ( .a(n37940), .o(n37941) );
ao12f01 g34150 ( .a(n37941), .b(n37933), .c(n37928), .o(n37942) );
in01f01 g34151 ( .a(n37942), .o(n37943) );
na02f01 g34152 ( .a(n37404), .b(n7712), .o(n37944) );
na02f01 g34153 ( .a(n37944), .b(n37814), .o(n37945) );
ao12f01 g34154 ( .a(n37818), .b(n37813), .c(n37812), .o(n37946) );
in01f01 g34155 ( .a(n37946), .o(n37947) );
no02f01 g34156 ( .a(n37947), .b(n37945), .o(n37948) );
in01f01 g34157 ( .a(n37945), .o(n37949) );
no02f01 g34158 ( .a(n37946), .b(n37949), .o(n37950) );
no02f01 g34159 ( .a(n17658), .b(n17510), .o(n37951) );
no02f01 g34160 ( .a(n37951), .b(n17797), .o(n37952) );
na02f01 g34161 ( .a(n37951), .b(n17797), .o(n37953) );
in01f01 g34162 ( .a(n37953), .o(n37954) );
no02f01 g34163 ( .a(n37954), .b(n37952), .o(n37955) );
no03f01 g34164 ( .a(n37955), .b(n37950), .c(n37948), .o(n37956) );
na02f01 g34165 ( .a(n37817), .b(n37813), .o(n37957) );
no03f01 g34166 ( .a(n37957), .b(n37887), .c(n37812), .o(n37958) );
no02f01 g34167 ( .a(n37888), .b(n37884), .o(n37959) );
ao12f01 g34168 ( .a(n37959), .b(n37816), .c(n37883), .o(n37960) );
no03f01 g34169 ( .a(n17655), .b(n17770), .c(n17523), .o(n37961) );
ao12f01 g34170 ( .a(n17652), .b(n17771), .c(n17736), .o(n37962) );
no02f01 g34171 ( .a(n37962), .b(n37961), .o(n37963) );
no03f01 g34172 ( .a(n37963), .b(n37960), .c(n37958), .o(n37964) );
in01f01 g34173 ( .a(n37964), .o(n37965) );
ao12f01 g34174 ( .a(n32685), .b(n32729), .c(n32567), .o(n37966) );
na03f01 g34175 ( .a(n37959), .b(n37816), .c(n37883), .o(n37967) );
in01f01 g34176 ( .a(n37960), .o(n37968) );
in01f01 g34177 ( .a(n37963), .o(n37969) );
ao12f01 g34178 ( .a(n37969), .b(n37968), .c(n37967), .o(n37970) );
oa12f01 g34179 ( .a(n37965), .b(n37970), .c(n37966), .o(n37971) );
oa12f01 g34180 ( .a(n37955), .b(n37950), .c(n37948), .o(n37972) );
ao12f01 g34181 ( .a(n37956), .b(n37972), .c(n37971), .o(n37973) );
na04f01 g34182 ( .a(n37828), .b(n37929), .c(n37819), .d(n37815), .o(n37974) );
oa12f01 g34183 ( .a(n37820), .b(n37895), .c(n37823), .o(n37975) );
na02f01 g34184 ( .a(n37975), .b(n37974), .o(n37976) );
no02f01 g34185 ( .a(n17778), .b(n17674), .o(n37977) );
no02f01 g34186 ( .a(n37977), .b(n17804), .o(n37978) );
na02f01 g34187 ( .a(n37977), .b(n17804), .o(n37979) );
in01f01 g34188 ( .a(n37979), .o(n37980) );
no02f01 g34189 ( .a(n37980), .b(n37978), .o(n37981) );
na02f01 g34190 ( .a(n37981), .b(n37976), .o(n37982) );
in01f01 g34191 ( .a(n37982), .o(n37983) );
ao12f01 g34192 ( .a(n37931), .b(n37932), .c(n37929), .o(n37984) );
no03f01 g34193 ( .a(n37927), .b(n37926), .c(n37823), .o(n37985) );
no03f01 g34194 ( .a(n37940), .b(n37985), .c(n37984), .o(n37986) );
in01f01 g34195 ( .a(n37981), .o(n37987) );
na03f01 g34196 ( .a(n37987), .b(n37975), .c(n37974), .o(n37988) );
in01f01 g34197 ( .a(n37988), .o(n37989) );
no02f01 g34198 ( .a(n37989), .b(n37986), .o(n37990) );
oa12f01 g34199 ( .a(n37990), .b(n37983), .c(n37973), .o(n37991) );
oa22f01 g34200 ( .a(n37831), .b(n37826), .c(n37829), .d(n37892), .o(n37992) );
na04f01 g34201 ( .a(n37830), .b(n37896), .c(n37893), .d(n37825), .o(n37993) );
ao12f01 g34202 ( .a(n17833), .b(n37993), .c(n37992), .o(n37994) );
in01f01 g34203 ( .a(n37994), .o(n37995) );
na03f01 g34204 ( .a(n37995), .b(n37991), .c(n37943), .o(n37996) );
ao12f01 g34205 ( .a(n37923), .b(n37922), .c(n37893), .o(n37997) );
no03f01 g34206 ( .a(n37920), .b(n37919), .c(n37826), .o(n37998) );
no03f01 g34207 ( .a(n37998), .b(n37997), .c(n17809), .o(n37999) );
na03f01 g34208 ( .a(n37993), .b(n37992), .c(n17833), .o(n38000) );
in01f01 g34209 ( .a(n38000), .o(n38001) );
no02f01 g34210 ( .a(n38001), .b(n37999), .o(n38002) );
ao12f01 g34211 ( .a(n37925), .b(n38002), .c(n37996), .o(n38003) );
no02f01 g34212 ( .a(n37911), .b(n37905), .o(n38004) );
in01f01 g34213 ( .a(n38004), .o(n38005) );
na04f01 g34214 ( .a(n38005), .b(n38003), .c(n37918), .d(n37877), .o(n38006) );
na02f01 g34215 ( .a(n38006), .b(n37915), .o(n38007) );
no02f01 g34216 ( .a(n37869), .b(n37868), .o(n38008) );
ao12f01 g34217 ( .a(n37864), .b(n37862), .c(n37859), .o(n38009) );
no02f01 g34218 ( .a(n38009), .b(n38008), .o(n38010) );
ao12f01 g34219 ( .a(n38010), .b(n26336), .c(n26332), .o(n38011) );
in01f01 g34220 ( .a(n38011), .o(n38012) );
ao12f01 g34221 ( .a(n37872), .b(n38012), .c(n38007), .o(n38013) );
no02f01 g34222 ( .a(n37871), .b(n26388), .o(n38014) );
no02f01 g34223 ( .a(n38010), .b(n26347), .o(n38015) );
no02f01 g34224 ( .a(n38015), .b(n38014), .o(n38016) );
na02f01 g34225 ( .a(n38016), .b(n38013), .o(n38017) );
in01f01 g34226 ( .a(n37872), .o(n38018) );
no02f01 g34227 ( .a(n37875), .b(n38010), .o(n38019) );
no03f01 g34228 ( .a(n37917), .b(n37916), .c(n37878), .o(n38020) );
na02f01 g34229 ( .a(n37907), .b(n37866), .o(n38021) );
na02f01 g34230 ( .a(n37908), .b(n37906), .o(n38022) );
na02f01 g34231 ( .a(n38022), .b(n38021), .o(n38023) );
no02f01 g34232 ( .a(n38023), .b(n37904), .o(n38024) );
oa12f01 g34233 ( .a(n37918), .b(n38024), .c(n38020), .o(n38025) );
in01f01 g34234 ( .a(n37873), .o(n38026) );
in01f01 g34235 ( .a(n37874), .o(n38027) );
oa12f01 g34236 ( .a(n38010), .b(n38027), .c(n38026), .o(n38028) );
ao12f01 g34237 ( .a(n38019), .b(n38028), .c(n38025), .o(n38029) );
in01f01 g34238 ( .a(n37925), .o(n38030) );
na02f01 g34239 ( .a(n37946), .b(n37949), .o(n38031) );
na02f01 g34240 ( .a(n37947), .b(n37945), .o(n38032) );
in01f01 g34241 ( .a(n37955), .o(n38033) );
na03f01 g34242 ( .a(n38033), .b(n38032), .c(n38031), .o(n38034) );
oa12f01 g34243 ( .a(n32564), .b(n32683), .c(n32686), .o(n38035) );
oa12f01 g34244 ( .a(n37963), .b(n37960), .c(n37958), .o(n38036) );
ao12f01 g34245 ( .a(n37964), .b(n38036), .c(n38035), .o(n38037) );
ao12f01 g34246 ( .a(n38033), .b(n38032), .c(n38031), .o(n38038) );
oa12f01 g34247 ( .a(n38034), .b(n38038), .c(n38037), .o(n38039) );
na03f01 g34248 ( .a(n37941), .b(n37933), .c(n37928), .o(n38040) );
na02f01 g34249 ( .a(n37988), .b(n38040), .o(n38041) );
ao12f01 g34250 ( .a(n38041), .b(n37982), .c(n38039), .o(n38042) );
no03f01 g34251 ( .a(n37994), .b(n38042), .c(n37942), .o(n38043) );
na03f01 g34252 ( .a(n37924), .b(n37921), .c(n17830), .o(n38044) );
na02f01 g34253 ( .a(n38000), .b(n38044), .o(n38045) );
oa12f01 g34254 ( .a(n38030), .b(n38045), .c(n38043), .o(n38046) );
no04f01 g34255 ( .a(n38004), .b(n38046), .c(n37902), .d(n38019), .o(n38047) );
no02f01 g34256 ( .a(n38047), .b(n38029), .o(n38048) );
oa12f01 g34257 ( .a(n38018), .b(n38011), .c(n38048), .o(n38049) );
in01f01 g34258 ( .a(n38016), .o(n38050) );
na02f01 g34259 ( .a(n38050), .b(n38049), .o(n38051) );
na03f01 g34260 ( .a(n38051), .b(n38017), .c(n1821), .o(n38052) );
na02f01 g34261 ( .a(n38051), .b(n38017), .o(n1845) );
na02f01 g34262 ( .a(n1845), .b(n8066), .o(n38054) );
na02f01 g34263 ( .a(n38054), .b(n38052), .o(n579) );
in01f01 g34264 ( .a(n11007), .o(n38056) );
in01f01 g34265 ( .a(n11008), .o(n38057) );
na03f01 g34266 ( .a(n38057), .b(n10995), .c(n10797), .o(n38058) );
ao12f01 g34267 ( .a(n10636), .b(n10658), .c(n10632), .o(n38059) );
in01f01 g34268 ( .a(n38059), .o(n38060) );
no02f01 g34269 ( .a(n38060), .b(n10681), .o(n38061) );
no02f01 g34270 ( .a(n10683), .b(n4088), .o(n38062) );
no02f01 g34271 ( .a(n38062), .b(n10677), .o(n38063) );
no02f01 g34272 ( .a(n38063), .b(n38061), .o(n38064) );
na02f01 g34273 ( .a(n38063), .b(n38061), .o(n38065) );
in01f01 g34274 ( .a(n38065), .o(n38066) );
no03f01 g34275 ( .a(n38066), .b(n38064), .c(n10735), .o(n38067) );
no02f01 g34276 ( .a(n38066), .b(n38064), .o(n38068) );
no02f01 g34277 ( .a(n38068), .b(n3521), .o(n38069) );
no02f01 g34278 ( .a(n38069), .b(n38067), .o(n38070) );
in01f01 g34279 ( .a(n38070), .o(n38071) );
na03f01 g34280 ( .a(n38071), .b(n38058), .c(n38056), .o(n38072) );
na02f01 g34281 ( .a(n38058), .b(n38056), .o(n38073) );
na02f01 g34282 ( .a(n38070), .b(n38073), .o(n38074) );
na02f01 g34283 ( .a(n38074), .b(n38072), .o(n584) );
na02f01 g34284 ( .a(n11717), .b(n11716), .o(n38076) );
in01f01 g34285 ( .a(n11735), .o(n38077) );
no02f01 g34286 ( .a(n38077), .b(n38076), .o(n38078) );
in01f01 g34287 ( .a(n38078), .o(n38079) );
no02f01 g34288 ( .a(n11762), .b(n11746), .o(n38080) );
na03f01 g34289 ( .a(n38080), .b(n11760), .c(n38079), .o(n38081) );
in01f01 g34290 ( .a(n38080), .o(n38082) );
oa12f01 g34291 ( .a(n38082), .b(n11761), .c(n38078), .o(n38083) );
na02f01 g34292 ( .a(n38083), .b(n38081), .o(n589) );
no02f01 g34293 ( .a(n6068), .b(n6056_1), .o(n38085) );
in01f01 g34294 ( .a(n38085), .o(n38086) );
in01f01 g34295 ( .a(n5895), .o(n38087) );
no02f01 g34296 ( .a(n38087), .b(n6037), .o(n38088) );
no03f01 g34297 ( .a(n38088), .b(n38086), .c(n34414), .o(n38089) );
in01f01 g34298 ( .a(n38089), .o(n38090) );
ao12f01 g34299 ( .a(n38090), .b(n6049), .c(n6046), .o(n38091) );
no02f01 g34300 ( .a(n5842), .b(n5818), .o(n38092) );
in01f01 g34301 ( .a(n38092), .o(n38093) );
no02f01 g34302 ( .a(n5858), .b(n5856), .o(n38094) );
oa12f01 g34303 ( .a(n38094), .b(n38093), .c(n5837), .o(n38095) );
no02f01 g34304 ( .a(n38095), .b(n5860), .o(n38096) );
no02f01 g34305 ( .a(n38096), .b(n5850), .o(n38097) );
no02f01 g34306 ( .a(n5854_1), .b(n5829_1), .o(n38098) );
in01f01 g34307 ( .a(n38098), .o(n38099) );
no02f01 g34308 ( .a(n38099), .b(n38097), .o(n38100) );
na02f01 g34309 ( .a(n38099), .b(n38097), .o(n38101) );
in01f01 g34310 ( .a(n38101), .o(n38102) );
no02f01 g34311 ( .a(n38102), .b(n38100), .o(n38103) );
in01f01 g34312 ( .a(n38103), .o(n38104) );
no02f01 g34313 ( .a(n38104), .b(n5873), .o(n38105) );
in01f01 g34314 ( .a(n5818), .o(n38106) );
no02f01 g34315 ( .a(n5858), .b(n5842), .o(n38107) );
in01f01 g34316 ( .a(n38107), .o(n38108) );
no02f01 g34317 ( .a(n38108), .b(n38106), .o(n38109) );
no02f01 g34318 ( .a(n38107), .b(n5818), .o(n38110) );
no02f01 g34319 ( .a(n38110), .b(n38109), .o(n38111) );
in01f01 g34320 ( .a(n38111), .o(n38112) );
no02f01 g34321 ( .a(n38112), .b(n5873), .o(n38113) );
no02f01 g34322 ( .a(n38092), .b(n5858), .o(n38114) );
no02f01 g34323 ( .a(n5856), .b(n5837), .o(n38115) );
no02f01 g34324 ( .a(n38115), .b(n38114), .o(n38116) );
na02f01 g34325 ( .a(n38115), .b(n38114), .o(n38117) );
in01f01 g34326 ( .a(n38117), .o(n38118) );
no03f01 g34327 ( .a(n38118), .b(n38116), .c(n5873), .o(n38119) );
no02f01 g34328 ( .a(n38119), .b(n38113), .o(n38120) );
in01f01 g34329 ( .a(n38120), .o(n38121) );
in01f01 g34330 ( .a(n38095), .o(n38122) );
no02f01 g34331 ( .a(n5860), .b(n5850), .o(n38123) );
no02f01 g34332 ( .a(n38123), .b(n38122), .o(n38124) );
na02f01 g34333 ( .a(n38123), .b(n38122), .o(n38125) );
in01f01 g34334 ( .a(n38125), .o(n38126) );
no03f01 g34335 ( .a(n38126), .b(n38124), .c(n5873), .o(n38127) );
no02f01 g34336 ( .a(n38127), .b(n38121), .o(n38128) );
in01f01 g34337 ( .a(n38128), .o(n38129) );
no02f01 g34338 ( .a(n38129), .b(n38105), .o(n38130) );
ao12f01 g34339 ( .a(n6037), .b(n6066_1), .c(n5883_1), .o(n38131) );
oa12f01 g34340 ( .a(n38085), .b(n38131), .c(n5896), .o(n38132) );
in01f01 g34341 ( .a(n38132), .o(n38133) );
no02f01 g34342 ( .a(n38126), .b(n38124), .o(n38134) );
no02f01 g34343 ( .a(n38134), .b(n6037), .o(n38135) );
oa12f01 g34344 ( .a(n5873), .b(n38135), .c(n38104), .o(n38136) );
no02f01 g34345 ( .a(n38118), .b(n38116), .o(n38137) );
ao12f01 g34346 ( .a(n6037), .b(n38137), .c(n38111), .o(n38138) );
in01f01 g34347 ( .a(n38138), .o(n38139) );
na02f01 g34348 ( .a(n38139), .b(n38136), .o(n38140) );
ao12f01 g34349 ( .a(n38140), .b(n38133), .c(n38130), .o(n38141) );
in01f01 g34350 ( .a(n38141), .o(n38142) );
ao12f01 g34351 ( .a(n38142), .b(n38130), .c(n38091), .o(n38143) );
in01f01 g34352 ( .a(n5863), .o(n38144) );
no02f01 g34353 ( .a(n38144), .b(n5543_1), .o(n38145) );
in01f01 g34354 ( .a(n38145), .o(n38146) );
no02f01 g34355 ( .a(n38146), .b(n5862), .o(n38147) );
in01f01 g34356 ( .a(n5862), .o(n38148) );
no02f01 g34357 ( .a(n38145), .b(n38148), .o(n38149) );
no02f01 g34358 ( .a(n38149), .b(n38147), .o(n38150) );
in01f01 g34359 ( .a(n38150), .o(n38151) );
no02f01 g34360 ( .a(n38151), .b(n5873), .o(n38152) );
no02f01 g34361 ( .a(n38150), .b(n6037), .o(n38153) );
no02f01 g34362 ( .a(n38153), .b(n38152), .o(n38154) );
na02f01 g34363 ( .a(n38154), .b(n38143), .o(n38155) );
na02f01 g34364 ( .a(n6025), .b(n6008), .o(n38156) );
na02f01 g34365 ( .a(n6045), .b(n6037_1), .o(n38157) );
no02f01 g34366 ( .a(n38157), .b(n38156), .o(n38158) );
in01f01 g34367 ( .a(n6049), .o(n38159) );
oa12f01 g34368 ( .a(n38089), .b(n38159), .c(n38158), .o(n38160) );
in01f01 g34369 ( .a(n38130), .o(n38161) );
oa12f01 g34370 ( .a(n38141), .b(n38161), .c(n38160), .o(n38162) );
in01f01 g34371 ( .a(n38154), .o(n38163) );
na02f01 g34372 ( .a(n38163), .b(n38162), .o(n38164) );
na02f01 g34373 ( .a(n38164), .b(n38155), .o(n594) );
in01f01 g34374 ( .a(n37384), .o(n38166) );
no03f01 g34375 ( .a(n9224), .b(n8899), .c(beta_31), .o(n38167) );
no02f01 g34376 ( .a(n38167), .b(n9602), .o(n38168) );
ao12f01 g34377 ( .a(n9596), .b(n38168), .c(n38166), .o(n38169) );
no02f01 g34378 ( .a(n38169), .b(n9610), .o(n38170) );
na02f01 g34379 ( .a(n38169), .b(n9610), .o(n38171) );
in01f01 g34380 ( .a(n38171), .o(n38172) );
no02f01 g34381 ( .a(n38172), .b(n38170), .o(n38173) );
in01f01 g34382 ( .a(n38173), .o(n599) );
in01f01 g34383 ( .a(n14208), .o(n38175) );
no02f01 g34384 ( .a(n38175), .b(n14035), .o(n38176) );
in01f01 g34385 ( .a(n14209), .o(n38177) );
no02f01 g34386 ( .a(n38177), .b(n14020), .o(n38178) );
in01f01 g34387 ( .a(n38178), .o(n38179) );
no02f01 g34388 ( .a(n38179), .b(n38176), .o(n38180) );
na02f01 g34389 ( .a(n38179), .b(n38176), .o(n38181) );
in01f01 g34390 ( .a(n38181), .o(n38182) );
no02f01 g34391 ( .a(n38182), .b(n38180), .o(n38183) );
in01f01 g34392 ( .a(n38183), .o(n604) );
in01f01 g34393 ( .a(n22334), .o(n38185) );
no02f01 g34394 ( .a(n22356), .b(n22347), .o(n38186) );
in01f01 g34395 ( .a(n38186), .o(n38187) );
no03f01 g34396 ( .a(n38187), .b(n22355), .c(n38185), .o(n38188) );
no02f01 g34397 ( .a(n22355), .b(n38185), .o(n38189) );
no02f01 g34398 ( .a(n38186), .b(n38189), .o(n38190) );
no02f01 g34399 ( .a(n38190), .b(n38188), .o(n38191) );
in01f01 g34400 ( .a(n38191), .o(n609) );
no02f01 g34401 ( .a(n15923), .b(n15866), .o(n38193) );
in01f01 g34402 ( .a(n38193), .o(n38194) );
no02f01 g34403 ( .a(n27395), .b(n38194), .o(n38195) );
no02f01 g34404 ( .a(n38195), .b(n27640), .o(n38196) );
in01f01 g34405 ( .a(n38196), .o(n38197) );
ao12f01 g34406 ( .a(n27367), .b(n15987), .c(n38193), .o(n38198) );
no03f01 g34407 ( .a(n38198), .b(n27677), .c(n27676), .o(n38199) );
no02f01 g34408 ( .a(n15990), .b(n15972), .o(n38200) );
in01f01 g34409 ( .a(n38200), .o(n38201) );
no02f01 g34410 ( .a(n27395), .b(n38201), .o(n38202) );
no02f01 g34411 ( .a(n27367), .b(n38200), .o(n38203) );
no02f01 g34412 ( .a(n38203), .b(n38202), .o(n38204) );
oa12f01 g34413 ( .a(n38204), .b(n38199), .c(n38197), .o(n38205) );
in01f01 g34414 ( .a(n38198), .o(n38206) );
na03f01 g34415 ( .a(n38206), .b(n27638), .c(n27624), .o(n38207) );
in01f01 g34416 ( .a(n38204), .o(n38208) );
na03f01 g34417 ( .a(n38208), .b(n38207), .c(n38196), .o(n38209) );
na02f01 g34418 ( .a(n38209), .b(n38205), .o(n614) );
na02f01 g34419 ( .a(n32037), .b(n_22641), .o(n38211) );
na02f01 g34420 ( .a(n32105), .b(n_22641), .o(n38212) );
oa12f01 g34421 ( .a(n_22641), .b(n32078), .c(n32423), .o(n38213) );
na02f01 g34422 ( .a(n32061), .b(n_22641), .o(n38214) );
na02f01 g34423 ( .a(n38214), .b(n38213), .o(n38215) );
no02f01 g34424 ( .a(n32092), .b(n32026), .o(n38216) );
no02f01 g34425 ( .a(n32090), .b(n31965), .o(n38217) );
no02f01 g34426 ( .a(n38217), .b(n38216), .o(n38218) );
no02f01 g34427 ( .a(n38218), .b(n6075), .o(n38219) );
no02f01 g34428 ( .a(n38219), .b(n38215), .o(n38220) );
na02f01 g34429 ( .a(n38220), .b(n38212), .o(n38221) );
no02f01 g34430 ( .a(n32128), .b(n6075), .o(n38222) );
no02f01 g34431 ( .a(n32117), .b(n6075), .o(n38223) );
no03f01 g34432 ( .a(n38223), .b(n38222), .c(n38221), .o(n38224) );
na02f01 g34433 ( .a(n38224), .b(n38211), .o(n38225) );
no02f01 g34434 ( .a(n32103), .b(n32101), .o(n38226) );
no02f01 g34435 ( .a(n32099), .b(n32097), .o(n38227) );
no02f01 g34436 ( .a(n38227), .b(n38226), .o(n38228) );
ao12f01 g34437 ( .a(n_22641), .b(n32117), .c(n38228), .o(n38229) );
ao12f01 g34438 ( .a(n_22641), .b(n32128), .c(n32033), .o(n38230) );
no02f01 g34439 ( .a(n38230), .b(n38229), .o(n38231) );
na02f01 g34440 ( .a(n36871), .b(n_22641), .o(n38232) );
in01f01 g34441 ( .a(n38232), .o(n38233) );
ao12f01 g34442 ( .a(n38233), .b(n38231), .c(n38225), .o(n38234) );
na02f01 g34443 ( .a(n36850), .b(n_22641), .o(n38235) );
na02f01 g34444 ( .a(n38235), .b(n38234), .o(n38236) );
no02f01 g34445 ( .a(n36882), .b(n6075), .o(n38237) );
no02f01 g34446 ( .a(n38237), .b(n38236), .o(n38238) );
ao12f01 g34447 ( .a(n_22641), .b(n36877), .c(n36880), .o(n38239) );
no02f01 g34448 ( .a(n36882), .b(n_22641), .o(n38240) );
no03f01 g34449 ( .a(n38240), .b(n38239), .c(n38238), .o(n38241) );
no02f01 g34450 ( .a(n36838), .b(n6075), .o(n38242) );
no02f01 g34451 ( .a(n36838), .b(n_22641), .o(n38243) );
no02f01 g34452 ( .a(n38243), .b(n38242), .o(n38244) );
no02f01 g34453 ( .a(n38244), .b(n38241), .o(n38245) );
no02f01 g34454 ( .a(n32033), .b(n6075), .o(n38246) );
no02f01 g34455 ( .a(n38228), .b(n6075), .o(n38247) );
no03f01 g34456 ( .a(n32076), .b(n32075), .c(n32064), .o(n38248) );
ao12f01 g34457 ( .a(n32069), .b(n32073), .c(n32065), .o(n38249) );
no02f01 g34458 ( .a(n38249), .b(n38248), .o(n38250) );
ao12f01 g34459 ( .a(n6075), .b(n38250), .c(n32050), .o(n38251) );
ao12f01 g34460 ( .a(n6075), .b(n32060), .c(n32056), .o(n38252) );
no02f01 g34461 ( .a(n38252), .b(n38251), .o(n38253) );
na02f01 g34462 ( .a(n32094), .b(n_22641), .o(n38254) );
na02f01 g34463 ( .a(n38254), .b(n38253), .o(n38255) );
no02f01 g34464 ( .a(n38255), .b(n38247), .o(n38256) );
in01f01 g34465 ( .a(n38222), .o(n38257) );
na02f01 g34466 ( .a(n32432), .b(n_22641), .o(n38258) );
na03f01 g34467 ( .a(n38258), .b(n38257), .c(n38256), .o(n38259) );
no02f01 g34468 ( .a(n38259), .b(n38246), .o(n38260) );
in01f01 g34469 ( .a(n38229), .o(n38261) );
no02f01 g34470 ( .a(n32128), .b(n_22641), .o(n38262) );
oa12f01 g34471 ( .a(n6075), .b(n38262), .c(n32037), .o(n38263) );
na02f01 g34472 ( .a(n38263), .b(n38261), .o(n38264) );
oa12f01 g34473 ( .a(n38232), .b(n38264), .c(n38260), .o(n38265) );
no02f01 g34474 ( .a(n36880), .b(n6075), .o(n38266) );
no02f01 g34475 ( .a(n38266), .b(n38265), .o(n38267) );
na02f01 g34476 ( .a(n36861), .b(n_22641), .o(n38268) );
na02f01 g34477 ( .a(n38268), .b(n38267), .o(n38269) );
in01f01 g34478 ( .a(n38239), .o(n38270) );
na02f01 g34479 ( .a(n36861), .b(n6075), .o(n38271) );
na03f01 g34480 ( .a(n38271), .b(n38270), .c(n38269), .o(n38272) );
in01f01 g34481 ( .a(n38244), .o(n38273) );
no02f01 g34482 ( .a(n38273), .b(n38272), .o(n38274) );
no02f01 g34483 ( .a(n31161), .b(n31010), .o(n38275) );
no02f01 g34484 ( .a(n31162), .b(n31000), .o(n38276) );
no02f01 g34485 ( .a(n38276), .b(n38275), .o(n38277) );
na02f01 g34486 ( .a(n38276), .b(n38275), .o(n38278) );
in01f01 g34487 ( .a(n38278), .o(n38279) );
no02f01 g34488 ( .a(n38279), .b(n38277), .o(n38280) );
in01f01 g34489 ( .a(n38280), .o(n38281) );
no03f01 g34490 ( .a(n38281), .b(n38274), .c(n38245), .o(n38282) );
no02f01 g34491 ( .a(n31157), .b(n31023), .o(n38283) );
no02f01 g34492 ( .a(n31160), .b(n31010), .o(n38284) );
in01f01 g34493 ( .a(n38284), .o(n38285) );
no02f01 g34494 ( .a(n38285), .b(n38283), .o(n38286) );
na02f01 g34495 ( .a(n38285), .b(n38283), .o(n38287) );
in01f01 g34496 ( .a(n38287), .o(n38288) );
no02f01 g34497 ( .a(n38288), .b(n38286), .o(n38289) );
na02f01 g34498 ( .a(n38270), .b(n38236), .o(n38290) );
na02f01 g34499 ( .a(n38271), .b(n38268), .o(n38291) );
na02f01 g34500 ( .a(n38291), .b(n38290), .o(n38292) );
no02f01 g34501 ( .a(n38239), .b(n38267), .o(n38293) );
no02f01 g34502 ( .a(n38240), .b(n38237), .o(n38294) );
na02f01 g34503 ( .a(n38294), .b(n38293), .o(n38295) );
ao12f01 g34504 ( .a(n38289), .b(n38295), .c(n38292), .o(n38296) );
na02f01 g34505 ( .a(n36871), .b(n6075), .o(n38297) );
no02f01 g34506 ( .a(n36880), .b(n_22641), .o(n38298) );
no02f01 g34507 ( .a(n38298), .b(n38266), .o(n38299) );
na03f01 g34508 ( .a(n38299), .b(n38297), .c(n38265), .o(n38300) );
in01f01 g34509 ( .a(n38297), .o(n38301) );
na02f01 g34510 ( .a(n36850), .b(n6075), .o(n38302) );
na02f01 g34511 ( .a(n38302), .b(n38235), .o(n38303) );
oa12f01 g34512 ( .a(n38303), .b(n38301), .c(n38234), .o(n38304) );
no04f01 g34513 ( .a(n31156), .b(n31154), .c(n31033), .d(n31023), .o(n38305) );
ao22f01 g34514 ( .a(n31440), .b(n31410), .c(n31439), .d(n31411), .o(n38306) );
no02f01 g34515 ( .a(n38306), .b(n38305), .o(n38307) );
na03f01 g34516 ( .a(n38307), .b(n38304), .c(n38300), .o(n38308) );
ao12f01 g34517 ( .a(n38307), .b(n38304), .c(n38300), .o(n38309) );
no02f01 g34518 ( .a(n38264), .b(n38260), .o(n38310) );
na02f01 g34519 ( .a(n38297), .b(n38232), .o(n38311) );
in01f01 g34520 ( .a(n38311), .o(n38312) );
na02f01 g34521 ( .a(n38312), .b(n38310), .o(n38313) );
in01f01 g34522 ( .a(n38310), .o(n38314) );
na02f01 g34523 ( .a(n38311), .b(n38314), .o(n38315) );
no02f01 g34524 ( .a(n31150), .b(n31045), .o(n38316) );
in01f01 g34525 ( .a(n38316), .o(n38317) );
no02f01 g34526 ( .a(n31153), .b(n31033), .o(n38318) );
no02f01 g34527 ( .a(n38318), .b(n38317), .o(n38319) );
na02f01 g34528 ( .a(n38318), .b(n38317), .o(n38320) );
in01f01 g34529 ( .a(n38320), .o(n38321) );
no02f01 g34530 ( .a(n38321), .b(n38319), .o(n38322) );
ao12f01 g34531 ( .a(n38322), .b(n38315), .c(n38313), .o(n38323) );
oa12f01 g34532 ( .a(n38308), .b(n38323), .c(n38309), .o(n38324) );
no02f01 g34533 ( .a(n38262), .b(n38229), .o(n38325) );
in01f01 g34534 ( .a(n38325), .o(n38326) );
na02f01 g34535 ( .a(n32037), .b(n6075), .o(n38327) );
na02f01 g34536 ( .a(n38327), .b(n38211), .o(n38328) );
no03f01 g34537 ( .a(n38328), .b(n38326), .c(n38224), .o(n38329) );
no02f01 g34538 ( .a(n32033), .b(n_22641), .o(n38330) );
no02f01 g34539 ( .a(n38330), .b(n38246), .o(n38331) );
ao12f01 g34540 ( .a(n38331), .b(n38325), .c(n38259), .o(n38332) );
no04f01 g34541 ( .a(n31149), .b(n31146), .c(n31056), .d(n31045), .o(n38333) );
ao22f01 g34542 ( .a(n31436), .b(n31412), .c(n31435), .d(n31413), .o(n38334) );
no02f01 g34543 ( .a(n38334), .b(n38333), .o(n38335) );
in01f01 g34544 ( .a(n38335), .o(n38336) );
no03f01 g34545 ( .a(n38336), .b(n38332), .c(n38329), .o(n38337) );
in01f01 g34546 ( .a(n38337), .o(n38338) );
no04f01 g34547 ( .a(n31141), .b(n31138), .c(n31091), .d(n31081), .o(n38339) );
ao22f01 g34548 ( .a(n31432), .b(n31414), .c(n31431), .d(n31415), .o(n38340) );
no02f01 g34549 ( .a(n38340), .b(n38339), .o(n38341) );
in01f01 g34550 ( .a(n38341), .o(n38342) );
no02f01 g34551 ( .a(n38228), .b(n_22641), .o(n38343) );
no02f01 g34552 ( .a(n32117), .b(n_22641), .o(n38344) );
no04f01 g34553 ( .a(n38344), .b(n38343), .c(n38223), .d(n38256), .o(n38345) );
in01f01 g34554 ( .a(n38343), .o(n38346) );
no02f01 g34555 ( .a(n38344), .b(n38223), .o(n38347) );
ao12f01 g34556 ( .a(n38347), .b(n38346), .c(n38221), .o(n38348) );
no03f01 g34557 ( .a(n38348), .b(n38345), .c(n38342), .o(n38349) );
in01f01 g34558 ( .a(n38349), .o(n38350) );
oa12f01 g34559 ( .a(n38220), .b(n38343), .c(n38247), .o(n38351) );
in01f01 g34560 ( .a(n38351), .o(n38352) );
no03f01 g34561 ( .a(n38343), .b(n38220), .c(n38247), .o(n38353) );
no02f01 g34562 ( .a(n31094), .b(n31091), .o(n38354) );
no02f01 g34563 ( .a(n38354), .b(n31137), .o(n38355) );
na02f01 g34564 ( .a(n38354), .b(n31137), .o(n38356) );
in01f01 g34565 ( .a(n38356), .o(n38357) );
no02f01 g34566 ( .a(n38357), .b(n38355), .o(n38358) );
in01f01 g34567 ( .a(n38358), .o(n38359) );
oa12f01 g34568 ( .a(n38359), .b(n38353), .c(n38352), .o(n38360) );
no02f01 g34569 ( .a(n38218), .b(n_22641), .o(n38361) );
no02f01 g34570 ( .a(n38361), .b(n38219), .o(n38362) );
na02f01 g34571 ( .a(n38362), .b(n38215), .o(n38363) );
na02f01 g34572 ( .a(n32094), .b(n6075), .o(n38364) );
na02f01 g34573 ( .a(n38364), .b(n38254), .o(n38365) );
na02f01 g34574 ( .a(n38365), .b(n38253), .o(n38366) );
no03f01 g34575 ( .a(n31429), .b(n31135), .c(n31102), .o(n38367) );
no02f01 g34576 ( .a(n31429), .b(n31102), .o(n38368) );
no02f01 g34577 ( .a(n38368), .b(n31426), .o(n38369) );
no02f01 g34578 ( .a(n38369), .b(n38367), .o(n38370) );
ao12f01 g34579 ( .a(n38370), .b(n38366), .c(n38363), .o(n38371) );
na03f01 g34580 ( .a(n32077), .b(n32074), .c(n_22641), .o(n38372) );
na03f01 g34581 ( .a(n32077), .b(n32074), .c(n6075), .o(n38373) );
in01f01 g34582 ( .a(n31117), .o(n38374) );
no02f01 g34583 ( .a(n38374), .b(n31114), .o(n38375) );
no02f01 g34584 ( .a(n31117), .b(n32070), .o(n38376) );
no02f01 g34585 ( .a(n38376), .b(n38375), .o(n38377) );
in01f01 g34586 ( .a(n38377), .o(n38378) );
na03f01 g34587 ( .a(n38378), .b(n38373), .c(n38372), .o(n38379) );
no02f01 g34588 ( .a(n31133), .b(n31127), .o(n38380) );
no02f01 g34589 ( .a(n31424), .b(n31125), .o(n38381) );
no03f01 g34590 ( .a(n38381), .b(n38380), .c(n31118), .o(n38382) );
no02f01 g34591 ( .a(n38381), .b(n38380), .o(n38383) );
no02f01 g34592 ( .a(n38383), .b(n31119), .o(n38384) );
no02f01 g34593 ( .a(n38384), .b(n38382), .o(n38385) );
no02f01 g34594 ( .a(n38385), .b(n38379), .o(n38386) );
na03f01 g34595 ( .a(n32078), .b(n32050), .c(n_22641), .o(n38387) );
oa12f01 g34596 ( .a(n32423), .b(n38250), .c(n6075), .o(n38388) );
na02f01 g34597 ( .a(n38388), .b(n38387), .o(n38389) );
na02f01 g34598 ( .a(n38385), .b(n38379), .o(n38390) );
ao12f01 g34599 ( .a(n38386), .b(n38390), .c(n38389), .o(n38391) );
ao12f01 g34600 ( .a(n_22641), .b(n32060), .c(n32056), .o(n38392) );
no03f01 g34601 ( .a(n38392), .b(n38252), .c(n38213), .o(n38393) );
na02f01 g34602 ( .a(n32061), .b(n6075), .o(n38394) );
ao12f01 g34603 ( .a(n38251), .b(n38394), .c(n38214), .o(n38395) );
no03f01 g34604 ( .a(n31425), .b(n31113), .c(n31419), .o(n38396) );
ao12f01 g34605 ( .a(n31134), .b(n31420), .c(n31112), .o(n38397) );
no02f01 g34606 ( .a(n38397), .b(n38396), .o(n38398) );
in01f01 g34607 ( .a(n38398), .o(n38399) );
no03f01 g34608 ( .a(n38399), .b(n38395), .c(n38393), .o(n38400) );
oa12f01 g34609 ( .a(n38399), .b(n38395), .c(n38393), .o(n38401) );
oa12f01 g34610 ( .a(n38401), .b(n38400), .c(n38391), .o(n38402) );
na03f01 g34611 ( .a(n38370), .b(n38366), .c(n38363), .o(n38403) );
ao12f01 g34612 ( .a(n38371), .b(n38403), .c(n38402), .o(n38404) );
no03f01 g34613 ( .a(n38359), .b(n38353), .c(n38352), .o(n38405) );
oa12f01 g34614 ( .a(n38360), .b(n38405), .c(n38404), .o(n38406) );
oa12f01 g34615 ( .a(n38342), .b(n38348), .c(n38345), .o(n38407) );
in01f01 g34616 ( .a(n38407), .o(n38408) );
oa12f01 g34617 ( .a(n38350), .b(n38408), .c(n38406), .o(n38409) );
no02f01 g34618 ( .a(n38223), .b(n38247), .o(n38410) );
ao12f01 g34619 ( .a(n38229), .b(n38410), .c(n38220), .o(n38411) );
no02f01 g34620 ( .a(n38262), .b(n38222), .o(n38412) );
no02f01 g34621 ( .a(n38412), .b(n38411), .o(n38413) );
na02f01 g34622 ( .a(n38258), .b(n38212), .o(n38414) );
oa12f01 g34623 ( .a(n38261), .b(n38414), .c(n38255), .o(n38415) );
in01f01 g34624 ( .a(n38412), .o(n38416) );
no02f01 g34625 ( .a(n38416), .b(n38415), .o(n38417) );
no02f01 g34626 ( .a(n38417), .b(n38413), .o(n38418) );
no02f01 g34627 ( .a(n31142), .b(n31081), .o(n38419) );
in01f01 g34628 ( .a(n38419), .o(n38420) );
no02f01 g34629 ( .a(n31145), .b(n31056), .o(n38421) );
no02f01 g34630 ( .a(n38421), .b(n38420), .o(n38422) );
na02f01 g34631 ( .a(n38421), .b(n38420), .o(n38423) );
in01f01 g34632 ( .a(n38423), .o(n38424) );
no02f01 g34633 ( .a(n38424), .b(n38422), .o(n38425) );
na02f01 g34634 ( .a(n38425), .b(n38418), .o(n38426) );
in01f01 g34635 ( .a(n38426), .o(n38427) );
na03f01 g34636 ( .a(n38331), .b(n38325), .c(n38259), .o(n38428) );
oa12f01 g34637 ( .a(n38328), .b(n38326), .c(n38224), .o(n38429) );
ao12f01 g34638 ( .a(n38335), .b(n38429), .c(n38428), .o(n38430) );
in01f01 g34639 ( .a(n38425), .o(n38431) );
oa12f01 g34640 ( .a(n38431), .b(n38417), .c(n38413), .o(n38432) );
in01f01 g34641 ( .a(n38432), .o(n38433) );
no02f01 g34642 ( .a(n38433), .b(n38430), .o(n38434) );
oa12f01 g34643 ( .a(n38434), .b(n38427), .c(n38409), .o(n38435) );
na03f01 g34644 ( .a(n38322), .b(n38315), .c(n38313), .o(n38436) );
na04f01 g34645 ( .a(n38436), .b(n38435), .c(n38338), .d(n38308), .o(n38437) );
in01f01 g34646 ( .a(n38289), .o(n38438) );
no02f01 g34647 ( .a(n38294), .b(n38293), .o(n38439) );
no02f01 g34648 ( .a(n38291), .b(n38290), .o(n38440) );
no03f01 g34649 ( .a(n38440), .b(n38439), .c(n38438), .o(n38441) );
ao12f01 g34650 ( .a(n38441), .b(n38437), .c(n38324), .o(n38442) );
na02f01 g34651 ( .a(n38273), .b(n38272), .o(n38443) );
na02f01 g34652 ( .a(n38244), .b(n38241), .o(n38444) );
ao12f01 g34653 ( .a(n38280), .b(n38444), .c(n38443), .o(n38445) );
no03f01 g34654 ( .a(n38445), .b(n38442), .c(n38296), .o(n38446) );
no02f01 g34655 ( .a(n38242), .b(n38269), .o(n38447) );
oa12f01 g34656 ( .a(n6075), .b(n36861), .c(n36839), .o(n38448) );
na02f01 g34657 ( .a(n38448), .b(n38270), .o(n38449) );
no02f01 g34658 ( .a(n38449), .b(n38447), .o(n38450) );
no02f01 g34659 ( .a(n36827), .b(n6075), .o(n38451) );
no02f01 g34660 ( .a(n36827), .b(n_22641), .o(n38452) );
no02f01 g34661 ( .a(n38452), .b(n38451), .o(n38453) );
na02f01 g34662 ( .a(n38453), .b(n38450), .o(n38454) );
in01f01 g34663 ( .a(n38242), .o(n38455) );
na02f01 g34664 ( .a(n38455), .b(n38238), .o(n38456) );
in01f01 g34665 ( .a(n38449), .o(n38457) );
na02f01 g34666 ( .a(n38457), .b(n38456), .o(n38458) );
in01f01 g34667 ( .a(n38453), .o(n38459) );
na02f01 g34668 ( .a(n38459), .b(n38458), .o(n38460) );
na02f01 g34669 ( .a(n38460), .b(n38454), .o(n38461) );
no02f01 g34670 ( .a(n31163), .b(n31000), .o(n38462) );
no03f01 g34671 ( .a(n31452), .b(n31174), .c(n38462), .o(n38463) );
in01f01 g34672 ( .a(n38462), .o(n38464) );
ao12f01 g34673 ( .a(n38464), .b(n31177), .c(n31448), .o(n38465) );
no02f01 g34674 ( .a(n38465), .b(n38463), .o(n38466) );
in01f01 g34675 ( .a(n38466), .o(n38467) );
no02f01 g34676 ( .a(n38467), .b(n38461), .o(n38468) );
no03f01 g34677 ( .a(n38468), .b(n38446), .c(n38282), .o(n38469) );
in01f01 g34678 ( .a(n38451), .o(n38470) );
na02f01 g34679 ( .a(n38470), .b(n38447), .o(n38471) );
no02f01 g34680 ( .a(n38452), .b(n38449), .o(n38472) );
no02f01 g34681 ( .a(n31666), .b(n30593), .o(n38473) );
no02f01 g34682 ( .a(n31664), .b(n30591), .o(n38474) );
no02f01 g34683 ( .a(n38474), .b(n38473), .o(n38475) );
in01f01 g34684 ( .a(n38475), .o(n38476) );
no03f01 g34685 ( .a(n36820), .b(n36819), .c(n36804), .o(n38477) );
in01f01 g34686 ( .a(n38477), .o(n38478) );
no02f01 g34687 ( .a(n36822), .b(n36803), .o(n38479) );
na02f01 g34688 ( .a(n38479), .b(n38478), .o(n38480) );
no02f01 g34689 ( .a(n38480), .b(n38476), .o(n38481) );
na02f01 g34690 ( .a(n38480), .b(n38476), .o(n38482) );
in01f01 g34691 ( .a(n38482), .o(n38483) );
no02f01 g34692 ( .a(n38483), .b(n38481), .o(n38484) );
no02f01 g34693 ( .a(n38484), .b(n6075), .o(n38485) );
no02f01 g34694 ( .a(n38484), .b(n_22641), .o(n38486) );
no02f01 g34695 ( .a(n38486), .b(n38485), .o(n38487) );
ao12f01 g34696 ( .a(n38487), .b(n38472), .c(n38471), .o(n38488) );
no02f01 g34697 ( .a(n38451), .b(n38456), .o(n38489) );
in01f01 g34698 ( .a(n38472), .o(n38490) );
in01f01 g34699 ( .a(n38481), .o(n38491) );
na02f01 g34700 ( .a(n38482), .b(n38491), .o(n38492) );
na02f01 g34701 ( .a(n38492), .b(n_22641), .o(n38493) );
na02f01 g34702 ( .a(n38492), .b(n6075), .o(n38494) );
na02f01 g34703 ( .a(n38494), .b(n38493), .o(n38495) );
no03f01 g34704 ( .a(n38495), .b(n38490), .c(n38489), .o(n38496) );
no02f01 g34705 ( .a(n38496), .b(n38488), .o(n38497) );
ao12f01 g34706 ( .a(n31174), .b(n31177), .c(n38464), .o(n38498) );
no02f01 g34707 ( .a(n31451), .b(n30987), .o(n38499) );
in01f01 g34708 ( .a(n38499), .o(n38500) );
no02f01 g34709 ( .a(n38500), .b(n38498), .o(n38501) );
na02f01 g34710 ( .a(n38500), .b(n38498), .o(n38502) );
in01f01 g34711 ( .a(n38502), .o(n38503) );
no02f01 g34712 ( .a(n38503), .b(n38501), .o(n38504) );
na02f01 g34713 ( .a(n38467), .b(n38461), .o(n38505) );
oa12f01 g34714 ( .a(n38505), .b(n38504), .c(n38497), .o(n38506) );
no02f01 g34715 ( .a(n38506), .b(n38469), .o(n38507) );
na02f01 g34716 ( .a(n38504), .b(n38497), .o(n38508) );
in01f01 g34717 ( .a(n38508), .o(n38509) );
no02f01 g34718 ( .a(n38509), .b(n38507), .o(n38510) );
in01f01 g34719 ( .a(n38510), .o(n38511) );
ao12f01 g34720 ( .a(n_22641), .b(n38484), .c(n36827), .o(n38512) );
no03f01 g34721 ( .a(n38485), .b(n38451), .c(n38450), .o(n38513) );
no02f01 g34722 ( .a(n31666), .b(n30619), .o(n38514) );
no02f01 g34723 ( .a(n31664), .b(n30616), .o(n38515) );
no02f01 g34724 ( .a(n38515), .b(n38514), .o(n38516) );
in01f01 g34725 ( .a(n38516), .o(n38517) );
no02f01 g34726 ( .a(n38480), .b(n30593), .o(n38518) );
oa22f01 g34727 ( .a(n38518), .b(n31664), .c(n38478), .d(n30591), .o(n38519) );
no02f01 g34728 ( .a(n38519), .b(n38517), .o(n38520) );
na02f01 g34729 ( .a(n38519), .b(n38517), .o(n38521) );
in01f01 g34730 ( .a(n38521), .o(n38522) );
oa12f01 g34731 ( .a(n_22641), .b(n38522), .c(n38520), .o(n38523) );
oa12f01 g34732 ( .a(n6075), .b(n38522), .c(n38520), .o(n38524) );
na02f01 g34733 ( .a(n38524), .b(n38523), .o(n38525) );
oa12f01 g34734 ( .a(n38525), .b(n38513), .c(n38512), .o(n38526) );
in01f01 g34735 ( .a(n38512), .o(n38527) );
na03f01 g34736 ( .a(n38493), .b(n38470), .c(n38458), .o(n38528) );
in01f01 g34737 ( .a(n38520), .o(n38529) );
ao12f01 g34738 ( .a(n6075), .b(n38521), .c(n38529), .o(n38530) );
ao12f01 g34739 ( .a(n_22641), .b(n38521), .c(n38529), .o(n38531) );
no02f01 g34740 ( .a(n38531), .b(n38530), .o(n38532) );
na03f01 g34741 ( .a(n38532), .b(n38528), .c(n38527), .o(n38533) );
no03f01 g34742 ( .a(n31212), .b(n31191), .c(n31454), .o(n38534) );
ao12f01 g34743 ( .a(n31179), .b(n31457), .c(n31455), .o(n38535) );
no02f01 g34744 ( .a(n38535), .b(n38534), .o(n38536) );
ao12f01 g34745 ( .a(n38536), .b(n38533), .c(n38526), .o(n38537) );
ao12f01 g34746 ( .a(n38532), .b(n38528), .c(n38527), .o(n38538) );
no03f01 g34747 ( .a(n38525), .b(n38513), .c(n38512), .o(n38539) );
in01f01 g34748 ( .a(n38536), .o(n38540) );
no03f01 g34749 ( .a(n38540), .b(n38539), .c(n38538), .o(n38541) );
no02f01 g34750 ( .a(n38541), .b(n38537), .o(n38542) );
na02f01 g34751 ( .a(n38542), .b(n38511), .o(n38543) );
in01f01 g34752 ( .a(n38542), .o(n38544) );
na02f01 g34753 ( .a(n38544), .b(n38510), .o(n38545) );
na02f01 g34754 ( .a(n38545), .b(n38543), .o(n619) );
no02f01 g34755 ( .a(n26836), .b(n26440), .o(n38547) );
in01f01 g34756 ( .a(n26836), .o(n38548) );
no02f01 g34757 ( .a(n38548), .b(n26441), .o(n38549) );
no02f01 g34758 ( .a(n38549), .b(n38547), .o(n38550) );
no02f01 g34759 ( .a(n26828), .b(n26440), .o(n38551) );
in01f01 g34760 ( .a(n38551), .o(n38552) );
na03f01 g34761 ( .a(n27111), .b(n27068), .c(n26870), .o(n38553) );
na02f01 g34762 ( .a(n27247), .b(n38553), .o(n38554) );
in01f01 g34763 ( .a(n26828), .o(n38555) );
no02f01 g34764 ( .a(n38555), .b(n26441), .o(n38556) );
in01f01 g34765 ( .a(n38556), .o(n38557) );
na02f01 g34766 ( .a(n38557), .b(n38554), .o(n38558) );
na03f01 g34767 ( .a(n38558), .b(n38552), .c(n38550), .o(n38559) );
in01f01 g34768 ( .a(n38550), .o(n38560) );
no03f01 g34769 ( .a(n27110), .b(n27238), .c(n26869), .o(n38561) );
no02f01 g34770 ( .a(n27119), .b(n38561), .o(n38562) );
oa12f01 g34771 ( .a(n38552), .b(n38556), .c(n38562), .o(n38563) );
na02f01 g34772 ( .a(n38563), .b(n38560), .o(n38564) );
na02f01 g34773 ( .a(n38564), .b(n38559), .o(n624) );
na03f01 g34774 ( .a(n32459), .b(n32323), .c(n32303), .o(n38566) );
oa12f01 g34775 ( .a(n32458), .b(n32324), .c(n32449), .o(n38567) );
na02f01 g34776 ( .a(n38567), .b(n38566), .o(n629) );
in01f01 g34777 ( .a(n22680), .o(n38569) );
in01f01 g34778 ( .a(n22683), .o(n38570) );
no02f01 g34779 ( .a(n22731), .b(n22693), .o(n38571) );
in01f01 g34780 ( .a(n38571), .o(n38572) );
oa12f01 g34781 ( .a(n38572), .b(n38570), .c(n38569), .o(n38573) );
no02f01 g34782 ( .a(n38570), .b(n38569), .o(n38574) );
na02f01 g34783 ( .a(n38571), .b(n38574), .o(n38575) );
na02f01 g34784 ( .a(n38575), .b(n38573), .o(n634) );
na02f01 g34785 ( .a(n36797), .b(n36793), .o(n639) );
in01f01 g34786 ( .a(n22239), .o(n38578) );
ao12f01 g34787 ( .a(n22246), .b(n22249), .c(n38578), .o(n38579) );
in01f01 g34788 ( .a(n38579), .o(n38580) );
in01f01 g34789 ( .a(n22155), .o(n38581) );
na02f01 g34790 ( .a(n22248), .b(n38581), .o(n38582) );
in01f01 g34791 ( .a(n38582), .o(n38583) );
no02f01 g34792 ( .a(n38583), .b(n38580), .o(n38584) );
no02f01 g34793 ( .a(n38582), .b(n38579), .o(n38585) );
no02f01 g34794 ( .a(n38585), .b(n38584), .o(n38586) );
na02f01 g34795 ( .a(n38586), .b(n2589), .o(n38587) );
in01f01 g34796 ( .a(n38586), .o(n3020) );
na02f01 g34797 ( .a(n3020), .b(n4116), .o(n38589) );
na02f01 g34798 ( .a(n38589), .b(n38587), .o(n644) );
na02f01 g34799 ( .a(n32732), .b(sin_out_11), .o(n38591) );
no04f01 g34800 ( .a(n36579), .b(n34393), .c(n34369), .d(n34348), .o(n38592) );
in01f01 g34801 ( .a(n36591), .o(n38593) );
in01f01 g34802 ( .a(n36594), .o(n38594) );
ao12f01 g34803 ( .a(n38594), .b(n38593), .c(n38592), .o(n38595) );
no02f01 g34804 ( .a(n36613), .b(n36597), .o(n38596) );
in01f01 g34805 ( .a(n38596), .o(n38597) );
no02f01 g34806 ( .a(n38597), .b(n38595), .o(n38598) );
ao12f01 g34807 ( .a(n35673), .b(n36544), .c(n35893), .o(n38599) );
no02f01 g34808 ( .a(n35667), .b(n34287), .o(n38600) );
no02f01 g34809 ( .a(n38600), .b(n35669), .o(n38601) );
no02f01 g34810 ( .a(n38601), .b(n38599), .o(n38602) );
na02f01 g34811 ( .a(n38601), .b(n38599), .o(n38603) );
in01f01 g34812 ( .a(n38603), .o(n38604) );
no02f01 g34813 ( .a(n38604), .b(n38602), .o(n38605) );
in01f01 g34814 ( .a(n38605), .o(n38606) );
no02f01 g34815 ( .a(n38606), .b(n34267), .o(n38607) );
in01f01 g34816 ( .a(n38607), .o(n38608) );
ao12f01 g34817 ( .a(n34307), .b(n36610), .c(n36552), .o(n38609) );
in01f01 g34818 ( .a(n38609), .o(n38610) );
no02f01 g34819 ( .a(n38605), .b(n34307), .o(n38611) );
in01f01 g34820 ( .a(n38611), .o(n38612) );
na02f01 g34821 ( .a(n38612), .b(n38610), .o(n38613) );
ao12f01 g34822 ( .a(n38613), .b(n38608), .c(n38598), .o(n38614) );
in01f01 g34823 ( .a(n38614), .o(n38615) );
no03f01 g34824 ( .a(n35669), .b(n36545), .c(n35618), .o(n38616) );
no02f01 g34825 ( .a(n38600), .b(n35673), .o(n38617) );
in01f01 g34826 ( .a(n38617), .o(n38618) );
no02f01 g34827 ( .a(n35659), .b(n34287), .o(n38619) );
no02f01 g34828 ( .a(n38619), .b(n35661), .o(n38620) );
in01f01 g34829 ( .a(n38620), .o(n38621) );
no03f01 g34830 ( .a(n38621), .b(n38618), .c(n38616), .o(n38622) );
no02f01 g34831 ( .a(n38618), .b(n38616), .o(n38623) );
no02f01 g34832 ( .a(n38620), .b(n38623), .o(n38624) );
no02f01 g34833 ( .a(n38624), .b(n38622), .o(n38625) );
no02f01 g34834 ( .a(n38625), .b(n34307), .o(n38626) );
in01f01 g34835 ( .a(n38625), .o(n38627) );
no02f01 g34836 ( .a(n38627), .b(n34267), .o(n38628) );
no02f01 g34837 ( .a(n38628), .b(n38626), .o(n38629) );
in01f01 g34838 ( .a(n38629), .o(n38630) );
no02f01 g34839 ( .a(n38630), .b(n38615), .o(n38631) );
no02f01 g34840 ( .a(n38629), .b(n38614), .o(n38632) );
oa12f01 g34841 ( .a(n32734), .b(n38632), .c(n38631), .o(n38633) );
na02f01 g34842 ( .a(n38633), .b(n38591), .o(n649) );
in01f01 g34843 ( .a(n5964), .o(n38635) );
na02f01 g34844 ( .a(n6003_1), .b(n38635), .o(n38636) );
no02f01 g34845 ( .a(n6013), .b(n5873), .o(n38637) );
no03f01 g34846 ( .a(n38637), .b(n6006), .c(n6005), .o(n38638) );
oa12f01 g34847 ( .a(n38638), .b(n6015), .c(n38636), .o(n38639) );
in01f01 g34848 ( .a(n38639), .o(n38640) );
no02f01 g34849 ( .a(n6022_1), .b(n5873), .o(n38641) );
no02f01 g34850 ( .a(n38641), .b(n6024), .o(n38642) );
na02f01 g34851 ( .a(n38642), .b(n38640), .o(n38643) );
in01f01 g34852 ( .a(n38642), .o(n38644) );
na02f01 g34853 ( .a(n38644), .b(n38639), .o(n38645) );
na02f01 g34854 ( .a(n38645), .b(n38643), .o(n653) );
na02f01 g34855 ( .a(n21186), .b(n21131), .o(n38647) );
no02f01 g34856 ( .a(n21189), .b(n21119), .o(n38648) );
in01f01 g34857 ( .a(n38648), .o(n38649) );
na02f01 g34858 ( .a(n38649), .b(n38647), .o(n38650) );
na03f01 g34859 ( .a(n38648), .b(n21186), .c(n21131), .o(n38651) );
na02f01 g34860 ( .a(n38651), .b(n38650), .o(n658) );
no02f01 g34861 ( .a(n22632), .b(n22501), .o(n38653) );
in01f01 g34862 ( .a(n22643), .o(n38654) );
ao12f01 g34863 ( .a(n22654), .b(n38654), .c(n38653), .o(n38655) );
no02f01 g34864 ( .a(n22655), .b(n22652), .o(n38656) );
na02f01 g34865 ( .a(n38656), .b(n38655), .o(n38657) );
in01f01 g34866 ( .a(n38655), .o(n38658) );
in01f01 g34867 ( .a(n38656), .o(n38659) );
na02f01 g34868 ( .a(n38659), .b(n38658), .o(n38660) );
na02f01 g34869 ( .a(n38660), .b(n38657), .o(n663) );
no02f01 g34870 ( .a(n37069), .b(n36963), .o(n38662) );
in01f01 g34871 ( .a(n38662), .o(n38663) );
no02f01 g34872 ( .a(n37070), .b(n36972), .o(n38664) );
ao12f01 g34873 ( .a(n38664), .b(n38663), .c(n37062), .o(n38665) );
in01f01 g34874 ( .a(n38665), .o(n38666) );
no02f01 g34875 ( .a(n37078), .b(n36963), .o(n38667) );
no02f01 g34876 ( .a(n37079), .b(n36972), .o(n38668) );
no02f01 g34877 ( .a(n38668), .b(n38667), .o(n38669) );
na02f01 g34878 ( .a(n38669), .b(n38666), .o(n38670) );
in01f01 g34879 ( .a(n38669), .o(n38671) );
na02f01 g34880 ( .a(n38671), .b(n38665), .o(n38672) );
na02f01 g34881 ( .a(n38672), .b(n38670), .o(n668) );
ao12f01 g34882 ( .a(n4635), .b(n4630), .c(n4697_1), .o(n38674) );
no02f01 g34883 ( .a(n4354_1), .b(n4344_1), .o(n38675) );
no02f01 g34884 ( .a(n4355), .b(n4340), .o(n38676) );
no02f01 g34885 ( .a(n38676), .b(n38675), .o(n38677) );
no02f01 g34886 ( .a(n38677), .b(n38674), .o(n38678) );
na02f01 g34887 ( .a(n38677), .b(n38674), .o(n38679) );
in01f01 g34888 ( .a(n38679), .o(n38680) );
no02f01 g34889 ( .a(n38680), .b(n38678), .o(n38681) );
in01f01 g34890 ( .a(n38681), .o(n38682) );
no02f01 g34891 ( .a(n38682), .b(n36038), .o(n38683) );
in01f01 g34892 ( .a(n38683), .o(n38684) );
ao12f01 g34893 ( .a(n36038), .b(n36200), .c(n36187), .o(n38685) );
no02f01 g34894 ( .a(n38685), .b(n36215), .o(n38686) );
na02f01 g34895 ( .a(n38686), .b(n38684), .o(n38687) );
in01f01 g34896 ( .a(n38687), .o(n38688) );
oa12f01 g34897 ( .a(n38688), .b(n36170), .c(n36166), .o(n38689) );
no02f01 g34898 ( .a(n38676), .b(n38674), .o(n38690) );
no02f01 g34899 ( .a(n38690), .b(n38675), .o(n38691) );
no02f01 g34900 ( .a(n4367), .b(n4340), .o(n38692) );
no02f01 g34901 ( .a(n4366), .b(n4344_1), .o(n38693) );
no02f01 g34902 ( .a(n38693), .b(n38692), .o(n38694) );
no02f01 g34903 ( .a(n38694), .b(n38691), .o(n38695) );
na02f01 g34904 ( .a(n38694), .b(n38691), .o(n38696) );
in01f01 g34905 ( .a(n38696), .o(n38697) );
no02f01 g34906 ( .a(n38697), .b(n38695), .o(n38698) );
in01f01 g34907 ( .a(n38698), .o(n38699) );
no02f01 g34908 ( .a(n38699), .b(n36038), .o(n38700) );
no02f01 g34909 ( .a(n4693), .b(n4692_1), .o(n38701) );
no02f01 g34910 ( .a(n4647), .b(n4643_1), .o(n38702) );
no02f01 g34911 ( .a(n38702), .b(n38701), .o(n38703) );
na02f01 g34912 ( .a(n38702), .b(n38701), .o(n38704) );
in01f01 g34913 ( .a(n38704), .o(n38705) );
no02f01 g34914 ( .a(n38705), .b(n38703), .o(n38706) );
in01f01 g34915 ( .a(n38706), .o(n38707) );
no02f01 g34916 ( .a(n38707), .b(n36038), .o(n38708) );
no02f01 g34917 ( .a(n36038), .b(n4927_1), .o(n38709) );
no02f01 g34918 ( .a(n38709), .b(n38708), .o(n38710) );
in01f01 g34919 ( .a(n38710), .o(n38711) );
no03f01 g34920 ( .a(n38711), .b(n38700), .c(n38689), .o(n38712) );
ao12f01 g34921 ( .a(n36122), .b(n36212), .c(n36196), .o(n38713) );
no02f01 g34922 ( .a(n38713), .b(n36198), .o(n38714) );
in01f01 g34923 ( .a(n38714), .o(n38715) );
ao12f01 g34924 ( .a(n36122), .b(n38698), .c(n38681), .o(n38716) );
no02f01 g34925 ( .a(n38716), .b(n38715), .o(n38717) );
ao12f01 g34926 ( .a(n36122), .b(n38706), .c(n4696), .o(n38718) );
in01f01 g34927 ( .a(n38718), .o(n38719) );
na02f01 g34928 ( .a(n38719), .b(n38717), .o(n38720) );
no02f01 g34929 ( .a(n4937_1), .b(n4751_1), .o(n38721) );
in01f01 g34930 ( .a(n38721), .o(n38722) );
no02f01 g34931 ( .a(n36038), .b(n38722), .o(n38723) );
no02f01 g34932 ( .a(n36038), .b(n4930), .o(n38724) );
no02f01 g34933 ( .a(n38724), .b(n38723), .o(n38725) );
no02f01 g34934 ( .a(n36038), .b(n4782), .o(n38726) );
no02f01 g34935 ( .a(n36038), .b(n4814), .o(n38727) );
no02f01 g34936 ( .a(n38727), .b(n38726), .o(n38728) );
na02f01 g34937 ( .a(n38728), .b(n38725), .o(n38729) );
in01f01 g34938 ( .a(n36937), .o(n38730) );
no02f01 g34939 ( .a(n38730), .b(n36038), .o(n38731) );
in01f01 g34940 ( .a(n36925), .o(n38732) );
no02f01 g34941 ( .a(n38732), .b(n36038), .o(n38733) );
no02f01 g34942 ( .a(n38733), .b(n38731), .o(n38734) );
in01f01 g34943 ( .a(n38734), .o(n38735) );
in01f01 g34944 ( .a(n36950), .o(n38736) );
no02f01 g34945 ( .a(n38736), .b(n36038), .o(n38737) );
no03f01 g34946 ( .a(n38737), .b(n38735), .c(n38729), .o(n38738) );
oa12f01 g34947 ( .a(n38738), .b(n38720), .c(n38712), .o(n38739) );
ao12f01 g34948 ( .a(n36122), .b(n38721), .c(n4729), .o(n38740) );
ao12f01 g34949 ( .a(n36122), .b(n4807), .c(n4785), .o(n38741) );
no02f01 g34950 ( .a(n38741), .b(n38740), .o(n38742) );
in01f01 g34951 ( .a(n38742), .o(n38743) );
no02f01 g34952 ( .a(n38730), .b(n38732), .o(n38744) );
ao12f01 g34953 ( .a(n36122), .b(n38744), .c(n36950), .o(n38745) );
no02f01 g34954 ( .a(n38745), .b(n38743), .o(n38746) );
no02f01 g34955 ( .a(n36913), .b(n36122), .o(n38747) );
na02f01 g34956 ( .a(n36913), .b(n36122), .o(n38748) );
in01f01 g34957 ( .a(n38748), .o(n38749) );
no02f01 g34958 ( .a(n38749), .b(n38747), .o(n38750) );
na03f01 g34959 ( .a(n38750), .b(n38746), .c(n38739), .o(n38751) );
ao12f01 g34960 ( .a(n38750), .b(n38746), .c(n38739), .o(n38752) );
in01f01 g34961 ( .a(n38752), .o(n38753) );
na03f01 g34962 ( .a(n38753), .b(n38751), .c(delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(n38754) );
na02f01 g34963 ( .a(n38753), .b(n38751), .o(n2687) );
na02f01 g34964 ( .a(n2687), .b(n37149), .o(n38756) );
no04f01 g34965 ( .a(n38724), .b(n38711), .c(n38700), .d(n38689), .o(n38757) );
no02f01 g34966 ( .a(n36122), .b(n4729), .o(n38758) );
no02f01 g34967 ( .a(n38758), .b(n38720), .o(n38759) );
in01f01 g34968 ( .a(n38759), .o(n38760) );
no02f01 g34969 ( .a(n36122), .b(n38721), .o(n38761) );
no02f01 g34970 ( .a(n38761), .b(n38723), .o(n38762) );
in01f01 g34971 ( .a(n38762), .o(n38763) );
oa12f01 g34972 ( .a(n38763), .b(n38760), .c(n38757), .o(n38764) );
in01f01 g34973 ( .a(n36057), .o(n38765) );
in01f01 g34974 ( .a(n36076), .o(n38766) );
ao12f01 g34975 ( .a(n7435), .b(n7521), .c(n7524), .o(n38767) );
oa12f01 g34976 ( .a(n36067), .b(n36066), .c(n36012), .o(n38768) );
na03f01 g34977 ( .a(n36064), .b(n36061), .c(n36060), .o(n38769) );
ao12f01 g34978 ( .a(n36074), .b(n38769), .c(n38768), .o(n38770) );
no02f01 g34979 ( .a(n36091), .b(n38770), .o(n38771) );
oa12f01 g34980 ( .a(n38771), .b(n36088), .c(n38767), .o(n38772) );
no03f01 g34981 ( .a(n36100), .b(n36099), .c(n36098), .o(n38773) );
ao12f01 g34982 ( .a(n36095), .b(n36035), .c(n36030), .o(n38774) );
no02f01 g34983 ( .a(n38774), .b(n38773), .o(n38775) );
na02f01 g34984 ( .a(n36105), .b(n38775), .o(n38776) );
na02f01 g34985 ( .a(n36113), .b(n36122), .o(n38777) );
na04f01 g34986 ( .a(n38777), .b(n38776), .c(n38772), .d(n38766), .o(n38778) );
no02f01 g34987 ( .a(n36105), .b(n38775), .o(n38779) );
no02f01 g34988 ( .a(n36113), .b(n36122), .o(n38780) );
oa12f01 g34989 ( .a(n38777), .b(n38780), .c(n38779), .o(n38781) );
in01f01 g34990 ( .a(n36123), .o(n38782) );
na03f01 g34991 ( .a(n38782), .b(n38781), .c(n38778), .o(n38783) );
in01f01 g34992 ( .a(n36142), .o(n38784) );
na04f01 g34993 ( .a(n36164), .b(n38784), .c(n38783), .d(n38765), .o(n38785) );
ao12f01 g34994 ( .a(n38687), .b(n36169), .c(n38785), .o(n38786) );
in01f01 g34995 ( .a(n38700), .o(n38787) );
in01f01 g34996 ( .a(n38724), .o(n38788) );
na04f01 g34997 ( .a(n38788), .b(n38710), .c(n38787), .d(n38786), .o(n38789) );
na03f01 g34998 ( .a(n38762), .b(n38759), .c(n38789), .o(n38790) );
ao12f01 g34999 ( .a(n37149), .b(n38790), .c(n38764), .o(n38791) );
no02f01 g35000 ( .a(n38758), .b(n38724), .o(n38792) );
in01f01 g35001 ( .a(n38792), .o(n38793) );
oa12f01 g35002 ( .a(n38793), .b(n38720), .c(n38712), .o(n38794) );
na03f01 g35003 ( .a(n38710), .b(n38787), .c(n38786), .o(n38795) );
in01f01 g35004 ( .a(n38720), .o(n38796) );
na03f01 g35005 ( .a(n38792), .b(n38796), .c(n38795), .o(n38797) );
ao12f01 g35006 ( .a(n37149), .b(n38797), .c(n38794), .o(n38798) );
na04f01 g35007 ( .a(n38725), .b(n38710), .c(n38787), .d(n38786), .o(n38799) );
no02f01 g35008 ( .a(n38740), .b(n38720), .o(n38800) );
no02f01 g35009 ( .a(n36122), .b(n4785), .o(n38801) );
no02f01 g35010 ( .a(n38801), .b(n38726), .o(n38802) );
na03f01 g35011 ( .a(n38802), .b(n38800), .c(n38799), .o(n38803) );
in01f01 g35012 ( .a(n38725), .o(n38804) );
no04f01 g35013 ( .a(n38804), .b(n38711), .c(n38700), .d(n38689), .o(n38805) );
in01f01 g35014 ( .a(n38800), .o(n38806) );
in01f01 g35015 ( .a(n38802), .o(n38807) );
oa12f01 g35016 ( .a(n38807), .b(n38806), .c(n38805), .o(n38808) );
ao12f01 g35017 ( .a(n37149), .b(n38808), .c(n38803), .o(n38809) );
no03f01 g35018 ( .a(n38809), .b(n38798), .c(n38791), .o(n38810) );
no02f01 g35019 ( .a(n36122), .b(n4807), .o(n38811) );
no02f01 g35020 ( .a(n38811), .b(n38727), .o(n38812) );
no03f01 g35021 ( .a(n38806), .b(n38805), .c(n38801), .o(n38813) );
no03f01 g35022 ( .a(n38813), .b(n38812), .c(n38726), .o(n38814) );
in01f01 g35023 ( .a(n38726), .o(n38815) );
in01f01 g35024 ( .a(n38812), .o(n38816) );
in01f01 g35025 ( .a(n38801), .o(n38817) );
na03f01 g35026 ( .a(n38800), .b(n38799), .c(n38817), .o(n38818) );
ao12f01 g35027 ( .a(n38816), .b(n38818), .c(n38815), .o(n38819) );
oa12f01 g35028 ( .a(delay_sub_ln23_0_unr23_stage8_stallmux_q), .b(n38819), .c(n38814), .o(n38820) );
no04f01 g35029 ( .a(n38729), .b(n38711), .c(n38700), .d(n38689), .o(n38821) );
no02f01 g35030 ( .a(n38743), .b(n38720), .o(n38822) );
in01f01 g35031 ( .a(n38822), .o(n38823) );
no02f01 g35032 ( .a(n38823), .b(n38821), .o(n38824) );
no02f01 g35033 ( .a(n36925), .b(n36122), .o(n38825) );
no02f01 g35034 ( .a(n38825), .b(n38733), .o(n38826) );
na02f01 g35035 ( .a(n38826), .b(n38824), .o(n38827) );
in01f01 g35036 ( .a(n38729), .o(n38828) );
na04f01 g35037 ( .a(n38828), .b(n38710), .c(n38787), .d(n38786), .o(n38829) );
na02f01 g35038 ( .a(n38822), .b(n38829), .o(n38830) );
in01f01 g35039 ( .a(n38826), .o(n38831) );
na02f01 g35040 ( .a(n38831), .b(n38830), .o(n38832) );
ao12f01 g35041 ( .a(n37149), .b(n38832), .c(n38827), .o(n38833) );
in01f01 g35042 ( .a(n38833), .o(n38834) );
no02f01 g35043 ( .a(n36937), .b(n36122), .o(n38835) );
no02f01 g35044 ( .a(n38835), .b(n38731), .o(n38836) );
no03f01 g35045 ( .a(n38825), .b(n38823), .c(n38821), .o(n38837) );
no03f01 g35046 ( .a(n38837), .b(n38836), .c(n38733), .o(n38838) );
in01f01 g35047 ( .a(n38733), .o(n38839) );
in01f01 g35048 ( .a(n38836), .o(n38840) );
in01f01 g35049 ( .a(n38825), .o(n38841) );
na03f01 g35050 ( .a(n38841), .b(n38822), .c(n38829), .o(n38842) );
ao12f01 g35051 ( .a(n38840), .b(n38842), .c(n38839), .o(n38843) );
oa12f01 g35052 ( .a(delay_sub_ln23_0_unr23_stage8_stallmux_q), .b(n38843), .c(n38838), .o(n38844) );
na04f01 g35053 ( .a(n38844), .b(n38834), .c(n38820), .d(n38810), .o(n38845) );
no02f01 g35054 ( .a(n36950), .b(n36122), .o(n38846) );
no02f01 g35055 ( .a(n38846), .b(n38737), .o(n38847) );
no02f01 g35056 ( .a(n38744), .b(n36122), .o(n38848) );
no02f01 g35057 ( .a(n38830), .b(n38848), .o(n38849) );
oa12f01 g35058 ( .a(n38847), .b(n38849), .c(n38735), .o(n38850) );
in01f01 g35059 ( .a(n38847), .o(n38851) );
in01f01 g35060 ( .a(n38848), .o(n38852) );
na02f01 g35061 ( .a(n38824), .b(n38852), .o(n38853) );
na03f01 g35062 ( .a(n38853), .b(n38851), .c(n38734), .o(n38854) );
ao12f01 g35063 ( .a(n37149), .b(n38854), .c(n38850), .o(n38855) );
no02f01 g35064 ( .a(n38855), .b(n38845), .o(n38856) );
ao22f01 g35065 ( .a(n38856), .b(delay_sub_ln23_0_unr23_stage8_stallmux_q), .c(n38756), .d(n38754), .o(n673) );
oa12f01 g35066 ( .a(n9232), .b(n9591), .c(n9228), .o(n38858) );
in01f01 g35067 ( .a(n38858), .o(n678) );
ao12f01 g35068 ( .a(n22302), .b(n22313), .c(n22296), .o(n38860) );
in01f01 g35069 ( .a(n38860), .o(n38861) );
no02f01 g35070 ( .a(n22317), .b(n22312), .o(n38862) );
no02f01 g35071 ( .a(n38862), .b(n38861), .o(n38863) );
na02f01 g35072 ( .a(n38862), .b(n38861), .o(n38864) );
in01f01 g35073 ( .a(n38864), .o(n38865) );
no02f01 g35074 ( .a(n38865), .b(n38863), .o(n38866) );
in01f01 g35075 ( .a(n38866), .o(n683) );
no02f01 g35076 ( .a(n37413), .b(n37407), .o(n38868) );
na02f01 g35077 ( .a(n38868), .b(n37418), .o(n38869) );
in01f01 g35078 ( .a(n38868), .o(n38870) );
na02f01 g35079 ( .a(n38870), .b(n37409), .o(n38871) );
na02f01 g35080 ( .a(n38871), .b(n38869), .o(n688) );
in01f01 g35081 ( .a(n36189), .o(n38873) );
na02f01 g35082 ( .a(n36201), .b(n36197), .o(n38874) );
in01f01 g35083 ( .a(n38874), .o(n38875) );
na03f01 g35084 ( .a(n38875), .b(n36199), .c(n38873), .o(n38876) );
oa12f01 g35085 ( .a(n38874), .b(n36198), .c(n36189), .o(n38877) );
na02f01 g35086 ( .a(n38877), .b(n38876), .o(n693) );
no02f01 g35087 ( .a(n21261), .b(n21004), .o(n38879) );
in01f01 g35088 ( .a(n38879), .o(n38880) );
ao12f01 g35089 ( .a(n20970), .b(n38880), .c(n20974), .o(n38881) );
no02f01 g35090 ( .a(n20953), .b(n20951), .o(n38882) );
no02f01 g35091 ( .a(n38882), .b(n38881), .o(n38883) );
in01f01 g35092 ( .a(n38883), .o(n38884) );
na02f01 g35093 ( .a(n38882), .b(n38881), .o(n38885) );
in01f01 g35094 ( .a(n29873), .o(n38886) );
no02f01 g35095 ( .a(n29874), .b(n29860), .o(n38887) );
oa12f01 g35096 ( .a(n38887), .b(n29858), .c(n29856), .o(n38888) );
no02f01 g35097 ( .a(n18393), .b(n29864), .o(n38889) );
no02f01 g35098 ( .a(n18450), .b(n18145), .o(n38890) );
no02f01 g35099 ( .a(n38890), .b(n18386), .o(n38891) );
in01f01 g35100 ( .a(n38891), .o(n38892) );
no03f01 g35101 ( .a(n38892), .b(n38889), .c(n29866), .o(n38893) );
no02f01 g35102 ( .a(n38889), .b(n29866), .o(n38894) );
no02f01 g35103 ( .a(n38891), .b(n38894), .o(n38895) );
no03f01 g35104 ( .a(n38895), .b(n38893), .c(n18459), .o(n38896) );
ao12f01 g35105 ( .a(n18452), .b(n18394), .c(n29865), .o(n38897) );
no02f01 g35106 ( .a(n18454), .b(n18145), .o(n38898) );
no02f01 g35107 ( .a(n38898), .b(n18412), .o(n38899) );
no02f01 g35108 ( .a(n38899), .b(n38897), .o(n38900) );
na02f01 g35109 ( .a(n38899), .b(n38897), .o(n38901) );
in01f01 g35110 ( .a(n38901), .o(n38902) );
no03f01 g35111 ( .a(n38902), .b(n38900), .c(n18459), .o(n38903) );
no02f01 g35112 ( .a(n38903), .b(n38896), .o(n38904) );
na03f01 g35113 ( .a(n38904), .b(n38888), .c(n38886), .o(n38905) );
no02f01 g35114 ( .a(n38895), .b(n38893), .o(n38906) );
no02f01 g35115 ( .a(n38906), .b(n18460), .o(n38907) );
in01f01 g35116 ( .a(n38900), .o(n38908) );
ao12f01 g35117 ( .a(n18460), .b(n38901), .c(n38908), .o(n38909) );
no02f01 g35118 ( .a(n38909), .b(n38907), .o(n38910) );
in01f01 g35119 ( .a(n38898), .o(n38911) );
ao12f01 g35120 ( .a(n18412), .b(n38897), .c(n38911), .o(n38912) );
no02f01 g35121 ( .a(n18453), .b(n18145), .o(n38913) );
no02f01 g35122 ( .a(n38913), .b(n18403), .o(n38914) );
in01f01 g35123 ( .a(n38914), .o(n38915) );
no02f01 g35124 ( .a(n38915), .b(n38912), .o(n38916) );
na02f01 g35125 ( .a(n38915), .b(n38912), .o(n38917) );
in01f01 g35126 ( .a(n38917), .o(n38918) );
no02f01 g35127 ( .a(n38918), .b(n38916), .o(n38919) );
in01f01 g35128 ( .a(n38919), .o(n38920) );
no02f01 g35129 ( .a(n38920), .b(n18459), .o(n38921) );
ao12f01 g35130 ( .a(n38921), .b(n38910), .c(n38905), .o(n38922) );
no02f01 g35131 ( .a(n38919), .b(n18460), .o(n38923) );
in01f01 g35132 ( .a(n18414), .o(n38924) );
no02f01 g35133 ( .a(n18457), .b(n38924), .o(n38925) );
in01f01 g35134 ( .a(n38925), .o(n38926) );
no02f01 g35135 ( .a(n18446), .b(n18145), .o(n38927) );
no02f01 g35136 ( .a(n38927), .b(n18430), .o(n38928) );
in01f01 g35137 ( .a(n38928), .o(n38929) );
no02f01 g35138 ( .a(n38929), .b(n38926), .o(n38930) );
no02f01 g35139 ( .a(n38928), .b(n38925), .o(n38931) );
no02f01 g35140 ( .a(n38931), .b(n38930), .o(n38932) );
no02f01 g35141 ( .a(n38932), .b(n18460), .o(n38933) );
no02f01 g35142 ( .a(n38933), .b(n38923), .o(n38934) );
in01f01 g35143 ( .a(n38934), .o(n38935) );
na02f01 g35144 ( .a(n38932), .b(n18460), .o(n38936) );
oa12f01 g35145 ( .a(n38936), .b(n38935), .c(n38922), .o(n38937) );
in01f01 g35146 ( .a(n38927), .o(n38938) );
ao12f01 g35147 ( .a(n18430), .b(n38925), .c(n38938), .o(n38939) );
no02f01 g35148 ( .a(n18445), .b(n18145), .o(n38940) );
no02f01 g35149 ( .a(n38940), .b(n18421), .o(n38941) );
in01f01 g35150 ( .a(n38941), .o(n38942) );
no02f01 g35151 ( .a(n38942), .b(n38939), .o(n38943) );
na02f01 g35152 ( .a(n38942), .b(n38939), .o(n38944) );
in01f01 g35153 ( .a(n38944), .o(n38945) );
no02f01 g35154 ( .a(n38945), .b(n38943), .o(n38946) );
in01f01 g35155 ( .a(n38946), .o(n38947) );
no02f01 g35156 ( .a(n38947), .b(n18459), .o(n38948) );
ao12f01 g35157 ( .a(n18447), .b(n38926), .c(n18431), .o(n38949) );
in01f01 g35158 ( .a(n38949), .o(n38950) );
no02f01 g35159 ( .a(n18444), .b(n18145), .o(n38951) );
no02f01 g35160 ( .a(n38951), .b(n18441), .o(n38952) );
in01f01 g35161 ( .a(n38952), .o(n38953) );
no02f01 g35162 ( .a(n38953), .b(n38950), .o(n38954) );
no02f01 g35163 ( .a(n38952), .b(n38949), .o(n38955) );
no03f01 g35164 ( .a(n38955), .b(n38954), .c(n18459), .o(n38956) );
no02f01 g35165 ( .a(n38956), .b(n38948), .o(n38957) );
in01f01 g35166 ( .a(n38957), .o(n38958) );
no02f01 g35167 ( .a(n38946), .b(n18460), .o(n38959) );
no02f01 g35168 ( .a(n38955), .b(n38954), .o(n38960) );
no02f01 g35169 ( .a(n38960), .b(n18460), .o(n38961) );
no02f01 g35170 ( .a(n38961), .b(n38959), .o(n38962) );
oa12f01 g35171 ( .a(n38962), .b(n38958), .c(n38937), .o(n911) );
in01f01 g35172 ( .a(n911), .o(n5799) );
na03f01 g35173 ( .a(n5799), .b(n38885), .c(n38884), .o(n38965) );
na02f01 g35174 ( .a(n38885), .b(n38884), .o(n5633) );
na02f01 g35175 ( .a(n911), .b(n5633), .o(n38967) );
na02f01 g35176 ( .a(n38967), .b(n38965), .o(n698) );
na03f01 g35177 ( .a(n38842), .b(n38840), .c(n38839), .o(n38969) );
oa12f01 g35178 ( .a(n38836), .b(n38837), .c(n38733), .o(n38970) );
na02f01 g35179 ( .a(n38970), .b(n38969), .o(n703) );
no02f01 g35180 ( .a(n9353), .b(n9352), .o(n38972) );
no02f01 g35181 ( .a(n9370), .b(n9224), .o(n38973) );
no02f01 g35182 ( .a(n9359), .b(n9225), .o(n38974) );
no02f01 g35183 ( .a(n38974), .b(n38973), .o(n38975) );
na02f01 g35184 ( .a(n38975), .b(n38972), .o(n38976) );
oa22f01 g35185 ( .a(n38974), .b(n38973), .c(n9353), .d(n9352), .o(n38977) );
na02f01 g35186 ( .a(n38977), .b(n38976), .o(n708) );
no02f01 g35187 ( .a(n35339), .b(n35271), .o(n38979) );
in01f01 g35188 ( .a(n38979), .o(n38980) );
no02f01 g35189 ( .a(n35360), .b(n38980), .o(n38981) );
in01f01 g35190 ( .a(n38981), .o(n38982) );
in01f01 g35191 ( .a(n35386), .o(n38983) );
no02f01 g35192 ( .a(n35368), .b(n4176), .o(n38984) );
no02f01 g35193 ( .a(n38984), .b(n35370), .o(n38985) );
na03f01 g35194 ( .a(n38985), .b(n38983), .c(n38982), .o(n38986) );
in01f01 g35195 ( .a(n38985), .o(n38987) );
oa12f01 g35196 ( .a(n38987), .b(n35386), .c(n38981), .o(n38988) );
na02f01 g35197 ( .a(n38988), .b(n38986), .o(n713) );
ao12f01 g35198 ( .a(n9591), .b(n9232), .c(n936), .o(n38990) );
ao12f01 g35199 ( .a(n4201), .b(n9231), .c(n936), .o(n38991) );
no02f01 g35200 ( .a(n38991), .b(n38990), .o(n38992) );
na03f01 g35201 ( .a(n38992), .b(n9590), .c(n9589), .o(n38993) );
in01f01 g35202 ( .a(n38992), .o(n732) );
oa12f01 g35203 ( .a(n732), .b(n9646), .c(n9645), .o(n38995) );
na02f01 g35204 ( .a(n38995), .b(n38993), .o(n718) );
na02f01 g35205 ( .a(n32732), .b(sin_out_6), .o(n38997) );
no03f01 g35206 ( .a(n34393), .b(n34369), .c(n34348), .o(n38998) );
no02f01 g35207 ( .a(n36577), .b(n34307), .o(n38999) );
no02f01 g35208 ( .a(n38999), .b(n36579), .o(n39000) );
in01f01 g35209 ( .a(n39000), .o(n39001) );
no03f01 g35210 ( .a(n39001), .b(n36593), .c(n38998), .o(n39002) );
no02f01 g35211 ( .a(n36593), .b(n38998), .o(n39003) );
no02f01 g35212 ( .a(n39000), .b(n39003), .o(n39004) );
oa12f01 g35213 ( .a(n32734), .b(n39004), .c(n39002), .o(n39005) );
na02f01 g35214 ( .a(n39005), .b(n38997), .o(n723) );
na02f01 g35215 ( .a(n8625), .b(n8604), .o(n39007) );
oa12f01 g35216 ( .a(n8670), .b(n8654), .c(n39007), .o(n39008) );
in01f01 g35217 ( .a(n39008), .o(n39009) );
no02f01 g35218 ( .a(n8673), .b(n5973), .o(n39010) );
no02f01 g35219 ( .a(n39010), .b(n8659), .o(n39011) );
na02f01 g35220 ( .a(n39011), .b(n39009), .o(n39012) );
in01f01 g35221 ( .a(n39011), .o(n39013) );
na02f01 g35222 ( .a(n39013), .b(n39008), .o(n39014) );
na02f01 g35223 ( .a(n39014), .b(n39012), .o(n727) );
no02f01 g35224 ( .a(n37142), .b(n37141), .o(n39016) );
oa12f01 g35225 ( .a(n25302), .b(n39016), .c(n25565), .o(n39017) );
oa12f01 g35226 ( .a(n25283), .b(n39017), .c(n25250), .o(n39018) );
in01f01 g35227 ( .a(n39018), .o(n39019) );
no02f01 g35228 ( .a(n25567), .b(n25230), .o(n39020) );
na02f01 g35229 ( .a(n39020), .b(n39019), .o(n39021) );
in01f01 g35230 ( .a(n39020), .o(n39022) );
na02f01 g35231 ( .a(n39022), .b(n39018), .o(n39023) );
na03f01 g35232 ( .a(n39023), .b(n39021), .c(n6037), .o(n39024) );
na02f01 g35233 ( .a(n39023), .b(n39021), .o(n5548) );
na02f01 g35234 ( .a(n5548), .b(n5873), .o(n39026) );
na02f01 g35235 ( .a(n39026), .b(n39024), .o(n737) );
in01f01 g35236 ( .a(n14213), .o(n39028) );
no02f01 g35237 ( .a(n39028), .b(n14006), .o(n39029) );
no02f01 g35238 ( .a(n14230), .b(n39029), .o(n39030) );
no02f01 g35239 ( .a(n39030), .b(n14226), .o(n39031) );
in01f01 g35240 ( .a(n39031), .o(n39032) );
no02f01 g35241 ( .a(n14229), .b(n13986), .o(n39033) );
no02f01 g35242 ( .a(n39033), .b(n39032), .o(n39034) );
na02f01 g35243 ( .a(n39033), .b(n39032), .o(n39035) );
in01f01 g35244 ( .a(n39035), .o(n39036) );
no02f01 g35245 ( .a(n39036), .b(n39034), .o(n39037) );
in01f01 g35246 ( .a(n39037), .o(n742) );
na03f01 g35247 ( .a(n9590), .b(n9589), .c(n9228), .o(n39039) );
oa12f01 g35248 ( .a(n936), .b(n9646), .c(n9645), .o(n39040) );
na02f01 g35249 ( .a(n39040), .b(n39039), .o(n747) );
na02f01 g35250 ( .a(n32732), .b(cos_out_12), .o(n39042) );
no02f01 g35251 ( .a(n36315), .b(n36269), .o(n39043) );
no02f01 g35252 ( .a(n36337), .b(n35944), .o(n39044) );
no02f01 g35253 ( .a(n39044), .b(n36339), .o(n39045) );
in01f01 g35254 ( .a(n39045), .o(n39046) );
no03f01 g35255 ( .a(n39046), .b(n36369), .c(n39043), .o(n39047) );
in01f01 g35256 ( .a(n39043), .o(n39048) );
ao12f01 g35257 ( .a(n39045), .b(n36368), .c(n39048), .o(n39049) );
oa12f01 g35258 ( .a(n32734), .b(n39049), .c(n39047), .o(n39050) );
na02f01 g35259 ( .a(n39050), .b(n39042), .o(n752) );
no02f01 g35260 ( .a(n38522), .b(n38520), .o(n39052) );
ao12f01 g35261 ( .a(n_22641), .b(n39052), .c(n38527), .o(n39053) );
no02f01 g35262 ( .a(n39053), .b(n38513), .o(n39054) );
na02f01 g35263 ( .a(n38521), .b(n38529), .o(n39055) );
oa12f01 g35264 ( .a(n6075), .b(n39055), .c(n38512), .o(n39056) );
na03f01 g35265 ( .a(n39056), .b(n38532), .c(n38528), .o(n39057) );
na02f01 g35266 ( .a(n39055), .b(n6075), .o(n39058) );
oa12f01 g35267 ( .a(n39057), .b(n39058), .c(n39054), .o(n39059) );
no02f01 g35268 ( .a(n31467), .b(n31471), .o(n39060) );
in01f01 g35269 ( .a(n39060), .o(n39061) );
ao12f01 g35270 ( .a(n39061), .b(n31219), .c(n31214), .o(n39062) );
no03f01 g35271 ( .a(n39060), .b(n31218), .c(n31459), .o(n39063) );
no02f01 g35272 ( .a(n39063), .b(n39062), .o(n39064) );
in01f01 g35273 ( .a(n39064), .o(n39065) );
ao12f01 g35274 ( .a(n39059), .b(n39065), .c(n31474), .o(n39066) );
ao12f01 g35275 ( .a(n31191), .b(n31457), .c(n31179), .o(n39067) );
no02f01 g35276 ( .a(n31218), .b(n31211), .o(n39068) );
in01f01 g35277 ( .a(n39068), .o(n39069) );
no02f01 g35278 ( .a(n39069), .b(n39067), .o(n39070) );
na02f01 g35279 ( .a(n39069), .b(n39067), .o(n39071) );
in01f01 g35280 ( .a(n39071), .o(n39072) );
no02f01 g35281 ( .a(n39072), .b(n39070), .o(n39073) );
in01f01 g35282 ( .a(n39073), .o(n39074) );
no02f01 g35283 ( .a(n39074), .b(n39059), .o(n39075) );
in01f01 g35284 ( .a(n38282), .o(n39076) );
in01f01 g35285 ( .a(n38296), .o(n39077) );
no03f01 g35286 ( .a(n38303), .b(n38301), .c(n38234), .o(n39078) );
ao12f01 g35287 ( .a(n38299), .b(n38297), .c(n38265), .o(n39079) );
in01f01 g35288 ( .a(n38307), .o(n39080) );
no03f01 g35289 ( .a(n39080), .b(n39079), .c(n39078), .o(n39081) );
oa12f01 g35290 ( .a(n39080), .b(n39079), .c(n39078), .o(n39082) );
no02f01 g35291 ( .a(n38311), .b(n38314), .o(n39083) );
no02f01 g35292 ( .a(n38312), .b(n38310), .o(n39084) );
in01f01 g35293 ( .a(n38322), .o(n39085) );
oa12f01 g35294 ( .a(n39085), .b(n39084), .c(n39083), .o(n39086) );
ao12f01 g35295 ( .a(n39081), .b(n39086), .c(n39082), .o(n39087) );
in01f01 g35296 ( .a(n38353), .o(n39088) );
ao12f01 g35297 ( .a(n38358), .b(n39088), .c(n38351), .o(n39089) );
no02f01 g35298 ( .a(n38365), .b(n38253), .o(n39090) );
no02f01 g35299 ( .a(n38362), .b(n38215), .o(n39091) );
in01f01 g35300 ( .a(n38370), .o(n39092) );
oa12f01 g35301 ( .a(n39092), .b(n39091), .c(n39090), .o(n39093) );
no03f01 g35302 ( .a(n38249), .b(n38248), .c(n6075), .o(n39094) );
no03f01 g35303 ( .a(n38249), .b(n38248), .c(n_22641), .o(n39095) );
no03f01 g35304 ( .a(n38377), .b(n39095), .c(n39094), .o(n39096) );
in01f01 g35305 ( .a(n38385), .o(n39097) );
na02f01 g35306 ( .a(n39097), .b(n39096), .o(n39098) );
no03f01 g35307 ( .a(n38250), .b(n32423), .c(n6075), .o(n39099) );
ao12f01 g35308 ( .a(n32050), .b(n32078), .c(n_22641), .o(n39100) );
no02f01 g35309 ( .a(n39100), .b(n39099), .o(n39101) );
no02f01 g35310 ( .a(n39097), .b(n39096), .o(n39102) );
oa12f01 g35311 ( .a(n39098), .b(n39102), .c(n39101), .o(n39103) );
na03f01 g35312 ( .a(n38394), .b(n38214), .c(n38251), .o(n39104) );
oa12f01 g35313 ( .a(n38213), .b(n38392), .c(n38252), .o(n39105) );
na03f01 g35314 ( .a(n38398), .b(n39105), .c(n39104), .o(n39106) );
ao12f01 g35315 ( .a(n38398), .b(n39105), .c(n39104), .o(n39107) );
ao12f01 g35316 ( .a(n39107), .b(n39106), .c(n39103), .o(n39108) );
no03f01 g35317 ( .a(n39092), .b(n39091), .c(n39090), .o(n39109) );
oa12f01 g35318 ( .a(n39093), .b(n39109), .c(n39108), .o(n39110) );
na03f01 g35319 ( .a(n38358), .b(n39088), .c(n38351), .o(n39111) );
ao12f01 g35320 ( .a(n39089), .b(n39111), .c(n39110), .o(n39112) );
ao12f01 g35321 ( .a(n38349), .b(n38407), .c(n39112), .o(n39113) );
oa12f01 g35322 ( .a(n38336), .b(n38332), .c(n38329), .o(n39114) );
na02f01 g35323 ( .a(n38432), .b(n39114), .o(n39115) );
ao12f01 g35324 ( .a(n39115), .b(n38426), .c(n39113), .o(n39116) );
no03f01 g35325 ( .a(n39085), .b(n39084), .c(n39083), .o(n39117) );
no04f01 g35326 ( .a(n39117), .b(n39116), .c(n38337), .d(n39081), .o(n39118) );
na03f01 g35327 ( .a(n38295), .b(n38292), .c(n38289), .o(n39119) );
oa12f01 g35328 ( .a(n39119), .b(n39118), .c(n39087), .o(n39120) );
oa12f01 g35329 ( .a(n38281), .b(n38274), .c(n38245), .o(n39121) );
na03f01 g35330 ( .a(n39121), .b(n39120), .c(n39077), .o(n39122) );
no02f01 g35331 ( .a(n38459), .b(n38458), .o(n39123) );
no02f01 g35332 ( .a(n38453), .b(n38450), .o(n39124) );
no02f01 g35333 ( .a(n39124), .b(n39123), .o(n39125) );
na02f01 g35334 ( .a(n38466), .b(n39125), .o(n39126) );
na03f01 g35335 ( .a(n39126), .b(n39122), .c(n39076), .o(n39127) );
no02f01 g35336 ( .a(n38504), .b(n38497), .o(n39128) );
no02f01 g35337 ( .a(n38466), .b(n39125), .o(n39129) );
no02f01 g35338 ( .a(n39129), .b(n39128), .o(n39130) );
na02f01 g35339 ( .a(n39130), .b(n39127), .o(n39131) );
no02f01 g35340 ( .a(n38541), .b(n38509), .o(n39132) );
oa12f01 g35341 ( .a(n38540), .b(n38539), .c(n38538), .o(n39133) );
ao12f01 g35342 ( .a(n39058), .b(n39056), .c(n38528), .o(n39134) );
ao12f01 g35343 ( .a(n39134), .b(n39054), .c(n38532), .o(n39135) );
oa12f01 g35344 ( .a(n39133), .b(n39073), .c(n39135), .o(n39136) );
ao12f01 g35345 ( .a(n39136), .b(n39132), .c(n39131), .o(n39137) );
no02f01 g35346 ( .a(n39059), .b(n32252), .o(n39138) );
no02f01 g35347 ( .a(n39059), .b(n31463), .o(n39139) );
no02f01 g35348 ( .a(n39139), .b(n39138), .o(n39140) );
in01f01 g35349 ( .a(n39140), .o(n39141) );
no04f01 g35350 ( .a(n39141), .b(n39137), .c(n39075), .d(n39066), .o(n39142) );
in01f01 g35351 ( .a(n31515), .o(n39143) );
no02f01 g35352 ( .a(n39059), .b(n39143), .o(n39144) );
no02f01 g35353 ( .a(n39059), .b(n32251), .o(n39145) );
no02f01 g35354 ( .a(n39145), .b(n39144), .o(n39146) );
in01f01 g35355 ( .a(n31502), .o(n39147) );
no02f01 g35356 ( .a(n39059), .b(n39147), .o(n39148) );
no02f01 g35357 ( .a(n39059), .b(n31518), .o(n39149) );
no02f01 g35358 ( .a(n39149), .b(n39148), .o(n39150) );
na02f01 g35359 ( .a(n39150), .b(n39146), .o(n39151) );
in01f01 g35360 ( .a(n39151), .o(n39152) );
na02f01 g35361 ( .a(n39152), .b(n39142), .o(n39153) );
ao12f01 g35362 ( .a(n39135), .b(n39064), .c(n32243), .o(n39154) );
ao12f01 g35363 ( .a(n39135), .b(n31485), .c(n32240), .o(n39155) );
no02f01 g35364 ( .a(n39155), .b(n39154), .o(n39156) );
ao12f01 g35365 ( .a(n39135), .b(n31515), .c(n31401), .o(n39157) );
in01f01 g35366 ( .a(n39157), .o(n39158) );
oa12f01 g35367 ( .a(n39059), .b(n39147), .c(n31518), .o(n39159) );
na03f01 g35368 ( .a(n39159), .b(n39158), .c(n39156), .o(n39160) );
in01f01 g35369 ( .a(n39160), .o(n39161) );
no02f01 g35370 ( .a(n39135), .b(n31511), .o(n39162) );
no02f01 g35371 ( .a(n39059), .b(n31519), .o(n39163) );
no02f01 g35372 ( .a(n39163), .b(n39162), .o(n39164) );
na03f01 g35373 ( .a(n39164), .b(n39161), .c(n39153), .o(n39165) );
in01f01 g35374 ( .a(n39066), .o(n39166) );
in01f01 g35375 ( .a(n39075), .o(n39167) );
na03f01 g35376 ( .a(n38536), .b(n38533), .c(n38526), .o(n39168) );
na02f01 g35377 ( .a(n39168), .b(n38508), .o(n39169) );
ao12f01 g35378 ( .a(n38537), .b(n39074), .c(n39059), .o(n39170) );
oa12f01 g35379 ( .a(n39170), .b(n39169), .c(n38507), .o(n39171) );
na04f01 g35380 ( .a(n39140), .b(n39171), .c(n39167), .d(n39166), .o(n39172) );
no02f01 g35381 ( .a(n39151), .b(n39172), .o(n39173) );
in01f01 g35382 ( .a(n39164), .o(n39174) );
oa12f01 g35383 ( .a(n39174), .b(n39160), .c(n39173), .o(n39175) );
na02f01 g35384 ( .a(n39175), .b(n39165), .o(n756) );
no02f01 g35385 ( .a(n38010), .b(n26336), .o(n39177) );
no02f01 g35386 ( .a(n37871), .b(n26327), .o(n39178) );
no02f01 g35387 ( .a(n39178), .b(n39177), .o(n39179) );
no02f01 g35388 ( .a(n38010), .b(n26332), .o(n39180) );
in01f01 g35389 ( .a(n39180), .o(n39181) );
no02f01 g35390 ( .a(n37871), .b(n26874), .o(n39182) );
ao12f01 g35391 ( .a(n39182), .b(n39181), .c(n38007), .o(n39183) );
na02f01 g35392 ( .a(n39183), .b(n39179), .o(n39184) );
in01f01 g35393 ( .a(n39179), .o(n39185) );
in01f01 g35394 ( .a(n39183), .o(n39186) );
na02f01 g35395 ( .a(n39186), .b(n39185), .o(n39187) );
na02f01 g35396 ( .a(n39187), .b(n39184), .o(n761) );
no02f01 g35397 ( .a(n38492), .b(n31606), .o(n39189) );
no02f01 g35398 ( .a(n38484), .b(n31607), .o(n39190) );
no02f01 g35399 ( .a(n39190), .b(n39189), .o(n39191) );
ao12f01 g35400 ( .a(n31607), .b(n36838), .c(n36827), .o(n39192) );
in01f01 g35401 ( .a(n39192), .o(n39193) );
no02f01 g35402 ( .a(n36838), .b(n36827), .o(n39194) );
no02f01 g35403 ( .a(n39194), .b(n31606), .o(n39195) );
in01f01 g35404 ( .a(n39195), .o(n39196) );
oa12f01 g35405 ( .a(n39196), .b(n36885), .c(n36891), .o(n39197) );
na03f01 g35406 ( .a(n39197), .b(n39193), .c(n39191), .o(n39198) );
in01f01 g35407 ( .a(n39191), .o(n39199) );
ao12f01 g35408 ( .a(n39195), .b(n36886), .c(n36876), .o(n39200) );
oa12f01 g35409 ( .a(n39199), .b(n39200), .c(n39192), .o(n39201) );
na03f01 g35410 ( .a(n39201), .b(n39198), .c(n3633), .o(n39202) );
no03f01 g35411 ( .a(n39200), .b(n39192), .c(n39199), .o(n39203) );
ao12f01 g35412 ( .a(n39191), .b(n39197), .c(n39193), .o(n39204) );
oa12f01 g35413 ( .a(n6203), .b(n39204), .c(n39203), .o(n39205) );
na02f01 g35414 ( .a(n39205), .b(n39202), .o(n770) );
no02f01 g35415 ( .a(n20872), .b(n20869), .o(n39207) );
in01f01 g35416 ( .a(n39207), .o(n39208) );
no02f01 g35417 ( .a(n21333), .b(n21006), .o(n39209) );
no02f01 g35418 ( .a(n39209), .b(n20931), .o(n39210) );
ao12f01 g35419 ( .a(n20921), .b(n39210), .c(n21318), .o(n39211) );
ao12f01 g35420 ( .a(n20930), .b(n39211), .c(n21312), .o(n39212) );
na02f01 g35421 ( .a(n39212), .b(n39208), .o(n39213) );
na02f01 g35422 ( .a(n21262), .b(n21007), .o(n39214) );
na03f01 g35423 ( .a(n39214), .b(n21328), .c(n21318), .o(n39215) );
na02f01 g35424 ( .a(n39215), .b(n21325), .o(n39216) );
oa12f01 g35425 ( .a(n20888), .b(n39216), .c(n20887), .o(n39217) );
na02f01 g35426 ( .a(n39217), .b(n39207), .o(n39218) );
na02f01 g35427 ( .a(n39218), .b(n39213), .o(n775) );
na03f01 g35428 ( .a(n36750), .b(n36747), .c(n36746), .o(n39220) );
oa12f01 g35429 ( .a(n36742), .b(n36744), .c(n36696), .o(n39221) );
ao12f01 g35430 ( .a(n_27014), .b(n39221), .c(n39220), .o(n39222) );
no03f01 g35431 ( .a(n36751), .b(n36745), .c(n27681), .o(n39223) );
no02f01 g35432 ( .a(n39223), .b(n39222), .o(n39224) );
ao12f01 g35433 ( .a(n27681), .b(n29661), .c(n29658), .o(n39225) );
no02f01 g35434 ( .a(n29649), .b(n27681), .o(n39226) );
oa12f01 g35435 ( .a(n36757), .b(n36698), .c(n36694), .o(n39227) );
na03f01 g35436 ( .a(n36755), .b(n36748), .c(n36714), .o(n39228) );
ao12f01 g35437 ( .a(n27681), .b(n39228), .c(n39227), .o(n39229) );
no03f01 g35438 ( .a(n39229), .b(n39226), .c(n39225), .o(n39230) );
no02f01 g35439 ( .a(n39230), .b(n27681), .o(n39231) );
ao12f01 g35440 ( .a(n_27014), .b(n39228), .c(n39227), .o(n39232) );
no02f01 g35441 ( .a(n39232), .b(n39230), .o(n39233) );
oa22f01 g35442 ( .a(n39233), .b(n_27014), .c(n39231), .d(n39224), .o(n39234) );
na02f01 g35443 ( .a(n36776), .b(n_27014), .o(n39235) );
na02f01 g35444 ( .a(n36771), .b(n_27014), .o(n39236) );
na02f01 g35445 ( .a(n36736), .b(n_27014), .o(n39237) );
na04f01 g35446 ( .a(n39237), .b(n39236), .c(n39235), .d(n39234), .o(n39238) );
no02f01 g35447 ( .a(n36726), .b(n_27014), .o(n39239) );
no02f01 g35448 ( .a(n36722), .b(n27681), .o(n39240) );
no02f01 g35449 ( .a(n36789), .b(n_27014), .o(n39241) );
no03f01 g35450 ( .a(n39241), .b(n39240), .c(n39239), .o(n39242) );
ao12f01 g35451 ( .a(n_27014), .b(n39242), .c(n39238), .o(n39243) );
in01f01 g35452 ( .a(n39243), .o(n39244) );
oa12f01 g35453 ( .a(n27681), .b(n36751), .c(n36745), .o(n39245) );
na03f01 g35454 ( .a(n39221), .b(n39220), .c(n_27014), .o(n39246) );
na02f01 g35455 ( .a(n39246), .b(n39245), .o(n39247) );
oa12f01 g35456 ( .a(n_27014), .b(n29665), .c(n29664), .o(n39248) );
na02f01 g35457 ( .a(n29635), .b(n_27014), .o(n39249) );
oa12f01 g35458 ( .a(n_27014), .b(n36758), .c(n36756), .o(n39250) );
na03f01 g35459 ( .a(n39250), .b(n39249), .c(n39248), .o(n39251) );
na02f01 g35460 ( .a(n39251), .b(n_27014), .o(n39252) );
oa12f01 g35461 ( .a(n27681), .b(n36758), .c(n36756), .o(n39253) );
na02f01 g35462 ( .a(n39253), .b(n39251), .o(n39254) );
ao22f01 g35463 ( .a(n39254), .b(n27681), .c(n39252), .d(n39247), .o(n39255) );
in01f01 g35464 ( .a(n36775), .o(n39256) );
no02f01 g35465 ( .a(n39256), .b(n36773), .o(n39257) );
no02f01 g35466 ( .a(n39257), .b(n27681), .o(n39258) );
in01f01 g35467 ( .a(n36770), .o(n39259) );
no02f01 g35468 ( .a(n39259), .b(n36768), .o(n39260) );
no02f01 g35469 ( .a(n39260), .b(n27681), .o(n39261) );
no02f01 g35470 ( .a(n36789), .b(n27681), .o(n39262) );
no04f01 g35471 ( .a(n39262), .b(n39261), .c(n39258), .d(n39255), .o(n39263) );
na02f01 g35472 ( .a(n36722), .b(n27681), .o(n39264) );
na02f01 g35473 ( .a(n36726), .b(n_27014), .o(n39265) );
na02f01 g35474 ( .a(n39265), .b(n39264), .o(n39266) );
ao12f01 g35475 ( .a(n_27014), .b(n39257), .c(n39260), .o(n39267) );
ao12f01 g35476 ( .a(n39267), .b(n39266), .c(n39263), .o(n39268) );
no02f01 g35477 ( .a(n36710), .b(n36688), .o(n39269) );
ao12f01 g35478 ( .a(n29460), .b(n28064), .c(n28461), .o(n39270) );
no02f01 g35479 ( .a(n39270), .b(n36691), .o(n39271) );
in01f01 g35480 ( .a(n39271), .o(n39272) );
ao12f01 g35481 ( .a(n39272), .b(n39269), .c(n36707), .o(n39273) );
no02f01 g35482 ( .a(n29491), .b(n28436), .o(n39274) );
no02f01 g35483 ( .a(n29460), .b(n28071), .o(n39275) );
no02f01 g35484 ( .a(n39275), .b(n39274), .o(n39276) );
no02f01 g35485 ( .a(n39276), .b(n39273), .o(n39277) );
na02f01 g35486 ( .a(n39276), .b(n39273), .o(n39278) );
in01f01 g35487 ( .a(n39278), .o(n39279) );
no02f01 g35488 ( .a(n39279), .b(n39277), .o(n39280) );
no02f01 g35489 ( .a(n39280), .b(n27681), .o(n39281) );
ao12f01 g35490 ( .a(n39281), .b(n39268), .c(n39244), .o(n39282) );
no02f01 g35491 ( .a(n39274), .b(n39273), .o(n39283) );
no02f01 g35492 ( .a(n39283), .b(n39275), .o(n39284) );
in01f01 g35493 ( .a(n39284), .o(n39285) );
no02f01 g35494 ( .a(n29491), .b(n28091), .o(n39286) );
no02f01 g35495 ( .a(n29460), .b(n28092), .o(n39287) );
no02f01 g35496 ( .a(n39287), .b(n39286), .o(n39288) );
in01f01 g35497 ( .a(n39288), .o(n39289) );
no02f01 g35498 ( .a(n39289), .b(n39285), .o(n39290) );
no02f01 g35499 ( .a(n39288), .b(n39284), .o(n39291) );
no02f01 g35500 ( .a(n39291), .b(n39290), .o(n39292) );
no02f01 g35501 ( .a(n39292), .b(n27681), .o(n39293) );
in01f01 g35502 ( .a(n39293), .o(n39294) );
na02f01 g35503 ( .a(n39294), .b(n39282), .o(n39295) );
ao12f01 g35504 ( .a(n_27014), .b(n39292), .c(n39280), .o(n39296) );
in01f01 g35505 ( .a(n39296), .o(n39297) );
na02f01 g35506 ( .a(n39297), .b(n39295), .o(n39298) );
no03f01 g35507 ( .a(n39286), .b(n39274), .c(n39273), .o(n39299) );
no03f01 g35508 ( .a(n39299), .b(n39287), .c(n39275), .o(n39300) );
no02f01 g35509 ( .a(n29491), .b(n28414), .o(n39301) );
no02f01 g35510 ( .a(n29460), .b(n28081), .o(n39302) );
no02f01 g35511 ( .a(n39302), .b(n39301), .o(n39303) );
no02f01 g35512 ( .a(n39303), .b(n39300), .o(n39304) );
na02f01 g35513 ( .a(n39303), .b(n39300), .o(n39305) );
in01f01 g35514 ( .a(n39305), .o(n39306) );
no02f01 g35515 ( .a(n39306), .b(n39304), .o(n39307) );
no02f01 g35516 ( .a(n39307), .b(n27681), .o(n39308) );
no02f01 g35517 ( .a(n39307), .b(n_27014), .o(n39309) );
no02f01 g35518 ( .a(n39309), .b(n39308), .o(n39310) );
in01f01 g35519 ( .a(n39310), .o(n39311) );
na02f01 g35520 ( .a(n39311), .b(n39298), .o(n39312) );
in01f01 g35521 ( .a(n39268), .o(n39313) );
in01f01 g35522 ( .a(n39281), .o(n39314) );
oa12f01 g35523 ( .a(n39314), .b(n39313), .c(n39243), .o(n39315) );
no02f01 g35524 ( .a(n39293), .b(n39315), .o(n39316) );
no02f01 g35525 ( .a(n39296), .b(n39316), .o(n39317) );
na02f01 g35526 ( .a(n39310), .b(n39317), .o(n39318) );
no02f01 g35527 ( .a(n28585), .b(n28871), .o(n39319) );
no02f01 g35528 ( .a(n28604), .b(n28598), .o(n39320) );
in01f01 g35529 ( .a(n39320), .o(n39321) );
no02f01 g35530 ( .a(n39321), .b(n39319), .o(n39322) );
na02f01 g35531 ( .a(n39321), .b(n39319), .o(n39323) );
in01f01 g35532 ( .a(n39323), .o(n39324) );
no02f01 g35533 ( .a(n39324), .b(n39322), .o(n39325) );
ao12f01 g35534 ( .a(n39325), .b(n39318), .c(n39312), .o(n39326) );
in01f01 g35535 ( .a(n39326), .o(n39327) );
na03f01 g35536 ( .a(n39325), .b(n39318), .c(n39312), .o(n39328) );
no02f01 g35537 ( .a(n39280), .b(n_27014), .o(n39329) );
in01f01 g35538 ( .a(n39329), .o(n39330) );
no02f01 g35539 ( .a(n39292), .b(n_27014), .o(n39331) );
no02f01 g35540 ( .a(n39331), .b(n39293), .o(n39332) );
na03f01 g35541 ( .a(n39332), .b(n39330), .c(n39315), .o(n39333) );
in01f01 g35542 ( .a(n39332), .o(n39334) );
oa12f01 g35543 ( .a(n39334), .b(n39329), .c(n39282), .o(n39335) );
ao22f01 g35544 ( .a(n28586), .b(n28446), .c(n28583), .d(n28460), .o(n39336) );
ao12f01 g35545 ( .a(n39336), .b(n28586), .c(n28871), .o(n39337) );
ao12f01 g35546 ( .a(n39337), .b(n39335), .c(n39333), .o(n39338) );
no03f01 g35547 ( .a(n39334), .b(n39329), .c(n39282), .o(n39339) );
ao12f01 g35548 ( .a(n39332), .b(n39330), .c(n39315), .o(n39340) );
in01f01 g35549 ( .a(n39337), .o(n39341) );
no03f01 g35550 ( .a(n39341), .b(n39340), .c(n39339), .o(n39342) );
no02f01 g35551 ( .a(n39329), .b(n39281), .o(n39343) );
na03f01 g35552 ( .a(n39343), .b(n39268), .c(n39244), .o(n39344) );
in01f01 g35553 ( .a(n39343), .o(n39345) );
oa12f01 g35554 ( .a(n39345), .b(n39313), .c(n39243), .o(n39346) );
no02f01 g35555 ( .a(n28865), .b(n28475), .o(n39347) );
no02f01 g35556 ( .a(n28869), .b(n28459), .o(n39348) );
in01f01 g35557 ( .a(n39348), .o(n39349) );
no02f01 g35558 ( .a(n39349), .b(n39347), .o(n39350) );
na02f01 g35559 ( .a(n39349), .b(n39347), .o(n39351) );
in01f01 g35560 ( .a(n39351), .o(n39352) );
no02f01 g35561 ( .a(n39352), .b(n39350), .o(n39353) );
ao12f01 g35562 ( .a(n39353), .b(n39346), .c(n39344), .o(n39354) );
in01f01 g35563 ( .a(n39354), .o(n39355) );
no02f01 g35564 ( .a(n39267), .b(n39241), .o(n39356) );
no02f01 g35565 ( .a(n36726), .b(n27681), .o(n39357) );
no02f01 g35566 ( .a(n36726), .b(n_27014), .o(n39358) );
no02f01 g35567 ( .a(n39358), .b(n39357), .o(n39359) );
ao12f01 g35568 ( .a(n39359), .b(n39356), .c(n39238), .o(n39360) );
in01f01 g35569 ( .a(n39241), .o(n39361) );
oa12f01 g35570 ( .a(n27681), .b(n36776), .c(n36771), .o(n39362) );
na02f01 g35571 ( .a(n39362), .b(n39361), .o(n39363) );
na02f01 g35572 ( .a(n36722), .b(n_27014), .o(n39364) );
na02f01 g35573 ( .a(n36722), .b(n27681), .o(n39365) );
na02f01 g35574 ( .a(n39365), .b(n39364), .o(n39366) );
no03f01 g35575 ( .a(n39366), .b(n39363), .c(n39263), .o(n39367) );
no04f01 g35576 ( .a(n28864), .b(n28862), .c(n28487), .d(n28475), .o(n39368) );
ao22f01 g35577 ( .a(n28580), .b(n28476), .c(n28579), .d(n28488), .o(n39369) );
no02f01 g35578 ( .a(n39369), .b(n39368), .o(n39370) );
in01f01 g35579 ( .a(n39370), .o(n39371) );
no03f01 g35580 ( .a(n39371), .b(n39367), .c(n39360), .o(n39372) );
in01f01 g35581 ( .a(n39372), .o(n39373) );
na02f01 g35582 ( .a(n39235), .b(n39234), .o(n39374) );
no02f01 g35583 ( .a(n39260), .b(n_27014), .o(n39375) );
no02f01 g35584 ( .a(n39375), .b(n39261), .o(n39376) );
na02f01 g35585 ( .a(n36776), .b(n27681), .o(n39377) );
na03f01 g35586 ( .a(n39377), .b(n39376), .c(n39374), .o(n39378) );
no02f01 g35587 ( .a(n39258), .b(n39255), .o(n39379) );
na02f01 g35588 ( .a(n36771), .b(n27681), .o(n39380) );
na02f01 g35589 ( .a(n39380), .b(n39236), .o(n39381) );
no02f01 g35590 ( .a(n39257), .b(n_27014), .o(n39382) );
oa12f01 g35591 ( .a(n39381), .b(n39382), .c(n39379), .o(n39383) );
ao22f01 g35592 ( .a(n28577), .b(n28574), .c(n28562), .d(n28512), .o(n39384) );
ao12f01 g35593 ( .a(n39384), .b(n28577), .c(n28858), .o(n39385) );
ao12f01 g35594 ( .a(n39385), .b(n39383), .c(n39378), .o(n39386) );
na02f01 g35595 ( .a(n39377), .b(n39235), .o(n39387) );
no02f01 g35596 ( .a(n39387), .b(n39234), .o(n39388) );
no02f01 g35597 ( .a(n39382), .b(n39258), .o(n39389) );
no02f01 g35598 ( .a(n39389), .b(n39255), .o(n39390) );
no02f01 g35599 ( .a(n28558), .b(n28522), .o(n39391) );
no02f01 g35600 ( .a(n28560), .b(n28511), .o(n39392) );
no02f01 g35601 ( .a(n39392), .b(n39391), .o(n39393) );
na02f01 g35602 ( .a(n39392), .b(n39391), .o(n39394) );
in01f01 g35603 ( .a(n39394), .o(n39395) );
no02f01 g35604 ( .a(n39395), .b(n39393), .o(n39396) );
in01f01 g35605 ( .a(n39396), .o(n39397) );
oa12f01 g35606 ( .a(n39397), .b(n39390), .c(n39388), .o(n39398) );
no03f01 g35607 ( .a(n39397), .b(n39390), .c(n39388), .o(n39399) );
oa12f01 g35608 ( .a(n_27014), .b(n36751), .c(n36745), .o(n39400) );
oa12f01 g35609 ( .a(n27681), .b(n36751), .c(n36745), .o(n39401) );
na04f01 g35610 ( .a(n39401), .b(n39400), .c(n39253), .d(n39251), .o(n39402) );
na02f01 g35611 ( .a(n39401), .b(n39400), .o(n39403) );
na02f01 g35612 ( .a(n39403), .b(n39254), .o(n39404) );
no02f01 g35613 ( .a(n28850), .b(n28842), .o(n39405) );
no02f01 g35614 ( .a(n28557), .b(n28522), .o(n39406) );
no02f01 g35615 ( .a(n39406), .b(n39405), .o(n39407) );
na02f01 g35616 ( .a(n39406), .b(n39405), .o(n39408) );
in01f01 g35617 ( .a(n39408), .o(n39409) );
no02f01 g35618 ( .a(n39409), .b(n39407), .o(n39410) );
ao12f01 g35619 ( .a(n39410), .b(n39404), .c(n39402), .o(n39411) );
na03f01 g35620 ( .a(n39410), .b(n39404), .c(n39402), .o(n39412) );
na02f01 g35621 ( .a(n39249), .b(n39248), .o(n39413) );
no02f01 g35622 ( .a(n39232), .b(n39229), .o(n39414) );
no02f01 g35623 ( .a(n39414), .b(n39413), .o(n39415) );
no02f01 g35624 ( .a(n39226), .b(n39225), .o(n39416) );
na02f01 g35625 ( .a(n39253), .b(n39250), .o(n39417) );
no02f01 g35626 ( .a(n39417), .b(n39416), .o(n39418) );
no02f01 g35627 ( .a(n28552), .b(n28549), .o(n39419) );
no02f01 g35628 ( .a(n28532), .b(n28525), .o(n39420) );
no02f01 g35629 ( .a(n39420), .b(n28842), .o(n39421) );
no02f01 g35630 ( .a(n39421), .b(n39419), .o(n39422) );
na02f01 g35631 ( .a(n39421), .b(n39419), .o(n39423) );
in01f01 g35632 ( .a(n39423), .o(n39424) );
no02f01 g35633 ( .a(n39424), .b(n39422), .o(n39425) );
in01f01 g35634 ( .a(n39425), .o(n39426) );
oa12f01 g35635 ( .a(n39426), .b(n39418), .c(n39415), .o(n39427) );
no03f01 g35636 ( .a(n39426), .b(n39418), .c(n39415), .o(n39428) );
no03f01 g35637 ( .a(n28848), .b(n28847), .c(n28846), .o(n39429) );
ao12f01 g35638 ( .a(n28548), .b(n28551), .c(n28550), .o(n39430) );
no03f01 g35639 ( .a(n39430), .b(n39429), .c(n28845), .o(n39431) );
no02f01 g35640 ( .a(n39430), .b(n39429), .o(n39432) );
no02f01 g35641 ( .a(n39432), .b(n28540), .o(n39433) );
no02f01 g35642 ( .a(n39433), .b(n39431), .o(n39434) );
na03f01 g35643 ( .a(n29634), .b(n29627), .c(n_27014), .o(n39435) );
na03f01 g35644 ( .a(n29634), .b(n29627), .c(n27681), .o(n39436) );
no02f01 g35645 ( .a(n28538), .b(n28534), .o(n39437) );
no02f01 g35646 ( .a(n28539), .b(n28844), .o(n39438) );
no02f01 g35647 ( .a(n39438), .b(n39437), .o(n39439) );
in01f01 g35648 ( .a(n39439), .o(n39440) );
na03f01 g35649 ( .a(n39440), .b(n39436), .c(n39435), .o(n39441) );
no02f01 g35650 ( .a(n39441), .b(n39434), .o(n39442) );
na02f01 g35651 ( .a(n39441), .b(n39434), .o(n39443) );
oa12f01 g35652 ( .a(n29662), .b(n29649), .c(n27681), .o(n39444) );
na03f01 g35653 ( .a(n29666), .b(n29635), .c(n_27014), .o(n39445) );
na02f01 g35654 ( .a(n39445), .b(n39444), .o(n39446) );
ao12f01 g35655 ( .a(n39442), .b(n39446), .c(n39443), .o(n39447) );
oa12f01 g35656 ( .a(n39427), .b(n39447), .c(n39428), .o(n39448) );
ao12f01 g35657 ( .a(n39411), .b(n39448), .c(n39412), .o(n39449) );
oa12f01 g35658 ( .a(n39398), .b(n39449), .c(n39399), .o(n39450) );
na03f01 g35659 ( .a(n39385), .b(n39383), .c(n39378), .o(n39451) );
oa12f01 g35660 ( .a(n39451), .b(n39450), .c(n39386), .o(n39452) );
na03f01 g35661 ( .a(n39236), .b(n39235), .c(n39234), .o(n39453) );
no02f01 g35662 ( .a(n39241), .b(n39262), .o(n39454) );
na03f01 g35663 ( .a(n39454), .b(n39362), .c(n39453), .o(n39455) );
in01f01 g35664 ( .a(n39455), .o(n39456) );
ao12f01 g35665 ( .a(n39454), .b(n39362), .c(n39453), .o(n39457) );
no02f01 g35666 ( .a(n28576), .b(n28858), .o(n39458) );
in01f01 g35667 ( .a(n39458), .o(n39459) );
no02f01 g35668 ( .a(n28861), .b(n28487), .o(n39460) );
no02f01 g35669 ( .a(n39460), .b(n39459), .o(n39461) );
na02f01 g35670 ( .a(n39460), .b(n39459), .o(n39462) );
in01f01 g35671 ( .a(n39462), .o(n39463) );
no02f01 g35672 ( .a(n39463), .b(n39461), .o(n39464) );
in01f01 g35673 ( .a(n39464), .o(n39465) );
no03f01 g35674 ( .a(n39465), .b(n39457), .c(n39456), .o(n39466) );
oa12f01 g35675 ( .a(n39366), .b(n39363), .c(n39263), .o(n39467) );
na03f01 g35676 ( .a(n39359), .b(n39356), .c(n39238), .o(n39468) );
ao12f01 g35677 ( .a(n39370), .b(n39468), .c(n39467), .o(n39469) );
no03f01 g35678 ( .a(n39261), .b(n39258), .c(n39255), .o(n39470) );
in01f01 g35679 ( .a(n39454), .o(n39471) );
oa12f01 g35680 ( .a(n39471), .b(n39267), .c(n39470), .o(n39472) );
ao12f01 g35681 ( .a(n39464), .b(n39472), .c(n39455), .o(n39473) );
no02f01 g35682 ( .a(n39473), .b(n39469), .o(n39474) );
oa12f01 g35683 ( .a(n39474), .b(n39466), .c(n39452), .o(n39475) );
na03f01 g35684 ( .a(n39353), .b(n39346), .c(n39344), .o(n39476) );
na03f01 g35685 ( .a(n39476), .b(n39475), .c(n39373), .o(n39477) );
ao12f01 g35686 ( .a(n39342), .b(n39477), .c(n39355), .o(n39478) );
no02f01 g35687 ( .a(n39478), .b(n39338), .o(n39479) );
na03f01 g35688 ( .a(n39479), .b(n39328), .c(n39327), .o(n39480) );
no02f01 g35689 ( .a(n39310), .b(n39317), .o(n39481) );
no02f01 g35690 ( .a(n39311), .b(n39298), .o(n39482) );
in01f01 g35691 ( .a(n39325), .o(n39483) );
no03f01 g35692 ( .a(n39483), .b(n39482), .c(n39481), .o(n39484) );
oa22f01 g35693 ( .a(n39478), .b(n39338), .c(n39484), .d(n39326), .o(n39485) );
na02f01 g35694 ( .a(n39485), .b(n39480), .o(n780) );
na02f01 g35695 ( .a(n14247), .b(n13890), .o(n39487) );
no02f01 g35696 ( .a(n39487), .b(n14242), .o(n39488) );
na02f01 g35697 ( .a(n39487), .b(n14242), .o(n39489) );
in01f01 g35698 ( .a(n39489), .o(n39490) );
no02f01 g35699 ( .a(n39490), .b(n39488), .o(n39491) );
in01f01 g35700 ( .a(n39491), .o(n785) );
na02f01 g35701 ( .a(n32732), .b(sin_out_12), .o(n39493) );
no03f01 g35702 ( .a(n38628), .b(n38607), .c(n38597), .o(n39494) );
in01f01 g35703 ( .a(n39494), .o(n39495) );
no02f01 g35704 ( .a(n39495), .b(n38595), .o(n39496) );
ao12f01 g35705 ( .a(n34307), .b(n38625), .c(n38605), .o(n39497) );
no02f01 g35706 ( .a(n39497), .b(n38609), .o(n39498) );
in01f01 g35707 ( .a(n39498), .o(n39499) );
no02f01 g35708 ( .a(n35676), .b(n35672), .o(n39500) );
in01f01 g35709 ( .a(n39500), .o(n39501) );
no02f01 g35710 ( .a(n35702), .b(n34287), .o(n39502) );
na02f01 g35711 ( .a(n35702), .b(n34287), .o(n39503) );
in01f01 g35712 ( .a(n39503), .o(n39504) );
no02f01 g35713 ( .a(n39504), .b(n39502), .o(n39505) );
in01f01 g35714 ( .a(n39505), .o(n39506) );
no02f01 g35715 ( .a(n39506), .b(n39501), .o(n39507) );
no02f01 g35716 ( .a(n39505), .b(n39500), .o(n39508) );
no02f01 g35717 ( .a(n39508), .b(n39507), .o(n39509) );
in01f01 g35718 ( .a(n39509), .o(n39510) );
no02f01 g35719 ( .a(n39510), .b(n34267), .o(n39511) );
no02f01 g35720 ( .a(n39509), .b(n34307), .o(n39512) );
no02f01 g35721 ( .a(n39512), .b(n39511), .o(n39513) );
in01f01 g35722 ( .a(n39513), .o(n39514) );
no03f01 g35723 ( .a(n39514), .b(n39499), .c(n39496), .o(n39515) );
in01f01 g35724 ( .a(n39496), .o(n39516) );
ao12f01 g35725 ( .a(n39513), .b(n39498), .c(n39516), .o(n39517) );
oa12f01 g35726 ( .a(n32734), .b(n39517), .c(n39515), .o(n39518) );
na02f01 g35727 ( .a(n39518), .b(n39493), .o(n790) );
in01f01 g35728 ( .a(n32086), .o(n39520) );
no02f01 g35729 ( .a(n32418), .b(n32139), .o(n39521) );
na02f01 g35730 ( .a(n32492), .b(n39521), .o(n39522) );
na02f01 g35731 ( .a(n32423), .b(n31606), .o(n39523) );
in01f01 g35732 ( .a(n39523), .o(n39524) );
no02f01 g35733 ( .a(n32424), .b(n39524), .o(n39525) );
na03f01 g35734 ( .a(n39525), .b(n39522), .c(n39520), .o(n39526) );
in01f01 g35735 ( .a(n39522), .o(n39527) );
in01f01 g35736 ( .a(n39525), .o(n39528) );
oa12f01 g35737 ( .a(n39528), .b(n39527), .c(n32086), .o(n39529) );
na03f01 g35738 ( .a(n39529), .b(n39526), .c(n3633), .o(n39530) );
na02f01 g35739 ( .a(n39529), .b(n39526), .o(n1719) );
na02f01 g35740 ( .a(n1719), .b(n6203), .o(n39532) );
na02f01 g35741 ( .a(n39532), .b(n39530), .o(n794) );
in01f01 g35742 ( .a(n21209), .o(n39534) );
in01f01 g35743 ( .a(n21210), .o(n39535) );
no02f01 g35744 ( .a(n39535), .b(n21066), .o(n39536) );
no02f01 g35745 ( .a(n39536), .b(n39534), .o(n39537) );
na02f01 g35746 ( .a(n39536), .b(n39534), .o(n39538) );
in01f01 g35747 ( .a(n39538), .o(n39539) );
no02f01 g35748 ( .a(n39539), .b(n39537), .o(n39540) );
in01f01 g35749 ( .a(n39540), .o(n799) );
na03f01 g35750 ( .a(n38858), .b(n9590), .c(n9589), .o(n39542) );
oa12f01 g35751 ( .a(n678), .b(n9646), .c(n9645), .o(n39543) );
na02f01 g35752 ( .a(n39543), .b(n39542), .o(n809) );
na02f01 g35753 ( .a(n32732), .b(sin_out_17), .o(n39545) );
no02f01 g35754 ( .a(n35905), .b(n35904), .o(n39546) );
no02f01 g35755 ( .a(n35761), .b(n34287), .o(n39547) );
no02f01 g35756 ( .a(n35762), .b(n34336), .o(n39548) );
no02f01 g35757 ( .a(n39548), .b(n39547), .o(n39549) );
no02f01 g35758 ( .a(n39549), .b(n39546), .o(n39550) );
na02f01 g35759 ( .a(n39549), .b(n39546), .o(n39551) );
in01f01 g35760 ( .a(n39551), .o(n39552) );
no02f01 g35761 ( .a(n39552), .b(n39550), .o(n39553) );
no02f01 g35762 ( .a(n39553), .b(n34307), .o(n39554) );
ao12f01 g35763 ( .a(n39502), .b(n39503), .c(n39501), .o(n39555) );
in01f01 g35764 ( .a(n39555), .o(n39556) );
in01f01 g35765 ( .a(n35696), .o(n39557) );
no02f01 g35766 ( .a(n39557), .b(n34336), .o(n39558) );
no02f01 g35767 ( .a(n35696), .b(n34287), .o(n39559) );
no02f01 g35768 ( .a(n39559), .b(n39558), .o(n39560) );
in01f01 g35769 ( .a(n39560), .o(n39561) );
no02f01 g35770 ( .a(n39561), .b(n39556), .o(n39562) );
no02f01 g35771 ( .a(n39560), .b(n39555), .o(n39563) );
no03f01 g35772 ( .a(n39563), .b(n39562), .c(n34267), .o(n39564) );
no02f01 g35773 ( .a(n39564), .b(n39511), .o(n39565) );
in01f01 g35774 ( .a(n39565), .o(n39566) );
no02f01 g35775 ( .a(n35718), .b(n35676), .o(n39567) );
oa12f01 g35776 ( .a(n39567), .b(n35704), .c(n35902), .o(n39568) );
in01f01 g35777 ( .a(n39568), .o(n39569) );
no02f01 g35778 ( .a(n35685), .b(n34287), .o(n39570) );
no02f01 g35779 ( .a(n39570), .b(n35687), .o(n39571) );
no02f01 g35780 ( .a(n39571), .b(n39569), .o(n39572) );
na02f01 g35781 ( .a(n39571), .b(n39569), .o(n39573) );
in01f01 g35782 ( .a(n39573), .o(n39574) );
no02f01 g35783 ( .a(n39574), .b(n39572), .o(n39575) );
in01f01 g35784 ( .a(n39575), .o(n39576) );
no02f01 g35785 ( .a(n39576), .b(n34267), .o(n39577) );
no02f01 g35786 ( .a(n39577), .b(n39566), .o(n39578) );
in01f01 g35787 ( .a(n39578), .o(n39579) );
no02f01 g35788 ( .a(n39568), .b(n39570), .o(n39580) );
no02f01 g35789 ( .a(n39580), .b(n35687), .o(n39581) );
no02f01 g35790 ( .a(n35713), .b(n34287), .o(n39582) );
no02f01 g35791 ( .a(n39582), .b(n35715), .o(n39583) );
in01f01 g35792 ( .a(n39583), .o(n39584) );
no02f01 g35793 ( .a(n39584), .b(n39581), .o(n39585) );
na02f01 g35794 ( .a(n39584), .b(n39581), .o(n39586) );
in01f01 g35795 ( .a(n39586), .o(n39587) );
no02f01 g35796 ( .a(n39587), .b(n39585), .o(n39588) );
in01f01 g35797 ( .a(n39588), .o(n39589) );
no02f01 g35798 ( .a(n39589), .b(n34267), .o(n39590) );
no04f01 g35799 ( .a(n39590), .b(n39579), .c(n39495), .d(n38595), .o(n39591) );
no02f01 g35800 ( .a(n39563), .b(n39562), .o(n39592) );
ao12f01 g35801 ( .a(n34307), .b(n39592), .c(n39509), .o(n39593) );
no02f01 g35802 ( .a(n39593), .b(n39499), .o(n39594) );
in01f01 g35803 ( .a(n39594), .o(n39595) );
ao12f01 g35804 ( .a(n34307), .b(n39588), .c(n39575), .o(n39596) );
no02f01 g35805 ( .a(n39596), .b(n39595), .o(n39597) );
in01f01 g35806 ( .a(n39597), .o(n39598) );
no02f01 g35807 ( .a(n39598), .b(n39591), .o(n39599) );
in01f01 g35808 ( .a(n39553), .o(n39600) );
no02f01 g35809 ( .a(n39600), .b(n34267), .o(n39601) );
no02f01 g35810 ( .a(n39601), .b(n39599), .o(n39602) );
no02f01 g35811 ( .a(n39548), .b(n39546), .o(n39603) );
no02f01 g35812 ( .a(n39603), .b(n39547), .o(n39604) );
no02f01 g35813 ( .a(n35754), .b(n34287), .o(n39605) );
no02f01 g35814 ( .a(n35755), .b(n34336), .o(n39606) );
no02f01 g35815 ( .a(n39606), .b(n39605), .o(n39607) );
no02f01 g35816 ( .a(n39607), .b(n39604), .o(n39608) );
na02f01 g35817 ( .a(n39607), .b(n39604), .o(n39609) );
in01f01 g35818 ( .a(n39609), .o(n39610) );
no03f01 g35819 ( .a(n39610), .b(n39608), .c(n34267), .o(n39611) );
no02f01 g35820 ( .a(n39610), .b(n39608), .o(n39612) );
no02f01 g35821 ( .a(n39612), .b(n34307), .o(n39613) );
no02f01 g35822 ( .a(n39613), .b(n39611), .o(n39614) );
in01f01 g35823 ( .a(n39614), .o(n39615) );
no03f01 g35824 ( .a(n39615), .b(n39602), .c(n39554), .o(n39616) );
no02f01 g35825 ( .a(n39602), .b(n39554), .o(n39617) );
no02f01 g35826 ( .a(n39614), .b(n39617), .o(n39618) );
oa12f01 g35827 ( .a(n32734), .b(n39618), .c(n39616), .o(n39619) );
na02f01 g35828 ( .a(n39619), .b(n39545), .o(n814) );
in01f01 g35829 ( .a(n37390), .o(n39621) );
no02f01 g35830 ( .a(n37389), .b(n9233), .o(n39622) );
oa12f01 g35831 ( .a(n39622), .b(n37385), .c(n9234), .o(n39623) );
na02f01 g35832 ( .a(n39623), .b(n39621), .o(n39624) );
in01f01 g35833 ( .a(n39624), .o(n39625) );
no03f01 g35834 ( .a(n9226), .b(n9224), .c(n8765), .o(n39626) );
no03f01 g35835 ( .a(n39624), .b(n9233), .c(n9227), .o(n39627) );
no03f01 g35836 ( .a(n39627), .b(n9234), .c(n9226), .o(n39628) );
no02f01 g35837 ( .a(n9224), .b(beta_31), .o(n39629) );
no02f01 g35838 ( .a(n9225), .b(n8765), .o(n39630) );
no02f01 g35839 ( .a(n39630), .b(n39629), .o(n39631) );
no02f01 g35840 ( .a(n39631), .b(n39628), .o(n39632) );
no02f01 g35841 ( .a(n39632), .b(n39626), .o(n39633) );
na03f01 g35842 ( .a(n39633), .b(n9590), .c(n9589), .o(n39634) );
in01f01 g35843 ( .a(n39633), .o(n3935) );
oa12f01 g35844 ( .a(n3935), .b(n9646), .c(n9645), .o(n39636) );
na02f01 g35845 ( .a(n39636), .b(n39634), .o(n823) );
na02f01 g35846 ( .a(n27253), .b(n27195), .o(n828) );
na03f01 g35847 ( .a(n9590), .b(n9589), .c(n9591), .o(n39639) );
oa12f01 g35848 ( .a(n4201), .b(n9646), .c(n9645), .o(n39640) );
na02f01 g35849 ( .a(n39640), .b(n39639), .o(n833) );
na03f01 g35850 ( .a(n9769), .b(n9746), .c(n36539), .o(n39642) );
in01f01 g35851 ( .a(n9816), .o(n39643) );
ao12f01 g35852 ( .a(n39643), .b(n9774), .c(n39642), .o(n39644) );
in01f01 g35853 ( .a(n9823), .o(n39645) );
in01f01 g35854 ( .a(n9831), .o(n39646) );
oa12f01 g35855 ( .a(n39646), .b(n39645), .c(n39644), .o(n39647) );
no04f01 g35856 ( .a(n9866), .b(n9854), .c(n9844), .d(n39647), .o(n39648) );
no03f01 g35857 ( .a(n9898), .b(n9873), .c(n39648), .o(n39649) );
no02f01 g35858 ( .a(n9897), .b(n9884), .o(n39650) );
oa12f01 g35859 ( .a(n39650), .b(n39649), .c(n9891), .o(n39651) );
in01f01 g35860 ( .a(n9891), .o(n39652) );
in01f01 g35861 ( .a(n9898), .o(n39653) );
na03f01 g35862 ( .a(n39653), .b(n9874), .c(n9868), .o(n39654) );
in01f01 g35863 ( .a(n39650), .o(n39655) );
na03f01 g35864 ( .a(n39655), .b(n39654), .c(n39652), .o(n39656) );
na02f01 g35865 ( .a(n39656), .b(n39651), .o(n838) );
na02f01 g35866 ( .a(n32732), .b(cos_out_20), .o(n39658) );
in01f01 g35867 ( .a(n35965), .o(n39659) );
na04f01 g35868 ( .a(n36264), .b(n36251), .c(n39659), .d(n35957), .o(n39660) );
na02f01 g35869 ( .a(n36267), .b(n39660), .o(n39661) );
na03f01 g35870 ( .a(n36363), .b(n36314), .c(n39661), .o(n39662) );
no02f01 g35871 ( .a(n36387), .b(n36230), .o(n39663) );
no02f01 g35872 ( .a(n39663), .b(n35912), .o(n39664) );
in01f01 g35873 ( .a(n34204), .o(n39665) );
ao12f01 g35874 ( .a(n34209), .b(n39665), .c(n34163), .o(n39666) );
no02f01 g35875 ( .a(n34171), .b(n33507), .o(n39667) );
no02f01 g35876 ( .a(n39667), .b(n34173), .o(n39668) );
no02f01 g35877 ( .a(n39668), .b(n39666), .o(n39669) );
na02f01 g35878 ( .a(n39668), .b(n39666), .o(n39670) );
in01f01 g35879 ( .a(n39670), .o(n39671) );
no02f01 g35880 ( .a(n39671), .b(n39669), .o(n39672) );
in01f01 g35881 ( .a(n39672), .o(n39673) );
no02f01 g35882 ( .a(n39673), .b(n35912), .o(n39674) );
no02f01 g35883 ( .a(n39674), .b(n39664), .o(n39675) );
in01f01 g35884 ( .a(n39675), .o(n39676) );
no03f01 g35885 ( .a(n34204), .b(n34173), .c(n34262), .o(n39677) );
no02f01 g35886 ( .a(n39667), .b(n34209), .o(n39678) );
in01f01 g35887 ( .a(n39678), .o(n39679) );
no02f01 g35888 ( .a(n34183), .b(n33507), .o(n39680) );
no02f01 g35889 ( .a(n39680), .b(n34185), .o(n39681) );
in01f01 g35890 ( .a(n39681), .o(n39682) );
no03f01 g35891 ( .a(n39682), .b(n39679), .c(n39677), .o(n39683) );
no02f01 g35892 ( .a(n39679), .b(n39677), .o(n39684) );
no02f01 g35893 ( .a(n39681), .b(n39684), .o(n39685) );
no02f01 g35894 ( .a(n39685), .b(n39683), .o(n39686) );
in01f01 g35895 ( .a(n39686), .o(n39687) );
no02f01 g35896 ( .a(n39687), .b(n35912), .o(n39688) );
no02f01 g35897 ( .a(n39688), .b(n39676), .o(n39689) );
in01f01 g35898 ( .a(n39689), .o(n39690) );
ao12f01 g35899 ( .a(n39690), .b(n36372), .c(n39662), .o(n39691) );
ao12f01 g35900 ( .a(n35944), .b(n36387), .c(n36230), .o(n39692) );
ao12f01 g35901 ( .a(n35944), .b(n39686), .c(n39672), .o(n39693) );
no02f01 g35902 ( .a(n39693), .b(n39692), .o(n39694) );
in01f01 g35903 ( .a(n39694), .o(n39695) );
no02f01 g35904 ( .a(n34263), .b(n34262), .o(n39696) );
in01f01 g35905 ( .a(n34211), .o(n39697) );
no02f01 g35906 ( .a(n33984), .b(n33507), .o(n39698) );
no02f01 g35907 ( .a(n33985), .b(n33508), .o(n39699) );
no02f01 g35908 ( .a(n39699), .b(n39698), .o(n39700) );
in01f01 g35909 ( .a(n39700), .o(n39701) );
no03f01 g35910 ( .a(n39701), .b(n39697), .c(n39696), .o(n39702) );
no02f01 g35911 ( .a(n39697), .b(n39696), .o(n39703) );
no02f01 g35912 ( .a(n39700), .b(n39703), .o(n39704) );
no02f01 g35913 ( .a(n39704), .b(n39702), .o(n39705) );
no02f01 g35914 ( .a(n39705), .b(n35944), .o(n39706) );
na02f01 g35915 ( .a(n39705), .b(n35944), .o(n39707) );
in01f01 g35916 ( .a(n39707), .o(n39708) );
no02f01 g35917 ( .a(n39708), .b(n39706), .o(n39709) );
in01f01 g35918 ( .a(n39709), .o(n39710) );
no03f01 g35919 ( .a(n39710), .b(n39695), .c(n39691), .o(n39711) );
oa12f01 g35920 ( .a(n39689), .b(n36373), .c(n36365), .o(n39712) );
ao12f01 g35921 ( .a(n39709), .b(n39694), .c(n39712), .o(n39713) );
oa12f01 g35922 ( .a(n32734), .b(n39713), .c(n39711), .o(n39714) );
na02f01 g35923 ( .a(n39714), .b(n39658), .o(n843) );
no03f01 g35924 ( .a(n9591), .b(n9232), .c(n936), .o(n39716) );
no02f01 g35925 ( .a(n4201), .b(n9238), .o(n39717) );
no02f01 g35926 ( .a(n39717), .b(n39716), .o(n39718) );
in01f01 g35927 ( .a(n39718), .o(n847) );
no02f01 g35928 ( .a(n37802), .b(n8534), .o(n39720) );
no02f01 g35929 ( .a(n8516), .b(n8471), .o(n39721) );
no02f01 g35930 ( .a(n39721), .b(n8518), .o(n39722) );
na02f01 g35931 ( .a(n39722), .b(n39720), .o(n39723) );
in01f01 g35932 ( .a(n39722), .o(n39724) );
oa12f01 g35933 ( .a(n39724), .b(n37802), .c(n8534), .o(n39725) );
na02f01 g35934 ( .a(n39725), .b(n39723), .o(n852) );
no02f01 g35935 ( .a(n8899), .b(beta_1), .o(n39727) );
no02f01 g35936 ( .a(n8862), .b(n8972), .o(n39728) );
oa12f01 g35937 ( .a(beta_0), .b(n39728), .c(n39727), .o(n39729) );
no02f01 g35938 ( .a(n39728), .b(n39727), .o(n39730) );
na02f01 g35939 ( .a(n39730), .b(n4932), .o(n39731) );
na02f01 g35940 ( .a(n39731), .b(n39729), .o(n857) );
in01f01 g35941 ( .a(n16232), .o(n39733) );
na03f01 g35942 ( .a(n39733), .b(n16149), .c(n16089), .o(n39734) );
oa12f01 g35943 ( .a(n21366), .b(n16232), .c(n16150), .o(n39735) );
na02f01 g35944 ( .a(n39735), .b(n39734), .o(n862) );
no02f01 g35945 ( .a(n38664), .b(n38662), .o(n39737) );
na02f01 g35946 ( .a(n39737), .b(n37062), .o(n39738) );
in01f01 g35947 ( .a(n39737), .o(n39739) );
na02f01 g35948 ( .a(n39739), .b(n37180), .o(n39740) );
na02f01 g35949 ( .a(n39740), .b(n39738), .o(n867) );
na02f01 g35950 ( .a(n32732), .b(cos_out_14), .o(n39742) );
no02f01 g35951 ( .a(n36370), .b(n36369), .o(n39743) );
in01f01 g35952 ( .a(n39743), .o(n39744) );
ao12f01 g35953 ( .a(n39744), .b(n36340), .c(n39043), .o(n39745) );
in01f01 g35954 ( .a(n39745), .o(n39746) );
no02f01 g35955 ( .a(n36360), .b(n35944), .o(n39747) );
no02f01 g35956 ( .a(n39747), .b(n36362), .o(n39748) );
in01f01 g35957 ( .a(n39748), .o(n39749) );
no02f01 g35958 ( .a(n39749), .b(n39746), .o(n39750) );
no02f01 g35959 ( .a(n39748), .b(n39745), .o(n39751) );
oa12f01 g35960 ( .a(n32734), .b(n39751), .c(n39750), .o(n39752) );
na02f01 g35961 ( .a(n39752), .b(n39742), .o(n872) );
no02f01 g35962 ( .a(n38556), .b(n38551), .o(n39754) );
na02f01 g35963 ( .a(n39754), .b(n38562), .o(n39755) );
in01f01 g35964 ( .a(n39754), .o(n39756) );
na02f01 g35965 ( .a(n39756), .b(n38554), .o(n39757) );
na03f01 g35966 ( .a(n39757), .b(n39755), .c(n1821), .o(n39758) );
na02f01 g35967 ( .a(n39757), .b(n39755), .o(n1889) );
na02f01 g35968 ( .a(n1889), .b(n8066), .o(n39760) );
na02f01 g35969 ( .a(n39760), .b(n39758), .o(n876) );
no02f01 g35970 ( .a(n20930), .b(n20887), .o(n39762) );
in01f01 g35971 ( .a(n39762), .o(n39763) );
na02f01 g35972 ( .a(n39763), .b(n39216), .o(n39764) );
na02f01 g35973 ( .a(n39762), .b(n39211), .o(n39765) );
na03f01 g35974 ( .a(n39765), .b(n39764), .c(n5799), .o(n39766) );
na02f01 g35975 ( .a(n39765), .b(n39764), .o(n2506) );
na02f01 g35976 ( .a(n2506), .b(n911), .o(n39768) );
na02f01 g35977 ( .a(n39768), .b(n39766), .o(n881) );
in01f01 g35978 ( .a(n14201), .o(n39770) );
no02f01 g35979 ( .a(n39770), .b(n14060), .o(n39771) );
in01f01 g35980 ( .a(n39771), .o(n39772) );
no02f01 g35981 ( .a(n14203), .b(n14048), .o(n39773) );
no02f01 g35982 ( .a(n39773), .b(n39772), .o(n39774) );
na02f01 g35983 ( .a(n39773), .b(n39772), .o(n39775) );
in01f01 g35984 ( .a(n39775), .o(n39776) );
no02f01 g35985 ( .a(n39776), .b(n39774), .o(n39777) );
in01f01 g35986 ( .a(n39777), .o(n4568) );
na02f01 g35987 ( .a(n4568), .b(n4116), .o(n39779) );
na02f01 g35988 ( .a(n39777), .b(n2589), .o(n39780) );
na02f01 g35989 ( .a(n39780), .b(n39779), .o(n886) );
in01f01 g35990 ( .a(n39162), .o(n39782) );
no02f01 g35991 ( .a(n39135), .b(n31532), .o(n39783) );
in01f01 g35992 ( .a(n31532), .o(n39784) );
no02f01 g35993 ( .a(n39059), .b(n39784), .o(n39785) );
no02f01 g35994 ( .a(n39785), .b(n39783), .o(n39786) );
in01f01 g35995 ( .a(n39163), .o(n39787) );
oa12f01 g35996 ( .a(n39787), .b(n39160), .c(n39173), .o(n39788) );
na03f01 g35997 ( .a(n39788), .b(n39786), .c(n39782), .o(n39789) );
in01f01 g35998 ( .a(n39786), .o(n39790) );
ao12f01 g35999 ( .a(n39163), .b(n39161), .c(n39153), .o(n39791) );
oa12f01 g36000 ( .a(n39790), .b(n39791), .c(n39162), .o(n39792) );
na02f01 g36001 ( .a(n39792), .b(n39789), .o(n891) );
no02f01 g36002 ( .a(n11814), .b(n11551), .o(n39794) );
na03f01 g36003 ( .a(n39794), .b(n11812), .c(n11801), .o(n39795) );
na02f01 g36004 ( .a(n11812), .b(n11801), .o(n39796) );
in01f01 g36005 ( .a(n39794), .o(n39797) );
na02f01 g36006 ( .a(n39797), .b(n39796), .o(n39798) );
na02f01 g36007 ( .a(n39798), .b(n39795), .o(n896) );
no02f01 g36008 ( .a(n27367), .b(n16153), .o(n39800) );
no02f01 g36009 ( .a(n27395), .b(n16152), .o(n39801) );
no02f01 g36010 ( .a(n39801), .b(n39800), .o(n39802) );
no02f01 g36011 ( .a(n38202), .b(n38197), .o(n39803) );
na02f01 g36012 ( .a(n39803), .b(n27676), .o(n39804) );
ao12f01 g36013 ( .a(n27367), .b(n38206), .c(n38200), .o(n39805) );
no02f01 g36014 ( .a(n39805), .b(n27677), .o(n39806) );
na03f01 g36015 ( .a(n39806), .b(n39804), .c(n39802), .o(n39807) );
in01f01 g36016 ( .a(n39802), .o(n39808) );
no03f01 g36017 ( .a(n38202), .b(n38197), .c(n27624), .o(n39809) );
in01f01 g36018 ( .a(n39806), .o(n39810) );
oa12f01 g36019 ( .a(n39808), .b(n39810), .c(n39809), .o(n39811) );
na02f01 g36020 ( .a(n39811), .b(n39807), .o(n901) );
in01f01 g36021 ( .a(n25328), .o(n39813) );
in01f01 g36022 ( .a(n25504), .o(n39814) );
oa12f01 g36023 ( .a(n39814), .b(n36666), .c(n25343), .o(n39815) );
in01f01 g36024 ( .a(n25516), .o(n39816) );
ao12f01 g36025 ( .a(n39813), .b(n39816), .c(n39815), .o(n39817) );
ao12f01 g36026 ( .a(n25515), .b(n25506), .c(n39815), .o(n39818) );
no04f01 g36027 ( .a(n25532), .b(n25527), .c(n39818), .d(n39817), .o(n39819) );
no02f01 g36028 ( .a(n39818), .b(n39817), .o(n39820) );
no02f01 g36029 ( .a(n25532), .b(n25527), .o(n39821) );
no02f01 g36030 ( .a(n39821), .b(n39820), .o(n39822) );
no02f01 g36031 ( .a(n39822), .b(n39819), .o(n39823) );
in01f01 g36032 ( .a(n39823), .o(n906) );
no02f01 g36033 ( .a(n39117), .b(n38323), .o(n39825) );
oa12f01 g36034 ( .a(n39825), .b(n39116), .c(n38337), .o(n39826) );
no02f01 g36035 ( .a(n39116), .b(n38337), .o(n39827) );
oa12f01 g36036 ( .a(n39827), .b(n39117), .c(n38323), .o(n39828) );
na02f01 g36037 ( .a(n39828), .b(n39826), .o(n916) );
in01f01 g36038 ( .a(n9600), .o(n39830) );
no02f01 g36039 ( .a(n39629), .b(n37389), .o(n39831) );
no02f01 g36040 ( .a(n39630), .b(n39831), .o(n39832) );
ao22f01 g36041 ( .a(n39832), .b(n39830), .c(n37384), .d(n9594), .o(n39833) );
in01f01 g36042 ( .a(n39833), .o(n39834) );
no02f01 g36043 ( .a(n39834), .b(n9591), .o(n39835) );
no02f01 g36044 ( .a(n39833), .b(n4201), .o(n39836) );
no02f01 g36045 ( .a(n39836), .b(n39835), .o(n39837) );
in01f01 g36046 ( .a(n39837), .o(n921) );
in01f01 g36047 ( .a(n28944), .o(n39839) );
in01f01 g36048 ( .a(n39308), .o(n39840) );
no02f01 g36049 ( .a(n39309), .b(n39296), .o(n39841) );
in01f01 g36050 ( .a(n39841), .o(n39842) );
ao12f01 g36051 ( .a(n39842), .b(n39840), .c(n39316), .o(n39843) );
in01f01 g36052 ( .a(n27964), .o(n39844) );
no02f01 g36053 ( .a(n29491), .b(n39844), .o(n39845) );
no02f01 g36054 ( .a(n29460), .b(n27964), .o(n39846) );
no02f01 g36055 ( .a(n39846), .b(n39845), .o(n39847) );
in01f01 g36056 ( .a(n39847), .o(n39848) );
in01f01 g36057 ( .a(n39299), .o(n39849) );
no02f01 g36058 ( .a(n39849), .b(n28081), .o(n39850) );
na02f01 g36059 ( .a(n39300), .b(n28081), .o(n39851) );
ao12f01 g36060 ( .a(n39850), .b(n39851), .c(n29491), .o(n39852) );
in01f01 g36061 ( .a(n39852), .o(n39853) );
no02f01 g36062 ( .a(n39853), .b(n39848), .o(n39854) );
no02f01 g36063 ( .a(n39852), .b(n39847), .o(n39855) );
no02f01 g36064 ( .a(n39855), .b(n39854), .o(n39856) );
no02f01 g36065 ( .a(n39856), .b(n_27014), .o(n39857) );
no02f01 g36066 ( .a(n39856), .b(n27681), .o(n39858) );
in01f01 g36067 ( .a(n39858), .o(n39859) );
oa12f01 g36068 ( .a(n39859), .b(n39857), .c(n39843), .o(n39860) );
in01f01 g36069 ( .a(n39860), .o(n39861) );
no02f01 g36070 ( .a(n39861), .b(n39839), .o(n39862) );
no02f01 g36071 ( .a(n39860), .b(n28944), .o(n39863) );
no02f01 g36072 ( .a(n39863), .b(n39862), .o(n39864) );
no02f01 g36073 ( .a(n28662), .b(n28383), .o(n39865) );
no02f01 g36074 ( .a(n28663), .b(n28102), .o(n39866) );
no02f01 g36075 ( .a(n39866), .b(n39865), .o(n39867) );
in01f01 g36076 ( .a(n39867), .o(n39868) );
ao12f01 g36077 ( .a(n39868), .b(n28633), .c(n28628), .o(n39869) );
na02f01 g36078 ( .a(n28633), .b(n28628), .o(n39870) );
no02f01 g36079 ( .a(n39867), .b(n39870), .o(n39871) );
no02f01 g36080 ( .a(n39871), .b(n39869), .o(n39872) );
in01f01 g36081 ( .a(n39872), .o(n39873) );
no02f01 g36082 ( .a(n39866), .b(n39870), .o(n39874) );
no02f01 g36083 ( .a(n39874), .b(n39865), .o(n39875) );
no02f01 g36084 ( .a(n28655), .b(n28383), .o(n39876) );
no02f01 g36085 ( .a(n28656), .b(n28102), .o(n39877) );
no02f01 g36086 ( .a(n39877), .b(n39876), .o(n39878) );
no02f01 g36087 ( .a(n39878), .b(n39875), .o(n39879) );
na02f01 g36088 ( .a(n39878), .b(n39875), .o(n39880) );
in01f01 g36089 ( .a(n39880), .o(n39881) );
no02f01 g36090 ( .a(n39881), .b(n39879), .o(n39882) );
in01f01 g36091 ( .a(n39882), .o(n39883) );
ao12f01 g36092 ( .a(n39861), .b(n39883), .c(n39873), .o(n39884) );
no02f01 g36093 ( .a(n39858), .b(n39857), .o(n39885) );
no02f01 g36094 ( .a(n39885), .b(n39843), .o(n39886) );
na02f01 g36095 ( .a(n39885), .b(n39843), .o(n39887) );
in01f01 g36096 ( .a(n39887), .o(n39888) );
no02f01 g36097 ( .a(n28604), .b(n28872), .o(n39889) );
no02f01 g36098 ( .a(n28602), .b(n28427), .o(n39890) );
no02f01 g36099 ( .a(n39890), .b(n39889), .o(n39891) );
na02f01 g36100 ( .a(n39890), .b(n39889), .o(n39892) );
in01f01 g36101 ( .a(n39892), .o(n39893) );
no02f01 g36102 ( .a(n39893), .b(n39891), .o(n39894) );
in01f01 g36103 ( .a(n39894), .o(n39895) );
no03f01 g36104 ( .a(n39895), .b(n39888), .c(n39886), .o(n39896) );
in01f01 g36105 ( .a(n39896), .o(n39897) );
oa12f01 g36106 ( .a(n39328), .b(n39478), .c(n39338), .o(n39898) );
oa12f01 g36107 ( .a(n39895), .b(n39888), .c(n39886), .o(n39899) );
na03f01 g36108 ( .a(n39899), .b(n39898), .c(n39327), .o(n39900) );
no02f01 g36109 ( .a(n28874), .b(n28427), .o(n39901) );
in01f01 g36110 ( .a(n39901), .o(n39902) );
in01f01 g36111 ( .a(n28400), .o(n39903) );
no02f01 g36112 ( .a(n28607), .b(n39903), .o(n39904) );
no02f01 g36113 ( .a(n39904), .b(n39902), .o(n39905) );
na02f01 g36114 ( .a(n39904), .b(n39902), .o(n39906) );
in01f01 g36115 ( .a(n39906), .o(n39907) );
no02f01 g36116 ( .a(n39907), .b(n39905), .o(n39908) );
in01f01 g36117 ( .a(n39908), .o(n39909) );
ao12f01 g36118 ( .a(n39903), .b(n28608), .c(n39901), .o(n39910) );
in01f01 g36119 ( .a(n28409), .o(n39911) );
no02f01 g36120 ( .a(n28410), .b(n39911), .o(n39912) );
no02f01 g36121 ( .a(n39912), .b(n39910), .o(n39913) );
na02f01 g36122 ( .a(n39912), .b(n39910), .o(n39914) );
in01f01 g36123 ( .a(n39914), .o(n39915) );
no02f01 g36124 ( .a(n39915), .b(n39913), .o(n39916) );
in01f01 g36125 ( .a(n39916), .o(n39917) );
ao12f01 g36126 ( .a(n39861), .b(n39917), .c(n39909), .o(n39918) );
in01f01 g36127 ( .a(n39918), .o(n39919) );
no02f01 g36128 ( .a(n28875), .b(n28411), .o(n39920) );
na02f01 g36129 ( .a(n28631), .b(n28102), .o(n39921) );
ao12f01 g36130 ( .a(n28632), .b(n39921), .c(n39920), .o(n39922) );
in01f01 g36131 ( .a(n39922), .o(n39923) );
no02f01 g36132 ( .a(n28620), .b(n28383), .o(n39924) );
no02f01 g36133 ( .a(n39924), .b(n28630), .o(n39925) );
no02f01 g36134 ( .a(n39925), .b(n39923), .o(n39926) );
na02f01 g36135 ( .a(n39925), .b(n39923), .o(n39927) );
in01f01 g36136 ( .a(n39927), .o(n39928) );
no02f01 g36137 ( .a(n39928), .b(n39926), .o(n39929) );
na02f01 g36138 ( .a(n39929), .b(n39860), .o(n39930) );
in01f01 g36139 ( .a(n39921), .o(n39931) );
no02f01 g36140 ( .a(n28632), .b(n39931), .o(n39932) );
no02f01 g36141 ( .a(n39932), .b(n39920), .o(n39933) );
na02f01 g36142 ( .a(n39932), .b(n39920), .o(n39934) );
in01f01 g36143 ( .a(n39934), .o(n39935) );
no02f01 g36144 ( .a(n39935), .b(n39933), .o(n39936) );
na02f01 g36145 ( .a(n39936), .b(n39860), .o(n39937) );
na02f01 g36146 ( .a(n39937), .b(n39930), .o(n39938) );
in01f01 g36147 ( .a(n39938), .o(n39939) );
na04f01 g36148 ( .a(n39939), .b(n39919), .c(n39900), .d(n39897), .o(n39940) );
no02f01 g36149 ( .a(n39917), .b(n39909), .o(n39941) );
no02f01 g36150 ( .a(n39941), .b(n39860), .o(n39942) );
ao12f01 g36151 ( .a(n39860), .b(n39936), .c(n39929), .o(n39943) );
no02f01 g36152 ( .a(n39943), .b(n39942), .o(n39944) );
ao12f01 g36153 ( .a(n39884), .b(n39944), .c(n39940), .o(n39945) );
no02f01 g36154 ( .a(n39870), .b(n28664), .o(n39946) );
in01f01 g36155 ( .a(n39946), .o(n39947) );
na02f01 g36156 ( .a(n28674), .b(n28102), .o(n39948) );
in01f01 g36157 ( .a(n39948), .o(n39949) );
no02f01 g36158 ( .a(n39949), .b(n28679), .o(n39950) );
oa12f01 g36159 ( .a(n39950), .b(n39947), .c(n28675), .o(n39951) );
no02f01 g36160 ( .a(n28681), .b(n28383), .o(n39952) );
no02f01 g36161 ( .a(n39952), .b(n28641), .o(n39953) );
in01f01 g36162 ( .a(n39953), .o(n39954) );
no02f01 g36163 ( .a(n39954), .b(n39951), .o(n39955) );
na02f01 g36164 ( .a(n39954), .b(n39951), .o(n39956) );
in01f01 g36165 ( .a(n39956), .o(n39957) );
no02f01 g36166 ( .a(n39957), .b(n39955), .o(n39958) );
in01f01 g36167 ( .a(n39958), .o(n39959) );
no02f01 g36168 ( .a(n39959), .b(n39861), .o(n39960) );
no02f01 g36169 ( .a(n39949), .b(n28675), .o(n39961) );
in01f01 g36170 ( .a(n39961), .o(n39962) );
no03f01 g36171 ( .a(n39962), .b(n39946), .c(n28679), .o(n39963) );
no02f01 g36172 ( .a(n39946), .b(n28679), .o(n39964) );
no02f01 g36173 ( .a(n39961), .b(n39964), .o(n39965) );
no02f01 g36174 ( .a(n39965), .b(n39963), .o(n39966) );
in01f01 g36175 ( .a(n39966), .o(n39967) );
no02f01 g36176 ( .a(n39967), .b(n39861), .o(n39968) );
no02f01 g36177 ( .a(n39968), .b(n39960), .o(n39969) );
no02f01 g36178 ( .a(n28902), .b(n28900), .o(n39970) );
in01f01 g36179 ( .a(n39970), .o(n39971) );
no02f01 g36180 ( .a(n28914), .b(n28909), .o(n39972) );
in01f01 g36181 ( .a(n39972), .o(n39973) );
ao12f01 g36182 ( .a(n39861), .b(n39973), .c(n39971), .o(n39974) );
in01f01 g36183 ( .a(n39974), .o(n39975) );
no02f01 g36184 ( .a(n39861), .b(n29296), .o(n39976) );
no02f01 g36185 ( .a(n39861), .b(n29295), .o(n39977) );
no02f01 g36186 ( .a(n39977), .b(n39976), .o(n39978) );
na02f01 g36187 ( .a(n39978), .b(n39975), .o(n39979) );
in01f01 g36188 ( .a(n39979), .o(n39980) );
ao12f01 g36189 ( .a(n39861), .b(n28934), .c(n28965), .o(n39981) );
in01f01 g36190 ( .a(n39981), .o(n39982) );
na04f01 g36191 ( .a(n39982), .b(n39980), .c(n39969), .d(n39945), .o(n39983) );
in01f01 g36192 ( .a(n28934), .o(n39984) );
ao12f01 g36193 ( .a(n39860), .b(n39984), .c(n28924), .o(n39985) );
in01f01 g36194 ( .a(n39985), .o(n39986) );
ao12f01 g36195 ( .a(n39860), .b(n39966), .c(n39958), .o(n39987) );
ao12f01 g36196 ( .a(n39860), .b(n39882), .c(n39872), .o(n39988) );
no02f01 g36197 ( .a(n39988), .b(n39987), .o(n39989) );
ao12f01 g36198 ( .a(n39860), .b(n28893), .c(n28888), .o(n39990) );
in01f01 g36199 ( .a(n39990), .o(n39991) );
na02f01 g36200 ( .a(n39991), .b(n39989), .o(n39992) );
ao12f01 g36201 ( .a(n39860), .b(n39972), .c(n39970), .o(n39993) );
no02f01 g36202 ( .a(n39993), .b(n39992), .o(n39994) );
na02f01 g36203 ( .a(n39994), .b(n39986), .o(n39995) );
in01f01 g36204 ( .a(n39995), .o(n39996) );
na03f01 g36205 ( .a(n39996), .b(n39983), .c(n39864), .o(n39997) );
in01f01 g36206 ( .a(n39864), .o(n39998) );
in01f01 g36207 ( .a(n39884), .o(n39999) );
in01f01 g36208 ( .a(n39338), .o(n40000) );
na03f01 g36209 ( .a(n39337), .b(n39335), .c(n39333), .o(n40001) );
no03f01 g36210 ( .a(n39382), .b(n39381), .c(n39379), .o(n40002) );
ao12f01 g36211 ( .a(n39376), .b(n39377), .c(n39374), .o(n40003) );
in01f01 g36212 ( .a(n39385), .o(n40004) );
oa12f01 g36213 ( .a(n40004), .b(n40003), .c(n40002), .o(n40005) );
na02f01 g36214 ( .a(n39389), .b(n39255), .o(n40006) );
na02f01 g36215 ( .a(n39387), .b(n39234), .o(n40007) );
ao12f01 g36216 ( .a(n39396), .b(n40007), .c(n40006), .o(n40008) );
na03f01 g36217 ( .a(n39396), .b(n40007), .c(n40006), .o(n40009) );
in01f01 g36218 ( .a(n39402), .o(n40010) );
ao12f01 g36219 ( .a(n39233), .b(n39401), .c(n39400), .o(n40011) );
in01f01 g36220 ( .a(n39410), .o(n40012) );
oa12f01 g36221 ( .a(n40012), .b(n40011), .c(n40010), .o(n40013) );
no03f01 g36222 ( .a(n40012), .b(n40011), .c(n40010), .o(n40014) );
na02f01 g36223 ( .a(n39417), .b(n39416), .o(n40015) );
na02f01 g36224 ( .a(n39414), .b(n39413), .o(n40016) );
ao12f01 g36225 ( .a(n39425), .b(n40016), .c(n40015), .o(n40017) );
na03f01 g36226 ( .a(n39425), .b(n40016), .c(n40015), .o(n40018) );
in01f01 g36227 ( .a(n39442), .o(n40019) );
in01f01 g36228 ( .a(n39443), .o(n40020) );
ao12f01 g36229 ( .a(n29666), .b(n29635), .c(n_27014), .o(n40021) );
no03f01 g36230 ( .a(n29662), .b(n29649), .c(n27681), .o(n40022) );
no02f01 g36231 ( .a(n40022), .b(n40021), .o(n40023) );
oa12f01 g36232 ( .a(n40019), .b(n40023), .c(n40020), .o(n40024) );
ao12f01 g36233 ( .a(n40017), .b(n40024), .c(n40018), .o(n40025) );
oa12f01 g36234 ( .a(n40013), .b(n40025), .c(n40014), .o(n40026) );
ao12f01 g36235 ( .a(n40008), .b(n40026), .c(n40009), .o(n40027) );
no03f01 g36236 ( .a(n40004), .b(n40003), .c(n40002), .o(n40028) );
ao12f01 g36237 ( .a(n40028), .b(n40027), .c(n40005), .o(n40029) );
in01f01 g36238 ( .a(n39466), .o(n40030) );
oa12f01 g36239 ( .a(n39371), .b(n39367), .c(n39360), .o(n40031) );
oa12f01 g36240 ( .a(n39465), .b(n39457), .c(n39456), .o(n40032) );
na02f01 g36241 ( .a(n40032), .b(n40031), .o(n40033) );
ao12f01 g36242 ( .a(n40033), .b(n40030), .c(n40029), .o(n40034) );
no03f01 g36243 ( .a(n39345), .b(n39313), .c(n39243), .o(n40035) );
ao12f01 g36244 ( .a(n39343), .b(n39268), .c(n39244), .o(n40036) );
in01f01 g36245 ( .a(n39353), .o(n40037) );
no03f01 g36246 ( .a(n40037), .b(n40036), .c(n40035), .o(n40038) );
no03f01 g36247 ( .a(n40038), .b(n40034), .c(n39372), .o(n40039) );
oa12f01 g36248 ( .a(n40001), .b(n40039), .c(n39354), .o(n40040) );
ao12f01 g36249 ( .a(n39484), .b(n40040), .c(n40000), .o(n40041) );
in01f01 g36250 ( .a(n39886), .o(n40042) );
ao12f01 g36251 ( .a(n39894), .b(n39887), .c(n40042), .o(n40043) );
no03f01 g36252 ( .a(n40043), .b(n40041), .c(n39326), .o(n40044) );
no04f01 g36253 ( .a(n39938), .b(n39918), .c(n40044), .d(n39896), .o(n40045) );
in01f01 g36254 ( .a(n39944), .o(n40046) );
oa12f01 g36255 ( .a(n39999), .b(n40046), .c(n40045), .o(n40047) );
in01f01 g36256 ( .a(n39969), .o(n40048) );
no04f01 g36257 ( .a(n39981), .b(n39979), .c(n40048), .d(n40047), .o(n40049) );
oa12f01 g36258 ( .a(n39998), .b(n39995), .c(n40049), .o(n40050) );
na02f01 g36259 ( .a(n40050), .b(n39997), .o(n926) );
no02f01 g36260 ( .a(n29938), .b(n24383), .o(n40052) );
no02f01 g36261 ( .a(n29937), .b(n24608), .o(n40053) );
no02f01 g36262 ( .a(n40053), .b(n40052), .o(n40054) );
no02f01 g36263 ( .a(n24576), .b(n24571), .o(n40055) );
ao12f01 g36264 ( .a(n29937), .b(n24602), .c(n40055), .o(n40056) );
in01f01 g36265 ( .a(n40056), .o(n40057) );
no02f01 g36266 ( .a(n24602), .b(n40055), .o(n40058) );
no02f01 g36267 ( .a(n40058), .b(n29938), .o(n40059) );
in01f01 g36268 ( .a(n40059), .o(n40060) );
oa12f01 g36269 ( .a(n40060), .b(n30046), .c(n30134), .o(n40061) );
na03f01 g36270 ( .a(n40061), .b(n40057), .c(n40054), .o(n40062) );
in01f01 g36271 ( .a(n40054), .o(n40063) );
ao12f01 g36272 ( .a(n40059), .b(n30047), .c(n30042), .o(n40064) );
oa12f01 g36273 ( .a(n40063), .b(n40064), .c(n40056), .o(n40065) );
na02f01 g36274 ( .a(n40065), .b(n40062), .o(n931) );
na03f01 g36275 ( .a(n40065), .b(n40062), .c(n6037), .o(n40067) );
no03f01 g36276 ( .a(n40064), .b(n40056), .c(n40063), .o(n40068) );
ao12f01 g36277 ( .a(n40054), .b(n40061), .c(n40057), .o(n40069) );
oa12f01 g36278 ( .a(n5873), .b(n40069), .c(n40068), .o(n40070) );
na02f01 g36279 ( .a(n40070), .b(n40067), .o(n941) );
no02f01 g36280 ( .a(n40044), .b(n39896), .o(n40072) );
no02f01 g36281 ( .a(n39908), .b(n39860), .o(n40073) );
no02f01 g36282 ( .a(n39909), .b(n39861), .o(n40074) );
in01f01 g36283 ( .a(n40074), .o(n40075) );
ao12f01 g36284 ( .a(n40073), .b(n40075), .c(n40072), .o(n40076) );
no02f01 g36285 ( .a(n39916), .b(n39860), .o(n40077) );
no02f01 g36286 ( .a(n39917), .b(n39861), .o(n40078) );
no02f01 g36287 ( .a(n40078), .b(n40077), .o(n40079) );
na02f01 g36288 ( .a(n40079), .b(n40076), .o(n40080) );
in01f01 g36289 ( .a(n40076), .o(n40081) );
in01f01 g36290 ( .a(n40079), .o(n40082) );
na02f01 g36291 ( .a(n40082), .b(n40081), .o(n40083) );
na02f01 g36292 ( .a(n40083), .b(n40080), .o(n946) );
na02f01 g36293 ( .a(n21025), .b(n18460), .o(n40085) );
in01f01 g36294 ( .a(n40085), .o(n40086) );
na02f01 g36295 ( .a(n29820), .b(n29817), .o(n40087) );
no02f01 g36296 ( .a(n21252), .b(n18459), .o(n40088) );
no02f01 g36297 ( .a(n40088), .b(n40087), .o(n40089) );
ao12f01 g36298 ( .a(n29747), .b(n21033), .c(n18459), .o(n40090) );
oa12f01 g36299 ( .a(n40090), .b(n21252), .c(n18460), .o(n40091) );
ao12f01 g36300 ( .a(n18460), .b(n21024), .c(n21023), .o(n40092) );
no03f01 g36301 ( .a(n40092), .b(n40091), .c(n40089), .o(n40093) );
no02f01 g36302 ( .a(n21001), .b(n18459), .o(n40094) );
no03f01 g36303 ( .a(n40094), .b(n40093), .c(n40086), .o(n40095) );
na02f01 g36304 ( .a(n20992), .b(n18460), .o(n40096) );
na02f01 g36305 ( .a(n40096), .b(n40095), .o(n40097) );
no02f01 g36306 ( .a(n20973), .b(n18459), .o(n40098) );
no02f01 g36307 ( .a(n40098), .b(n40097), .o(n40099) );
na02f01 g36308 ( .a(n20968), .b(n18459), .o(n40100) );
no02f01 g36309 ( .a(n20987), .b(n18460), .o(n40101) );
no02f01 g36310 ( .a(n21001), .b(n18460), .o(n40102) );
no02f01 g36311 ( .a(n40102), .b(n40101), .o(n40103) );
na02f01 g36312 ( .a(n40103), .b(n40100), .o(n40104) );
ao12f01 g36313 ( .a(n18460), .b(n20947), .c(n20945), .o(n40105) );
no02f01 g36314 ( .a(n20949), .b(n18459), .o(n40106) );
no04f01 g36315 ( .a(n40106), .b(n40105), .c(n40104), .d(n40099), .o(n40107) );
in01f01 g36316 ( .a(n40099), .o(n40108) );
in01f01 g36317 ( .a(n40104), .o(n40109) );
in01f01 g36318 ( .a(n40105), .o(n40110) );
in01f01 g36319 ( .a(n40106), .o(n40111) );
ao22f01 g36320 ( .a(n40111), .b(n40110), .c(n40109), .d(n40108), .o(n40112) );
no02f01 g36321 ( .a(n40112), .b(n40107), .o(n40113) );
no02f01 g36322 ( .a(n40113), .b(n20379), .o(n40114) );
in01f01 g36323 ( .a(n40103), .o(n40115) );
ao12f01 g36324 ( .a(n40115), .b(n40096), .c(n40095), .o(n40116) );
in01f01 g36325 ( .a(n40100), .o(n40117) );
no02f01 g36326 ( .a(n40117), .b(n40098), .o(n40118) );
no02f01 g36327 ( .a(n40118), .b(n40116), .o(n40119) );
na02f01 g36328 ( .a(n40118), .b(n40116), .o(n40120) );
in01f01 g36329 ( .a(n40120), .o(n40121) );
no02f01 g36330 ( .a(n40121), .b(n40119), .o(n40122) );
no02f01 g36331 ( .a(n40122), .b(n20221), .o(n40123) );
in01f01 g36332 ( .a(n40123), .o(n40124) );
no02f01 g36333 ( .a(n40102), .b(n40095), .o(n40125) );
in01f01 g36334 ( .a(n40096), .o(n40126) );
no02f01 g36335 ( .a(n40101), .b(n40126), .o(n40127) );
no02f01 g36336 ( .a(n40127), .b(n40125), .o(n40128) );
na02f01 g36337 ( .a(n40127), .b(n40125), .o(n40129) );
in01f01 g36338 ( .a(n40129), .o(n40130) );
no02f01 g36339 ( .a(n40130), .b(n40128), .o(n40131) );
na02f01 g36340 ( .a(n40131), .b(n20214), .o(n40132) );
no02f01 g36341 ( .a(n40093), .b(n40086), .o(n40133) );
in01f01 g36342 ( .a(n40133), .o(n40134) );
no02f01 g36343 ( .a(n40102), .b(n40094), .o(n40135) );
no02f01 g36344 ( .a(n40135), .b(n40134), .o(n40136) );
in01f01 g36345 ( .a(n40136), .o(n40137) );
na02f01 g36346 ( .a(n40135), .b(n40134), .o(n40138) );
na02f01 g36347 ( .a(n40138), .b(n40137), .o(n40139) );
na02f01 g36348 ( .a(n40139), .b(n21154), .o(n40140) );
no02f01 g36349 ( .a(n40091), .b(n40089), .o(n40141) );
in01f01 g36350 ( .a(n40092), .o(n40142) );
ao12f01 g36351 ( .a(n40141), .b(n40142), .c(n40085), .o(n40143) );
no04f01 g36352 ( .a(n40092), .b(n40091), .c(n40089), .d(n40086), .o(n40144) );
no02f01 g36353 ( .a(n40144), .b(n40143), .o(n40145) );
in01f01 g36354 ( .a(n40145), .o(n40146) );
no02f01 g36355 ( .a(n20055), .b(n19763), .o(n40147) );
ao12f01 g36356 ( .a(n19833), .b(n40147), .c(n20044), .o(n40148) );
no02f01 g36357 ( .a(n19836), .b(n19739), .o(n40149) );
in01f01 g36358 ( .a(n40149), .o(n40150) );
no02f01 g36359 ( .a(n40150), .b(n40148), .o(n40151) );
na02f01 g36360 ( .a(n40150), .b(n40148), .o(n40152) );
in01f01 g36361 ( .a(n40152), .o(n40153) );
no02f01 g36362 ( .a(n40153), .b(n40151), .o(n40154) );
in01f01 g36363 ( .a(n40154), .o(n40155) );
no02f01 g36364 ( .a(n40155), .b(n40146), .o(n40156) );
in01f01 g36365 ( .a(n40156), .o(n40157) );
oa12f01 g36366 ( .a(n29829), .b(n29828), .c(n29816), .o(n40158) );
no02f01 g36367 ( .a(n21252), .b(n18460), .o(n40159) );
na02f01 g36368 ( .a(n40090), .b(n40087), .o(n40160) );
no03f01 g36369 ( .a(n40160), .b(n40159), .c(n40088), .o(n40161) );
no02f01 g36370 ( .a(n40159), .b(n40088), .o(n40162) );
ao12f01 g36371 ( .a(n40162), .b(n40090), .c(n40087), .o(n40163) );
no04f01 g36372 ( .a(n19833), .b(n20055), .c(n19763), .d(n19752), .o(n40164) );
ao12f01 g36373 ( .a(n40147), .b(n20056), .c(n20044), .o(n40165) );
no02f01 g36374 ( .a(n40165), .b(n40164), .o(n40166) );
in01f01 g36375 ( .a(n40166), .o(n40167) );
no03f01 g36376 ( .a(n40167), .b(n40163), .c(n40161), .o(n40168) );
no02f01 g36377 ( .a(n40154), .b(n40145), .o(n40169) );
no02f01 g36378 ( .a(n40163), .b(n40161), .o(n40170) );
no02f01 g36379 ( .a(n40166), .b(n40170), .o(n40171) );
no02f01 g36380 ( .a(n40171), .b(n40169), .o(n40172) );
oa12f01 g36381 ( .a(n40172), .b(n40168), .c(n40158), .o(n40173) );
na02f01 g36382 ( .a(n40173), .b(n40157), .o(n40174) );
no02f01 g36383 ( .a(n40139), .b(n21154), .o(n40175) );
oa12f01 g36384 ( .a(n40140), .b(n40175), .c(n40174), .o(n40176) );
no02f01 g36385 ( .a(n40131), .b(n20214), .o(n40177) );
oa12f01 g36386 ( .a(n40132), .b(n40177), .c(n40176), .o(n40178) );
na02f01 g36387 ( .a(n40122), .b(n20221), .o(n40179) );
in01f01 g36388 ( .a(n40179), .o(n40180) );
oa12f01 g36389 ( .a(n40124), .b(n40180), .c(n40178), .o(n40181) );
na02f01 g36390 ( .a(n40113), .b(n20379), .o(n40182) );
ao12f01 g36391 ( .a(n40114), .b(n40182), .c(n40181), .o(n40183) );
no03f01 g36392 ( .a(n40105), .b(n40104), .c(n40099), .o(n40184) );
no02f01 g36393 ( .a(n40184), .b(n40106), .o(n40185) );
no02f01 g36394 ( .a(n21323), .b(n18460), .o(n40186) );
ao12f01 g36395 ( .a(n18459), .b(n20918), .c(n20917), .o(n40187) );
no03f01 g36396 ( .a(n40187), .b(n40186), .c(n40185), .o(n40188) );
in01f01 g36397 ( .a(n40185), .o(n40189) );
no02f01 g36398 ( .a(n40187), .b(n40186), .o(n40190) );
no02f01 g36399 ( .a(n40190), .b(n40189), .o(n40191) );
no02f01 g36400 ( .a(n40191), .b(n40188), .o(n40192) );
no02f01 g36401 ( .a(n40192), .b(n20236), .o(n40193) );
na02f01 g36402 ( .a(n40192), .b(n20236), .o(n40194) );
in01f01 g36403 ( .a(n40194), .o(n40195) );
no02f01 g36404 ( .a(n40195), .b(n40193), .o(n40196) );
no02f01 g36405 ( .a(n40196), .b(n40183), .o(n40197) );
na02f01 g36406 ( .a(n40196), .b(n40183), .o(n40198) );
in01f01 g36407 ( .a(n40198), .o(n40199) );
no02f01 g36408 ( .a(n40199), .b(n40197), .o(n40200) );
in01f01 g36409 ( .a(n40200), .o(n951) );
in01f01 g36410 ( .a(n40072), .o(n40202) );
in01f01 g36411 ( .a(n39942), .o(n40203) );
ao12f01 g36412 ( .a(n39918), .b(n40203), .c(n40202), .o(n40204) );
in01f01 g36413 ( .a(n39937), .o(n40205) );
no02f01 g36414 ( .a(n39936), .b(n39860), .o(n40206) );
no02f01 g36415 ( .a(n40206), .b(n40205), .o(n40207) );
in01f01 g36416 ( .a(n40207), .o(n40208) );
na02f01 g36417 ( .a(n40208), .b(n40204), .o(n40209) );
in01f01 g36418 ( .a(n40204), .o(n40210) );
na02f01 g36419 ( .a(n40207), .b(n40210), .o(n40211) );
na02f01 g36420 ( .a(n40211), .b(n40209), .o(n956) );
na02f01 g36421 ( .a(n30037), .b(n29944), .o(n40213) );
no02f01 g36422 ( .a(n36521), .b(n36518), .o(n40214) );
na02f01 g36423 ( .a(n40214), .b(n40213), .o(n40215) );
in01f01 g36424 ( .a(n40214), .o(n40216) );
na02f01 g36425 ( .a(n40216), .b(n36520), .o(n40217) );
na03f01 g36426 ( .a(n40217), .b(n40215), .c(n6037), .o(n40218) );
na02f01 g36427 ( .a(n40217), .b(n40215), .o(n2003) );
na02f01 g36428 ( .a(n2003), .b(n5873), .o(n40220) );
na02f01 g36429 ( .a(n40220), .b(n40218), .o(n961) );
oa12f01 g36430 ( .a(n7506), .b(n7532), .c(n7531), .o(n40222) );
na03f01 g36431 ( .a(n7505), .b(n7501), .c(n7500), .o(n40223) );
na02f01 g36432 ( .a(n40223), .b(n40222), .o(n966) );
na02f01 g36433 ( .a(n37323), .b(n37319), .o(n971) );
no02f01 g36434 ( .a(n30123), .b(n29967), .o(n40226) );
no02f01 g36435 ( .a(n40226), .b(n30014), .o(n40227) );
na02f01 g36436 ( .a(n40226), .b(n30014), .o(n40228) );
in01f01 g36437 ( .a(n40228), .o(n40229) );
no02f01 g36438 ( .a(n40229), .b(n40227), .o(n40230) );
in01f01 g36439 ( .a(n40230), .o(n976) );
no02f01 g36440 ( .a(n9631), .b(n9287), .o(n40232) );
in01f01 g36441 ( .a(n40232), .o(n40233) );
na02f01 g36442 ( .a(n40233), .b(n9426), .o(n40234) );
na02f01 g36443 ( .a(n40232), .b(n9630), .o(n40235) );
na02f01 g36444 ( .a(n40235), .b(n40234), .o(n981) );
no02f01 g36445 ( .a(n36483), .b(n36504), .o(n40237) );
in01f01 g36446 ( .a(n40237), .o(n40238) );
no02f01 g36447 ( .a(n40238), .b(n36501), .o(n40239) );
no02f01 g36448 ( .a(n40237), .b(n36461), .o(n40240) );
no02f01 g36449 ( .a(n40240), .b(n40239), .o(n40241) );
na02f01 g36450 ( .a(n40241), .b(n2589), .o(n40242) );
in01f01 g36451 ( .a(n40241), .o(n5730) );
na02f01 g36452 ( .a(n5730), .b(n4116), .o(n40244) );
na02f01 g36453 ( .a(n40244), .b(n40242), .o(n986) );
no02f01 g36454 ( .a(n38144), .b(n38148), .o(n40246) );
in01f01 g36455 ( .a(n40246), .o(n40247) );
in01f01 g36456 ( .a(n5870), .o(n40248) );
oa12f01 g36457 ( .a(n5563_1), .b(n40248), .c(n40247), .o(n40249) );
no02f01 g36458 ( .a(n40249), .b(n5585), .o(n40250) );
no02f01 g36459 ( .a(n40250), .b(n5578_1), .o(n40251) );
in01f01 g36460 ( .a(n40251), .o(n40252) );
no02f01 g36461 ( .a(n5583_1), .b(n5569), .o(n40253) );
no02f01 g36462 ( .a(n40253), .b(n40252), .o(n40254) );
na02f01 g36463 ( .a(n40253), .b(n40252), .o(n40255) );
in01f01 g36464 ( .a(n40255), .o(n40256) );
no03f01 g36465 ( .a(n40256), .b(n40254), .c(n5873), .o(n40257) );
in01f01 g36466 ( .a(n40249), .o(n40258) );
no02f01 g36467 ( .a(n5585), .b(n5578_1), .o(n40259) );
no02f01 g36468 ( .a(n40259), .b(n40258), .o(n40260) );
na02f01 g36469 ( .a(n40259), .b(n40258), .o(n40261) );
in01f01 g36470 ( .a(n40261), .o(n40262) );
no02f01 g36471 ( .a(n40262), .b(n40260), .o(n40263) );
in01f01 g36472 ( .a(n40263), .o(n40264) );
no02f01 g36473 ( .a(n40264), .b(n5873), .o(n40265) );
no02f01 g36474 ( .a(n40265), .b(n40257), .o(n40266) );
in01f01 g36475 ( .a(n40266), .o(n40267) );
ao12f01 g36476 ( .a(n5587), .b(n40249), .c(n5579), .o(n40268) );
in01f01 g36477 ( .a(n40268), .o(n40269) );
no02f01 g36478 ( .a(n5589), .b(n5528_1), .o(n40270) );
in01f01 g36479 ( .a(n40270), .o(n40271) );
no02f01 g36480 ( .a(n40271), .b(n40269), .o(n40272) );
no02f01 g36481 ( .a(n40270), .b(n40268), .o(n40273) );
no03f01 g36482 ( .a(n40273), .b(n40272), .c(n5873), .o(n40274) );
in01f01 g36483 ( .a(n5554), .o(n40275) );
ao12f01 g36484 ( .a(n5545), .b(n5866), .c(n40246), .o(n40276) );
ao12f01 g36485 ( .a(n5865), .b(n40276), .c(n40275), .o(n40277) );
in01f01 g36486 ( .a(n40277), .o(n40278) );
no02f01 g36487 ( .a(n5869_1), .b(n5562), .o(n40279) );
no02f01 g36488 ( .a(n40279), .b(n40278), .o(n40280) );
na02f01 g36489 ( .a(n40279), .b(n40278), .o(n40281) );
in01f01 g36490 ( .a(n40281), .o(n40282) );
no02f01 g36491 ( .a(n40282), .b(n40280), .o(n40283) );
in01f01 g36492 ( .a(n40283), .o(n40284) );
no02f01 g36493 ( .a(n40284), .b(n5873), .o(n40285) );
in01f01 g36494 ( .a(n40276), .o(n40286) );
no02f01 g36495 ( .a(n5865), .b(n5554), .o(n40287) );
in01f01 g36496 ( .a(n40287), .o(n40288) );
no02f01 g36497 ( .a(n40288), .b(n40286), .o(n40289) );
no02f01 g36498 ( .a(n40287), .b(n40276), .o(n40290) );
no02f01 g36499 ( .a(n40290), .b(n40289), .o(n40291) );
in01f01 g36500 ( .a(n40291), .o(n40292) );
no02f01 g36501 ( .a(n40292), .b(n5873), .o(n40293) );
no02f01 g36502 ( .a(n5867), .b(n5537), .o(n40294) );
in01f01 g36503 ( .a(n40294), .o(n40295) );
no03f01 g36504 ( .a(n40295), .b(n40246), .c(n5543_1), .o(n40296) );
no02f01 g36505 ( .a(n40246), .b(n5543_1), .o(n40297) );
no02f01 g36506 ( .a(n40294), .b(n40297), .o(n40298) );
no03f01 g36507 ( .a(n40298), .b(n40296), .c(n5873), .o(n40299) );
no02f01 g36508 ( .a(n40299), .b(n38152), .o(n40300) );
in01f01 g36509 ( .a(n40300), .o(n40301) );
no03f01 g36510 ( .a(n40301), .b(n40293), .c(n40285), .o(n40302) );
in01f01 g36511 ( .a(n40302), .o(n40303) );
no03f01 g36512 ( .a(n40303), .b(n40274), .c(n40267), .o(n40304) );
in01f01 g36513 ( .a(n40304), .o(n40305) );
no02f01 g36514 ( .a(n40298), .b(n40296), .o(n40306) );
ao12f01 g36515 ( .a(n6037), .b(n40306), .c(n38150), .o(n40307) );
in01f01 g36516 ( .a(n40307), .o(n40308) );
oa12f01 g36517 ( .a(n5873), .b(n40292), .c(n40284), .o(n40309) );
na02f01 g36518 ( .a(n40309), .b(n40308), .o(n40310) );
no02f01 g36519 ( .a(n40273), .b(n40272), .o(n40311) );
no02f01 g36520 ( .a(n40256), .b(n40254), .o(n40312) );
no02f01 g36521 ( .a(n40263), .b(n6037), .o(n40313) );
in01f01 g36522 ( .a(n40313), .o(n40314) );
ao12f01 g36523 ( .a(n6037), .b(n40314), .c(n40312), .o(n40315) );
in01f01 g36524 ( .a(n40315), .o(n40316) );
ao12f01 g36525 ( .a(n6037), .b(n40316), .c(n40311), .o(n40317) );
no02f01 g36526 ( .a(n40317), .b(n40310), .o(n40318) );
oa12f01 g36527 ( .a(n40318), .b(n40305), .c(n38143), .o(n2861) );
in01f01 g36528 ( .a(n2861), .o(n991) );
na03f01 g36529 ( .a(n39980), .b(n39969), .c(n39945), .o(n40321) );
no02f01 g36530 ( .a(n39860), .b(n28924), .o(n40322) );
no02f01 g36531 ( .a(n39861), .b(n28965), .o(n40323) );
no02f01 g36532 ( .a(n40323), .b(n40322), .o(n40324) );
na03f01 g36533 ( .a(n40324), .b(n39994), .c(n40321), .o(n40325) );
no03f01 g36534 ( .a(n39979), .b(n40048), .c(n40047), .o(n40326) );
in01f01 g36535 ( .a(n39994), .o(n40327) );
in01f01 g36536 ( .a(n40324), .o(n40328) );
oa12f01 g36537 ( .a(n40328), .b(n40327), .c(n40326), .o(n40329) );
na02f01 g36538 ( .a(n40329), .b(n40325), .o(n996) );
in01f01 g36539 ( .a(n39029), .o(n40331) );
no02f01 g36540 ( .a(n14230), .b(n14226), .o(n40332) );
no02f01 g36541 ( .a(n40332), .b(n40331), .o(n40333) );
na02f01 g36542 ( .a(n40332), .b(n40331), .o(n40334) );
in01f01 g36543 ( .a(n40334), .o(n40335) );
no02f01 g36544 ( .a(n40335), .b(n40333), .o(n40336) );
in01f01 g36545 ( .a(n40336), .o(n5036) );
na02f01 g36546 ( .a(n5036), .b(n4116), .o(n40338) );
na02f01 g36547 ( .a(n40336), .b(n2589), .o(n40339) );
na02f01 g36548 ( .a(n40339), .b(n40338), .o(n1001) );
no02f01 g36549 ( .a(n9775), .b(n9771), .o(n40341) );
no02f01 g36550 ( .a(n9793), .b(n5001), .o(n40342) );
no02f01 g36551 ( .a(n40342), .b(n9795), .o(n40343) );
na02f01 g36552 ( .a(n40343), .b(n40341), .o(n40344) );
in01f01 g36553 ( .a(n40343), .o(n40345) );
oa12f01 g36554 ( .a(n40345), .b(n9775), .c(n9771), .o(n40346) );
na02f01 g36555 ( .a(n40346), .b(n40344), .o(n1006) );
no02f01 g36556 ( .a(n11815), .b(n11551), .o(n40348) );
no02f01 g36557 ( .a(n11816), .b(n11535), .o(n40349) );
na02f01 g36558 ( .a(n40349), .b(n40348), .o(n40350) );
in01f01 g36559 ( .a(n40349), .o(n40351) );
oa12f01 g36560 ( .a(n40351), .b(n11815), .c(n11551), .o(n40352) );
na02f01 g36561 ( .a(n40352), .b(n40350), .o(n1011) );
in01f01 g36562 ( .a(n27167), .o(n40354) );
in01f01 g36563 ( .a(n27146), .o(n40355) );
oa12f01 g36564 ( .a(n40355), .b(n27248), .c(n27239), .o(n40356) );
no02f01 g36565 ( .a(n27169), .b(n26440), .o(n40357) );
no02f01 g36566 ( .a(n40357), .b(n27154), .o(n40358) );
na03f01 g36567 ( .a(n40358), .b(n40356), .c(n40354), .o(n40359) );
ao12f01 g36568 ( .a(n27146), .b(n27124), .c(n27112), .o(n40360) );
in01f01 g36569 ( .a(n40358), .o(n40361) );
oa12f01 g36570 ( .a(n40361), .b(n40360), .c(n27167), .o(n40362) );
na03f01 g36571 ( .a(n40362), .b(n40359), .c(n1821), .o(n40363) );
na02f01 g36572 ( .a(n40362), .b(n40359), .o(n5385) );
na02f01 g36573 ( .a(n5385), .b(n8066), .o(n40365) );
na02f01 g36574 ( .a(n40365), .b(n40363), .o(n1016) );
no02f01 g36575 ( .a(n9591), .b(n9232), .o(n40367) );
no03f01 g36576 ( .a(n40367), .b(n4201), .c(n936), .o(n40368) );
ao12f01 g36577 ( .a(n9591), .b(n9232), .c(n9228), .o(n40369) );
no02f01 g36578 ( .a(n40369), .b(n40368), .o(n40370) );
in01f01 g36579 ( .a(n40370), .o(n1021) );
na02f01 g36580 ( .a(n40200), .b(n5799), .o(n40372) );
na02f01 g36581 ( .a(n951), .b(n911), .o(n40373) );
na02f01 g36582 ( .a(n40373), .b(n40372), .o(n1026) );
na02f01 g36583 ( .a(n32732), .b(sin_out_3), .o(n40375) );
no02f01 g36584 ( .a(n34344), .b(n34267), .o(n40376) );
no02f01 g36585 ( .a(n34343), .b(n34307), .o(n40377) );
no02f01 g36586 ( .a(n40377), .b(n40376), .o(n40378) );
in01f01 g36587 ( .a(n40378), .o(n40379) );
no03f01 g36588 ( .a(n40379), .b(n34345), .c(n34328), .o(n40380) );
in01f01 g36589 ( .a(n34345), .o(n40381) );
ao12f01 g36590 ( .a(n40378), .b(n40381), .c(n36563), .o(n40382) );
oa12f01 g36591 ( .a(n32734), .b(n40382), .c(n40380), .o(n40383) );
na02f01 g36592 ( .a(n40383), .b(n40375), .o(n1031) );
na02f01 g36593 ( .a(n39919), .b(n40072), .o(n40385) );
no02f01 g36594 ( .a(n40206), .b(n39942), .o(n40386) );
ao12f01 g36595 ( .a(n40205), .b(n40386), .c(n40385), .o(n40387) );
in01f01 g36596 ( .a(n39930), .o(n40388) );
no02f01 g36597 ( .a(n39929), .b(n39860), .o(n40389) );
no02f01 g36598 ( .a(n40389), .b(n40388), .o(n40390) );
in01f01 g36599 ( .a(n40390), .o(n40391) );
na02f01 g36600 ( .a(n40391), .b(n40387), .o(n40392) );
in01f01 g36601 ( .a(n40387), .o(n40393) );
na02f01 g36602 ( .a(n40390), .b(n40393), .o(n40394) );
na02f01 g36603 ( .a(n40394), .b(n40392), .o(n1035) );
in01f01 g36604 ( .a(n11854), .o(n40396) );
in01f01 g36605 ( .a(n11862), .o(n40397) );
na02f01 g36606 ( .a(n40397), .b(n30140), .o(n40398) );
no02f01 g36607 ( .a(n11864), .b(n11859), .o(n40399) );
in01f01 g36608 ( .a(n40399), .o(n40400) );
na03f01 g36609 ( .a(n40400), .b(n40398), .c(n40396), .o(n40401) );
na02f01 g36610 ( .a(n40398), .b(n40396), .o(n40402) );
na02f01 g36611 ( .a(n40399), .b(n40402), .o(n40403) );
na02f01 g36612 ( .a(n40403), .b(n40401), .o(n1040) );
no02f01 g36613 ( .a(n9720), .b(n9697), .o(n40405) );
no02f01 g36614 ( .a(n9705), .b(n5001), .o(n40406) );
no02f01 g36615 ( .a(n40406), .b(n9707), .o(n40407) );
na02f01 g36616 ( .a(n40407), .b(n40405), .o(n40408) );
in01f01 g36617 ( .a(n40407), .o(n40409) );
oa12f01 g36618 ( .a(n40409), .b(n9720), .c(n9697), .o(n40410) );
na02f01 g36619 ( .a(n40410), .b(n40408), .o(n1045) );
ao12f01 g36620 ( .a(n9234), .b(n37382), .c(n8899), .o(n40412) );
in01f01 g36621 ( .a(n40412), .o(n40413) );
no02f01 g36622 ( .a(n40413), .b(n3623), .o(n40414) );
no02f01 g36623 ( .a(n40412), .b(n37391), .o(n40415) );
no02f01 g36624 ( .a(n40415), .b(n40414), .o(n40416) );
in01f01 g36625 ( .a(n40416), .o(n1050) );
in01f01 g36626 ( .a(n39988), .o(n40418) );
no02f01 g36627 ( .a(n39966), .b(n39860), .o(n40419) );
no02f01 g36628 ( .a(n40419), .b(n39968), .o(n40420) );
na03f01 g36629 ( .a(n40420), .b(n40418), .c(n40047), .o(n40421) );
in01f01 g36630 ( .a(n40420), .o(n40422) );
oa12f01 g36631 ( .a(n40422), .b(n39988), .c(n39945), .o(n40423) );
na02f01 g36632 ( .a(n40423), .b(n40421), .o(n1055) );
in01f01 g36633 ( .a(n5900), .o(n40425) );
oa22f01 g36634 ( .a(n5912), .b(n5910), .c(n5901), .d(n40425), .o(n40426) );
no02f01 g36635 ( .a(n5912), .b(n5910), .o(n40427) );
na03f01 g36636 ( .a(n40427), .b(n5902), .c(n5900), .o(n40428) );
na02f01 g36637 ( .a(n40428), .b(n40426), .o(n1060) );
no02f01 g36638 ( .a(n38681), .b(n36122), .o(n40430) );
no02f01 g36639 ( .a(n40430), .b(n38715), .o(n40431) );
no02f01 g36640 ( .a(n38698), .b(n36122), .o(n40432) );
no02f01 g36641 ( .a(n40432), .b(n38700), .o(n40433) );
na03f01 g36642 ( .a(n40433), .b(n40431), .c(n38689), .o(n40434) );
in01f01 g36643 ( .a(n40431), .o(n40435) );
in01f01 g36644 ( .a(n40433), .o(n40436) );
oa12f01 g36645 ( .a(n40436), .b(n40435), .c(n38786), .o(n40437) );
na02f01 g36646 ( .a(n40437), .b(n40434), .o(n1065) );
no02f01 g36647 ( .a(n16486), .b(n16329), .o(n40439) );
no02f01 g36648 ( .a(n16487), .b(n16155), .o(n40440) );
no02f01 g36649 ( .a(n40440), .b(n40439), .o(n40441) );
na02f01 g36650 ( .a(n40441), .b(n16441), .o(n40442) );
in01f01 g36651 ( .a(n40441), .o(n40443) );
na02f01 g36652 ( .a(n40443), .b(n21374), .o(n40444) );
na02f01 g36653 ( .a(n40444), .b(n40442), .o(n1070) );
na03f01 g36654 ( .a(n36762), .b(n29614), .c(n29721), .o(n40446) );
no02f01 g36655 ( .a(n39257), .b(n29639), .o(n40447) );
no02f01 g36656 ( .a(n36776), .b(n29430), .o(n40448) );
no02f01 g36657 ( .a(n40448), .b(n40447), .o(n40449) );
na03f01 g36658 ( .a(n40449), .b(n36783), .c(n40446), .o(n40450) );
no03f01 g36659 ( .a(n36794), .b(n29615), .c(n29578), .o(n40451) );
in01f01 g36660 ( .a(n36783), .o(n40452) );
in01f01 g36661 ( .a(n40449), .o(n40453) );
oa12f01 g36662 ( .a(n40453), .b(n40452), .c(n40451), .o(n40454) );
na02f01 g36663 ( .a(n40454), .b(n40450), .o(n1075) );
in01f01 g36664 ( .a(n22267), .o(n40456) );
no02f01 g36665 ( .a(n22254), .b(n22148), .o(n40457) );
ao12f01 g36666 ( .a(n40457), .b(n40456), .c(n22264), .o(n40458) );
ao12f01 g36667 ( .a(n40458), .b(n40456), .c(n22266), .o(n40459) );
in01f01 g36668 ( .a(n40459), .o(n1080) );
no03f01 g36669 ( .a(n37390), .b(n39630), .c(n37389), .o(n40461) );
ao12f01 g36670 ( .a(n37390), .b(n39630), .c(n37389), .o(n40462) );
in01f01 g36671 ( .a(n40462), .o(n40463) );
no02f01 g36672 ( .a(n40463), .b(n40461), .o(n40464) );
na03f01 g36673 ( .a(n40464), .b(n9590), .c(n9589), .o(n40465) );
in01f01 g36674 ( .a(n40464), .o(n3065) );
oa12f01 g36675 ( .a(n3065), .b(n9646), .c(n9645), .o(n40467) );
na02f01 g36676 ( .a(n40467), .b(n40465), .o(n1085) );
ao12f01 g36677 ( .a(n36483), .b(n36480), .c(n36501), .o(n40469) );
in01f01 g36678 ( .a(n40469), .o(n40470) );
no02f01 g36679 ( .a(n36482), .b(n36472), .o(n40471) );
in01f01 g36680 ( .a(n40471), .o(n40472) );
na02f01 g36681 ( .a(n40472), .b(n40470), .o(n40473) );
na02f01 g36682 ( .a(n40471), .b(n40469), .o(n40474) );
na02f01 g36683 ( .a(n40474), .b(n40473), .o(n1090) );
no02f01 g36684 ( .a(n37110), .b(n36971), .o(n40476) );
na02f01 g36685 ( .a(n40476), .b(n37182), .o(n40477) );
in01f01 g36686 ( .a(n40476), .o(n40478) );
na02f01 g36687 ( .a(n40478), .b(n37108), .o(n40479) );
na02f01 g36688 ( .a(n40479), .b(n40477), .o(n1095) );
ao12f01 g36689 ( .a(n37162), .b(n37161), .c(n37156), .o(n40481) );
in01f01 g36690 ( .a(n40481), .o(n40482) );
na03f01 g36691 ( .a(n40482), .b(n37164), .c(n36987), .o(n40483) );
oa12f01 g36692 ( .a(n40481), .b(n37016), .c(n36986), .o(n40484) );
na02f01 g36693 ( .a(n40484), .b(n40483), .o(n1100) );
no02f01 g36694 ( .a(n22436), .b(n22050), .o(n40486) );
no02f01 g36695 ( .a(n22435), .b(n21993), .o(n40487) );
no02f01 g36696 ( .a(n40487), .b(n40486), .o(n40488) );
na02f01 g36697 ( .a(n40488), .b(n22426), .o(n40489) );
in01f01 g36698 ( .a(n40488), .o(n40490) );
na02f01 g36699 ( .a(n40490), .b(n22484), .o(n40491) );
na02f01 g36700 ( .a(n40491), .b(n40489), .o(n1105) );
oa22f01 g36701 ( .a(n36659), .b(n25363), .c(n25485), .d(n25377), .o(n40493) );
na04f01 g36702 ( .a(n25486), .b(n36655), .c(n36621), .d(n25364), .o(n40494) );
na02f01 g36703 ( .a(n40494), .b(n40493), .o(n1110) );
na03f01 g36704 ( .a(n37988), .b(n37982), .c(n37973), .o(n40496) );
oa12f01 g36705 ( .a(n38039), .b(n37989), .c(n37983), .o(n40497) );
na02f01 g36706 ( .a(n40497), .b(n40496), .o(n1115) );
na04f01 g36707 ( .a(n25493), .b(n36662), .c(n36620), .d(n25344), .o(n40499) );
oa22f01 g36708 ( .a(n36665), .b(n25343), .c(n25492), .d(n25355), .o(n40500) );
na02f01 g36709 ( .a(n40500), .b(n40499), .o(n1120) );
no02f01 g36710 ( .a(n27161), .b(n26440), .o(n40502) );
no02f01 g36711 ( .a(n40502), .b(n27163), .o(n40503) );
no03f01 g36712 ( .a(n40360), .b(n40357), .c(n27167), .o(n40504) );
oa12f01 g36713 ( .a(n40503), .b(n40504), .c(n27154), .o(n40505) );
in01f01 g36714 ( .a(n27154), .o(n40506) );
in01f01 g36715 ( .a(n40503), .o(n40507) );
in01f01 g36716 ( .a(n40357), .o(n40508) );
na03f01 g36717 ( .a(n40356), .b(n40508), .c(n40354), .o(n40509) );
na03f01 g36718 ( .a(n40509), .b(n40507), .c(n40506), .o(n40510) );
na03f01 g36719 ( .a(n40510), .b(n40505), .c(n1821), .o(n40511) );
ao12f01 g36720 ( .a(n40507), .b(n40509), .c(n40506), .o(n40512) );
no03f01 g36721 ( .a(n40504), .b(n40503), .c(n27154), .o(n40513) );
oa12f01 g36722 ( .a(n8066), .b(n40513), .c(n40512), .o(n40514) );
na02f01 g36723 ( .a(n40514), .b(n40511), .o(n1125) );
no02f01 g36724 ( .a(n6056_1), .b(n5884), .o(n40516) );
na02f01 g36725 ( .a(n40516), .b(n6054), .o(n40517) );
no02f01 g36726 ( .a(n6052), .b(n34411), .o(n40518) );
in01f01 g36727 ( .a(n40516), .o(n40519) );
oa12f01 g36728 ( .a(n40519), .b(n40518), .c(n5896), .o(n40520) );
na02f01 g36729 ( .a(n40520), .b(n40517), .o(n1130) );
in01f01 g36730 ( .a(n9659), .o(n40522) );
oa12f01 g36731 ( .a(n9892), .b(n9873), .c(n39648), .o(n40523) );
na02f01 g36732 ( .a(n40523), .b(n5001), .o(n40524) );
na02f01 g36733 ( .a(n9899), .b(n40523), .o(n40525) );
ao22f01 g36734 ( .a(n40525), .b(n6934), .c(n40524), .d(n40522), .o(n1135) );
in01f01 g36735 ( .a(n27600), .o(n40527) );
no02f01 g36736 ( .a(n27598), .b(n27367), .o(n40528) );
in01f01 g36737 ( .a(n40528), .o(n40529) );
na02f01 g36738 ( .a(n40529), .b(n27633), .o(n40530) );
ao12f01 g36739 ( .a(n40530), .b(n40527), .c(n27588), .o(n40531) );
no02f01 g36740 ( .a(n27609), .b(n27367), .o(n40532) );
no02f01 g36741 ( .a(n40532), .b(n27611), .o(n40533) );
na02f01 g36742 ( .a(n40533), .b(n40531), .o(n40534) );
in01f01 g36743 ( .a(n40531), .o(n40535) );
in01f01 g36744 ( .a(n40533), .o(n40536) );
na02f01 g36745 ( .a(n40536), .b(n40535), .o(n40537) );
na02f01 g36746 ( .a(n40537), .b(n40534), .o(n1140) );
no02f01 g36747 ( .a(n10896), .b(n3521), .o(n40539) );
no02f01 g36748 ( .a(n40539), .b(n10898), .o(n40540) );
in01f01 g36749 ( .a(n40540), .o(n40541) );
na02f01 g36750 ( .a(n40541), .b(n25630), .o(n40542) );
na02f01 g36751 ( .a(n40540), .b(n25629), .o(n40543) );
na02f01 g36752 ( .a(n40543), .b(n40542), .o(n1145) );
ao12f01 g36753 ( .a(n25527), .b(n25531), .c(n39820), .o(n40545) );
in01f01 g36754 ( .a(n40545), .o(n40546) );
no02f01 g36755 ( .a(n25530), .b(n25322), .o(n40547) );
no02f01 g36756 ( .a(n40547), .b(n40546), .o(n40548) );
na02f01 g36757 ( .a(n40547), .b(n40546), .o(n40549) );
in01f01 g36758 ( .a(n40549), .o(n40550) );
no02f01 g36759 ( .a(n40550), .b(n40548), .o(n40551) );
in01f01 g36760 ( .a(n40551), .o(n1150) );
oa12f01 g36761 ( .a(n25835), .b(n25829), .c(n25828), .o(n40553) );
na02f01 g36762 ( .a(n25834), .b(n25830), .o(n40554) );
na02f01 g36763 ( .a(n40554), .b(n40553), .o(n1155) );
no02f01 g36764 ( .a(n9591), .b(n936), .o(n40556) );
no02f01 g36765 ( .a(n4201), .b(n9228), .o(n40557) );
no02f01 g36766 ( .a(n40557), .b(n40556), .o(n3707) );
na03f01 g36767 ( .a(n3707), .b(n9590), .c(n9589), .o(n40559) );
in01f01 g36768 ( .a(n3707), .o(n5716) );
oa12f01 g36769 ( .a(n5716), .b(n9646), .c(n9645), .o(n40561) );
na02f01 g36770 ( .a(n40561), .b(n40559), .o(n1160) );
in01f01 g36771 ( .a(n28973), .o(n40563) );
no02f01 g36772 ( .a(n39861), .b(n40563), .o(n40564) );
in01f01 g36773 ( .a(n28982), .o(n40565) );
no02f01 g36774 ( .a(n39861), .b(n40565), .o(n40566) );
no02f01 g36775 ( .a(n40566), .b(n40564), .o(n40567) );
no02f01 g36776 ( .a(n40565), .b(n40563), .o(n40568) );
no02f01 g36777 ( .a(n40568), .b(n39860), .o(n40569) );
in01f01 g36778 ( .a(n40569), .o(n40570) );
no02f01 g36779 ( .a(n28956), .b(n28954), .o(n40571) );
in01f01 g36780 ( .a(n40571), .o(n40572) );
no02f01 g36781 ( .a(n39861), .b(n40572), .o(n40573) );
in01f01 g36782 ( .a(n40573), .o(n40574) );
no02f01 g36783 ( .a(n39981), .b(n39862), .o(n40575) );
na02f01 g36784 ( .a(n40575), .b(n40574), .o(n40576) );
in01f01 g36785 ( .a(n40576), .o(n40577) );
na04f01 g36786 ( .a(n40577), .b(n39980), .c(n39969), .d(n39945), .o(n40578) );
ao12f01 g36787 ( .a(n39860), .b(n40571), .c(n28944), .o(n40579) );
no02f01 g36788 ( .a(n40579), .b(n39985), .o(n40580) );
na02f01 g36789 ( .a(n40580), .b(n39994), .o(n40581) );
in01f01 g36790 ( .a(n40581), .o(n40582) );
na03f01 g36791 ( .a(n40582), .b(n40578), .c(n40570), .o(n40583) );
in01f01 g36792 ( .a(n28833), .o(n40584) );
no02f01 g36793 ( .a(n39861), .b(n40584), .o(n40585) );
no02f01 g36794 ( .a(n39860), .b(n28833), .o(n40586) );
no02f01 g36795 ( .a(n40586), .b(n40585), .o(n40587) );
in01f01 g36796 ( .a(n40587), .o(n40588) );
na03f01 g36797 ( .a(n40588), .b(n40583), .c(n40567), .o(n40589) );
in01f01 g36798 ( .a(n40567), .o(n40590) );
no04f01 g36799 ( .a(n40576), .b(n39979), .c(n40048), .d(n40047), .o(n40591) );
no03f01 g36800 ( .a(n40581), .b(n40591), .c(n40569), .o(n40592) );
oa12f01 g36801 ( .a(n40587), .b(n40592), .c(n40590), .o(n40593) );
na03f01 g36802 ( .a(n40593), .b(n40589), .c(n_27923), .o(n40594) );
no03f01 g36803 ( .a(n40587), .b(n40592), .c(n40590), .o(n40595) );
ao12f01 g36804 ( .a(n40588), .b(n40583), .c(n40567), .o(n40596) );
oa12f01 g36805 ( .a(n34420), .b(n40596), .c(n40595), .o(n40597) );
na02f01 g36806 ( .a(n40597), .b(n40594), .o(n1165) );
no02f01 g36807 ( .a(n37384), .b(n9596), .o(n40599) );
no02f01 g36808 ( .a(n40599), .b(n38168), .o(n40600) );
na02f01 g36809 ( .a(n40599), .b(n38168), .o(n40601) );
in01f01 g36810 ( .a(n40601), .o(n40602) );
no02f01 g36811 ( .a(n40602), .b(n40600), .o(n40603) );
na03f01 g36812 ( .a(n40603), .b(n9590), .c(n9589), .o(n40604) );
in01f01 g36813 ( .a(n40603), .o(n3287) );
oa12f01 g36814 ( .a(n3287), .b(n9646), .c(n9645), .o(n40606) );
na02f01 g36815 ( .a(n40606), .b(n40604), .o(n1170) );
na02f01 g36816 ( .a(n11866), .b(n11860), .o(n40608) );
no02f01 g36817 ( .a(n11867), .b(n11526), .o(n40609) );
na03f01 g36818 ( .a(n40609), .b(n40608), .c(n11861), .o(n40610) );
na02f01 g36819 ( .a(n40608), .b(n11861), .o(n40611) );
in01f01 g36820 ( .a(n40609), .o(n40612) );
na02f01 g36821 ( .a(n40612), .b(n40611), .o(n40613) );
na02f01 g36822 ( .a(n40613), .b(n40610), .o(n1175) );
na02f01 g36823 ( .a(n29366), .b(n29365), .o(n40615) );
na02f01 g36824 ( .a(n29370), .b(n40615), .o(n40616) );
na02f01 g36825 ( .a(n40616), .b(n29372), .o(n1180) );
ao12f01 g36826 ( .a(n21279), .b(n21274), .c(n21278), .o(n40618) );
in01f01 g36827 ( .a(n40618), .o(n40619) );
no02f01 g36828 ( .a(n40619), .b(n18868), .o(n40620) );
no02f01 g36829 ( .a(n40618), .b(n19114), .o(n40621) );
no02f01 g36830 ( .a(n40621), .b(n40620), .o(n40622) );
in01f01 g36831 ( .a(n40622), .o(n40623) );
no02f01 g36832 ( .a(n40618), .b(n19068), .o(n40624) );
in01f01 g36833 ( .a(n40624), .o(n40625) );
oa12f01 g36834 ( .a(n21295), .b(n21292), .c(n21284), .o(n40626) );
no02f01 g36835 ( .a(n40619), .b(n19067), .o(n40627) );
oa12f01 g36836 ( .a(n40625), .b(n40627), .c(n40626), .o(n40628) );
no02f01 g36837 ( .a(n40619), .b(n19074), .o(n40629) );
in01f01 g36838 ( .a(n40629), .o(n40630) );
na03f01 g36839 ( .a(n40630), .b(n40628), .c(n19108), .o(n40631) );
oa12f01 g36840 ( .a(n40619), .b(n40628), .c(n19108), .o(n40632) );
na02f01 g36841 ( .a(n40619), .b(n19074), .o(n40633) );
ao12f01 g36842 ( .a(n40618), .b(n19106), .c(n19102), .o(n40634) );
in01f01 g36843 ( .a(n40634), .o(n40635) );
na04f01 g36844 ( .a(n40635), .b(n40633), .c(n40632), .d(n40631), .o(n40636) );
in01f01 g36845 ( .a(n18896), .o(n40637) );
ao12f01 g36846 ( .a(n21288), .b(n21299), .c(n21294), .o(n40638) );
in01f01 g36847 ( .a(n40627), .o(n40639) );
ao12f01 g36848 ( .a(n40624), .b(n40639), .c(n40638), .o(n40640) );
no03f01 g36849 ( .a(n40629), .b(n40640), .c(n19090), .o(n40641) );
ao12f01 g36850 ( .a(n40618), .b(n40640), .c(n19090), .o(n40642) );
in01f01 g36851 ( .a(n40633), .o(n40643) );
no04f01 g36852 ( .a(n40634), .b(n40643), .c(n40642), .d(n40641), .o(n40644) );
ao12f01 g36853 ( .a(n40619), .b(n19096), .c(n18882), .o(n40645) );
no03f01 g36854 ( .a(n40645), .b(n40644), .c(n40637), .o(n40646) );
oa22f01 g36855 ( .a(n40646), .b(n40619), .c(n40636), .d(n18896), .o(n40647) );
no02f01 g36856 ( .a(n40647), .b(n40623), .o(n40648) );
in01f01 g36857 ( .a(n40645), .o(n40649) );
na03f01 g36858 ( .a(n40649), .b(n40636), .c(n18896), .o(n40650) );
ao22f01 g36859 ( .a(n40650), .b(n40618), .c(n40644), .d(n40637), .o(n40651) );
no02f01 g36860 ( .a(n40651), .b(n40622), .o(n40652) );
oa12f01 g36861 ( .a(n18460), .b(n40652), .c(n40648), .o(n40653) );
no02f01 g36862 ( .a(n40618), .b(n19106), .o(n40654) );
in01f01 g36863 ( .a(n40654), .o(n40655) );
na04f01 g36864 ( .a(n40655), .b(n40633), .c(n40632), .d(n40631), .o(n40656) );
no02f01 g36865 ( .a(n40619), .b(n19096), .o(n40657) );
in01f01 g36866 ( .a(n40657), .o(n40658) );
no02f01 g36867 ( .a(n40619), .b(n18882), .o(n40659) );
no02f01 g36868 ( .a(n40618), .b(n19102), .o(n40660) );
no02f01 g36869 ( .a(n40660), .b(n40659), .o(n40661) );
na03f01 g36870 ( .a(n40661), .b(n40658), .c(n40656), .o(n40662) );
no04f01 g36871 ( .a(n40654), .b(n40643), .c(n40642), .d(n40641), .o(n40663) );
in01f01 g36872 ( .a(n40661), .o(n40664) );
oa12f01 g36873 ( .a(n40664), .b(n40657), .c(n40663), .o(n40665) );
ao12f01 g36874 ( .a(n18459), .b(n40665), .c(n40662), .o(n40666) );
na02f01 g36875 ( .a(n21298), .b(n21297), .o(n40667) );
na03f01 g36876 ( .a(n40667), .b(n21294), .c(n20547), .o(n40668) );
na03f01 g36877 ( .a(n40639), .b(n40668), .c(n21295), .o(n40669) );
ao12f01 g36878 ( .a(n40629), .b(n40669), .c(n40625), .o(n40670) );
no02f01 g36879 ( .a(n40618), .b(n19090), .o(n40671) );
no02f01 g36880 ( .a(n40619), .b(n19108), .o(n40672) );
no02f01 g36881 ( .a(n40672), .b(n40671), .o(n40673) );
oa12f01 g36882 ( .a(n40673), .b(n40643), .c(n40670), .o(n40674) );
no02f01 g36883 ( .a(n21291), .b(n21290), .o(n40675) );
no03f01 g36884 ( .a(n40675), .b(n21284), .c(n20789), .o(n40676) );
no03f01 g36885 ( .a(n40627), .b(n40676), .c(n21288), .o(n40677) );
oa12f01 g36886 ( .a(n40630), .b(n40677), .c(n40624), .o(n40678) );
in01f01 g36887 ( .a(n40673), .o(n40679) );
na03f01 g36888 ( .a(n40679), .b(n40633), .c(n40678), .o(n40680) );
na02f01 g36889 ( .a(n40680), .b(n40674), .o(n40681) );
no02f01 g36890 ( .a(n40643), .b(n40629), .o(n40682) );
no02f01 g36891 ( .a(n40682), .b(n40628), .o(n40683) );
in01f01 g36892 ( .a(n40682), .o(n40684) );
no02f01 g36893 ( .a(n40684), .b(n40640), .o(n40685) );
oa12f01 g36894 ( .a(n18460), .b(n40685), .c(n40683), .o(n40686) );
no02f01 g36895 ( .a(n40627), .b(n40624), .o(n40687) );
na02f01 g36896 ( .a(n40687), .b(n40638), .o(n40688) );
in01f01 g36897 ( .a(n40687), .o(n40689) );
na02f01 g36898 ( .a(n40689), .b(n40626), .o(n40690) );
ao12f01 g36899 ( .a(n18459), .b(n40690), .c(n40688), .o(n40691) );
no02f01 g36900 ( .a(n20867), .b(n18459), .o(n40692) );
oa12f01 g36901 ( .a(n18460), .b(n20885), .c(n20882), .o(n40693) );
oa12f01 g36902 ( .a(n18460), .b(n21316), .c(n21315), .o(n40694) );
no03f01 g36903 ( .a(n40187), .b(n40184), .c(n40106), .o(n40695) );
na03f01 g36904 ( .a(n40695), .b(n40694), .c(n40693), .o(n40696) );
no02f01 g36905 ( .a(n40696), .b(n40692), .o(n40697) );
oa12f01 g36906 ( .a(n18459), .b(n20866), .c(n20787), .o(n40698) );
na02f01 g36907 ( .a(n20929), .b(n18459), .o(n40699) );
oa12f01 g36908 ( .a(n18459), .b(n20919), .c(n20903), .o(n40700) );
na03f01 g36909 ( .a(n40700), .b(n40699), .c(n40698), .o(n40701) );
no02f01 g36910 ( .a(n40701), .b(n40697), .o(n40702) );
no02f01 g36911 ( .a(n21301), .b(n18459), .o(n40703) );
no03f01 g36912 ( .a(n40703), .b(n40702), .c(n40691), .o(n40704) );
na02f01 g36913 ( .a(n40704), .b(n40686), .o(n40705) );
ao12f01 g36914 ( .a(n40705), .b(n40681), .c(n18460), .o(n40706) );
ao12f01 g36915 ( .a(n40679), .b(n40633), .c(n40678), .o(n40707) );
no03f01 g36916 ( .a(n40673), .b(n40643), .c(n40670), .o(n40708) );
no02f01 g36917 ( .a(n40708), .b(n40707), .o(n40709) );
na02f01 g36918 ( .a(n40684), .b(n40640), .o(n40710) );
na02f01 g36919 ( .a(n40682), .b(n40628), .o(n40711) );
na02f01 g36920 ( .a(n40711), .b(n40710), .o(n40712) );
no02f01 g36921 ( .a(n40689), .b(n40626), .o(n40713) );
no02f01 g36922 ( .a(n40687), .b(n40638), .o(n40714) );
no02f01 g36923 ( .a(n40714), .b(n40713), .o(n40715) );
ao12f01 g36924 ( .a(n18460), .b(n40715), .c(n21301), .o(n40716) );
ao12f01 g36925 ( .a(n40716), .b(n40712), .c(n18459), .o(n40717) );
oa12f01 g36926 ( .a(n40717), .b(n40709), .c(n18460), .o(n40718) );
no02f01 g36927 ( .a(n40657), .b(n40654), .o(n40719) );
in01f01 g36928 ( .a(n40719), .o(n40720) );
na04f01 g36929 ( .a(n40720), .b(n40633), .c(n40632), .d(n40631), .o(n40721) );
in01f01 g36930 ( .a(n40721), .o(n40722) );
no03f01 g36931 ( .a(n40643), .b(n40642), .c(n40641), .o(n40723) );
no02f01 g36932 ( .a(n40720), .b(n40723), .o(n40724) );
no02f01 g36933 ( .a(n40724), .b(n40722), .o(n40725) );
oa22f01 g36934 ( .a(n40725), .b(n18459), .c(n40718), .d(n40706), .o(n40726) );
no02f01 g36935 ( .a(n40726), .b(n40666), .o(n40727) );
na02f01 g36936 ( .a(n40649), .b(n40636), .o(n40728) );
no02f01 g36937 ( .a(n40619), .b(n18896), .o(n40729) );
no02f01 g36938 ( .a(n40618), .b(n40637), .o(n40730) );
no02f01 g36939 ( .a(n40730), .b(n40729), .o(n40731) );
in01f01 g36940 ( .a(n40731), .o(n40732) );
na02f01 g36941 ( .a(n40732), .b(n40728), .o(n40733) );
no02f01 g36942 ( .a(n40645), .b(n40644), .o(n40734) );
na02f01 g36943 ( .a(n40731), .b(n40734), .o(n40735) );
na02f01 g36944 ( .a(n40735), .b(n40733), .o(n40736) );
na02f01 g36945 ( .a(n40736), .b(n18460), .o(n40737) );
na03f01 g36946 ( .a(n40737), .b(n40727), .c(n40653), .o(n40738) );
na02f01 g36947 ( .a(n40651), .b(n40622), .o(n40739) );
na02f01 g36948 ( .a(n40647), .b(n40623), .o(n40740) );
ao12f01 g36949 ( .a(n18460), .b(n40740), .c(n40739), .o(n40741) );
no03f01 g36950 ( .a(n40664), .b(n40657), .c(n40663), .o(n40742) );
ao12f01 g36951 ( .a(n40661), .b(n40658), .c(n40656), .o(n40743) );
no02f01 g36952 ( .a(n40743), .b(n40742), .o(n40744) );
ao12f01 g36953 ( .a(n18460), .b(n40725), .c(n40744), .o(n40745) );
no02f01 g36954 ( .a(n40731), .b(n40734), .o(n40746) );
no02f01 g36955 ( .a(n40732), .b(n40728), .o(n40747) );
no02f01 g36956 ( .a(n40747), .b(n40746), .o(n40748) );
no02f01 g36957 ( .a(n40748), .b(n18460), .o(n40749) );
no03f01 g36958 ( .a(n40749), .b(n40745), .c(n40741), .o(n40750) );
na02f01 g36959 ( .a(n40750), .b(n40738), .o(n40751) );
oa12f01 g36960 ( .a(n18459), .b(n40652), .c(n40648), .o(n40752) );
na02f01 g36961 ( .a(n40752), .b(n40653), .o(n40753) );
no02f01 g36962 ( .a(n40753), .b(n40751), .o(n40754) );
ao12f01 g36963 ( .a(n18459), .b(n40740), .c(n40739), .o(n40755) );
oa12f01 g36964 ( .a(n18460), .b(n40743), .c(n40742), .o(n40756) );
ao12f01 g36965 ( .a(n18459), .b(n40711), .c(n40710), .o(n40757) );
oa12f01 g36966 ( .a(n18460), .b(n40714), .c(n40713), .o(n40758) );
oa12f01 g36967 ( .a(n20790), .b(n20865), .c(n20791), .o(n40759) );
na03f01 g36968 ( .a(n20786), .b(n20553), .c(n20548), .o(n40760) );
ao12f01 g36969 ( .a(n18460), .b(n40760), .c(n40759), .o(n40761) );
no02f01 g36970 ( .a(n20886), .b(n18460), .o(n40762) );
ao12f01 g36971 ( .a(n18460), .b(n21323), .c(n21317), .o(n40763) );
no03f01 g36972 ( .a(n40763), .b(n40762), .c(n40761), .o(n40764) );
oa12f01 g36973 ( .a(n40764), .b(n40696), .c(n40692), .o(n40765) );
na02f01 g36974 ( .a(n21308), .b(n18460), .o(n40766) );
na03f01 g36975 ( .a(n40766), .b(n40765), .c(n40758), .o(n40767) );
no02f01 g36976 ( .a(n40767), .b(n40757), .o(n40768) );
oa12f01 g36977 ( .a(n40768), .b(n40709), .c(n18459), .o(n40769) );
no02f01 g36978 ( .a(n40685), .b(n40683), .o(n40770) );
na02f01 g36979 ( .a(n40690), .b(n40688), .o(n40771) );
no02f01 g36980 ( .a(n21301), .b(n18460), .o(n40772) );
ao12f01 g36981 ( .a(n40772), .b(n40771), .c(n18459), .o(n40773) );
oa12f01 g36982 ( .a(n40773), .b(n40770), .c(n18460), .o(n40774) );
ao12f01 g36983 ( .a(n40774), .b(n40681), .c(n18459), .o(n40775) );
no03f01 g36984 ( .a(n40677), .b(n40624), .c(n19108), .o(n40776) );
oa12f01 g36985 ( .a(n40633), .b(n40776), .c(n40618), .o(n40777) );
oa12f01 g36986 ( .a(n40719), .b(n40777), .c(n40641), .o(n40778) );
na02f01 g36987 ( .a(n40778), .b(n40721), .o(n40779) );
ao22f01 g36988 ( .a(n40779), .b(n18460), .c(n40775), .d(n40769), .o(n40780) );
na02f01 g36989 ( .a(n40780), .b(n40756), .o(n40781) );
no02f01 g36990 ( .a(n40748), .b(n18459), .o(n40782) );
no03f01 g36991 ( .a(n40782), .b(n40781), .c(n40755), .o(n40783) );
na02f01 g36992 ( .a(n40665), .b(n40662), .o(n40784) );
oa12f01 g36993 ( .a(n18459), .b(n40779), .c(n40784), .o(n40785) );
na02f01 g36994 ( .a(n40736), .b(n18459), .o(n40786) );
na03f01 g36995 ( .a(n40786), .b(n40785), .c(n40752), .o(n40787) );
no02f01 g36996 ( .a(n40787), .b(n40783), .o(n40788) );
no02f01 g36997 ( .a(n40741), .b(n40755), .o(n40789) );
no02f01 g36998 ( .a(n40789), .b(n40788), .o(n40790) );
no02f01 g36999 ( .a(n40790), .b(n40754), .o(n40791) );
no02f01 g37000 ( .a(n40791), .b(n20164), .o(n40792) );
in01f01 g37001 ( .a(n20164), .o(n40793) );
in01f01 g37002 ( .a(n40791), .o(n40794) );
no02f01 g37003 ( .a(n40794), .b(n40793), .o(n40795) );
no02f01 g37004 ( .a(n40795), .b(n40792), .o(n40796) );
na03f01 g37005 ( .a(n40786), .b(n40785), .c(n40781), .o(n40797) );
na02f01 g37006 ( .a(n40797), .b(n40737), .o(n40798) );
no02f01 g37007 ( .a(n40798), .b(n40789), .o(n40799) );
ao12f01 g37008 ( .a(n40753), .b(n40797), .c(n40737), .o(n40800) );
no03f01 g37009 ( .a(n40800), .b(n40799), .c(n20300), .o(n40801) );
no02f01 g37010 ( .a(n20311), .b(n20310), .o(n40802) );
in01f01 g37011 ( .a(n40802), .o(n40803) );
no02f01 g37012 ( .a(n40745), .b(n40727), .o(n40804) );
no02f01 g37013 ( .a(n40749), .b(n40782), .o(n40805) );
no02f01 g37014 ( .a(n40805), .b(n40804), .o(n40806) );
na02f01 g37015 ( .a(n40785), .b(n40781), .o(n40807) );
na02f01 g37016 ( .a(n40786), .b(n40737), .o(n40808) );
no02f01 g37017 ( .a(n40808), .b(n40807), .o(n40809) );
no03f01 g37018 ( .a(n40809), .b(n40806), .c(n40803), .o(n40810) );
no02f01 g37019 ( .a(n40744), .b(n18460), .o(n40811) );
no02f01 g37020 ( .a(n40725), .b(n18460), .o(n40812) );
no04f01 g37021 ( .a(n40812), .b(n40811), .c(n40780), .d(n40666), .o(n40813) );
na02f01 g37022 ( .a(n40784), .b(n18459), .o(n40814) );
in01f01 g37023 ( .a(n40812), .o(n40815) );
ao22f01 g37024 ( .a(n40815), .b(n40726), .c(n40814), .d(n40756), .o(n40816) );
no03f01 g37025 ( .a(n40816), .b(n40813), .c(n20303), .o(n40817) );
na04f01 g37026 ( .a(n40815), .b(n40814), .c(n40726), .d(n40756), .o(n40818) );
oa22f01 g37027 ( .a(n40812), .b(n40780), .c(n40811), .d(n40666), .o(n40819) );
ao12f01 g37028 ( .a(n20179), .b(n40819), .c(n40818), .o(n40820) );
no02f01 g37029 ( .a(n40718), .b(n40706), .o(n40821) );
in01f01 g37030 ( .a(n40821), .o(n40822) );
no02f01 g37031 ( .a(n40725), .b(n18459), .o(n40823) );
oa12f01 g37032 ( .a(n40822), .b(n40812), .c(n40823), .o(n40824) );
no02f01 g37033 ( .a(n40812), .b(n40823), .o(n40825) );
na02f01 g37034 ( .a(n40825), .b(n40821), .o(n40826) );
ao12f01 g37035 ( .a(n20307), .b(n40826), .c(n40824), .o(n40827) );
no02f01 g37036 ( .a(n40827), .b(n40820), .o(n40828) );
no03f01 g37037 ( .a(n40828), .b(n40817), .c(n40810), .o(n40829) );
na03f01 g37038 ( .a(n40797), .b(n40753), .c(n40737), .o(n40830) );
na02f01 g37039 ( .a(n40798), .b(n40789), .o(n40831) );
ao12f01 g37040 ( .a(n20172), .b(n40831), .c(n40830), .o(n40832) );
na02f01 g37041 ( .a(n40808), .b(n40807), .o(n40833) );
na02f01 g37042 ( .a(n40805), .b(n40804), .o(n40834) );
ao12f01 g37043 ( .a(n40802), .b(n40834), .c(n40833), .o(n40835) );
no03f01 g37044 ( .a(n40835), .b(n40832), .c(n40829), .o(n40836) );
no02f01 g37045 ( .a(n40836), .b(n40801), .o(n40837) );
na03f01 g37046 ( .a(n40831), .b(n40830), .c(n20172), .o(n40838) );
no02f01 g37047 ( .a(n40825), .b(n40821), .o(n40839) );
no03f01 g37048 ( .a(n40812), .b(n40823), .c(n40822), .o(n40840) );
no02f01 g37049 ( .a(n40840), .b(n40839), .o(n40841) );
na02f01 g37050 ( .a(n40841), .b(n20307), .o(n40842) );
in01f01 g37051 ( .a(n40842), .o(n40843) );
no03f01 g37052 ( .a(n40843), .b(n40817), .c(n40810), .o(n40844) );
na02f01 g37053 ( .a(n40844), .b(n40838), .o(n40845) );
no02f01 g37054 ( .a(n40709), .b(n18459), .o(n40846) );
no02f01 g37055 ( .a(n40709), .b(n18460), .o(n40847) );
no02f01 g37056 ( .a(n40847), .b(n40846), .o(n40848) );
no02f01 g37057 ( .a(n40774), .b(n40768), .o(n40849) );
na02f01 g37058 ( .a(n40849), .b(n40848), .o(n40850) );
in01f01 g37059 ( .a(n40850), .o(n40851) );
no02f01 g37060 ( .a(n40849), .b(n40848), .o(n40852) );
no02f01 g37061 ( .a(n40852), .b(n40851), .o(n40853) );
na02f01 g37062 ( .a(n40853), .b(n20185), .o(n40854) );
in01f01 g37063 ( .a(n40854), .o(n40855) );
in01f01 g37064 ( .a(n20185), .o(n40856) );
oa12f01 g37065 ( .a(n40856), .b(n40852), .c(n40851), .o(n40857) );
no02f01 g37066 ( .a(n20191), .b(n20189), .o(n40858) );
no02f01 g37067 ( .a(n40770), .b(n18460), .o(n40859) );
no02f01 g37068 ( .a(n40859), .b(n40757), .o(n40860) );
ao12f01 g37069 ( .a(n40860), .b(n40773), .c(n40767), .o(n40861) );
no04f01 g37070 ( .a(n40716), .b(n40859), .c(n40704), .d(n40757), .o(n40862) );
no02f01 g37071 ( .a(n40862), .b(n40861), .o(n40863) );
na02f01 g37072 ( .a(n40863), .b(n40858), .o(n40864) );
no02f01 g37073 ( .a(n20274), .b(n20272), .o(n40865) );
in01f01 g37074 ( .a(n40865), .o(n40866) );
no02f01 g37075 ( .a(n40715), .b(n18460), .o(n40867) );
no02f01 g37076 ( .a(n40867), .b(n40691), .o(n40868) );
ao12f01 g37077 ( .a(n40772), .b(n40766), .c(n40765), .o(n40869) );
na02f01 g37078 ( .a(n40869), .b(n40868), .o(n40870) );
in01f01 g37079 ( .a(n40870), .o(n40871) );
no02f01 g37080 ( .a(n40869), .b(n40868), .o(n40872) );
no02f01 g37081 ( .a(n40872), .b(n40871), .o(n40873) );
in01f01 g37082 ( .a(n40873), .o(n40874) );
no02f01 g37083 ( .a(n40874), .b(n40866), .o(n40875) );
na02f01 g37084 ( .a(n40874), .b(n40866), .o(n40876) );
no02f01 g37085 ( .a(n40772), .b(n40703), .o(n40877) );
no02f01 g37086 ( .a(n40877), .b(n40702), .o(n40878) );
na02f01 g37087 ( .a(n40877), .b(n40702), .o(n40879) );
in01f01 g37088 ( .a(n40879), .o(n40880) );
no02f01 g37089 ( .a(n40880), .b(n40878), .o(n40881) );
no02f01 g37090 ( .a(n40881), .b(n20266), .o(n40882) );
in01f01 g37091 ( .a(n40882), .o(n40883) );
ao12f01 g37092 ( .a(n40875), .b(n40883), .c(n40876), .o(n40884) );
no02f01 g37093 ( .a(n40863), .b(n40858), .o(n40885) );
ao12f01 g37094 ( .a(n40885), .b(n40884), .c(n40864), .o(n40886) );
ao12f01 g37095 ( .a(n40855), .b(n40886), .c(n40857), .o(n40887) );
in01f01 g37096 ( .a(n40887), .o(n40888) );
no02f01 g37097 ( .a(n40761), .b(n40692), .o(n40889) );
ao12f01 g37098 ( .a(n40763), .b(n40695), .c(n40694), .o(n40890) );
na02f01 g37099 ( .a(n40890), .b(n40699), .o(n40891) );
na02f01 g37100 ( .a(n40891), .b(n40693), .o(n40892) );
na02f01 g37101 ( .a(n40892), .b(n40889), .o(n40893) );
no02f01 g37102 ( .a(n40892), .b(n40889), .o(n40894) );
in01f01 g37103 ( .a(n40894), .o(n40895) );
na02f01 g37104 ( .a(n40895), .b(n40893), .o(n40896) );
no02f01 g37105 ( .a(n40896), .b(n20377), .o(n40897) );
in01f01 g37106 ( .a(n40897), .o(n40898) );
in01f01 g37107 ( .a(n20247), .o(n40899) );
in01f01 g37108 ( .a(n40186), .o(n40900) );
ao12f01 g37109 ( .a(n40187), .b(n40900), .c(n40189), .o(n40901) );
in01f01 g37110 ( .a(n40901), .o(n40902) );
no02f01 g37111 ( .a(n21317), .b(n18460), .o(n40903) );
in01f01 g37112 ( .a(n40903), .o(n40904) );
na02f01 g37113 ( .a(n40904), .b(n40694), .o(n40905) );
in01f01 g37114 ( .a(n40905), .o(n40906) );
no02f01 g37115 ( .a(n40906), .b(n40902), .o(n40907) );
no02f01 g37116 ( .a(n40905), .b(n40901), .o(n40908) );
no02f01 g37117 ( .a(n40908), .b(n40907), .o(n40909) );
in01f01 g37118 ( .a(n40909), .o(n40910) );
no02f01 g37119 ( .a(n40910), .b(n40899), .o(n40911) );
in01f01 g37120 ( .a(n40911), .o(n40912) );
in01f01 g37121 ( .a(n40193), .o(n40913) );
oa12f01 g37122 ( .a(n40913), .b(n40195), .c(n40183), .o(n40914) );
no02f01 g37123 ( .a(n40909), .b(n20247), .o(n40915) );
oa12f01 g37124 ( .a(n40912), .b(n40915), .c(n40914), .o(n40916) );
na02f01 g37125 ( .a(n40699), .b(n40693), .o(n40917) );
in01f01 g37126 ( .a(n40917), .o(n40918) );
no02f01 g37127 ( .a(n40918), .b(n40890), .o(n40919) );
na02f01 g37128 ( .a(n40918), .b(n40890), .o(n40920) );
in01f01 g37129 ( .a(n40920), .o(n40921) );
no02f01 g37130 ( .a(n40921), .b(n40919), .o(n40922) );
in01f01 g37131 ( .a(n40922), .o(n40923) );
no02f01 g37132 ( .a(n40923), .b(n20391), .o(n40924) );
ao12f01 g37133 ( .a(n20199), .b(n40895), .c(n40893), .o(n40925) );
no02f01 g37134 ( .a(n40922), .b(n20255), .o(n40926) );
no02f01 g37135 ( .a(n40926), .b(n40925), .o(n40927) );
oa12f01 g37136 ( .a(n40927), .b(n40924), .c(n40916), .o(n40928) );
na02f01 g37137 ( .a(n40928), .b(n40898), .o(n40929) );
na02f01 g37138 ( .a(n40881), .b(n20266), .o(n40930) );
in01f01 g37139 ( .a(n40930), .o(n40931) );
na02f01 g37140 ( .a(n40864), .b(n40854), .o(n40932) );
no04f01 g37141 ( .a(n40932), .b(n40931), .c(n40929), .d(n40875), .o(n40933) );
in01f01 g37142 ( .a(n40933), .o(n40934) );
ao12f01 g37143 ( .a(n40845), .b(n40934), .c(n40888), .o(n40935) );
no02f01 g37144 ( .a(n40935), .b(n40837), .o(n40936) );
na02f01 g37145 ( .a(n40936), .b(n40796), .o(n40937) );
na03f01 g37146 ( .a(n40834), .b(n40833), .c(n40802), .o(n40938) );
in01f01 g37147 ( .a(n40817), .o(n40939) );
no02f01 g37148 ( .a(n40816), .b(n40813), .o(n40940) );
oa22f01 g37149 ( .a(n40841), .b(n20307), .c(n40940), .d(n20179), .o(n40941) );
na03f01 g37150 ( .a(n40941), .b(n40939), .c(n40938), .o(n40942) );
oa12f01 g37151 ( .a(n20300), .b(n40800), .c(n40799), .o(n40943) );
in01f01 g37152 ( .a(n40835), .o(n40944) );
na03f01 g37153 ( .a(n40944), .b(n40943), .c(n40942), .o(n40945) );
na02f01 g37154 ( .a(n40945), .b(n40838), .o(n40946) );
na03f01 g37155 ( .a(n40842), .b(n40939), .c(n40938), .o(n40947) );
no02f01 g37156 ( .a(n40947), .b(n40801), .o(n40948) );
oa12f01 g37157 ( .a(n40948), .b(n40933), .c(n40887), .o(n40949) );
na02f01 g37158 ( .a(n40949), .b(n40946), .o(n40950) );
oa12f01 g37159 ( .a(n40950), .b(n40795), .c(n40792), .o(n40951) );
na03f01 g37160 ( .a(n40951), .b(n40937), .c(n5799), .o(n40952) );
na02f01 g37161 ( .a(n40951), .b(n40937), .o(n5195) );
na02f01 g37162 ( .a(n5195), .b(n911), .o(n40954) );
na02f01 g37163 ( .a(n40954), .b(n40952), .o(n1185) );
no02f01 g37164 ( .a(n6042_1), .b(n5873), .o(n40956) );
in01f01 g37165 ( .a(n40956), .o(n40957) );
ao12f01 g37166 ( .a(n6047_1), .b(n6025), .c(n6008), .o(n40958) );
ao12f01 g37167 ( .a(n6044), .b(n40958), .c(n40957), .o(n40959) );
in01f01 g37168 ( .a(n40959), .o(n40960) );
no02f01 g37169 ( .a(n6034), .b(n5873), .o(n40961) );
no02f01 g37170 ( .a(n40961), .b(n6036), .o(n40962) );
na02f01 g37171 ( .a(n40962), .b(n40960), .o(n40963) );
in01f01 g37172 ( .a(n40962), .o(n40964) );
na02f01 g37173 ( .a(n40964), .b(n40959), .o(n40965) );
na02f01 g37174 ( .a(n40965), .b(n40963), .o(n1190) );
no03f01 g37175 ( .a(n37386), .b(n37383), .c(n9591), .o(n40967) );
no02f01 g37176 ( .a(n37387), .b(n4201), .o(n40968) );
no02f01 g37177 ( .a(n40968), .b(n40967), .o(n40969) );
in01f01 g37178 ( .a(n40969), .o(n1195) );
no02f01 g37179 ( .a(n40926), .b(n40924), .o(n40971) );
no02f01 g37180 ( .a(n40971), .b(n40916), .o(n40972) );
na02f01 g37181 ( .a(n40971), .b(n40916), .o(n40973) );
in01f01 g37182 ( .a(n40973), .o(n40974) );
no02f01 g37183 ( .a(n40974), .b(n40972), .o(n40975) );
na02f01 g37184 ( .a(n40975), .b(n5799), .o(n40976) );
in01f01 g37185 ( .a(n40975), .o(n2048) );
na02f01 g37186 ( .a(n2048), .b(n911), .o(n40978) );
na02f01 g37187 ( .a(n40978), .b(n40976), .o(n1200) );
no02f01 g37188 ( .a(n38923), .b(n38921), .o(n40980) );
na03f01 g37189 ( .a(n40980), .b(n38910), .c(n38905), .o(n40981) );
na02f01 g37190 ( .a(n38910), .b(n38905), .o(n40982) );
in01f01 g37191 ( .a(n40980), .o(n40983) );
na02f01 g37192 ( .a(n40983), .b(n40982), .o(n40984) );
na02f01 g37193 ( .a(n40984), .b(n40981), .o(n1205) );
no02f01 g37194 ( .a(n38010), .b(n26393), .o(n40986) );
no03f01 g37195 ( .a(n40986), .b(n38015), .c(n38011), .o(n40987) );
oa12f01 g37196 ( .a(n40987), .b(n38047), .c(n38029), .o(n40988) );
ao12f01 g37197 ( .a(n37871), .b(n26361), .c(n26388), .o(n40989) );
no02f01 g37198 ( .a(n40989), .b(n37872), .o(n40990) );
no02f01 g37199 ( .a(n38010), .b(n26396), .o(n40991) );
no02f01 g37200 ( .a(n37871), .b(n26373), .o(n40992) );
no02f01 g37201 ( .a(n40992), .b(n40991), .o(n40993) );
na03f01 g37202 ( .a(n40993), .b(n40990), .c(n40988), .o(n40994) );
na02f01 g37203 ( .a(n40990), .b(n40988), .o(n40995) );
in01f01 g37204 ( .a(n40993), .o(n40996) );
na02f01 g37205 ( .a(n40996), .b(n40995), .o(n40997) );
na02f01 g37206 ( .a(n40997), .b(n40994), .o(n1210) );
na03f01 g37207 ( .a(n36399), .b(n9590), .c(n9589), .o(n40999) );
oa12f01 g37208 ( .a(n5638), .b(n9646), .c(n9645), .o(n41000) );
na02f01 g37209 ( .a(n41000), .b(n40999), .o(n1215) );
na03f01 g37210 ( .a(n5799), .b(n21337), .c(n21311), .o(n41002) );
na02f01 g37211 ( .a(n911), .b(n273), .o(n41003) );
na02f01 g37212 ( .a(n41003), .b(n41002), .o(n1220) );
no02f01 g37213 ( .a(n39135), .b(n31381), .o(n41005) );
na02f01 g37214 ( .a(n39135), .b(n31381), .o(n41006) );
in01f01 g37215 ( .a(n41006), .o(n41007) );
no02f01 g37216 ( .a(n41007), .b(n41005), .o(n41008) );
in01f01 g37217 ( .a(n31545), .o(n41009) );
no02f01 g37218 ( .a(n39059), .b(n41009), .o(n41010) );
no02f01 g37219 ( .a(n31532), .b(n31511), .o(n41011) );
no02f01 g37220 ( .a(n41011), .b(n39059), .o(n41012) );
in01f01 g37221 ( .a(n31557), .o(n41013) );
no02f01 g37222 ( .a(n39059), .b(n41013), .o(n41014) );
no03f01 g37223 ( .a(n41014), .b(n41012), .c(n41010), .o(n41015) );
in01f01 g37224 ( .a(n41015), .o(n41016) );
in01f01 g37225 ( .a(n31596), .o(n41017) );
no02f01 g37226 ( .a(n39059), .b(n41017), .o(n41018) );
no02f01 g37227 ( .a(n31586), .b(n31569), .o(n41019) );
no02f01 g37228 ( .a(n41019), .b(n39059), .o(n41020) );
no03f01 g37229 ( .a(n41020), .b(n41018), .c(n41016), .o(n41021) );
oa12f01 g37230 ( .a(n41021), .b(n39160), .c(n39173), .o(n41022) );
ao12f01 g37231 ( .a(n39135), .b(n31532), .c(n31511), .o(n41023) );
in01f01 g37232 ( .a(n41023), .o(n41024) );
oa12f01 g37233 ( .a(n39059), .b(n41013), .c(n41009), .o(n41025) );
na02f01 g37234 ( .a(n41025), .b(n41024), .o(n41026) );
ao12f01 g37235 ( .a(n39135), .b(n31586), .c(n31569), .o(n41027) );
in01f01 g37236 ( .a(n41027), .o(n41028) );
na02f01 g37237 ( .a(n41028), .b(n31596), .o(n41029) );
ao12f01 g37238 ( .a(n41026), .b(n41029), .c(n39059), .o(n41030) );
na03f01 g37239 ( .a(n41030), .b(n41022), .c(n41008), .o(n41031) );
in01f01 g37240 ( .a(n41008), .o(n41032) );
in01f01 g37241 ( .a(n41021), .o(n41033) );
ao12f01 g37242 ( .a(n41033), .b(n39161), .c(n39153), .o(n41034) );
in01f01 g37243 ( .a(n41030), .o(n41035) );
oa12f01 g37244 ( .a(n41032), .b(n41035), .c(n41034), .o(n41036) );
na03f01 g37245 ( .a(n41036), .b(n41031), .c(n3633), .o(n41037) );
no03f01 g37246 ( .a(n41035), .b(n41034), .c(n41032), .o(n41038) );
ao12f01 g37247 ( .a(n41008), .b(n41030), .c(n41022), .o(n41039) );
oa12f01 g37248 ( .a(n6203), .b(n41039), .c(n41038), .o(n41040) );
na02f01 g37249 ( .a(n41040), .b(n41037), .o(n1225) );
no02f01 g37250 ( .a(n38700), .b(n38689), .o(n41042) );
in01f01 g37251 ( .a(n38708), .o(n41043) );
no02f01 g37252 ( .a(n38706), .b(n36122), .o(n41044) );
in01f01 g37253 ( .a(n41044), .o(n41045) );
na02f01 g37254 ( .a(n41045), .b(n38717), .o(n41046) );
ao12f01 g37255 ( .a(n41046), .b(n41043), .c(n41042), .o(n41047) );
no02f01 g37256 ( .a(n36122), .b(n4696), .o(n41048) );
no02f01 g37257 ( .a(n41048), .b(n38709), .o(n41049) );
na02f01 g37258 ( .a(n41049), .b(n41047), .o(n41050) );
in01f01 g37259 ( .a(n41047), .o(n41051) );
in01f01 g37260 ( .a(n41049), .o(n41052) );
na02f01 g37261 ( .a(n41052), .b(n41051), .o(n41053) );
na02f01 g37262 ( .a(n41053), .b(n41050), .o(n1230) );
no02f01 g37263 ( .a(n9898), .b(n9891), .o(n41055) );
na03f01 g37264 ( .a(n41055), .b(n9874), .c(n9868), .o(n41056) );
in01f01 g37265 ( .a(n41055), .o(n41057) );
oa12f01 g37266 ( .a(n41057), .b(n9873), .c(n39648), .o(n41058) );
na02f01 g37267 ( .a(n41058), .b(n41056), .o(n1235) );
ao12f01 g37268 ( .a(n25504), .b(n25506), .c(n36667), .o(n41060) );
no02f01 g37269 ( .a(n25519), .b(n25328), .o(n41061) );
no02f01 g37270 ( .a(n25515), .b(n39813), .o(n41062) );
no02f01 g37271 ( .a(n41062), .b(n41061), .o(n41063) );
in01f01 g37272 ( .a(n41063), .o(n41064) );
no02f01 g37273 ( .a(n41064), .b(n41060), .o(n41065) );
na02f01 g37274 ( .a(n41064), .b(n41060), .o(n41066) );
in01f01 g37275 ( .a(n41066), .o(n41067) );
no02f01 g37276 ( .a(n41067), .b(n41065), .o(n41068) );
na02f01 g37277 ( .a(n41068), .b(n6037), .o(n41069) );
in01f01 g37278 ( .a(n41068), .o(n3865) );
na02f01 g37279 ( .a(n3865), .b(n5873), .o(n41071) );
na02f01 g37280 ( .a(n41071), .b(n41069), .o(n1240) );
no02f01 g37281 ( .a(n29937), .b(n24547), .o(n41073) );
no02f01 g37282 ( .a(n29938), .b(n24532), .o(n41074) );
no02f01 g37283 ( .a(n41074), .b(n41073), .o(n41075) );
in01f01 g37284 ( .a(n41075), .o(n41076) );
no02f01 g37285 ( .a(n29937), .b(n24405), .o(n41077) );
in01f01 g37286 ( .a(n41077), .o(n41078) );
no02f01 g37287 ( .a(n30131), .b(n30129), .o(n41079) );
no02f01 g37288 ( .a(n29938), .b(n24512), .o(n41080) );
ao12f01 g37289 ( .a(n41080), .b(n41079), .c(n41078), .o(n41081) );
na02f01 g37290 ( .a(n41081), .b(n41076), .o(n41082) );
in01f01 g37291 ( .a(n41081), .o(n41083) );
na02f01 g37292 ( .a(n41083), .b(n41075), .o(n41084) );
na03f01 g37293 ( .a(n41084), .b(n41082), .c(n6037), .o(n41085) );
na02f01 g37294 ( .a(n41084), .b(n41082), .o(n4786) );
na02f01 g37295 ( .a(n4786), .b(n5873), .o(n41087) );
na02f01 g37296 ( .a(n41087), .b(n41085), .o(n1245) );
no02f01 g37297 ( .a(n36963), .b(n35998), .o(n41089) );
na02f01 g37298 ( .a(n36963), .b(n35998), .o(n41090) );
in01f01 g37299 ( .a(n41090), .o(n41091) );
no02f01 g37300 ( .a(n41091), .b(n41089), .o(n41092) );
in01f01 g37301 ( .a(n41092), .o(n41093) );
in01f01 g37302 ( .a(n37150), .o(n41094) );
na02f01 g37303 ( .a(n37270), .b(n41094), .o(n41095) );
no02f01 g37304 ( .a(n41095), .b(n37325), .o(n41096) );
ao12f01 g37305 ( .a(n36963), .b(n37273), .c(n36023), .o(n41097) );
no02f01 g37306 ( .a(n41097), .b(n37263), .o(n41098) );
in01f01 g37307 ( .a(n41098), .o(n41099) );
ao12f01 g37308 ( .a(n41099), .b(n41096), .c(n37309), .o(n41100) );
in01f01 g37309 ( .a(n41100), .o(n41101) );
na02f01 g37310 ( .a(n41101), .b(n41093), .o(n41102) );
na02f01 g37311 ( .a(n41100), .b(n41092), .o(n41103) );
na02f01 g37312 ( .a(n41103), .b(n41102), .o(n1250) );
no03f01 g37313 ( .a(n9591), .b(n9232), .c(n936), .o(n41105) );
no02f01 g37314 ( .a(n40367), .b(n9228), .o(n41106) );
no02f01 g37315 ( .a(n41106), .b(n41105), .o(n41107) );
in01f01 g37316 ( .a(n41107), .o(n1255) );
in01f01 g37317 ( .a(n22559), .o(n41109) );
na03f01 g37318 ( .a(n22565), .b(n4448), .c(n41109), .o(n41110) );
in01f01 g37319 ( .a(n4448), .o(n41111) );
in01f01 g37320 ( .a(n22565), .o(n41112) );
oa12f01 g37321 ( .a(n41111), .b(n41112), .c(n22559), .o(n41113) );
na02f01 g37322 ( .a(n41113), .b(n41110), .o(n1260) );
no02f01 g37323 ( .a(n22654), .b(n22643), .o(n41115) );
in01f01 g37324 ( .a(n41115), .o(n41116) );
na02f01 g37325 ( .a(n41116), .b(n38653), .o(n41117) );
oa12f01 g37326 ( .a(n41115), .b(n22632), .c(n22501), .o(n41118) );
na02f01 g37327 ( .a(n41118), .b(n41117), .o(n1265) );
no02f01 g37328 ( .a(n27401), .b(n27394), .o(n41120) );
no02f01 g37329 ( .a(n27430), .b(n27367), .o(n41121) );
in01f01 g37330 ( .a(n27430), .o(n41122) );
no02f01 g37331 ( .a(n41122), .b(n27395), .o(n41123) );
in01f01 g37332 ( .a(n41123), .o(n41124) );
ao12f01 g37333 ( .a(n41121), .b(n41124), .c(n41120), .o(n41125) );
in01f01 g37334 ( .a(n27439), .o(n41126) );
no02f01 g37335 ( .a(n41126), .b(n27395), .o(n41127) );
no02f01 g37336 ( .a(n27439), .b(n27367), .o(n41128) );
no02f01 g37337 ( .a(n41128), .b(n41127), .o(n41129) );
na02f01 g37338 ( .a(n41129), .b(n41125), .o(n41130) );
in01f01 g37339 ( .a(n41125), .o(n41131) );
in01f01 g37340 ( .a(n41129), .o(n41132) );
na02f01 g37341 ( .a(n41132), .b(n41131), .o(n41133) );
na02f01 g37342 ( .a(n41133), .b(n41130), .o(n1270) );
in01f01 g37343 ( .a(n38921), .o(n41135) );
oa12f01 g37344 ( .a(n41135), .b(n38923), .c(n40982), .o(n41136) );
in01f01 g37345 ( .a(n38936), .o(n41137) );
no02f01 g37346 ( .a(n41137), .b(n38933), .o(n41138) );
na02f01 g37347 ( .a(n41138), .b(n41136), .o(n41139) );
in01f01 g37348 ( .a(n41136), .o(n41140) );
in01f01 g37349 ( .a(n41138), .o(n41141) );
na02f01 g37350 ( .a(n41141), .b(n41140), .o(n41142) );
na02f01 g37351 ( .a(n41142), .b(n41139), .o(n1275) );
in01f01 g37352 ( .a(n8667), .o(n41144) );
in01f01 g37353 ( .a(n8644), .o(n41145) );
na02f01 g37354 ( .a(n8665), .b(n39007), .o(n41146) );
na02f01 g37355 ( .a(n41146), .b(n41145), .o(n41147) );
no02f01 g37356 ( .a(n8669), .b(n8652), .o(n41148) );
na03f01 g37357 ( .a(n41148), .b(n41147), .c(n41144), .o(n41149) );
na02f01 g37358 ( .a(n41147), .b(n41144), .o(n41150) );
in01f01 g37359 ( .a(n41148), .o(n41151) );
na02f01 g37360 ( .a(n41151), .b(n41150), .o(n41152) );
na02f01 g37361 ( .a(n41152), .b(n41149), .o(n1280) );
in01f01 g37362 ( .a(n14232), .o(n41154) );
no02f01 g37363 ( .a(n14235), .b(n41154), .o(n41155) );
no02f01 g37364 ( .a(n41155), .b(n13960), .o(n41156) );
in01f01 g37365 ( .a(n13944), .o(n41157) );
no02f01 g37366 ( .a(n41157), .b(n13943), .o(n41158) );
no02f01 g37367 ( .a(n41158), .b(n41156), .o(n41159) );
na02f01 g37368 ( .a(n41158), .b(n41156), .o(n41160) );
in01f01 g37369 ( .a(n41160), .o(n41161) );
no02f01 g37370 ( .a(n41161), .b(n41159), .o(n41162) );
in01f01 g37371 ( .a(n41162), .o(n1290) );
no02f01 g37372 ( .a(n39135), .b(n31557), .o(n41164) );
no02f01 g37373 ( .a(n41164), .b(n41014), .o(n41165) );
no02f01 g37374 ( .a(n39135), .b(n31545), .o(n41166) );
no03f01 g37375 ( .a(n41012), .b(n39151), .c(n39172), .o(n41167) );
no02f01 g37376 ( .a(n41023), .b(n39160), .o(n41168) );
in01f01 g37377 ( .a(n41168), .o(n41169) );
no03f01 g37378 ( .a(n41169), .b(n41167), .c(n41166), .o(n41170) );
oa12f01 g37379 ( .a(n41165), .b(n41170), .c(n41010), .o(n41171) );
in01f01 g37380 ( .a(n41010), .o(n41172) );
in01f01 g37381 ( .a(n41165), .o(n41173) );
in01f01 g37382 ( .a(n41166), .o(n41174) );
in01f01 g37383 ( .a(n41012), .o(n41175) );
na03f01 g37384 ( .a(n41175), .b(n39152), .c(n39142), .o(n41176) );
na03f01 g37385 ( .a(n41168), .b(n41176), .c(n41174), .o(n41177) );
na03f01 g37386 ( .a(n41177), .b(n41173), .c(n41172), .o(n41178) );
na02f01 g37387 ( .a(n41178), .b(n41171), .o(n1295) );
no02f01 g37388 ( .a(n40794), .b(n20360), .o(n41180) );
no02f01 g37389 ( .a(n40791), .b(n20436), .o(n41181) );
no02f01 g37390 ( .a(n41181), .b(n41180), .o(n41182) );
ao12f01 g37391 ( .a(n40791), .b(n20349), .c(n20431), .o(n41183) );
in01f01 g37392 ( .a(n41183), .o(n41184) );
na02f01 g37393 ( .a(n40789), .b(n40788), .o(n41185) );
na02f01 g37394 ( .a(n40753), .b(n40751), .o(n41186) );
no02f01 g37395 ( .a(n20424), .b(n20164), .o(n41187) );
in01f01 g37396 ( .a(n41187), .o(n41188) );
na03f01 g37397 ( .a(n41188), .b(n41186), .c(n41185), .o(n41189) );
na03f01 g37398 ( .a(n41186), .b(n41185), .c(n20334), .o(n41190) );
na03f01 g37399 ( .a(n41186), .b(n41185), .c(n20159), .o(n41191) );
na03f01 g37400 ( .a(n41191), .b(n41190), .c(n41189), .o(n41192) );
ao12f01 g37401 ( .a(n41192), .b(n40949), .c(n40946), .o(n41193) );
ao12f01 g37402 ( .a(n40791), .b(n20334), .c(n20159), .o(n41194) );
ao12f01 g37403 ( .a(n40791), .b(n20424), .c(n20164), .o(n41195) );
no02f01 g37404 ( .a(n41195), .b(n41194), .o(n41196) );
in01f01 g37405 ( .a(n41196), .o(n41197) );
na02f01 g37406 ( .a(n40791), .b(n20431), .o(n41198) );
na02f01 g37407 ( .a(n40791), .b(n20349), .o(n41199) );
na02f01 g37408 ( .a(n41199), .b(n41198), .o(n41200) );
in01f01 g37409 ( .a(n41200), .o(n41201) );
oa12f01 g37410 ( .a(n41201), .b(n41197), .c(n41193), .o(n41202) );
na03f01 g37411 ( .a(n41202), .b(n41184), .c(n41182), .o(n41203) );
in01f01 g37412 ( .a(n41182), .o(n41204) );
no03f01 g37413 ( .a(n41187), .b(n40790), .c(n40754), .o(n41205) );
no03f01 g37414 ( .a(n40790), .b(n40754), .c(n20326), .o(n41206) );
no03f01 g37415 ( .a(n40790), .b(n40754), .c(n20331), .o(n41207) );
no03f01 g37416 ( .a(n41207), .b(n41206), .c(n41205), .o(n41208) );
oa12f01 g37417 ( .a(n41208), .b(n40935), .c(n40837), .o(n41209) );
ao12f01 g37418 ( .a(n41200), .b(n41196), .c(n41209), .o(n41210) );
oa12f01 g37419 ( .a(n41204), .b(n41210), .c(n41183), .o(n41211) );
na03f01 g37420 ( .a(n41211), .b(n41203), .c(n5799), .o(n41212) );
no03f01 g37421 ( .a(n41210), .b(n41183), .c(n41204), .o(n41213) );
ao12f01 g37422 ( .a(n41182), .b(n41202), .c(n41184), .o(n41214) );
oa12f01 g37423 ( .a(n911), .b(n41214), .c(n41213), .o(n41215) );
na02f01 g37424 ( .a(n41215), .b(n41212), .o(n1300) );
no02f01 g37425 ( .a(n37871), .b(n26232), .o(n41217) );
in01f01 g37426 ( .a(n26232), .o(n41218) );
no02f01 g37427 ( .a(n38010), .b(n41218), .o(n41219) );
no02f01 g37428 ( .a(n41219), .b(n41217), .o(n41220) );
no02f01 g37429 ( .a(n38010), .b(n26413), .o(n41221) );
no02f01 g37430 ( .a(n38010), .b(n26411), .o(n41222) );
no02f01 g37431 ( .a(n26399), .b(n26398), .o(n41223) );
no02f01 g37432 ( .a(n41223), .b(n26373), .o(n41224) );
no02f01 g37433 ( .a(n41224), .b(n38010), .o(n41225) );
no03f01 g37434 ( .a(n41225), .b(n41222), .c(n41221), .o(n41226) );
in01f01 g37435 ( .a(n41226), .o(n41227) );
ao12f01 g37436 ( .a(n41227), .b(n40990), .c(n40988), .o(n41228) );
no02f01 g37437 ( .a(n38010), .b(n26428), .o(n41229) );
no02f01 g37438 ( .a(n26256), .b(n26250), .o(n41230) );
no02f01 g37439 ( .a(n41230), .b(n38010), .o(n41231) );
no02f01 g37440 ( .a(n41231), .b(n41229), .o(n41232) );
na02f01 g37441 ( .a(n41232), .b(n41228), .o(n41233) );
ao12f01 g37442 ( .a(n37871), .b(n26256), .c(n26250), .o(n41234) );
in01f01 g37443 ( .a(n41234), .o(n41235) );
ao12f01 g37444 ( .a(n37871), .b(n41235), .c(n26438), .o(n41236) );
ao12f01 g37445 ( .a(n37871), .b(n41223), .c(n26373), .o(n41237) );
ao12f01 g37446 ( .a(n37871), .b(n26407), .c(n26272), .o(n41238) );
no02f01 g37447 ( .a(n41238), .b(n41237), .o(n41239) );
in01f01 g37448 ( .a(n41239), .o(n41240) );
no02f01 g37449 ( .a(n41240), .b(n41236), .o(n41241) );
na03f01 g37450 ( .a(n41241), .b(n41233), .c(n41220), .o(n41242) );
in01f01 g37451 ( .a(n41220), .o(n41243) );
no02f01 g37452 ( .a(n40986), .b(n38015), .o(n41244) );
na02f01 g37453 ( .a(n41244), .b(n38012), .o(n41245) );
ao12f01 g37454 ( .a(n41245), .b(n38006), .c(n37915), .o(n41246) );
in01f01 g37455 ( .a(n40990), .o(n41247) );
oa12f01 g37456 ( .a(n41226), .b(n41247), .c(n41246), .o(n41248) );
no03f01 g37457 ( .a(n41231), .b(n41229), .c(n41248), .o(n41249) );
in01f01 g37458 ( .a(n41241), .o(n41250) );
oa12f01 g37459 ( .a(n41243), .b(n41250), .c(n41249), .o(n41251) );
na03f01 g37460 ( .a(n41251), .b(n41242), .c(n1821), .o(n41252) );
no03f01 g37461 ( .a(n41250), .b(n41249), .c(n41243), .o(n41253) );
ao12f01 g37462 ( .a(n41220), .b(n41241), .c(n41233), .o(n41254) );
oa12f01 g37463 ( .a(n8066), .b(n41254), .c(n41253), .o(n41255) );
na02f01 g37464 ( .a(n41255), .b(n41252), .o(n1305) );
no02f01 g37465 ( .a(n30020), .b(n30052), .o(n41257) );
no02f01 g37466 ( .a(n41257), .b(n30019), .o(n41258) );
na02f01 g37467 ( .a(n41257), .b(n30019), .o(n41259) );
in01f01 g37468 ( .a(n41259), .o(n41260) );
no02f01 g37469 ( .a(n41260), .b(n41258), .o(n41261) );
na02f01 g37470 ( .a(n41261), .b(n6037), .o(n41262) );
in01f01 g37471 ( .a(n41261), .o(n5493) );
na02f01 g37472 ( .a(n5493), .b(n5873), .o(n41264) );
na02f01 g37473 ( .a(n41264), .b(n41262), .o(n1310) );
na02f01 g37474 ( .a(n32732), .b(sin_out_25), .o(n41266) );
no02f01 g37475 ( .a(n35818), .b(n35807), .o(n41267) );
in01f01 g37476 ( .a(n41267), .o(n41268) );
no02f01 g37477 ( .a(n35845), .b(n34287), .o(n41269) );
no02f01 g37478 ( .a(n35846), .b(n34336), .o(n41270) );
in01f01 g37479 ( .a(n41270), .o(n41271) );
ao12f01 g37480 ( .a(n41269), .b(n41271), .c(n41268), .o(n41272) );
in01f01 g37481 ( .a(n41272), .o(n41273) );
no02f01 g37482 ( .a(n35839), .b(n34287), .o(n41274) );
no02f01 g37483 ( .a(n35840), .b(n34336), .o(n41275) );
no02f01 g37484 ( .a(n41275), .b(n41274), .o(n41276) );
in01f01 g37485 ( .a(n41276), .o(n41277) );
no02f01 g37486 ( .a(n41277), .b(n41273), .o(n41278) );
no02f01 g37487 ( .a(n41276), .b(n41272), .o(n41279) );
no03f01 g37488 ( .a(n41279), .b(n41278), .c(n34267), .o(n41280) );
no02f01 g37489 ( .a(n41279), .b(n41278), .o(n41281) );
no02f01 g37490 ( .a(n41281), .b(n34307), .o(n41282) );
no02f01 g37491 ( .a(n41282), .b(n41280), .o(n41283) );
in01f01 g37492 ( .a(n41283), .o(n41284) );
no02f01 g37493 ( .a(n41270), .b(n41269), .o(n41285) );
in01f01 g37494 ( .a(n41285), .o(n41286) );
no02f01 g37495 ( .a(n41286), .b(n41268), .o(n41287) );
no02f01 g37496 ( .a(n41285), .b(n41267), .o(n41288) );
no02f01 g37497 ( .a(n41288), .b(n41287), .o(n41289) );
in01f01 g37498 ( .a(n41289), .o(n41290) );
no02f01 g37499 ( .a(n41290), .b(n34267), .o(n41291) );
in01f01 g37500 ( .a(n39590), .o(n41292) );
na04f01 g37501 ( .a(n41292), .b(n39578), .c(n39494), .d(n36595), .o(n41293) );
na02f01 g37502 ( .a(n39597), .b(n41293), .o(n41294) );
no02f01 g37503 ( .a(n39611), .b(n39601), .o(n41295) );
in01f01 g37504 ( .a(n41295), .o(n41296) );
no02f01 g37505 ( .a(n35763), .b(n39546), .o(n41297) );
in01f01 g37506 ( .a(n41297), .o(n41298) );
no02f01 g37507 ( .a(n35730), .b(n34287), .o(n41299) );
no02f01 g37508 ( .a(n41299), .b(n35808), .o(n41300) );
oa12f01 g37509 ( .a(n41300), .b(n41298), .c(n35732), .o(n41301) );
no02f01 g37510 ( .a(n35744), .b(n34287), .o(n41302) );
no02f01 g37511 ( .a(n41302), .b(n35746), .o(n41303) );
in01f01 g37512 ( .a(n41303), .o(n41304) );
no02f01 g37513 ( .a(n41304), .b(n41301), .o(n41305) );
na02f01 g37514 ( .a(n41304), .b(n41301), .o(n41306) );
in01f01 g37515 ( .a(n41306), .o(n41307) );
no03f01 g37516 ( .a(n41307), .b(n41305), .c(n34267), .o(n41308) );
no02f01 g37517 ( .a(n41299), .b(n35732), .o(n41309) );
in01f01 g37518 ( .a(n41309), .o(n41310) );
no03f01 g37519 ( .a(n41310), .b(n41297), .c(n35808), .o(n41311) );
no02f01 g37520 ( .a(n41297), .b(n35808), .o(n41312) );
no02f01 g37521 ( .a(n41309), .b(n41312), .o(n41313) );
no03f01 g37522 ( .a(n41313), .b(n41311), .c(n34267), .o(n41314) );
no03f01 g37523 ( .a(n41314), .b(n41308), .c(n41296), .o(n41315) );
oa12f01 g37524 ( .a(n35810), .b(n35765), .c(n39546), .o(n41316) );
na02f01 g37525 ( .a(n35802), .b(n34287), .o(n41317) );
in01f01 g37526 ( .a(n41317), .o(n41318) );
no02f01 g37527 ( .a(n41318), .b(n35812), .o(n41319) );
in01f01 g37528 ( .a(n41319), .o(n41320) );
no02f01 g37529 ( .a(n41320), .b(n41316), .o(n41321) );
in01f01 g37530 ( .a(n41316), .o(n41322) );
no02f01 g37531 ( .a(n41319), .b(n41322), .o(n41323) );
no03f01 g37532 ( .a(n41323), .b(n41321), .c(n34267), .o(n41324) );
ao12f01 g37533 ( .a(n35812), .b(n41317), .c(n41316), .o(n41325) );
na02f01 g37534 ( .a(n35797), .b(n34287), .o(n41326) );
in01f01 g37535 ( .a(n41326), .o(n41327) );
no02f01 g37536 ( .a(n41327), .b(n35811), .o(n41328) );
no02f01 g37537 ( .a(n41328), .b(n41325), .o(n41329) );
na02f01 g37538 ( .a(n41328), .b(n41325), .o(n41330) );
in01f01 g37539 ( .a(n41330), .o(n41331) );
no03f01 g37540 ( .a(n41331), .b(n41329), .c(n34267), .o(n41332) );
no02f01 g37541 ( .a(n41332), .b(n41324), .o(n41333) );
in01f01 g37542 ( .a(n41333), .o(n41334) );
no02f01 g37543 ( .a(n35776), .b(n34287), .o(n41335) );
in01f01 g37544 ( .a(n41335), .o(n41336) );
no03f01 g37545 ( .a(n35804), .b(n35765), .c(n39546), .o(n41337) );
no02f01 g37546 ( .a(n41337), .b(n35814), .o(n41338) );
ao12f01 g37547 ( .a(n35778), .b(n41338), .c(n41336), .o(n41339) );
in01f01 g37548 ( .a(n41339), .o(n41340) );
no02f01 g37549 ( .a(n35815), .b(n34287), .o(n41341) );
no02f01 g37550 ( .a(n41341), .b(n35787), .o(n41342) );
no02f01 g37551 ( .a(n41342), .b(n41340), .o(n41343) );
na02f01 g37552 ( .a(n41342), .b(n41340), .o(n41344) );
in01f01 g37553 ( .a(n41344), .o(n41345) );
no03f01 g37554 ( .a(n41345), .b(n41343), .c(n34267), .o(n41346) );
no02f01 g37555 ( .a(n41335), .b(n35778), .o(n41347) );
no02f01 g37556 ( .a(n41347), .b(n41338), .o(n41348) );
na02f01 g37557 ( .a(n41347), .b(n41338), .o(n41349) );
in01f01 g37558 ( .a(n41349), .o(n41350) );
no03f01 g37559 ( .a(n41350), .b(n41348), .c(n34267), .o(n41351) );
no03f01 g37560 ( .a(n41351), .b(n41346), .c(n41334), .o(n41352) );
na03f01 g37561 ( .a(n41352), .b(n41315), .c(n41294), .o(n41353) );
no02f01 g37562 ( .a(n41353), .b(n41291), .o(n41354) );
no02f01 g37563 ( .a(n41289), .b(n34307), .o(n41355) );
in01f01 g37564 ( .a(n41355), .o(n41356) );
no02f01 g37565 ( .a(n41307), .b(n41305), .o(n41357) );
no02f01 g37566 ( .a(n41313), .b(n41311), .o(n41358) );
ao12f01 g37567 ( .a(n34307), .b(n41358), .c(n41357), .o(n41359) );
ao12f01 g37568 ( .a(n34307), .b(n39612), .c(n39553), .o(n41360) );
no02f01 g37569 ( .a(n41360), .b(n41359), .o(n41361) );
in01f01 g37570 ( .a(n41361), .o(n41362) );
no02f01 g37571 ( .a(n41323), .b(n41321), .o(n41363) );
no02f01 g37572 ( .a(n41331), .b(n41329), .o(n41364) );
ao12f01 g37573 ( .a(n34307), .b(n41364), .c(n41363), .o(n41365) );
no02f01 g37574 ( .a(n41365), .b(n41362), .o(n41366) );
in01f01 g37575 ( .a(n41366), .o(n41367) );
no02f01 g37576 ( .a(n41345), .b(n41343), .o(n41368) );
no02f01 g37577 ( .a(n41350), .b(n41348), .o(n41369) );
ao12f01 g37578 ( .a(n34307), .b(n41369), .c(n41368), .o(n41370) );
no02f01 g37579 ( .a(n41370), .b(n41367), .o(n41371) );
na02f01 g37580 ( .a(n41371), .b(n41356), .o(n41372) );
no03f01 g37581 ( .a(n41372), .b(n41354), .c(n41284), .o(n41373) );
no02f01 g37582 ( .a(n41372), .b(n41354), .o(n41374) );
no02f01 g37583 ( .a(n41374), .b(n41283), .o(n41375) );
oa12f01 g37584 ( .a(n32734), .b(n41375), .c(n41373), .o(n41376) );
na02f01 g37585 ( .a(n41376), .b(n41266), .o(n1315) );
ao12f01 g37586 ( .a(n21305), .b(n40771), .c(n21308), .o(n41378) );
no02f01 g37587 ( .a(n40712), .b(n21305), .o(n41379) );
no02f01 g37588 ( .a(n40681), .b(n21305), .o(n41380) );
no03f01 g37589 ( .a(n41380), .b(n41379), .c(n41378), .o(n41381) );
oa12f01 g37590 ( .a(n41381), .b(n21263), .c(n20923), .o(n41382) );
ao12f01 g37591 ( .a(n21270), .b(n40770), .c(n40709), .o(n41383) );
ao12f01 g37592 ( .a(n21270), .b(n40715), .c(n21301), .o(n41384) );
no02f01 g37593 ( .a(n41384), .b(n41383), .o(n41385) );
no02f01 g37594 ( .a(n40779), .b(n21305), .o(n41386) );
no02f01 g37595 ( .a(n40725), .b(n21270), .o(n41387) );
no02f01 g37596 ( .a(n41387), .b(n41386), .o(n41388) );
na03f01 g37597 ( .a(n41388), .b(n41385), .c(n41382), .o(n41389) );
oa12f01 g37598 ( .a(n21270), .b(n40715), .c(n21301), .o(n41390) );
oa12f01 g37599 ( .a(n21270), .b(n40770), .c(n40709), .o(n41391) );
na02f01 g37600 ( .a(n41391), .b(n41390), .o(n41392) );
ao12f01 g37601 ( .a(n41392), .b(n21334), .c(n21327), .o(n41393) );
in01f01 g37602 ( .a(n41385), .o(n41394) );
in01f01 g37603 ( .a(n41388), .o(n41395) );
oa12f01 g37604 ( .a(n41395), .b(n41394), .c(n41393), .o(n41396) );
na03f01 g37605 ( .a(n41396), .b(n41389), .c(n5799), .o(n41397) );
na02f01 g37606 ( .a(n41396), .b(n41389), .o(n5425) );
na02f01 g37607 ( .a(n5425), .b(n911), .o(n41399) );
na02f01 g37608 ( .a(n41399), .b(n41397), .o(n1319) );
oa12f01 g37609 ( .a(n37012), .b(n37162), .c(n36997), .o(n41401) );
na03f01 g37610 ( .a(n37013), .b(n37161), .c(n37156), .o(n41402) );
na02f01 g37611 ( .a(n41402), .b(n41401), .o(n1324) );
in01f01 g37612 ( .a(n8506), .o(n41404) );
no02f01 g37613 ( .a(n8504), .b(n8471), .o(n41405) );
ao12f01 g37614 ( .a(n41405), .b(n41404), .c(n37800), .o(n41406) );
no02f01 g37615 ( .a(n8496), .b(n8471), .o(n41407) );
no02f01 g37616 ( .a(n41407), .b(n8498), .o(n41408) );
na02f01 g37617 ( .a(n41408), .b(n41406), .o(n41409) );
in01f01 g37618 ( .a(n41406), .o(n41410) );
in01f01 g37619 ( .a(n41408), .o(n41411) );
na02f01 g37620 ( .a(n41411), .b(n41410), .o(n41412) );
na02f01 g37621 ( .a(n41412), .b(n41409), .o(n1329) );
in01f01 g37622 ( .a(rst), .o(n41414) );
in01f01 g37623 ( .a(mux_while_ln12_psv_q_6_), .o(n41415) );
in01f01 g37624 ( .a(state_cordic_1_), .o(n41416) );
no03f01 g37625 ( .a(n41416), .b(n41415), .c(n41414), .o(n1334) );
no02f01 g37626 ( .a(n36186), .b(n36122), .o(n41418) );
in01f01 g37627 ( .a(n36186), .o(n41419) );
no02f01 g37628 ( .a(n41419), .b(n36038), .o(n41420) );
no02f01 g37629 ( .a(n41420), .b(n41418), .o(n41421) );
na02f01 g37630 ( .a(n41421), .b(n36171), .o(n41422) );
na02f01 g37631 ( .a(n36169), .b(n38785), .o(n41423) );
in01f01 g37632 ( .a(n41421), .o(n41424) );
na02f01 g37633 ( .a(n41424), .b(n41423), .o(n41425) );
na02f01 g37634 ( .a(n41425), .b(n41422), .o(n1339) );
na02f01 g37635 ( .a(n32732), .b(cos_out_2), .o(n41427) );
no02f01 g37636 ( .a(n35940), .b(n35944), .o(n41428) );
no03f01 g37637 ( .a(n41428), .b(n35942), .c(n35933), .o(n41429) );
no02f01 g37638 ( .a(n41428), .b(n35942), .o(n41430) );
no02f01 g37639 ( .a(n41430), .b(n35976), .o(n41431) );
oa12f01 g37640 ( .a(n32734), .b(n41431), .c(n41429), .o(n41432) );
na02f01 g37641 ( .a(n41432), .b(n41427), .o(n1344) );
no02f01 g37642 ( .a(n29841), .b(n9238), .o(n41434) );
na03f01 g37643 ( .a(n41434), .b(n9590), .c(n9589), .o(n41435) );
in01f01 g37644 ( .a(n41434), .o(n5643) );
oa12f01 g37645 ( .a(n5643), .b(n9646), .c(n9645), .o(n41437) );
na02f01 g37646 ( .a(n41437), .b(n41435), .o(n1348) );
na03f01 g37647 ( .a(n39451), .b(n40027), .c(n40005), .o(n41439) );
oa12f01 g37648 ( .a(n39450), .b(n40028), .c(n39386), .o(n41440) );
na02f01 g37649 ( .a(n41440), .b(n41439), .o(n1353) );
no02f01 g37650 ( .a(n16300), .b(n16329), .o(n41442) );
no02f01 g37651 ( .a(n16430), .b(n16155), .o(n41443) );
in01f01 g37652 ( .a(n41443), .o(n41444) );
ao12f01 g37653 ( .a(n41442), .b(n41444), .c(n21371), .o(n41445) );
no02f01 g37654 ( .a(n16295), .b(n16329), .o(n41446) );
no02f01 g37655 ( .a(n16429), .b(n16155), .o(n41447) );
no02f01 g37656 ( .a(n41447), .b(n41446), .o(n41448) );
na02f01 g37657 ( .a(n41448), .b(n41445), .o(n41449) );
in01f01 g37658 ( .a(n41445), .o(n41450) );
in01f01 g37659 ( .a(n41448), .o(n41451) );
na02f01 g37660 ( .a(n41451), .b(n41450), .o(n41452) );
na02f01 g37661 ( .a(n41452), .b(n41449), .o(n1358) );
in01f01 g37662 ( .a(n9599), .o(n41454) );
no02f01 g37663 ( .a(n9595), .b(beta_31), .o(n41455) );
no02f01 g37664 ( .a(n41455), .b(n9600), .o(n41456) );
in01f01 g37665 ( .a(n41456), .o(n41457) );
no02f01 g37666 ( .a(n41457), .b(n41454), .o(n41458) );
no02f01 g37667 ( .a(n41456), .b(n9599), .o(n41459) );
no02f01 g37668 ( .a(n41459), .b(n41458), .o(n41460) );
na03f01 g37669 ( .a(n41460), .b(n9590), .c(n9589), .o(n41461) );
in01f01 g37670 ( .a(n41460), .o(n1645) );
oa12f01 g37671 ( .a(n1645), .b(n9646), .c(n9645), .o(n41463) );
na02f01 g37672 ( .a(n41463), .b(n41461), .o(n1363) );
na03f01 g37673 ( .a(n25864), .b(n30087), .c(n30076), .o(n41465) );
oa12f01 g37674 ( .a(n25863), .b(n30088), .c(n25818), .o(n41466) );
na02f01 g37675 ( .a(n41466), .b(n41465), .o(n1368) );
na02f01 g37676 ( .a(n32732), .b(cos_out_22), .o(n41468) );
no02f01 g37677 ( .a(n39699), .b(n39703), .o(n41469) );
no02f01 g37678 ( .a(n33979), .b(n33508), .o(n41470) );
no02f01 g37679 ( .a(n33978), .b(n33507), .o(n41471) );
no02f01 g37680 ( .a(n41471), .b(n41470), .o(n41472) );
in01f01 g37681 ( .a(n41472), .o(n41473) );
no03f01 g37682 ( .a(n41473), .b(n41469), .c(n39698), .o(n41474) );
no02f01 g37683 ( .a(n41469), .b(n39698), .o(n41475) );
no02f01 g37684 ( .a(n41472), .b(n41475), .o(n41476) );
no02f01 g37685 ( .a(n41476), .b(n41474), .o(n41477) );
ao12f01 g37686 ( .a(n35944), .b(n41477), .c(n39705), .o(n41478) );
no02f01 g37687 ( .a(n41478), .b(n39695), .o(n41479) );
in01f01 g37688 ( .a(n41479), .o(n41480) );
na02f01 g37689 ( .a(n41477), .b(n35944), .o(n41481) );
na02f01 g37690 ( .a(n41481), .b(n39707), .o(n41482) );
no02f01 g37691 ( .a(n41482), .b(n39712), .o(n41483) );
no02f01 g37692 ( .a(n39703), .b(n33986), .o(n41484) );
no02f01 g37693 ( .a(n33957), .b(n33507), .o(n41485) );
no02f01 g37694 ( .a(n41485), .b(n33959), .o(n41486) );
in01f01 g37695 ( .a(n41486), .o(n41487) );
no03f01 g37696 ( .a(n41487), .b(n41484), .c(n34212), .o(n41488) );
no02f01 g37697 ( .a(n41484), .b(n34212), .o(n41489) );
no02f01 g37698 ( .a(n41486), .b(n41489), .o(n41490) );
no02f01 g37699 ( .a(n41490), .b(n41488), .o(n41491) );
no02f01 g37700 ( .a(n41491), .b(n35944), .o(n41492) );
na02f01 g37701 ( .a(n41491), .b(n35944), .o(n41493) );
in01f01 g37702 ( .a(n41493), .o(n41494) );
no02f01 g37703 ( .a(n41494), .b(n41492), .o(n41495) );
in01f01 g37704 ( .a(n41495), .o(n41496) );
no03f01 g37705 ( .a(n41496), .b(n41483), .c(n41480), .o(n41497) );
in01f01 g37706 ( .a(n41482), .o(n41498) );
ao12f01 g37707 ( .a(n41480), .b(n41498), .c(n39691), .o(n41499) );
no02f01 g37708 ( .a(n41495), .b(n41499), .o(n41500) );
oa12f01 g37709 ( .a(n32734), .b(n41500), .c(n41497), .o(n41501) );
na02f01 g37710 ( .a(n41501), .b(n41468), .o(n1373) );
na03f01 g37711 ( .a(n38403), .b(n39108), .c(n39093), .o(n41503) );
oa12f01 g37712 ( .a(n38402), .b(n39109), .c(n38371), .o(n41504) );
na02f01 g37713 ( .a(n41504), .b(n41503), .o(n1377) );
no02f01 g37714 ( .a(n25179), .b(n25023), .o(n41506) );
no02f01 g37715 ( .a(n41506), .b(n25181), .o(n41507) );
no02f01 g37716 ( .a(n25543), .b(n25023), .o(n41508) );
na02f01 g37717 ( .a(n37144), .b(n25562), .o(n41509) );
na03f01 g37718 ( .a(n41509), .b(n25574), .c(n25570), .o(n41510) );
no02f01 g37719 ( .a(n41510), .b(n41508), .o(n41511) );
oa12f01 g37720 ( .a(n41507), .b(n41511), .c(n25159), .o(n41512) );
in01f01 g37721 ( .a(n25159), .o(n41513) );
in01f01 g37722 ( .a(n41507), .o(n41514) );
in01f01 g37723 ( .a(n41508), .o(n41515) );
no03f01 g37724 ( .a(n25538), .b(n25300), .c(n25287), .o(n41516) );
na02f01 g37725 ( .a(n41516), .b(n41515), .o(n41517) );
na03f01 g37726 ( .a(n41517), .b(n41514), .c(n41513), .o(n41518) );
na02f01 g37727 ( .a(n41518), .b(n41512), .o(n1382) );
no02f01 g37728 ( .a(n22480), .b(n22381), .o(n41520) );
no02f01 g37729 ( .a(n41520), .b(n22366), .o(n41521) );
na02f01 g37730 ( .a(n41520), .b(n22366), .o(n41522) );
in01f01 g37731 ( .a(n41522), .o(n41523) );
no02f01 g37732 ( .a(n41523), .b(n41521), .o(n41524) );
na02f01 g37733 ( .a(n41524), .b(n2589), .o(n41525) );
in01f01 g37734 ( .a(n41524), .o(n5160) );
na02f01 g37735 ( .a(n5160), .b(n4116), .o(n41527) );
na02f01 g37736 ( .a(n41527), .b(n41525), .o(n1387) );
na02f01 g37737 ( .a(n32732), .b(cos_out_31), .o(n41529) );
no02f01 g37738 ( .a(n34306), .b(n34305), .o(n41530) );
in01f01 g37739 ( .a(n41530), .o(n41531) );
no02f01 g37740 ( .a(n35912), .b(n41531), .o(n41532) );
no02f01 g37741 ( .a(n35944), .b(n41530), .o(n41533) );
no02f01 g37742 ( .a(n41533), .b(n41532), .o(n41534) );
in01f01 g37743 ( .a(n41534), .o(n41535) );
in01f01 g37744 ( .a(n41485), .o(n41536) );
ao12f01 g37745 ( .a(n33959), .b(n41489), .c(n41536), .o(n41537) );
no02f01 g37746 ( .a(n34213), .b(n33507), .o(n41538) );
no02f01 g37747 ( .a(n41538), .b(n33968), .o(n41539) );
in01f01 g37748 ( .a(n41539), .o(n41540) );
na02f01 g37749 ( .a(n41540), .b(n41537), .o(n41541) );
no02f01 g37750 ( .a(n41540), .b(n41537), .o(n41542) );
in01f01 g37751 ( .a(n41542), .o(n41543) );
na02f01 g37752 ( .a(n41543), .b(n41541), .o(n41544) );
no02f01 g37753 ( .a(n41544), .b(n35912), .o(n41545) );
no03f01 g37754 ( .a(n41545), .b(n41494), .c(n41482), .o(n41546) );
in01f01 g37755 ( .a(n41546), .o(n41547) );
no02f01 g37756 ( .a(n33890), .b(n33507), .o(n41548) );
ao12f01 g37757 ( .a(n34216), .b(n39696), .c(n33987), .o(n41549) );
in01f01 g37758 ( .a(n41549), .o(n41550) );
no02f01 g37759 ( .a(n33891), .b(n33508), .o(n41551) );
in01f01 g37760 ( .a(n41551), .o(n41552) );
ao12f01 g37761 ( .a(n41548), .b(n41552), .c(n41550), .o(n41553) );
in01f01 g37762 ( .a(n41553), .o(n41554) );
no02f01 g37763 ( .a(n33884), .b(n33508), .o(n41555) );
no02f01 g37764 ( .a(n33883), .b(n33507), .o(n41556) );
no02f01 g37765 ( .a(n41556), .b(n41555), .o(n41557) );
in01f01 g37766 ( .a(n41557), .o(n41558) );
no02f01 g37767 ( .a(n41558), .b(n41554), .o(n41559) );
no02f01 g37768 ( .a(n41557), .b(n41553), .o(n41560) );
no03f01 g37769 ( .a(n41560), .b(n41559), .c(n35912), .o(n41561) );
no02f01 g37770 ( .a(n41551), .b(n41548), .o(n41562) );
in01f01 g37771 ( .a(n41562), .o(n41563) );
no02f01 g37772 ( .a(n41563), .b(n41550), .o(n41564) );
no02f01 g37773 ( .a(n41562), .b(n41549), .o(n41565) );
no02f01 g37774 ( .a(n41565), .b(n41564), .o(n41566) );
in01f01 g37775 ( .a(n41566), .o(n41567) );
no02f01 g37776 ( .a(n41567), .b(n35912), .o(n41568) );
no02f01 g37777 ( .a(n41568), .b(n41561), .o(n41569) );
in01f01 g37778 ( .a(n41569), .o(n41570) );
no02f01 g37779 ( .a(n41549), .b(n33892), .o(n41571) );
no02f01 g37780 ( .a(n34220), .b(n33851), .o(n41572) );
in01f01 g37781 ( .a(n41572), .o(n41573) );
no03f01 g37782 ( .a(n41573), .b(n41571), .c(n34218), .o(n41574) );
no02f01 g37783 ( .a(n41571), .b(n34218), .o(n41575) );
no02f01 g37784 ( .a(n41572), .b(n41575), .o(n41576) );
no02f01 g37785 ( .a(n41576), .b(n41574), .o(n41577) );
in01f01 g37786 ( .a(n41577), .o(n41578) );
no02f01 g37787 ( .a(n41578), .b(n35912), .o(n41579) );
ao12f01 g37788 ( .a(n33851), .b(n41575), .c(n34221), .o(n41580) );
no02f01 g37789 ( .a(n34219), .b(n33507), .o(n41581) );
no02f01 g37790 ( .a(n41581), .b(n33874), .o(n41582) );
in01f01 g37791 ( .a(n41582), .o(n41583) );
no02f01 g37792 ( .a(n41583), .b(n41580), .o(n41584) );
na02f01 g37793 ( .a(n41583), .b(n41580), .o(n41585) );
in01f01 g37794 ( .a(n41585), .o(n41586) );
no03f01 g37795 ( .a(n41586), .b(n41584), .c(n35912), .o(n41587) );
no03f01 g37796 ( .a(n41587), .b(n41579), .c(n41570), .o(n41588) );
in01f01 g37797 ( .a(n41588), .o(n41589) );
no02f01 g37798 ( .a(n33929), .b(n33507), .o(n41590) );
no02f01 g37799 ( .a(n34222), .b(n34218), .o(n41591) );
oa12f01 g37800 ( .a(n41591), .b(n41549), .c(n33894), .o(n41592) );
no02f01 g37801 ( .a(n33930), .b(n33508), .o(n41593) );
in01f01 g37802 ( .a(n41593), .o(n41594) );
ao12f01 g37803 ( .a(n41590), .b(n41594), .c(n41592), .o(n41595) );
in01f01 g37804 ( .a(n41595), .o(n41596) );
no02f01 g37805 ( .a(n33923), .b(n33508), .o(n41597) );
no02f01 g37806 ( .a(n33922), .b(n33507), .o(n41598) );
no02f01 g37807 ( .a(n41598), .b(n41597), .o(n41599) );
in01f01 g37808 ( .a(n41599), .o(n41600) );
no02f01 g37809 ( .a(n41600), .b(n41596), .o(n41601) );
no02f01 g37810 ( .a(n41599), .b(n41595), .o(n41602) );
no03f01 g37811 ( .a(n41602), .b(n41601), .c(n35912), .o(n41603) );
no02f01 g37812 ( .a(n41593), .b(n41590), .o(n41604) );
in01f01 g37813 ( .a(n41604), .o(n41605) );
no02f01 g37814 ( .a(n41605), .b(n41592), .o(n41606) );
in01f01 g37815 ( .a(n41592), .o(n41607) );
no02f01 g37816 ( .a(n41604), .b(n41607), .o(n41608) );
no02f01 g37817 ( .a(n41608), .b(n41606), .o(n41609) );
in01f01 g37818 ( .a(n41609), .o(n41610) );
no02f01 g37819 ( .a(n41610), .b(n35912), .o(n41611) );
no02f01 g37820 ( .a(n41611), .b(n41603), .o(n41612) );
in01f01 g37821 ( .a(n41612), .o(n41613) );
oa12f01 g37822 ( .a(n34224), .b(n41607), .c(n33931), .o(n41614) );
no02f01 g37823 ( .a(n33943), .b(n33507), .o(n41615) );
no02f01 g37824 ( .a(n41615), .b(n33945), .o(n41616) );
in01f01 g37825 ( .a(n41616), .o(n41617) );
no02f01 g37826 ( .a(n41617), .b(n41614), .o(n41618) );
na02f01 g37827 ( .a(n41617), .b(n41614), .o(n41619) );
in01f01 g37828 ( .a(n41619), .o(n41620) );
no03f01 g37829 ( .a(n41620), .b(n41618), .c(n35912), .o(n41621) );
no02f01 g37830 ( .a(n41621), .b(n41613), .o(n41622) );
in01f01 g37831 ( .a(n41622), .o(n41623) );
no04f01 g37832 ( .a(n41623), .b(n41589), .c(n41547), .d(n39712), .o(n41624) );
ao12f01 g37833 ( .a(n41478), .b(n41546), .c(n39695), .o(n41625) );
in01f01 g37834 ( .a(n41544), .o(n41626) );
ao12f01 g37835 ( .a(n35944), .b(n41626), .c(n41491), .o(n41627) );
in01f01 g37836 ( .a(n41627), .o(n41628) );
na02f01 g37837 ( .a(n41628), .b(n41625), .o(n41629) );
no02f01 g37838 ( .a(n41560), .b(n41559), .o(n41630) );
ao12f01 g37839 ( .a(n35944), .b(n41566), .c(n41630), .o(n41631) );
no02f01 g37840 ( .a(n41631), .b(n41629), .o(n41632) );
no02f01 g37841 ( .a(n41586), .b(n41584), .o(n41633) );
ao12f01 g37842 ( .a(n35944), .b(n41633), .c(n41577), .o(n41634) );
in01f01 g37843 ( .a(n41634), .o(n41635) );
na02f01 g37844 ( .a(n41635), .b(n41632), .o(n41636) );
no02f01 g37845 ( .a(n41620), .b(n41618), .o(n41637) );
no02f01 g37846 ( .a(n41602), .b(n41601), .o(n41638) );
ao12f01 g37847 ( .a(n35944), .b(n41609), .c(n41638), .o(n41639) );
in01f01 g37848 ( .a(n41639), .o(n41640) );
ao12f01 g37849 ( .a(n35944), .b(n41640), .c(n41637), .o(n41641) );
no02f01 g37850 ( .a(n41641), .b(n41636), .o(n41642) );
in01f01 g37851 ( .a(n41642), .o(n41643) );
no03f01 g37852 ( .a(n41643), .b(n41624), .c(n41535), .o(n41644) );
na04f01 g37853 ( .a(n41622), .b(n41588), .c(n41546), .d(n39691), .o(n41645) );
ao12f01 g37854 ( .a(n41534), .b(n41642), .c(n41645), .o(n41646) );
oa12f01 g37855 ( .a(n32734), .b(n41646), .c(n41644), .o(n41647) );
na02f01 g37856 ( .a(n41647), .b(n41529), .o(n1392) );
in01f01 g37857 ( .a(n36872), .o(n41649) );
na04f01 g37858 ( .a(n41649), .b(n32436), .c(n32430), .d(n32427), .o(n41650) );
no02f01 g37859 ( .a(n36878), .b(n32440), .o(n41651) );
na02f01 g37860 ( .a(n36850), .b(n31606), .o(n41652) );
in01f01 g37861 ( .a(n41652), .o(n41653) );
no02f01 g37862 ( .a(n41653), .b(n36851), .o(n41654) );
na03f01 g37863 ( .a(n41654), .b(n41651), .c(n41650), .o(n41655) );
no04f01 g37864 ( .a(n36872), .b(n32495), .c(n32494), .d(n32493), .o(n41656) );
in01f01 g37865 ( .a(n41651), .o(n41657) );
in01f01 g37866 ( .a(n41654), .o(n41658) );
oa12f01 g37867 ( .a(n41658), .b(n41657), .c(n41656), .o(n41659) );
na02f01 g37868 ( .a(n41659), .b(n41655), .o(n1396) );
na03f01 g37869 ( .a(n16086), .b(n21354), .c(n16069), .o(n41661) );
oa12f01 g37870 ( .a(n21363), .b(n16070), .c(n21353), .o(n41662) );
na02f01 g37871 ( .a(n41662), .b(n41661), .o(n1401) );
no02f01 g37872 ( .a(n38133), .b(n38091), .o(n41664) );
no02f01 g37873 ( .a(n41664), .b(n38129), .o(n41665) );
oa12f01 g37874 ( .a(n38139), .b(n38134), .c(n6037), .o(n41666) );
no02f01 g37875 ( .a(n41666), .b(n41665), .o(n41667) );
no02f01 g37876 ( .a(n38103), .b(n6037), .o(n41668) );
no02f01 g37877 ( .a(n41668), .b(n38105), .o(n41669) );
na02f01 g37878 ( .a(n41669), .b(n41667), .o(n41670) );
in01f01 g37879 ( .a(n41669), .o(n41671) );
oa12f01 g37880 ( .a(n41671), .b(n41666), .c(n41665), .o(n41672) );
na02f01 g37881 ( .a(n41672), .b(n41670), .o(n1406) );
no02f01 g37882 ( .a(n21823), .b(n21816), .o(n41674) );
no02f01 g37883 ( .a(n36432), .b(n41674), .o(n41675) );
na02f01 g37884 ( .a(n36432), .b(n41674), .o(n41676) );
in01f01 g37885 ( .a(n41676), .o(n41677) );
no02f01 g37886 ( .a(n41677), .b(n41675), .o(n41678) );
in01f01 g37887 ( .a(n41678), .o(n41679) );
no02f01 g37888 ( .a(n22384), .b(n22383), .o(n41680) );
in01f01 g37889 ( .a(n41680), .o(n41681) );
no02f01 g37890 ( .a(n36447), .b(n41681), .o(n41682) );
in01f01 g37891 ( .a(n41682), .o(n41683) );
ao12f01 g37892 ( .a(n36432), .b(n21959), .c(n21835), .o(n41684) );
oa12f01 g37893 ( .a(n36447), .b(n41684), .c(n41681), .o(n41685) );
no03f01 g37894 ( .a(n36494), .b(n36481), .c(n36448), .o(n41686) );
no02f01 g37895 ( .a(n21959), .b(n21835), .o(n41687) );
no02f01 g37896 ( .a(n41687), .b(n36447), .o(n41688) );
in01f01 g37897 ( .a(n41688), .o(n41689) );
na03f01 g37898 ( .a(n41689), .b(n41686), .c(n36501), .o(n41690) );
no03f01 g37899 ( .a(n36494), .b(n36484), .c(n36472), .o(n41691) );
oa12f01 g37900 ( .a(n36510), .b(n36432), .c(n21954), .o(n41692) );
no02f01 g37901 ( .a(n41688), .b(n36448), .o(n41693) );
oa12f01 g37902 ( .a(n41693), .b(n41692), .c(n41691), .o(n41694) );
na03f01 g37903 ( .a(n41694), .b(n41690), .c(n41685), .o(n41695) );
na03f01 g37904 ( .a(n41695), .b(n41683), .c(n41679), .o(n41696) );
in01f01 g37905 ( .a(n41685), .o(n41697) );
na02f01 g37906 ( .a(n36432), .b(n21954), .o(n41698) );
na03f01 g37907 ( .a(n36512), .b(n36505), .c(n41698), .o(n41699) );
no03f01 g37908 ( .a(n41688), .b(n41699), .c(n36461), .o(n41700) );
na03f01 g37909 ( .a(n36512), .b(n36508), .c(n36475), .o(n41701) );
no02f01 g37910 ( .a(n36490), .b(n36433), .o(n41702) );
in01f01 g37911 ( .a(n41693), .o(n41703) );
ao12f01 g37912 ( .a(n41703), .b(n41702), .c(n41701), .o(n41704) );
no03f01 g37913 ( .a(n41704), .b(n41700), .c(n41697), .o(n41705) );
oa12f01 g37914 ( .a(n41678), .b(n41705), .c(n41682), .o(n41706) );
na03f01 g37915 ( .a(n41706), .b(n41696), .c(n2589), .o(n41707) );
no03f01 g37916 ( .a(n41705), .b(n41682), .c(n41678), .o(n41708) );
ao12f01 g37917 ( .a(n41679), .b(n41695), .c(n41683), .o(n41709) );
oa12f01 g37918 ( .a(n4116), .b(n41709), .c(n41708), .o(n41710) );
na02f01 g37919 ( .a(n41710), .b(n41707), .o(n1411) );
no02f01 g37920 ( .a(n5979), .b(n5873), .o(n41712) );
no02f01 g37921 ( .a(n41712), .b(n5981), .o(n41713) );
in01f01 g37922 ( .a(n41713), .o(n41714) );
na02f01 g37923 ( .a(n41714), .b(n38635), .o(n41715) );
na02f01 g37924 ( .a(n41713), .b(n5964), .o(n41716) );
na02f01 g37925 ( .a(n41716), .b(n41715), .o(n1416) );
no02f01 g37926 ( .a(n39856), .b(n29639), .o(n41718) );
in01f01 g37927 ( .a(n39856), .o(n41719) );
no02f01 g37928 ( .a(n41719), .b(n29430), .o(n41720) );
no02f01 g37929 ( .a(n41720), .b(n41718), .o(n41721) );
no03f01 g37930 ( .a(n36777), .b(n36737), .c(n36723), .o(n41722) );
in01f01 g37931 ( .a(n39280), .o(n41723) );
no02f01 g37932 ( .a(n41723), .b(n29430), .o(n41724) );
in01f01 g37933 ( .a(n39292), .o(n41725) );
no02f01 g37934 ( .a(n41725), .b(n29430), .o(n41726) );
no02f01 g37935 ( .a(n41726), .b(n41724), .o(n41727) );
in01f01 g37936 ( .a(n39307), .o(n41728) );
no02f01 g37937 ( .a(n41728), .b(n29430), .o(n41729) );
in01f01 g37938 ( .a(n41729), .o(n41730) );
na03f01 g37939 ( .a(n41730), .b(n41727), .c(n41722), .o(n41731) );
in01f01 g37940 ( .a(n41731), .o(n41732) );
oa12f01 g37941 ( .a(n41732), .b(n40452), .c(n40451), .o(n41733) );
oa12f01 g37942 ( .a(n29430), .b(n36736), .c(n36722), .o(n41734) );
na02f01 g37943 ( .a(n41734), .b(n36784), .o(n41735) );
no02f01 g37944 ( .a(n41725), .b(n41723), .o(n41736) );
ao12f01 g37945 ( .a(n29639), .b(n41736), .c(n39307), .o(n41737) );
no02f01 g37946 ( .a(n41737), .b(n41735), .o(n41738) );
na03f01 g37947 ( .a(n41738), .b(n41733), .c(n41721), .o(n41739) );
in01f01 g37948 ( .a(n41721), .o(n41740) );
ao12f01 g37949 ( .a(n41731), .b(n36783), .c(n40446), .o(n41741) );
in01f01 g37950 ( .a(n41738), .o(n41742) );
oa12f01 g37951 ( .a(n41740), .b(n41742), .c(n41741), .o(n41743) );
na03f01 g37952 ( .a(n41743), .b(n41739), .c(n_27923), .o(n41744) );
no03f01 g37953 ( .a(n41742), .b(n41741), .c(n41740), .o(n41745) );
ao12f01 g37954 ( .a(n41721), .b(n41738), .c(n41733), .o(n41746) );
oa12f01 g37955 ( .a(n34420), .b(n41746), .c(n41745), .o(n41747) );
na02f01 g37956 ( .a(n41747), .b(n41744), .o(n1421) );
no02f01 g37957 ( .a(n38389), .b(n39097), .o(n41749) );
no02f01 g37958 ( .a(n39101), .b(n38385), .o(n41750) );
no02f01 g37959 ( .a(n41750), .b(n41749), .o(n41751) );
na02f01 g37960 ( .a(n41751), .b(n38379), .o(n41752) );
oa12f01 g37961 ( .a(n39096), .b(n41750), .c(n41749), .o(n41753) );
na02f01 g37962 ( .a(n41753), .b(n41752), .o(n1426) );
in01f01 g37963 ( .a(n11632), .o(n41755) );
no02f01 g37964 ( .a(n11633), .b(n11598), .o(n41756) );
in01f01 g37965 ( .a(n41756), .o(n41757) );
na02f01 g37966 ( .a(n41757), .b(n41755), .o(n41758) );
na02f01 g37967 ( .a(n41756), .b(n11632), .o(n41759) );
na02f01 g37968 ( .a(n41759), .b(n41758), .o(n1431) );
no02f01 g37969 ( .a(n36119), .b(n36116), .o(n41761) );
in01f01 g37970 ( .a(n41761), .o(n41762) );
no02f01 g37971 ( .a(n36055), .b(n36122), .o(n41763) );
no02f01 g37972 ( .a(n36056), .b(n36038), .o(n41764) );
in01f01 g37973 ( .a(n41764), .o(n41765) );
ao12f01 g37974 ( .a(n41763), .b(n41765), .c(n41762), .o(n41766) );
no02f01 g37975 ( .a(n36048), .b(n36122), .o(n41767) );
no02f01 g37976 ( .a(n36049), .b(n36038), .o(n41768) );
no02f01 g37977 ( .a(n41768), .b(n41767), .o(n41769) );
na02f01 g37978 ( .a(n41769), .b(n41766), .o(n41770) );
in01f01 g37979 ( .a(n41766), .o(n41771) );
in01f01 g37980 ( .a(n41769), .o(n41772) );
na02f01 g37981 ( .a(n41772), .b(n41771), .o(n41773) );
na02f01 g37982 ( .a(n41773), .b(n41770), .o(n1436) );
in01f01 g37983 ( .a(n9607), .o(n41775) );
oa12f01 g37984 ( .a(n41775), .b(n9608), .c(n9606), .o(n41776) );
no02f01 g37985 ( .a(n41776), .b(n4201), .o(n41777) );
na02f01 g37986 ( .a(n41776), .b(n4201), .o(n41778) );
in01f01 g37987 ( .a(n41778), .o(n41779) );
no02f01 g37988 ( .a(n41779), .b(n41777), .o(n41780) );
na03f01 g37989 ( .a(n41780), .b(n9590), .c(n9589), .o(n41781) );
in01f01 g37990 ( .a(n41780), .o(n5215) );
oa12f01 g37991 ( .a(n5215), .b(n9646), .c(n9645), .o(n41783) );
na02f01 g37992 ( .a(n41783), .b(n41781), .o(n1441) );
na03f01 g37993 ( .a(n9855), .b(n9845), .c(n9832), .o(n41785) );
no02f01 g37994 ( .a(n9871), .b(n9869), .o(n41786) );
no02f01 g37995 ( .a(n9864), .b(n5001), .o(n41787) );
no02f01 g37996 ( .a(n41787), .b(n9866), .o(n41788) );
na03f01 g37997 ( .a(n41788), .b(n41786), .c(n41785), .o(n41789) );
na02f01 g37998 ( .a(n41786), .b(n41785), .o(n41790) );
in01f01 g37999 ( .a(n41788), .o(n41791) );
na02f01 g38000 ( .a(n41791), .b(n41790), .o(n41792) );
na02f01 g38001 ( .a(n41792), .b(n41789), .o(n1446) );
na02f01 g38002 ( .a(n1080), .b(n4116), .o(n41794) );
na02f01 g38003 ( .a(n40459), .b(n2589), .o(n41795) );
na02f01 g38004 ( .a(n41795), .b(n41794), .o(n1451) );
in01f01 g38005 ( .a(n26846), .o(n41797) );
in01f01 g38006 ( .a(n26756), .o(n41798) );
no02f01 g38007 ( .a(n26755), .b(n26440), .o(n41799) );
no02f01 g38008 ( .a(n41799), .b(n41798), .o(n41800) );
no02f01 g38009 ( .a(n26845), .b(n26440), .o(n41801) );
in01f01 g38010 ( .a(n26839), .o(n41802) );
ao12f01 g38011 ( .a(n41802), .b(n27247), .c(n38553), .o(n41803) );
no03f01 g38012 ( .a(n41803), .b(n27121), .c(n41801), .o(n41804) );
oa12f01 g38013 ( .a(n41800), .b(n41804), .c(n41797), .o(n41805) );
in01f01 g38014 ( .a(n41800), .o(n41806) );
in01f01 g38015 ( .a(n41801), .o(n41807) );
in01f01 g38016 ( .a(n27121), .o(n41808) );
oa12f01 g38017 ( .a(n26839), .b(n27119), .c(n38561), .o(n41809) );
na03f01 g38018 ( .a(n41809), .b(n41808), .c(n41807), .o(n41810) );
na03f01 g38019 ( .a(n41810), .b(n41806), .c(n26846), .o(n41811) );
na03f01 g38020 ( .a(n41811), .b(n41805), .c(n1821), .o(n41812) );
ao12f01 g38021 ( .a(n41806), .b(n41810), .c(n26846), .o(n41813) );
no03f01 g38022 ( .a(n41804), .b(n41800), .c(n41797), .o(n41814) );
oa12f01 g38023 ( .a(n8066), .b(n41814), .c(n41813), .o(n41815) );
na02f01 g38024 ( .a(n41815), .b(n41812), .o(n1456) );
no02f01 g38025 ( .a(n32382), .b(n32473), .o(n41817) );
oa12f01 g38026 ( .a(n41817), .b(n32476), .c(n32234), .o(n41818) );
in01f01 g38027 ( .a(n41817), .o(n41819) );
na03f01 g38028 ( .a(n32384), .b(n41819), .c(n32235), .o(n41820) );
na02f01 g38029 ( .a(n41820), .b(n41818), .o(n1461) );
no02f01 g38030 ( .a(n7512), .b(n7530), .o(n41822) );
no02f01 g38031 ( .a(n7538), .b(n7499), .o(n41823) );
oa12f01 g38032 ( .a(n7533), .b(n41823), .c(n41822), .o(n41824) );
no02f01 g38033 ( .a(n41823), .b(n41822), .o(n41825) );
na02f01 g38034 ( .a(n41825), .b(n7507), .o(n41826) );
na02f01 g38035 ( .a(n41826), .b(n41824), .o(n1466) );
na03f01 g38036 ( .a(n41015), .b(n39152), .c(n39142), .o(n41828) );
no02f01 g38037 ( .a(n41026), .b(n39160), .o(n41829) );
no02f01 g38038 ( .a(n39135), .b(n31569), .o(n41830) );
in01f01 g38039 ( .a(n31569), .o(n41831) );
no02f01 g38040 ( .a(n39059), .b(n41831), .o(n41832) );
no02f01 g38041 ( .a(n41832), .b(n41830), .o(n41833) );
na03f01 g38042 ( .a(n41833), .b(n41829), .c(n41828), .o(n41834) );
no03f01 g38043 ( .a(n41016), .b(n39151), .c(n39172), .o(n41835) );
in01f01 g38044 ( .a(n41829), .o(n41836) );
in01f01 g38045 ( .a(n41833), .o(n41837) );
oa12f01 g38046 ( .a(n41837), .b(n41836), .c(n41835), .o(n41838) );
na03f01 g38047 ( .a(n41838), .b(n41834), .c(n3633), .o(n41839) );
na02f01 g38048 ( .a(n41838), .b(n41834), .o(n5330) );
na02f01 g38049 ( .a(n5330), .b(n6203), .o(n41841) );
na02f01 g38050 ( .a(n41841), .b(n41839), .o(n1471) );
in01f01 g38051 ( .a(n8614), .o(n41843) );
in01f01 g38052 ( .a(n8662), .o(n41844) );
no02f01 g38053 ( .a(n8612), .b(n5973), .o(n41845) );
in01f01 g38054 ( .a(n41845), .o(n41846) );
na02f01 g38055 ( .a(n41846), .b(n41844), .o(n41847) );
ao12f01 g38056 ( .a(n41847), .b(n41843), .c(n8604), .o(n41848) );
no02f01 g38057 ( .a(n8663), .b(n5973), .o(n41849) );
no02f01 g38058 ( .a(n41849), .b(n8624), .o(n41850) );
na02f01 g38059 ( .a(n41850), .b(n41848), .o(n41851) );
in01f01 g38060 ( .a(n41848), .o(n41852) );
in01f01 g38061 ( .a(n41850), .o(n41853) );
na02f01 g38062 ( .a(n41853), .b(n41852), .o(n41854) );
na02f01 g38063 ( .a(n41854), .b(n41851), .o(n1476) );
in01f01 g38064 ( .a(n11765), .o(n41856) );
no02f01 g38065 ( .a(n11775), .b(n41856), .o(n41857) );
in01f01 g38066 ( .a(n41857), .o(n41858) );
in01f01 g38067 ( .a(n11802), .o(n41859) );
no02f01 g38068 ( .a(n11803), .b(n11785), .o(n41860) );
na03f01 g38069 ( .a(n41860), .b(n41859), .c(n41858), .o(n41861) );
in01f01 g38070 ( .a(n41860), .o(n41862) );
oa12f01 g38071 ( .a(n41862), .b(n11802), .c(n41857), .o(n41863) );
na02f01 g38072 ( .a(n41863), .b(n41861), .o(n1481) );
no02f01 g38073 ( .a(n17935), .b(n17930), .o(n41865) );
no02f01 g38074 ( .a(n17954), .b(n17931), .o(n41866) );
no02f01 g38075 ( .a(n41866), .b(n41865), .o(n41867) );
na02f01 g38076 ( .a(n41867), .b(n17950), .o(n41868) );
oa12f01 g38077 ( .a(n17923), .b(n41866), .c(n41865), .o(n41869) );
na02f01 g38078 ( .a(n41869), .b(n41868), .o(n1486) );
no02f01 g38079 ( .a(n39135), .b(n31596), .o(n41871) );
no02f01 g38080 ( .a(n41871), .b(n41018), .o(n41872) );
no03f01 g38081 ( .a(n41836), .b(n41835), .c(n41027), .o(n41873) );
oa12f01 g38082 ( .a(n41872), .b(n41873), .c(n41020), .o(n41874) );
in01f01 g38083 ( .a(n41020), .o(n41875) );
in01f01 g38084 ( .a(n41872), .o(n41876) );
na03f01 g38085 ( .a(n41829), .b(n41828), .c(n41028), .o(n41877) );
na03f01 g38086 ( .a(n41877), .b(n41876), .c(n41875), .o(n41878) );
na03f01 g38087 ( .a(n41878), .b(n41874), .c(n3633), .o(n41879) );
ao12f01 g38088 ( .a(n41876), .b(n41877), .c(n41875), .o(n41880) );
no03f01 g38089 ( .a(n41873), .b(n41872), .c(n41020), .o(n41881) );
oa12f01 g38090 ( .a(n6203), .b(n41881), .c(n41880), .o(n41882) );
na02f01 g38091 ( .a(n41882), .b(n41879), .o(n1491) );
no03f01 g38092 ( .a(n40303), .b(n38161), .c(n38160), .o(n41884) );
ao12f01 g38093 ( .a(n40310), .b(n40302), .c(n38142), .o(n41885) );
in01f01 g38094 ( .a(n41885), .o(n41886) );
no03f01 g38095 ( .a(n41886), .b(n41884), .c(n40313), .o(n41887) );
no02f01 g38096 ( .a(n40312), .b(n6037), .o(n41888) );
no02f01 g38097 ( .a(n41888), .b(n40257), .o(n41889) );
oa12f01 g38098 ( .a(n41889), .b(n41887), .c(n40265), .o(n41890) );
in01f01 g38099 ( .a(n40265), .o(n41891) );
na03f01 g38100 ( .a(n40302), .b(n38130), .c(n38091), .o(n41892) );
na03f01 g38101 ( .a(n41885), .b(n41892), .c(n40314), .o(n41893) );
in01f01 g38102 ( .a(n41889), .o(n41894) );
na03f01 g38103 ( .a(n41894), .b(n41893), .c(n41891), .o(n41895) );
na02f01 g38104 ( .a(n41895), .b(n41890), .o(n1496) );
ao12f01 g38105 ( .a(n6005), .b(n5982), .c(n38635), .o(n41897) );
no02f01 g38106 ( .a(n6000), .b(n5873), .o(n41898) );
no02f01 g38107 ( .a(n41898), .b(n6002), .o(n41899) );
na02f01 g38108 ( .a(n41899), .b(n41897), .o(n41900) );
in01f01 g38109 ( .a(n41897), .o(n41901) );
in01f01 g38110 ( .a(n41899), .o(n41902) );
na02f01 g38111 ( .a(n41902), .b(n41901), .o(n41903) );
na02f01 g38112 ( .a(n41903), .b(n41900), .o(n1501) );
in01f01 g38113 ( .a(n14210), .o(n41905) );
no02f01 g38114 ( .a(n14211), .b(n14006), .o(n41906) );
in01f01 g38115 ( .a(n41906), .o(n41907) );
no03f01 g38116 ( .a(n41907), .b(n41905), .c(n14020), .o(n41908) );
ao12f01 g38117 ( .a(n41906), .b(n14210), .c(n14021), .o(n41909) );
no02f01 g38118 ( .a(n41909), .b(n41908), .o(n41910) );
na02f01 g38119 ( .a(n41910), .b(n2589), .o(n41911) );
in01f01 g38120 ( .a(n41910), .o(n5430) );
na02f01 g38121 ( .a(n5430), .b(n4116), .o(n41913) );
na02f01 g38122 ( .a(n41913), .b(n41911), .o(n1506) );
in01f01 g38123 ( .a(n27192), .o(n41915) );
in01f01 g38124 ( .a(n27193), .o(n41916) );
no02f01 g38125 ( .a(n27183), .b(n26440), .o(n41917) );
no02f01 g38126 ( .a(n41917), .b(n41916), .o(n41918) );
no02f01 g38127 ( .a(n27189), .b(n26440), .o(n41919) );
no03f01 g38128 ( .a(n41919), .b(n27172), .c(n27166), .o(n41920) );
oa12f01 g38129 ( .a(n41918), .b(n41920), .c(n41915), .o(n41921) );
in01f01 g38130 ( .a(n41918), .o(n41922) );
in01f01 g38131 ( .a(n41919), .o(n41923) );
na03f01 g38132 ( .a(n41923), .b(n27171), .c(n27249), .o(n41924) );
na03f01 g38133 ( .a(n41924), .b(n41922), .c(n27192), .o(n41925) );
na02f01 g38134 ( .a(n41925), .b(n41921), .o(n1511) );
no02f01 g38135 ( .a(n8667), .b(n8644), .o(n41927) );
na03f01 g38136 ( .a(n41927), .b(n8665), .c(n39007), .o(n41928) );
in01f01 g38137 ( .a(n41927), .o(n41929) );
na02f01 g38138 ( .a(n41929), .b(n41146), .o(n41930) );
na02f01 g38139 ( .a(n41930), .b(n41928), .o(n1516) );
in01f01 g38140 ( .a(n22195), .o(n41932) );
na03f01 g38141 ( .a(n22235), .b(n22234), .c(n41932), .o(n41933) );
in01f01 g38142 ( .a(n22234), .o(n41934) );
in01f01 g38143 ( .a(n22235), .o(n41935) );
oa12f01 g38144 ( .a(n41934), .b(n41935), .c(n22195), .o(n41936) );
na02f01 g38145 ( .a(n41936), .b(n41933), .o(n1521) );
no02f01 g38146 ( .a(n21190), .b(n21119), .o(n41938) );
in01f01 g38147 ( .a(n21199), .o(n41939) );
in01f01 g38148 ( .a(n21203), .o(n41940) );
ao12f01 g38149 ( .a(n41939), .b(n41940), .c(n41938), .o(n41941) );
in01f01 g38150 ( .a(n41941), .o(n41942) );
no02f01 g38151 ( .a(n21202), .b(n21107), .o(n41943) );
na02f01 g38152 ( .a(n41943), .b(n41942), .o(n41944) );
in01f01 g38153 ( .a(n41943), .o(n41945) );
na02f01 g38154 ( .a(n41945), .b(n41941), .o(n41946) );
na02f01 g38155 ( .a(n41946), .b(n41944), .o(n1531) );
no02f01 g38156 ( .a(n35433), .b(n4176), .o(n41948) );
no02f01 g38157 ( .a(n35435), .b(n35414), .o(n41949) );
no03f01 g38158 ( .a(n41949), .b(n35439), .c(n41948), .o(n41950) );
no02f01 g38159 ( .a(n35426), .b(n4176), .o(n41951) );
no02f01 g38160 ( .a(n41951), .b(n35428), .o(n41952) );
na02f01 g38161 ( .a(n41952), .b(n41950), .o(n41953) );
in01f01 g38162 ( .a(n41950), .o(n41954) );
in01f01 g38163 ( .a(n41952), .o(n41955) );
na02f01 g38164 ( .a(n41955), .b(n41954), .o(n41956) );
na02f01 g38165 ( .a(n41956), .b(n41953), .o(n1536) );
in01f01 g38166 ( .a(n35370), .o(n41958) );
in01f01 g38167 ( .a(n38984), .o(n41959) );
na02f01 g38168 ( .a(n41959), .b(n38983), .o(n41960) );
ao12f01 g38169 ( .a(n41960), .b(n41958), .c(n38981), .o(n41961) );
no02f01 g38170 ( .a(n35380), .b(n4176), .o(n41962) );
no02f01 g38171 ( .a(n41962), .b(n35382), .o(n41963) );
na02f01 g38172 ( .a(n41963), .b(n41961), .o(n41964) );
in01f01 g38173 ( .a(n41961), .o(n41965) );
in01f01 g38174 ( .a(n41963), .o(n41966) );
na02f01 g38175 ( .a(n41966), .b(n41965), .o(n41967) );
na02f01 g38176 ( .a(n41967), .b(n41964), .o(n1545) );
in01f01 g38177 ( .a(n22049), .o(n41969) );
no02f01 g38178 ( .a(n36419), .b(n36418), .o(n41970) );
no02f01 g38179 ( .a(n41970), .b(n22050), .o(n41971) );
na02f01 g38180 ( .a(n41970), .b(n22050), .o(n41972) );
in01f01 g38181 ( .a(n41972), .o(n41973) );
no02f01 g38182 ( .a(n41973), .b(n41971), .o(n41974) );
in01f01 g38183 ( .a(n41974), .o(n41975) );
ao12f01 g38184 ( .a(n22050), .b(n22448), .c(n22053), .o(n41976) );
in01f01 g38185 ( .a(n41976), .o(n41977) );
oa12f01 g38186 ( .a(n41977), .b(n22453), .c(n22426), .o(n41978) );
ao12f01 g38187 ( .a(n41975), .b(n41978), .c(n41969), .o(n41979) );
ao12f01 g38188 ( .a(n41976), .b(n22454), .c(n22484), .o(n41980) );
no03f01 g38189 ( .a(n41980), .b(n41974), .c(n22049), .o(n41981) );
oa12f01 g38190 ( .a(n4116), .b(n41981), .c(n41979), .o(n41982) );
oa12f01 g38191 ( .a(n41974), .b(n41980), .c(n22049), .o(n41983) );
na03f01 g38192 ( .a(n41978), .b(n41975), .c(n41969), .o(n41984) );
na03f01 g38193 ( .a(n41984), .b(n41983), .c(n2589), .o(n41985) );
na02f01 g38194 ( .a(n41985), .b(n41982), .o(n1550) );
in01f01 g38195 ( .a(n10994), .o(n41987) );
no03f01 g38196 ( .a(n38067), .b(n11007), .c(n41987), .o(n41988) );
in01f01 g38197 ( .a(n41988), .o(n41989) );
no02f01 g38198 ( .a(n38062), .b(n10681), .o(n41990) );
oa12f01 g38199 ( .a(n41990), .b(n38059), .c(n10677), .o(n41991) );
in01f01 g38200 ( .a(n41991), .o(n41992) );
no02f01 g38201 ( .a(n10682), .b(n4088), .o(n41993) );
no02f01 g38202 ( .a(n41993), .b(n10668), .o(n41994) );
no02f01 g38203 ( .a(n41994), .b(n41992), .o(n41995) );
na02f01 g38204 ( .a(n41994), .b(n41992), .o(n41996) );
in01f01 g38205 ( .a(n41996), .o(n41997) );
no02f01 g38206 ( .a(n41997), .b(n41995), .o(n41998) );
in01f01 g38207 ( .a(n41998), .o(n41999) );
no02f01 g38208 ( .a(n10696), .b(n4088), .o(n42000) );
no02f01 g38209 ( .a(n42000), .b(n10698), .o(n42001) );
in01f01 g38210 ( .a(n42001), .o(n42002) );
no02f01 g38211 ( .a(n42002), .b(n10686), .o(n42003) );
in01f01 g38212 ( .a(n10686), .o(n42004) );
no02f01 g38213 ( .a(n42001), .b(n42004), .o(n42005) );
no02f01 g38214 ( .a(n42005), .b(n42003), .o(n42006) );
in01f01 g38215 ( .a(n42006), .o(n42007) );
ao12f01 g38216 ( .a(n10735), .b(n42007), .c(n41999), .o(n42008) );
no04f01 g38217 ( .a(n42008), .b(n41989), .c(n10988), .d(n10976), .o(n42009) );
in01f01 g38218 ( .a(n42009), .o(n42010) );
ao12f01 g38219 ( .a(n3521), .b(n38068), .c(n11005), .o(n42011) );
no02f01 g38220 ( .a(n42011), .b(n10796), .o(n42012) );
in01f01 g38221 ( .a(n42012), .o(n42013) );
ao12f01 g38222 ( .a(n3521), .b(n42006), .c(n41998), .o(n42014) );
no02f01 g38223 ( .a(n42014), .b(n42013), .o(n42015) );
no02f01 g38224 ( .a(n10698), .b(n42004), .o(n42016) );
no02f01 g38225 ( .a(n10707), .b(n4088), .o(n42017) );
no02f01 g38226 ( .a(n42017), .b(n10709), .o(n42018) );
in01f01 g38227 ( .a(n42018), .o(n42019) );
no03f01 g38228 ( .a(n42019), .b(n42000), .c(n42016), .o(n42020) );
no02f01 g38229 ( .a(n42000), .b(n42016), .o(n42021) );
no02f01 g38230 ( .a(n42018), .b(n42021), .o(n42022) );
no03f01 g38231 ( .a(n42022), .b(n42020), .c(n10735), .o(n42023) );
no02f01 g38232 ( .a(n42022), .b(n42020), .o(n42024) );
no02f01 g38233 ( .a(n42024), .b(n3521), .o(n42025) );
no02f01 g38234 ( .a(n42025), .b(n42023), .o(n42026) );
na03f01 g38235 ( .a(n42026), .b(n42015), .c(n42010), .o(n42027) );
in01f01 g38236 ( .a(n42015), .o(n42028) );
in01f01 g38237 ( .a(n42026), .o(n42029) );
oa12f01 g38238 ( .a(n42029), .b(n42028), .c(n42009), .o(n42030) );
na02f01 g38239 ( .a(n42030), .b(n42027), .o(n1555) );
in01f01 g38240 ( .a(n8532), .o(n42032) );
in01f01 g38241 ( .a(n8536), .o(n42033) );
no02f01 g38242 ( .a(n8558), .b(n8544), .o(n42034) );
in01f01 g38243 ( .a(n42034), .o(n42035) );
oa12f01 g38244 ( .a(n42035), .b(n42033), .c(n42032), .o(n42036) );
no02f01 g38245 ( .a(n42033), .b(n42032), .o(n42037) );
na02f01 g38246 ( .a(n42034), .b(n42037), .o(n42038) );
na02f01 g38247 ( .a(n42038), .b(n42036), .o(n1560) );
na02f01 g38248 ( .a(n25420), .b(n25419), .o(n42040) );
na02f01 g38249 ( .a(n25424), .b(n42040), .o(n42041) );
na02f01 g38250 ( .a(n42041), .b(n25426), .o(n1565) );
in01f01 g38251 ( .a(n37250), .o(n42043) );
no02f01 g38252 ( .a(n37184), .b(n37182), .o(n42044) );
in01f01 g38253 ( .a(n42044), .o(n42045) );
no02f01 g38254 ( .a(n37192), .b(n36963), .o(n42046) );
no02f01 g38255 ( .a(n42046), .b(n37194), .o(n42047) );
na03f01 g38256 ( .a(n42047), .b(n42045), .c(n42043), .o(n42048) );
in01f01 g38257 ( .a(n42047), .o(n42049) );
oa12f01 g38258 ( .a(n42049), .b(n42044), .c(n37250), .o(n42050) );
na02f01 g38259 ( .a(n42050), .b(n42048), .o(n1570) );
in01f01 g38260 ( .a(n14129), .o(n42052) );
in01f01 g38261 ( .a(n14152), .o(n42053) );
na03f01 g38262 ( .a(n42053), .b(n14130), .c(n42052), .o(n42054) );
in01f01 g38263 ( .a(n14130), .o(n42055) );
oa12f01 g38264 ( .a(n14152), .b(n42055), .c(n14129), .o(n42056) );
na02f01 g38265 ( .a(n42056), .b(n42054), .o(n1575) );
no03f01 g38266 ( .a(n40931), .b(n40929), .c(n40875), .o(n42058) );
no02f01 g38267 ( .a(n42058), .b(n40884), .o(n42059) );
in01f01 g38268 ( .a(n40864), .o(n42060) );
no02f01 g38269 ( .a(n40885), .b(n42060), .o(n42061) );
no02f01 g38270 ( .a(n42061), .b(n42059), .o(n42062) );
na02f01 g38271 ( .a(n42061), .b(n42059), .o(n42063) );
in01f01 g38272 ( .a(n42063), .o(n42064) );
no02f01 g38273 ( .a(n42064), .b(n42062), .o(n42065) );
in01f01 g38274 ( .a(n42065), .o(n1580) );
na04f01 g38275 ( .a(n39119), .b(n38437), .c(n38324), .d(n39077), .o(n42067) );
oa22f01 g38276 ( .a(n38441), .b(n38296), .c(n39118), .d(n39087), .o(n42068) );
na02f01 g38277 ( .a(n42068), .b(n42067), .o(n1585) );
no02f01 g38278 ( .a(n37208), .b(n37182), .o(n42070) );
in01f01 g38279 ( .a(n37228), .o(n42071) );
no02f01 g38280 ( .a(n37226), .b(n36963), .o(n42072) );
in01f01 g38281 ( .a(n42072), .o(n42073) );
na02f01 g38282 ( .a(n42073), .b(n37252), .o(n42074) );
ao12f01 g38283 ( .a(n42074), .b(n42071), .c(n42070), .o(n42075) );
no02f01 g38284 ( .a(n37219), .b(n36963), .o(n42076) );
no02f01 g38285 ( .a(n42076), .b(n37221), .o(n42077) );
na02f01 g38286 ( .a(n42077), .b(n42075), .o(n42078) );
in01f01 g38287 ( .a(n42075), .o(n42079) );
in01f01 g38288 ( .a(n42077), .o(n42080) );
na02f01 g38289 ( .a(n42080), .b(n42079), .o(n42081) );
na02f01 g38290 ( .a(n42081), .b(n42078), .o(n1590) );
na02f01 g38291 ( .a(n37343), .b(n37341), .o(n1595) );
oa12f01 g38292 ( .a(n27024), .b(n27222), .c(n27012), .o(n42084) );
na03f01 g38293 ( .a(n27025), .b(n27221), .c(n27213), .o(n42085) );
na02f01 g38294 ( .a(n42085), .b(n42084), .o(n1600) );
in01f01 g38295 ( .a(n14195), .o(n42087) );
no02f01 g38296 ( .a(n14197), .b(n14071), .o(n42088) );
no02f01 g38297 ( .a(n42088), .b(n42087), .o(n42089) );
na02f01 g38298 ( .a(n42088), .b(n42087), .o(n42090) );
in01f01 g38299 ( .a(n42090), .o(n42091) );
no02f01 g38300 ( .a(n42091), .b(n42089), .o(n42092) );
in01f01 g38301 ( .a(n42092), .o(n1729) );
na02f01 g38302 ( .a(n1729), .b(n4116), .o(n42094) );
na02f01 g38303 ( .a(n42092), .b(n2589), .o(n42095) );
na02f01 g38304 ( .a(n42095), .b(n42094), .o(n1605) );
in01f01 g38305 ( .a(n38015), .o(n42097) );
no02f01 g38306 ( .a(n37871), .b(n26361), .o(n42098) );
no02f01 g38307 ( .a(n42098), .b(n40986), .o(n42099) );
in01f01 g38308 ( .a(n42099), .o(n42100) );
oa12f01 g38309 ( .a(n38013), .b(n37871), .c(n26388), .o(n42101) );
na03f01 g38310 ( .a(n42101), .b(n42100), .c(n42097), .o(n42102) );
no02f01 g38311 ( .a(n38014), .b(n38049), .o(n42103) );
oa12f01 g38312 ( .a(n42099), .b(n42103), .c(n38015), .o(n42104) );
na02f01 g38313 ( .a(n42104), .b(n42102), .o(n1610) );
na03f01 g38314 ( .a(n36641), .b(n25462), .c(n25402), .o(n42106) );
oa12f01 g38315 ( .a(n36638), .b(n25463), .c(n36630), .o(n42107) );
na02f01 g38316 ( .a(n42107), .b(n42106), .o(n1615) );
no02f01 g38317 ( .a(n29917), .b(n25023), .o(n42109) );
no02f01 g38318 ( .a(n42109), .b(n25171), .o(n42110) );
in01f01 g38319 ( .a(n42110), .o(n42111) );
in01f01 g38320 ( .a(n25544), .o(n42112) );
oa12f01 g38321 ( .a(n42112), .b(n41516), .c(n25159), .o(n42113) );
na03f01 g38322 ( .a(n42113), .b(n42111), .c(n25180), .o(n42114) );
ao12f01 g38323 ( .a(n25544), .b(n41510), .c(n41513), .o(n42115) );
oa12f01 g38324 ( .a(n42110), .b(n42115), .c(n25181), .o(n42116) );
na02f01 g38325 ( .a(n42116), .b(n42114), .o(n1620) );
no02f01 g38326 ( .a(n37871), .b(n41223), .o(n42118) );
na02f01 g38327 ( .a(n37871), .b(n41223), .o(n42119) );
in01f01 g38328 ( .a(n42119), .o(n42120) );
no02f01 g38329 ( .a(n42120), .b(n42118), .o(n42121) );
in01f01 g38330 ( .a(n40991), .o(n42122) );
oa12f01 g38331 ( .a(n42122), .b(n40992), .c(n40995), .o(n42123) );
na02f01 g38332 ( .a(n42123), .b(n42121), .o(n42124) );
no02f01 g38333 ( .a(n42123), .b(n42121), .o(n42125) );
in01f01 g38334 ( .a(n42125), .o(n42126) );
na02f01 g38335 ( .a(n42126), .b(n42124), .o(n1625) );
in01f01 g38336 ( .a(n29772), .o(n42128) );
in01f01 g38337 ( .a(n29811), .o(n42129) );
na03f01 g38338 ( .a(n29812), .b(n42129), .c(n42128), .o(n42130) );
in01f01 g38339 ( .a(n29812), .o(n42131) );
oa12f01 g38340 ( .a(n29811), .b(n42131), .c(n29772), .o(n42132) );
na02f01 g38341 ( .a(n42132), .b(n42130), .o(n1630) );
no02f01 g38342 ( .a(n29611), .b(n29639), .o(n42134) );
no02f01 g38343 ( .a(n42134), .b(n29613), .o(n42135) );
in01f01 g38344 ( .a(n29600), .o(n42136) );
ao12f01 g38345 ( .a(n29639), .b(n29643), .c(n29598), .o(n42137) );
ao12f01 g38346 ( .a(n42137), .b(n42136), .c(n29721), .o(n42138) );
na02f01 g38347 ( .a(n42138), .b(n42135), .o(n42139) );
in01f01 g38348 ( .a(n42135), .o(n42140) );
in01f01 g38349 ( .a(n42138), .o(n42141) );
na02f01 g38350 ( .a(n42141), .b(n42140), .o(n42142) );
na02f01 g38351 ( .a(n42142), .b(n42139), .o(n1635) );
no02f01 g38352 ( .a(n35389), .b(n35385), .o(n42144) );
in01f01 g38353 ( .a(n42144), .o(n42145) );
in01f01 g38354 ( .a(n35412), .o(n42146) );
no02f01 g38355 ( .a(n35410), .b(n4176), .o(n42147) );
ao12f01 g38356 ( .a(n42147), .b(n42146), .c(n42145), .o(n42148) );
no02f01 g38357 ( .a(n35402), .b(n4176), .o(n42149) );
no02f01 g38358 ( .a(n42149), .b(n35404), .o(n42150) );
na02f01 g38359 ( .a(n42150), .b(n42148), .o(n42151) );
in01f01 g38360 ( .a(n42148), .o(n42152) );
in01f01 g38361 ( .a(n42150), .o(n42153) );
na02f01 g38362 ( .a(n42153), .b(n42152), .o(n42154) );
na02f01 g38363 ( .a(n42154), .b(n42151), .o(n1640) );
in01f01 g38364 ( .a(mux_while_ln12_psv_q_7_), .o(n42156) );
no03f01 g38365 ( .a(n41416), .b(n42156), .c(n41414), .o(n1650) );
no02f01 g38366 ( .a(n40931), .b(n40882), .o(n42158) );
in01f01 g38367 ( .a(n42158), .o(n42159) );
ao12f01 g38368 ( .a(n42159), .b(n40928), .c(n40898), .o(n42160) );
no02f01 g38369 ( .a(n42158), .b(n40929), .o(n42161) );
no02f01 g38370 ( .a(n42161), .b(n42160), .o(n42162) );
na02f01 g38371 ( .a(n42162), .b(n5799), .o(n42163) );
in01f01 g38372 ( .a(n42162), .o(n4488) );
na02f01 g38373 ( .a(n4488), .b(n911), .o(n42165) );
na02f01 g38374 ( .a(n42165), .b(n42163), .o(n1655) );
no02f01 g38375 ( .a(n9646), .b(n9587), .o(n42167) );
na03f01 g38376 ( .a(n42167), .b(n9644), .c(n9643), .o(n42168) );
in01f01 g38377 ( .a(n42167), .o(n42169) );
oa12f01 g38378 ( .a(n42169), .b(n9585), .c(n9578), .o(n42170) );
na02f01 g38379 ( .a(n42170), .b(n42168), .o(n1660) );
in01f01 g38380 ( .a(n10776), .o(n42172) );
no02f01 g38381 ( .a(n10989), .b(n42172), .o(n42173) );
no02f01 g38382 ( .a(n42173), .b(n10991), .o(n42174) );
no02f01 g38383 ( .a(n42174), .b(n10787), .o(n42175) );
no02f01 g38384 ( .a(n10993), .b(n10794), .o(n42176) );
na02f01 g38385 ( .a(n42176), .b(n42175), .o(n42177) );
in01f01 g38386 ( .a(n42176), .o(n42178) );
oa12f01 g38387 ( .a(n42178), .b(n42174), .c(n10787), .o(n42179) );
na02f01 g38388 ( .a(n42179), .b(n42177), .o(n1669) );
ao12f01 g38389 ( .a(n30091), .b(n25890), .c(n30090), .o(n42181) );
in01f01 g38390 ( .a(n42181), .o(n42182) );
no02f01 g38391 ( .a(n25883), .b(n25800), .o(n42183) );
no02f01 g38392 ( .a(n25884), .b(n30068), .o(n42184) );
no02f01 g38393 ( .a(n42184), .b(n42183), .o(n42185) );
na02f01 g38394 ( .a(n42185), .b(n42182), .o(n42186) );
oa12f01 g38395 ( .a(n42181), .b(n42184), .c(n42183), .o(n42187) );
na02f01 g38396 ( .a(n42187), .b(n42186), .o(n1674) );
in01f01 g38397 ( .a(n37278), .o(n42189) );
ao12f01 g38398 ( .a(delay_sub_ln23_0_unr23_stage8_stallmux_q), .b(n41103), .c(n41102), .o(n42190) );
ao12f01 g38399 ( .a(n37149), .b(n41103), .c(n41102), .o(n42191) );
no02f01 g38400 ( .a(n42191), .b(n42190), .o(n42192) );
in01f01 g38401 ( .a(n42192), .o(n42193) );
na03f01 g38402 ( .a(n42193), .b(n37345), .c(n42189), .o(n42194) );
oa12f01 g38403 ( .a(n42192), .b(n37366), .c(n37278), .o(n42195) );
na02f01 g38404 ( .a(n42195), .b(n42194), .o(n1679) );
no04f01 g38405 ( .a(n40933), .b(n40887), .c(n40843), .d(n40827), .o(n42197) );
no02f01 g38406 ( .a(n40933), .b(n40887), .o(n42198) );
no02f01 g38407 ( .a(n40843), .b(n40827), .o(n42199) );
no02f01 g38408 ( .a(n42199), .b(n42198), .o(n42200) );
no02f01 g38409 ( .a(n42200), .b(n42197), .o(n42201) );
na02f01 g38410 ( .a(n42201), .b(n5799), .o(n42202) );
in01f01 g38411 ( .a(n42201), .o(n5474) );
na02f01 g38412 ( .a(n5474), .b(n911), .o(n42204) );
na02f01 g38413 ( .a(n42204), .b(n42202), .o(n1684) );
ao12f01 g38414 ( .a(n25723), .b(n25922), .c(n30109), .o(n42206) );
no02f01 g38415 ( .a(n29998), .b(n29994), .o(n42207) );
in01f01 g38416 ( .a(n42207), .o(n42208) );
no02f01 g38417 ( .a(n42208), .b(n42206), .o(n42209) );
na02f01 g38418 ( .a(n42208), .b(n42206), .o(n42210) );
in01f01 g38419 ( .a(n42210), .o(n42211) );
no02f01 g38420 ( .a(n42211), .b(n42209), .o(n42212) );
in01f01 g38421 ( .a(n42212), .o(n1689) );
no02f01 g38422 ( .a(n10768), .b(n3521), .o(n42214) );
in01f01 g38423 ( .a(n42214), .o(n42215) );
oa12f01 g38424 ( .a(n42215), .b(n10980), .c(n10976), .o(n42216) );
in01f01 g38425 ( .a(n42216), .o(n42217) );
no02f01 g38426 ( .a(n10774), .b(n3521), .o(n42218) );
no02f01 g38427 ( .a(n42218), .b(n10978), .o(n42219) );
na02f01 g38428 ( .a(n42219), .b(n42217), .o(n42220) );
in01f01 g38429 ( .a(n42219), .o(n42221) );
na02f01 g38430 ( .a(n42221), .b(n42216), .o(n42222) );
na02f01 g38431 ( .a(n42222), .b(n42220), .o(n1694) );
in01f01 g38432 ( .a(n9240), .o(n42224) );
no02f01 g38433 ( .a(n40556), .b(n42224), .o(n42225) );
na02f01 g38434 ( .a(n40556), .b(n42224), .o(n42226) );
in01f01 g38435 ( .a(n42226), .o(n42227) );
no02f01 g38436 ( .a(n42227), .b(n42225), .o(n42228) );
na03f01 g38437 ( .a(n42228), .b(n9590), .c(n9589), .o(n42229) );
in01f01 g38438 ( .a(n42228), .o(n2063) );
oa12f01 g38439 ( .a(n2063), .b(n9646), .c(n9645), .o(n42231) );
na02f01 g38440 ( .a(n42231), .b(n42229), .o(n1699) );
no02f01 g38441 ( .a(n21522), .b(n16329), .o(n42233) );
no02f01 g38442 ( .a(n42233), .b(n21524), .o(n42234) );
na02f01 g38443 ( .a(n21474), .b(n21615), .o(n42235) );
in01f01 g38444 ( .a(n42235), .o(n42236) );
in01f01 g38445 ( .a(n21502), .o(n42237) );
na02f01 g38446 ( .a(n42237), .b(n42236), .o(n42238) );
no02f01 g38447 ( .a(n21500), .b(n16329), .o(n42239) );
no02f01 g38448 ( .a(n42239), .b(n21585), .o(n42240) );
na03f01 g38449 ( .a(n42240), .b(n42238), .c(n42234), .o(n42241) );
in01f01 g38450 ( .a(n42234), .o(n42242) );
oa12f01 g38451 ( .a(n42240), .b(n21502), .c(n42235), .o(n42243) );
na02f01 g38452 ( .a(n42243), .b(n42242), .o(n42244) );
na02f01 g38453 ( .a(n42244), .b(n42241), .o(n1704) );
ao12f01 g38454 ( .a(n38715), .b(n38686), .c(n41423), .o(n42246) );
no02f01 g38455 ( .a(n40430), .b(n38683), .o(n42247) );
na02f01 g38456 ( .a(n42247), .b(n42246), .o(n42248) );
in01f01 g38457 ( .a(n42246), .o(n42249) );
in01f01 g38458 ( .a(n42247), .o(n42250) );
na02f01 g38459 ( .a(n42250), .b(n42249), .o(n42251) );
na02f01 g38460 ( .a(n42251), .b(n42248), .o(n1709) );
no02f01 g38461 ( .a(n30044), .b(n30040), .o(n42253) );
no02f01 g38462 ( .a(n30043), .b(n36520), .o(n42254) );
oa12f01 g38463 ( .a(n42253), .b(n42254), .c(n30039), .o(n42255) );
no03f01 g38464 ( .a(n42254), .b(n42253), .c(n30039), .o(n42256) );
in01f01 g38465 ( .a(n42256), .o(n42257) );
na02f01 g38466 ( .a(n42257), .b(n42255), .o(n1714) );
no02f01 g38467 ( .a(n5928_1), .b(n5873), .o(n42259) );
no02f01 g38468 ( .a(n42259), .b(n5930), .o(n42260) );
in01f01 g38469 ( .a(n42260), .o(n42261) );
na02f01 g38470 ( .a(n42261), .b(n5923_1), .o(n42262) );
in01f01 g38471 ( .a(n5923_1), .o(n42263) );
na02f01 g38472 ( .a(n42260), .b(n42263), .o(n42264) );
na02f01 g38473 ( .a(n42264), .b(n42262), .o(n1724) );
no02f01 g38474 ( .a(n9747), .b(n9724), .o(n42266) );
in01f01 g38475 ( .a(n42266), .o(n42267) );
in01f01 g38476 ( .a(n9773), .o(n42268) );
no02f01 g38477 ( .a(n9766), .b(n5001), .o(n42269) );
no02f01 g38478 ( .a(n42269), .b(n9768), .o(n42270) );
na03f01 g38479 ( .a(n42270), .b(n42268), .c(n42267), .o(n42271) );
in01f01 g38480 ( .a(n42270), .o(n42272) );
oa12f01 g38481 ( .a(n42272), .b(n9773), .c(n42266), .o(n42273) );
na02f01 g38482 ( .a(n42273), .b(n42271), .o(n1734) );
ao12f01 g38483 ( .a(n14174), .b(n14191), .c(n36677), .o(n42275) );
in01f01 g38484 ( .a(n14194), .o(n42276) );
na02f01 g38485 ( .a(n42276), .b(n14189), .o(n42277) );
no02f01 g38486 ( .a(n42277), .b(n42275), .o(n42278) );
na02f01 g38487 ( .a(n42277), .b(n42275), .o(n42279) );
in01f01 g38488 ( .a(n42279), .o(n42280) );
no02f01 g38489 ( .a(n42280), .b(n42278), .o(n42281) );
in01f01 g38490 ( .a(n42281), .o(n1739) );
no02f01 g38491 ( .a(n25553), .b(n24958), .o(n42283) );
na02f01 g38492 ( .a(n42283), .b(n25182), .o(n42284) );
no02f01 g38493 ( .a(n42284), .b(n41516), .o(n42285) );
in01f01 g38494 ( .a(n25545), .o(n42286) );
ao12f01 g38495 ( .a(n25023), .b(n25548), .c(n24956), .o(n42287) );
no02f01 g38496 ( .a(n42287), .b(n42286), .o(n42288) );
in01f01 g38497 ( .a(n42288), .o(n42289) );
in01f01 g38498 ( .a(n29898), .o(n42290) );
no02f01 g38499 ( .a(n42290), .b(n24613), .o(n42291) );
no02f01 g38500 ( .a(n29898), .b(n25023), .o(n42292) );
no02f01 g38501 ( .a(n42292), .b(n42291), .o(n42293) );
in01f01 g38502 ( .a(n42293), .o(n42294) );
no03f01 g38503 ( .a(n42294), .b(n42289), .c(n42285), .o(n42295) );
in01f01 g38504 ( .a(n42295), .o(n42296) );
oa12f01 g38505 ( .a(n42294), .b(n42289), .c(n42285), .o(n42297) );
na03f01 g38506 ( .a(n42297), .b(n42296), .c(n6037), .o(n42298) );
na03f01 g38507 ( .a(n42283), .b(n41510), .c(n25182), .o(n42299) );
ao12f01 g38508 ( .a(n42293), .b(n42288), .c(n42299), .o(n42300) );
oa12f01 g38509 ( .a(n5873), .b(n42300), .c(n42295), .o(n42301) );
na02f01 g38510 ( .a(n42301), .b(n42298), .o(n1744) );
in01f01 g38511 ( .a(n39434), .o(n42303) );
no02f01 g38512 ( .a(n39446), .b(n42303), .o(n42304) );
no02f01 g38513 ( .a(n40023), .b(n39434), .o(n42305) );
no02f01 g38514 ( .a(n42305), .b(n42304), .o(n42306) );
na02f01 g38515 ( .a(n42306), .b(n39441), .o(n42307) );
in01f01 g38516 ( .a(n39441), .o(n42308) );
oa12f01 g38517 ( .a(n42308), .b(n42305), .c(n42304), .o(n42309) );
na02f01 g38518 ( .a(n42309), .b(n42307), .o(n1749) );
no02f01 g38519 ( .a(n22274), .b(n22133), .o(n42311) );
in01f01 g38520 ( .a(n42311), .o(n42312) );
ao12f01 g38521 ( .a(n22281), .b(n22291), .c(n42312), .o(n42313) );
in01f01 g38522 ( .a(n22295), .o(n42314) );
no02f01 g38523 ( .a(n42314), .b(n22290), .o(n42315) );
in01f01 g38524 ( .a(n42315), .o(n42316) );
no02f01 g38525 ( .a(n42316), .b(n42313), .o(n42317) );
na02f01 g38526 ( .a(n42316), .b(n42313), .o(n42318) );
in01f01 g38527 ( .a(n42318), .o(n42319) );
no02f01 g38528 ( .a(n42319), .b(n42317), .o(n42320) );
in01f01 g38529 ( .a(n42320), .o(n1754) );
na02f01 g38530 ( .a(n40551), .b(n6037), .o(n42322) );
na02f01 g38531 ( .a(n1150), .b(n5873), .o(n42323) );
na02f01 g38532 ( .a(n42323), .b(n42322), .o(n1759) );
in01f01 g38533 ( .a(n8604), .o(n42325) );
no02f01 g38534 ( .a(n41845), .b(n8614), .o(n42326) );
na03f01 g38535 ( .a(n42326), .b(n41844), .c(n42325), .o(n42327) );
in01f01 g38536 ( .a(n42326), .o(n42328) );
oa12f01 g38537 ( .a(n42328), .b(n8662), .c(n8604), .o(n42329) );
na02f01 g38538 ( .a(n42329), .b(n42327), .o(n1767) );
na03f01 g38539 ( .a(n27033), .b(n27229), .c(n27200), .o(n42331) );
oa12f01 g38540 ( .a(n27032), .b(n27230), .c(n26957), .o(n42332) );
na02f01 g38541 ( .a(n42332), .b(n42331), .o(n1772) );
na03f01 g38542 ( .a(n32497), .b(n32438), .c(n3633), .o(n42334) );
na02f01 g38543 ( .a(n403), .b(n6203), .o(n42335) );
na02f01 g38544 ( .a(n42335), .b(n42334), .o(n1777) );
in01f01 g38545 ( .a(n35485), .o(n42337) );
in01f01 g38546 ( .a(n35441), .o(n42338) );
no02f01 g38547 ( .a(n35465), .b(n42338), .o(n42339) );
na02f01 g38548 ( .a(n42339), .b(n42337), .o(n42340) );
no02f01 g38549 ( .a(n35483), .b(n4176), .o(n42341) );
no02f01 g38550 ( .a(n35535), .b(n42341), .o(n42342) );
no02f01 g38551 ( .a(n35533), .b(n4176), .o(n42343) );
no02f01 g38552 ( .a(n42343), .b(n35477), .o(n42344) );
na03f01 g38553 ( .a(n42344), .b(n42342), .c(n42340), .o(n42345) );
na02f01 g38554 ( .a(n42342), .b(n42340), .o(n42346) );
in01f01 g38555 ( .a(n42344), .o(n42347) );
na02f01 g38556 ( .a(n42347), .b(n42346), .o(n42348) );
na02f01 g38557 ( .a(n42348), .b(n42345), .o(n1782) );
na02f01 g38558 ( .a(n27667), .b(n41120), .o(n42350) );
in01f01 g38559 ( .a(n27465), .o(n42351) );
no02f01 g38560 ( .a(n42351), .b(n42350), .o(n42352) );
in01f01 g38561 ( .a(n42352), .o(n42353) );
in01f01 g38562 ( .a(n27490), .o(n42354) );
no02f01 g38563 ( .a(n27491), .b(n42354), .o(n42355) );
in01f01 g38564 ( .a(n27485), .o(n42356) );
no02f01 g38565 ( .a(n27484), .b(n27367), .o(n42357) );
no02f01 g38566 ( .a(n42357), .b(n42356), .o(n42358) );
na03f01 g38567 ( .a(n42358), .b(n42355), .c(n42353), .o(n42359) );
in01f01 g38568 ( .a(n42355), .o(n42360) );
in01f01 g38569 ( .a(n42358), .o(n42361) );
oa12f01 g38570 ( .a(n42361), .b(n42360), .c(n42352), .o(n42362) );
na02f01 g38571 ( .a(n42362), .b(n42359), .o(n1787) );
na02f01 g38572 ( .a(n32732), .b(cos_out_26), .o(n42364) );
in01f01 g38573 ( .a(n41632), .o(n42365) );
na03f01 g38574 ( .a(n41569), .b(n41546), .c(n39691), .o(n42366) );
in01f01 g38575 ( .a(n42366), .o(n42367) );
no02f01 g38576 ( .a(n41577), .b(n35944), .o(n42368) );
no02f01 g38577 ( .a(n42368), .b(n41579), .o(n42369) );
in01f01 g38578 ( .a(n42369), .o(n42370) );
no03f01 g38579 ( .a(n42370), .b(n42367), .c(n42365), .o(n42371) );
ao12f01 g38580 ( .a(n42369), .b(n42366), .c(n41632), .o(n42372) );
oa12f01 g38581 ( .a(n32734), .b(n42372), .c(n42371), .o(n42373) );
na02f01 g38582 ( .a(n42373), .b(n42364), .o(n1792) );
na02f01 g38583 ( .a(n38832), .b(n38827), .o(n1796) );
in01f01 g38584 ( .a(n41724), .o(n42376) );
no02f01 g38585 ( .a(n39292), .b(n29639), .o(n42377) );
no02f01 g38586 ( .a(n42377), .b(n41726), .o(n42378) );
in01f01 g38587 ( .a(n42378), .o(n42379) );
na04f01 g38588 ( .a(n41722), .b(n36762), .c(n29614), .d(n29721), .o(n42380) );
in01f01 g38589 ( .a(n41735), .o(n42381) );
na02f01 g38590 ( .a(n42381), .b(n36783), .o(n42382) );
in01f01 g38591 ( .a(n42382), .o(n42383) );
no02f01 g38592 ( .a(n39280), .b(n29639), .o(n42384) );
in01f01 g38593 ( .a(n42384), .o(n42385) );
na03f01 g38594 ( .a(n42385), .b(n42383), .c(n42380), .o(n42386) );
na03f01 g38595 ( .a(n42386), .b(n42379), .c(n42376), .o(n42387) );
in01f01 g38596 ( .a(n41722), .o(n42388) );
no04f01 g38597 ( .a(n42388), .b(n36794), .c(n29615), .d(n29578), .o(n42389) );
no03f01 g38598 ( .a(n42384), .b(n42382), .c(n42389), .o(n42390) );
oa12f01 g38599 ( .a(n42378), .b(n42390), .c(n41724), .o(n42391) );
na02f01 g38600 ( .a(n42391), .b(n42387), .o(n1801) );
in01f01 g38601 ( .a(n25146), .o(n42393) );
in01f01 g38602 ( .a(n25158), .o(n42394) );
no02f01 g38603 ( .a(n25157), .b(n25023), .o(n42395) );
no02f01 g38604 ( .a(n42395), .b(n42394), .o(n42396) );
no02f01 g38605 ( .a(n25145), .b(n25023), .o(n42397) );
no02f01 g38606 ( .a(n42397), .b(n41510), .o(n42398) );
oa12f01 g38607 ( .a(n42396), .b(n42398), .c(n42393), .o(n42399) );
in01f01 g38608 ( .a(n42396), .o(n42400) );
in01f01 g38609 ( .a(n42397), .o(n42401) );
na02f01 g38610 ( .a(n42401), .b(n41516), .o(n42402) );
na03f01 g38611 ( .a(n42402), .b(n42400), .c(n25146), .o(n42403) );
na02f01 g38612 ( .a(n42403), .b(n42399), .o(n1806) );
ao12f01 g38613 ( .a(n9224), .b(n9556), .c(n9545), .o(n42405) );
no02f01 g38614 ( .a(n42405), .b(n9536), .o(n42406) );
in01f01 g38615 ( .a(n42406), .o(n42407) );
no02f01 g38616 ( .a(n9581), .b(n9573), .o(n42408) );
na03f01 g38617 ( .a(n42408), .b(n42407), .c(n9580), .o(n42409) );
in01f01 g38618 ( .a(n42408), .o(n42410) );
oa12f01 g38619 ( .a(n42410), .b(n42406), .c(n9579), .o(n42411) );
na02f01 g38620 ( .a(n42411), .b(n42409), .o(n1811) );
no02f01 g38621 ( .a(n37142), .b(n25277), .o(n42413) );
no02f01 g38622 ( .a(n42413), .b(n37141), .o(n42414) );
na02f01 g38623 ( .a(n42413), .b(n37141), .o(n42415) );
in01f01 g38624 ( .a(n42415), .o(n42416) );
no02f01 g38625 ( .a(n42416), .b(n42414), .o(n42417) );
in01f01 g38626 ( .a(n42417), .o(n1816) );
in01f01 g38627 ( .a(n29810), .o(n42419) );
na03f01 g38628 ( .a(n42419), .b(n29809), .c(n29786), .o(n42420) );
in01f01 g38629 ( .a(n29786), .o(n42421) );
in01f01 g38630 ( .a(n29809), .o(n42422) );
oa12f01 g38631 ( .a(n42422), .b(n29810), .c(n42421), .o(n42423) );
na02f01 g38632 ( .a(n42423), .b(n42420), .o(n1826) );
na02f01 g38633 ( .a(n32732), .b(sin_out_10), .o(n42425) );
no02f01 g38634 ( .a(n38611), .b(n38607), .o(n42426) );
in01f01 g38635 ( .a(n42426), .o(n42427) );
no03f01 g38636 ( .a(n42427), .b(n38609), .c(n38598), .o(n42428) );
no02f01 g38637 ( .a(n38609), .b(n38598), .o(n42429) );
no02f01 g38638 ( .a(n42426), .b(n42429), .o(n42430) );
oa12f01 g38639 ( .a(n32734), .b(n42430), .c(n42428), .o(n42431) );
na02f01 g38640 ( .a(n42431), .b(n42425), .o(n1831) );
na03f01 g38641 ( .a(n21558), .b(n21474), .c(n21615), .o(n42433) );
no02f01 g38642 ( .a(n21596), .b(n21576), .o(n42434) );
na03f01 g38643 ( .a(n42434), .b(n21593), .c(n42433), .o(n42435) );
no03f01 g38644 ( .a(n21559), .b(n21475), .c(n21428), .o(n42436) );
in01f01 g38645 ( .a(n21593), .o(n42437) );
in01f01 g38646 ( .a(n42434), .o(n42438) );
oa12f01 g38647 ( .a(n42438), .b(n42437), .c(n42436), .o(n42439) );
na02f01 g38648 ( .a(n42439), .b(n42435), .o(n1835) );
ao12f01 g38649 ( .a(n38762), .b(n38759), .c(n38789), .o(n42441) );
no03f01 g38650 ( .a(n38763), .b(n38760), .c(n38757), .o(n42442) );
oa12f01 g38651 ( .a(delay_sub_ln23_0_unr23_stage8_stallmux_q), .b(n42442), .c(n42441), .o(n42443) );
ao12f01 g38652 ( .a(n38792), .b(n38796), .c(n38795), .o(n42444) );
no03f01 g38653 ( .a(n38793), .b(n38720), .c(n38712), .o(n42445) );
oa12f01 g38654 ( .a(delay_sub_ln23_0_unr23_stage8_stallmux_q), .b(n42445), .c(n42444), .o(n42446) );
no03f01 g38655 ( .a(n38807), .b(n38806), .c(n38805), .o(n42447) );
ao12f01 g38656 ( .a(n38802), .b(n38800), .c(n38799), .o(n42448) );
oa12f01 g38657 ( .a(delay_sub_ln23_0_unr23_stage8_stallmux_q), .b(n42448), .c(n42447), .o(n42449) );
na03f01 g38658 ( .a(n42449), .b(n42446), .c(n42443), .o(n42450) );
na03f01 g38659 ( .a(n38818), .b(n38816), .c(n38815), .o(n42451) );
oa12f01 g38660 ( .a(n38812), .b(n38813), .c(n38726), .o(n42452) );
ao12f01 g38661 ( .a(n37149), .b(n42452), .c(n42451), .o(n42453) );
ao12f01 g38662 ( .a(n37149), .b(n38970), .c(n38969), .o(n42454) );
no04f01 g38663 ( .a(n42454), .b(n38833), .c(n42453), .d(n42450), .o(n42455) );
ao12f01 g38664 ( .a(delay_sub_ln23_0_unr23_stage8_stallmux_q), .b(n38854), .c(n38850), .o(n42456) );
oa12f01 g38665 ( .a(n42455), .b(n42456), .c(n38855), .o(n42457) );
no02f01 g38666 ( .a(n42456), .b(n38855), .o(n42458) );
na02f01 g38667 ( .a(n42458), .b(n38845), .o(n42459) );
na02f01 g38668 ( .a(n42459), .b(n42457), .o(n1840) );
no02f01 g38669 ( .a(n27552), .b(n27495), .o(n42461) );
no03f01 g38670 ( .a(n29732), .b(n27628), .c(n42461), .o(n42462) );
no02f01 g38671 ( .a(n27561), .b(n27367), .o(n42463) );
no02f01 g38672 ( .a(n42463), .b(n27563), .o(n42464) );
na02f01 g38673 ( .a(n42464), .b(n42462), .o(n42465) );
in01f01 g38674 ( .a(n42462), .o(n42466) );
in01f01 g38675 ( .a(n42464), .o(n42467) );
na02f01 g38676 ( .a(n42467), .b(n42466), .o(n42468) );
na02f01 g38677 ( .a(n42468), .b(n42465), .o(n1850) );
ao12f01 g38678 ( .a(n9234), .b(n37382), .c(n8862), .o(n42470) );
in01f01 g38679 ( .a(n42470), .o(n42471) );
no02f01 g38680 ( .a(n42471), .b(n40599), .o(n42472) );
in01f01 g38681 ( .a(n40599), .o(n42473) );
no02f01 g38682 ( .a(n42470), .b(n42473), .o(n42474) );
no02f01 g38683 ( .a(n42474), .b(n42472), .o(n42475) );
na03f01 g38684 ( .a(n42475), .b(n9590), .c(n9589), .o(n42476) );
in01f01 g38685 ( .a(n42475), .o(n5051) );
oa12f01 g38686 ( .a(n5051), .b(n9646), .c(n9645), .o(n42478) );
na02f01 g38687 ( .a(n42478), .b(n42476), .o(n1855) );
no02f01 g38688 ( .a(n40828), .b(n40817), .o(n42480) );
no02f01 g38689 ( .a(n42198), .b(n40843), .o(n42481) );
ao12f01 g38690 ( .a(n42480), .b(n42481), .c(n40939), .o(n42482) );
in01f01 g38691 ( .a(n42482), .o(n42483) );
no02f01 g38692 ( .a(n40835), .b(n40810), .o(n42484) );
in01f01 g38693 ( .a(n42484), .o(n42485) );
na02f01 g38694 ( .a(n42485), .b(n42483), .o(n42486) );
na02f01 g38695 ( .a(n42484), .b(n42482), .o(n42487) );
na03f01 g38696 ( .a(n42487), .b(n42486), .c(n5799), .o(n42488) );
na02f01 g38697 ( .a(n42487), .b(n42486), .o(n3199) );
na02f01 g38698 ( .a(n3199), .b(n911), .o(n42490) );
na02f01 g38699 ( .a(n42490), .b(n42488), .o(n1860) );
na02f01 g38700 ( .a(n32732), .b(cos_out_30), .o(n42492) );
no04f01 g38701 ( .a(n41613), .b(n41589), .c(n41547), .d(n39712), .o(n42493) );
no02f01 g38702 ( .a(n41639), .b(n41636), .o(n42494) );
in01f01 g38703 ( .a(n42494), .o(n42495) );
no02f01 g38704 ( .a(n41637), .b(n35944), .o(n42496) );
no02f01 g38705 ( .a(n42496), .b(n41621), .o(n42497) );
in01f01 g38706 ( .a(n42497), .o(n42498) );
no03f01 g38707 ( .a(n42498), .b(n42495), .c(n42493), .o(n42499) );
na04f01 g38708 ( .a(n41612), .b(n41588), .c(n41546), .d(n39691), .o(n42500) );
ao12f01 g38709 ( .a(n42497), .b(n42494), .c(n42500), .o(n42501) );
oa12f01 g38710 ( .a(n32734), .b(n42501), .c(n42499), .o(n42502) );
na02f01 g38711 ( .a(n42502), .b(n42492), .o(n1865) );
oa12f01 g38712 ( .a(n4965), .b(n4961), .c(n4960), .o(n42504) );
na02f01 g38713 ( .a(n42504), .b(n4989), .o(n1869) );
in01f01 g38714 ( .a(n21213), .o(n42506) );
ao12f01 g38715 ( .a(n21227), .b(n21229), .c(n42506), .o(n42507) );
in01f01 g38716 ( .a(n42507), .o(n42508) );
no02f01 g38717 ( .a(n21239), .b(n21034), .o(n42509) );
no02f01 g38718 ( .a(n21238), .b(n21033), .o(n42510) );
no02f01 g38719 ( .a(n42510), .b(n42509), .o(n42511) );
no02f01 g38720 ( .a(n42511), .b(n42508), .o(n42512) );
na02f01 g38721 ( .a(n42511), .b(n42508), .o(n42513) );
in01f01 g38722 ( .a(n42513), .o(n42514) );
no02f01 g38723 ( .a(n42514), .b(n42512), .o(n42515) );
in01f01 g38724 ( .a(n42515), .o(n1874) );
oa12f01 g38725 ( .a(n9224), .b(n8899), .c(n8765), .o(n42517) );
in01f01 g38726 ( .a(n42517), .o(n42518) );
no02f01 g38727 ( .a(n42518), .b(n8899), .o(n42519) );
no02f01 g38728 ( .a(n9225), .b(n8862), .o(n42520) );
no02f01 g38729 ( .a(n42520), .b(n42519), .o(n42521) );
no02f01 g38730 ( .a(n42521), .b(n9232), .o(n42522) );
na02f01 g38731 ( .a(n42521), .b(n9232), .o(n42523) );
in01f01 g38732 ( .a(n42523), .o(n42524) );
no03f01 g38733 ( .a(n9224), .b(n8862), .c(beta_31), .o(n42525) );
in01f01 g38734 ( .a(n42525), .o(n42526) );
oa12f01 g38735 ( .a(n42526), .b(n42524), .c(n42522), .o(n42527) );
in01f01 g38736 ( .a(n42527), .o(n42528) );
no03f01 g38737 ( .a(n9224), .b(n8862), .c(beta_31), .o(n42529) );
no02f01 g38738 ( .a(n42529), .b(n42528), .o(n42530) );
in01f01 g38739 ( .a(n42530), .o(n1879) );
no02f01 g38740 ( .a(n9544), .b(n9225), .o(n42532) );
no02f01 g38741 ( .a(n42532), .b(n9546), .o(n42533) );
na02f01 g38742 ( .a(n42533), .b(n9536), .o(n42534) );
in01f01 g38743 ( .a(n42533), .o(n42535) );
na02f01 g38744 ( .a(n42535), .b(n9641), .o(n42536) );
na02f01 g38745 ( .a(n42536), .b(n42534), .o(n1884) );
in01f01 g38746 ( .a(n32087), .o(n42538) );
no02f01 g38747 ( .a(n38218), .b(n31607), .o(n42539) );
no02f01 g38748 ( .a(n32428), .b(n42539), .o(n42540) );
in01f01 g38749 ( .a(n42540), .o(n42541) );
oa12f01 g38750 ( .a(n42541), .b(n32427), .c(n42538), .o(n42542) );
na03f01 g38751 ( .a(n42540), .b(n32493), .c(n32087), .o(n42543) );
na02f01 g38752 ( .a(n42543), .b(n42542), .o(n1894) );
no02f01 g38753 ( .a(n11707), .b(n11706), .o(n42545) );
na02f01 g38754 ( .a(n42545), .b(n11696), .o(n42546) );
in01f01 g38755 ( .a(n11696), .o(n42547) );
in01f01 g38756 ( .a(n42545), .o(n42548) );
na02f01 g38757 ( .a(n42548), .b(n42547), .o(n42549) );
na02f01 g38758 ( .a(n42549), .b(n42546), .o(n1899) );
oa12f01 g38759 ( .a(n25866), .b(n25874), .c(n30091), .o(n42551) );
na03f01 g38760 ( .a(n25890), .b(n25872), .c(n30090), .o(n42552) );
na02f01 g38761 ( .a(n42552), .b(n42551), .o(n1904) );
no02f01 g38762 ( .a(n25546), .b(n25023), .o(n42554) );
no02f01 g38763 ( .a(n42554), .b(n25035), .o(n42555) );
in01f01 g38764 ( .a(n42555), .o(n42556) );
na02f01 g38765 ( .a(n41516), .b(n25545), .o(n42557) );
na03f01 g38766 ( .a(n42557), .b(n42556), .c(n25182), .o(n42558) );
no02f01 g38767 ( .a(n41510), .b(n42286), .o(n42559) );
oa12f01 g38768 ( .a(n42555), .b(n42559), .c(n25183), .o(n42560) );
na03f01 g38769 ( .a(n42560), .b(n42558), .c(n6037), .o(n42561) );
no03f01 g38770 ( .a(n42559), .b(n42555), .c(n25183), .o(n42562) );
ao12f01 g38771 ( .a(n42556), .b(n42557), .c(n25182), .o(n42563) );
oa12f01 g38772 ( .a(n5873), .b(n42563), .c(n42562), .o(n42564) );
na02f01 g38773 ( .a(n42564), .b(n42561), .o(n1909) );
in01f01 g38774 ( .a(n40914), .o(n42566) );
no02f01 g38775 ( .a(n40915), .b(n40911), .o(n42567) );
no02f01 g38776 ( .a(n42567), .b(n42566), .o(n42568) );
na02f01 g38777 ( .a(n42567), .b(n42566), .o(n42569) );
in01f01 g38778 ( .a(n42569), .o(n42570) );
no02f01 g38779 ( .a(n42570), .b(n42568), .o(n42571) );
in01f01 g38780 ( .a(n42571), .o(n1914) );
no02f01 g38781 ( .a(n6922), .b(n5001), .o(n42573) );
oa22f01 g38782 ( .a(n6935), .b(n42573), .c(n6914), .d(n6912), .o(n42574) );
no02f01 g38783 ( .a(n6914), .b(n6912), .o(n42575) );
in01f01 g38784 ( .a(n42573), .o(n42576) );
na03f01 g38785 ( .a(n6936), .b(n42576), .c(n42575), .o(n42577) );
na02f01 g38786 ( .a(n42577), .b(n42574), .o(n1919) );
no02f01 g38787 ( .a(n40048), .b(n40047), .o(n42579) );
in01f01 g38788 ( .a(n39976), .o(n42580) );
na02f01 g38789 ( .a(n42580), .b(n42579), .o(n42581) );
in01f01 g38790 ( .a(n39989), .o(n42582) );
no02f01 g38791 ( .a(n39860), .b(n28893), .o(n42583) );
no02f01 g38792 ( .a(n42583), .b(n42582), .o(n42584) );
no02f01 g38793 ( .a(n39860), .b(n28888), .o(n42585) );
no02f01 g38794 ( .a(n42585), .b(n39977), .o(n42586) );
na03f01 g38795 ( .a(n42586), .b(n42584), .c(n42581), .o(n42587) );
na02f01 g38796 ( .a(n39969), .b(n39945), .o(n42588) );
oa12f01 g38797 ( .a(n42584), .b(n39976), .c(n42588), .o(n42589) );
in01f01 g38798 ( .a(n42586), .o(n42590) );
na02f01 g38799 ( .a(n42590), .b(n42589), .o(n42591) );
na03f01 g38800 ( .a(n42591), .b(n42587), .c(n_27923), .o(n42592) );
na02f01 g38801 ( .a(n42591), .b(n42587), .o(n3233) );
na02f01 g38802 ( .a(n3233), .b(n34420), .o(n42594) );
na02f01 g38803 ( .a(n42594), .b(n42592), .o(n1924) );
ao12f01 g38804 ( .a(n35439), .b(n35413), .c(n42145), .o(n42596) );
no02f01 g38805 ( .a(n41948), .b(n35435), .o(n42597) );
na02f01 g38806 ( .a(n42597), .b(n42596), .o(n42598) );
in01f01 g38807 ( .a(n42596), .o(n42599) );
in01f01 g38808 ( .a(n42597), .o(n42600) );
na02f01 g38809 ( .a(n42600), .b(n42599), .o(n42601) );
na02f01 g38810 ( .a(n42601), .b(n42598), .o(n1929) );
no02f01 g38811 ( .a(n40832), .b(n40801), .o(n42603) );
in01f01 g38812 ( .a(n42603), .o(n42604) );
ao12f01 g38813 ( .a(n40810), .b(n42482), .c(n40944), .o(n42605) );
na02f01 g38814 ( .a(n42605), .b(n42604), .o(n42606) );
no02f01 g38815 ( .a(n42605), .b(n42604), .o(n42607) );
in01f01 g38816 ( .a(n42607), .o(n42608) );
na02f01 g38817 ( .a(n42608), .b(n42606), .o(n1934) );
no02f01 g38818 ( .a(n11746), .b(n38079), .o(n42610) );
no03f01 g38819 ( .a(n42610), .b(n11762), .c(n11761), .o(n42611) );
in01f01 g38820 ( .a(n42611), .o(n42612) );
no02f01 g38821 ( .a(n11763), .b(n11755), .o(n42613) );
in01f01 g38822 ( .a(n42613), .o(n42614) );
na02f01 g38823 ( .a(n42614), .b(n42612), .o(n42615) );
na02f01 g38824 ( .a(n42613), .b(n42611), .o(n42616) );
na02f01 g38825 ( .a(n42616), .b(n42615), .o(n1939) );
na02f01 g38826 ( .a(n9845), .b(n9832), .o(n42618) );
no02f01 g38827 ( .a(n9871), .b(n9854), .o(n42619) );
na03f01 g38828 ( .a(n42619), .b(n9870), .c(n42618), .o(n42620) );
na02f01 g38829 ( .a(n9870), .b(n42618), .o(n42621) );
in01f01 g38830 ( .a(n42619), .o(n42622) );
na02f01 g38831 ( .a(n42622), .b(n42621), .o(n42623) );
na02f01 g38832 ( .a(n42623), .b(n42620), .o(n1944) );
na03f01 g38833 ( .a(n41925), .b(n41921), .c(n1821), .o(n42625) );
ao12f01 g38834 ( .a(n41922), .b(n41924), .c(n27192), .o(n42626) );
no03f01 g38835 ( .a(n41920), .b(n41918), .c(n41915), .o(n42627) );
oa12f01 g38836 ( .a(n8066), .b(n42627), .c(n42626), .o(n42628) );
na02f01 g38837 ( .a(n42628), .b(n42625), .o(n1949) );
in01f01 g38838 ( .a(n42350), .o(n42630) );
no02f01 g38839 ( .a(n27451), .b(n27367), .o(n42631) );
in01f01 g38840 ( .a(n42631), .o(n42632) );
na02f01 g38841 ( .a(n42632), .b(n27490), .o(n42633) );
ao12f01 g38842 ( .a(n42633), .b(n27452), .c(n42630), .o(n42634) );
no02f01 g38843 ( .a(n27462), .b(n27367), .o(n42635) );
no02f01 g38844 ( .a(n42635), .b(n27464), .o(n42636) );
na02f01 g38845 ( .a(n42636), .b(n42634), .o(n42637) );
in01f01 g38846 ( .a(n42634), .o(n42638) );
in01f01 g38847 ( .a(n42636), .o(n42639) );
na02f01 g38848 ( .a(n42639), .b(n42638), .o(n42640) );
na02f01 g38849 ( .a(n42640), .b(n42637), .o(n1954) );
no02f01 g38850 ( .a(n8584), .b(n8578), .o(n42642) );
no02f01 g38851 ( .a(n8601), .b(n5973), .o(n42643) );
no02f01 g38852 ( .a(n8602), .b(n8471), .o(n42644) );
in01f01 g38853 ( .a(n42644), .o(n42645) );
ao12f01 g38854 ( .a(n42643), .b(n42645), .c(n42642), .o(n42646) );
no02f01 g38855 ( .a(n8596), .b(n8471), .o(n42647) );
no02f01 g38856 ( .a(n8595), .b(n5973), .o(n42648) );
no02f01 g38857 ( .a(n42648), .b(n42647), .o(n42649) );
na02f01 g38858 ( .a(n42649), .b(n42646), .o(n42650) );
in01f01 g38859 ( .a(n42646), .o(n42651) );
in01f01 g38860 ( .a(n42649), .o(n42652) );
na02f01 g38861 ( .a(n42652), .b(n42651), .o(n42653) );
na02f01 g38862 ( .a(n42653), .b(n42650), .o(n1959) );
ao12f01 g38863 ( .a(n29403), .b(n29406), .c(n29701), .o(n42655) );
in01f01 g38864 ( .a(n42655), .o(n42656) );
no02f01 g38865 ( .a(n29704), .b(n29327), .o(n42657) );
na02f01 g38866 ( .a(n42657), .b(n42656), .o(n42658) );
in01f01 g38867 ( .a(n42657), .o(n42659) );
na02f01 g38868 ( .a(n42659), .b(n42655), .o(n42660) );
na02f01 g38869 ( .a(n42660), .b(n42658), .o(n1964) );
no02f01 g38870 ( .a(n38446), .b(n38282), .o(n42662) );
in01f01 g38871 ( .a(n42662), .o(n42663) );
ao12f01 g38872 ( .a(n38468), .b(n38505), .c(n42663), .o(n42664) );
no02f01 g38873 ( .a(n38509), .b(n39128), .o(n42665) );
in01f01 g38874 ( .a(n42665), .o(n42666) );
na02f01 g38875 ( .a(n42666), .b(n42664), .o(n42667) );
in01f01 g38876 ( .a(n42664), .o(n42668) );
na02f01 g38877 ( .a(n42665), .b(n42668), .o(n42669) );
na02f01 g38878 ( .a(n42669), .b(n42667), .o(n1969) );
no02f01 g38879 ( .a(n37871), .b(n26256), .o(n42671) );
in01f01 g38880 ( .a(n26256), .o(n42672) );
no02f01 g38881 ( .a(n38010), .b(n42672), .o(n42673) );
no02f01 g38882 ( .a(n42673), .b(n42671), .o(n42674) );
na03f01 g38883 ( .a(n42674), .b(n41239), .c(n41248), .o(n42675) );
in01f01 g38884 ( .a(n42674), .o(n42676) );
oa12f01 g38885 ( .a(n42676), .b(n41240), .c(n41228), .o(n42677) );
na03f01 g38886 ( .a(n42677), .b(n42675), .c(n1821), .o(n42678) );
na02f01 g38887 ( .a(n42677), .b(n42675), .o(n3332) );
na02f01 g38888 ( .a(n3332), .b(n8066), .o(n42680) );
na02f01 g38889 ( .a(n42680), .b(n42678), .o(n1974) );
na02f01 g38890 ( .a(n32732), .b(sin_out_1), .o(n42682) );
ao12f01 g38891 ( .a(n36560), .b(n34326), .c(n36556), .o(n42683) );
no03f01 g38892 ( .a(n36561), .b(n34325), .c(n34317), .o(n42684) );
oa12f01 g38893 ( .a(n32734), .b(n42684), .c(n42683), .o(n42685) );
na02f01 g38894 ( .a(n42685), .b(n42682), .o(n1979) );
no02f01 g38895 ( .a(n39182), .b(n39180), .o(n42687) );
in01f01 g38896 ( .a(n42687), .o(n42688) );
no02f01 g38897 ( .a(n42688), .b(n38007), .o(n42689) );
no02f01 g38898 ( .a(n42687), .b(n38048), .o(n42690) );
no02f01 g38899 ( .a(n42690), .b(n42689), .o(n42691) );
in01f01 g38900 ( .a(n42691), .o(n1983) );
no02f01 g38901 ( .a(n40709), .b(n21270), .o(n42693) );
no02f01 g38902 ( .a(n42693), .b(n41380), .o(n42694) );
na02f01 g38903 ( .a(n40712), .b(n21305), .o(n42695) );
in01f01 g38904 ( .a(n42695), .o(n42696) );
ao12f01 g38905 ( .a(n41378), .b(n21334), .c(n21327), .o(n42697) );
no03f01 g38906 ( .a(n42697), .b(n41384), .c(n42696), .o(n42698) );
oa12f01 g38907 ( .a(n42694), .b(n42698), .c(n41379), .o(n42699) );
in01f01 g38908 ( .a(n41379), .o(n42700) );
in01f01 g38909 ( .a(n42694), .o(n42701) );
in01f01 g38910 ( .a(n41384), .o(n42702) );
oa12f01 g38911 ( .a(n41390), .b(n21263), .c(n20923), .o(n42703) );
na03f01 g38912 ( .a(n42703), .b(n42702), .c(n42695), .o(n42704) );
na03f01 g38913 ( .a(n42704), .b(n42701), .c(n42700), .o(n42705) );
na03f01 g38914 ( .a(n42705), .b(n42699), .c(n5799), .o(n42706) );
ao12f01 g38915 ( .a(n42701), .b(n42704), .c(n42700), .o(n42707) );
no03f01 g38916 ( .a(n42698), .b(n42694), .c(n41379), .o(n42708) );
oa12f01 g38917 ( .a(n911), .b(n42708), .c(n42707), .o(n42709) );
na02f01 g38918 ( .a(n42709), .b(n42706), .o(n1988) );
no02f01 g38919 ( .a(n9628), .b(n9307), .o(n42711) );
in01f01 g38920 ( .a(n42711), .o(n42712) );
na02f01 g38921 ( .a(n42712), .b(n9421), .o(n42713) );
na02f01 g38922 ( .a(n42711), .b(n9627), .o(n42714) );
na02f01 g38923 ( .a(n42714), .b(n42713), .o(n1993) );
na02f01 g38924 ( .a(n32432), .b(n31606), .o(n42716) );
in01f01 g38925 ( .a(n42716), .o(n42717) );
in01f01 g38926 ( .a(n32107), .o(n42718) );
oa12f01 g38927 ( .a(n42718), .b(n32494), .c(n32493), .o(n42719) );
no02f01 g38928 ( .a(n42719), .b(n42717), .o(n42720) );
no02f01 g38929 ( .a(n32128), .b(n31607), .o(n42721) );
no02f01 g38930 ( .a(n42721), .b(n32435), .o(n42722) );
no03f01 g38931 ( .a(n42722), .b(n42720), .c(n32433), .o(n42723) );
in01f01 g38932 ( .a(n42723), .o(n42724) );
oa12f01 g38933 ( .a(n42722), .b(n42720), .c(n32433), .o(n42725) );
na03f01 g38934 ( .a(n42725), .b(n42724), .c(n3633), .o(n42726) );
no02f01 g38935 ( .a(n42720), .b(n32433), .o(n42727) );
in01f01 g38936 ( .a(n42722), .o(n42728) );
no02f01 g38937 ( .a(n42728), .b(n42727), .o(n42729) );
oa12f01 g38938 ( .a(n6203), .b(n42729), .c(n42723), .o(n42730) );
na02f01 g38939 ( .a(n42730), .b(n42726), .o(n1998) );
oa22f01 g38940 ( .a(n27664), .b(n27373), .c(n27662), .d(n27310), .o(n42732) );
oa12f01 g38941 ( .a(n42732), .b(n27664), .c(n27375), .o(n2008) );
na02f01 g38942 ( .a(n22363), .b(n22466), .o(n42734) );
in01f01 g38943 ( .a(n42734), .o(n42735) );
no02f01 g38944 ( .a(n22467), .b(n22077), .o(n42736) );
no02f01 g38945 ( .a(n42736), .b(n42735), .o(n42737) );
na02f01 g38946 ( .a(n42736), .b(n42735), .o(n42738) );
in01f01 g38947 ( .a(n42738), .o(n42739) );
no02f01 g38948 ( .a(n42739), .b(n42737), .o(n42740) );
in01f01 g38949 ( .a(n42740), .o(n2013) );
na02f01 g38950 ( .a(n40593), .b(n40589), .o(n2018) );
na02f01 g38951 ( .a(n27440), .b(n41120), .o(n42743) );
in01f01 g38952 ( .a(n42743), .o(n42744) );
in01f01 g38953 ( .a(n27488), .o(n42745) );
in01f01 g38954 ( .a(n27411), .o(n42746) );
na02f01 g38955 ( .a(n42746), .b(n27395), .o(n42747) );
na02f01 g38956 ( .a(n42747), .b(n42745), .o(n42748) );
ao12f01 g38957 ( .a(n42748), .b(n42744), .c(n27412), .o(n42749) );
in01f01 g38958 ( .a(n27423), .o(n42750) );
no02f01 g38959 ( .a(n27422), .b(n27367), .o(n42751) );
no02f01 g38960 ( .a(n42751), .b(n42750), .o(n42752) );
na02f01 g38961 ( .a(n42752), .b(n42749), .o(n42753) );
in01f01 g38962 ( .a(n42749), .o(n42754) );
in01f01 g38963 ( .a(n42752), .o(n42755) );
na02f01 g38964 ( .a(n42755), .b(n42754), .o(n42756) );
na02f01 g38965 ( .a(n42756), .b(n42753), .o(n2023) );
in01f01 g38966 ( .a(n11628), .o(n42758) );
no02f01 g38967 ( .a(n42758), .b(n11611), .o(n42759) );
in01f01 g38968 ( .a(n42759), .o(n42760) );
na02f01 g38969 ( .a(n42760), .b(n11627), .o(n42761) );
na02f01 g38970 ( .a(n42759), .b(n11626), .o(n42762) );
na02f01 g38971 ( .a(n42762), .b(n42761), .o(n2028) );
no02f01 g38972 ( .a(n32084), .b(n31606), .o(n42764) );
no02f01 g38973 ( .a(n32083), .b(n31607), .o(n42765) );
no02f01 g38974 ( .a(n42765), .b(n42764), .o(n42766) );
oa12f01 g38975 ( .a(n42766), .b(n32418), .c(n32139), .o(n42767) );
in01f01 g38976 ( .a(n42766), .o(n42768) );
na02f01 g38977 ( .a(n42768), .b(n39521), .o(n42769) );
na02f01 g38978 ( .a(n42769), .b(n42767), .o(n2033) );
no02f01 g38979 ( .a(n35334), .b(n4176), .o(n42771) );
ao12f01 g38980 ( .a(n42771), .b(n35337), .c(n35327), .o(n42772) );
no02f01 g38981 ( .a(n35269), .b(n4176), .o(n42773) );
no02f01 g38982 ( .a(n42773), .b(n35271), .o(n42774) );
na02f01 g38983 ( .a(n42774), .b(n42772), .o(n42775) );
in01f01 g38984 ( .a(n42772), .o(n42776) );
in01f01 g38985 ( .a(n42774), .o(n42777) );
na02f01 g38986 ( .a(n42777), .b(n42776), .o(n42778) );
na02f01 g38987 ( .a(n42778), .b(n42775), .o(n2038) );
no02f01 g38988 ( .a(n39625), .b(n9591), .o(n42780) );
no02f01 g38989 ( .a(n39624), .b(n4201), .o(n42781) );
no02f01 g38990 ( .a(n42781), .b(n42780), .o(n42782) );
na03f01 g38991 ( .a(n42782), .b(n9590), .c(n9589), .o(n42783) );
in01f01 g38992 ( .a(n42782), .o(n3228) );
oa12f01 g38993 ( .a(n3228), .b(n9646), .c(n9645), .o(n42785) );
na02f01 g38994 ( .a(n42785), .b(n42783), .o(n2043) );
na02f01 g38995 ( .a(n38820), .b(n38810), .o(n42787) );
in01f01 g38996 ( .a(n42787), .o(n42788) );
ao12f01 g38997 ( .a(delay_sub_ln23_0_unr23_stage8_stallmux_q), .b(n38970), .c(n38969), .o(n42789) );
no02f01 g38998 ( .a(n42789), .b(n42454), .o(n42790) );
in01f01 g38999 ( .a(n42790), .o(n42791) );
na03f01 g39000 ( .a(n42791), .b(n38834), .c(n42788), .o(n42792) );
oa12f01 g39001 ( .a(n42790), .b(n38833), .c(n42787), .o(n42793) );
na02f01 g39002 ( .a(n42793), .b(n42792), .o(n2053) );
no02f01 g39003 ( .a(n30112), .b(n29994), .o(n42795) );
in01f01 g39004 ( .a(n42795), .o(n42796) );
no02f01 g39005 ( .a(n30010), .b(n30115), .o(n42797) );
no02f01 g39006 ( .a(n42797), .b(n42796), .o(n42798) );
na02f01 g39007 ( .a(n42797), .b(n42796), .o(n42799) );
in01f01 g39008 ( .a(n42799), .o(n42800) );
no02f01 g39009 ( .a(n42800), .b(n42798), .o(n42801) );
in01f01 g39010 ( .a(n42801), .o(n2058) );
na02f01 g39011 ( .a(n11651), .b(n11650), .o(n42803) );
in01f01 g39012 ( .a(n42803), .o(n42804) );
no02f01 g39013 ( .a(n11660), .b(n11515), .o(n42805) );
ao12f01 g39014 ( .a(n42805), .b(n11663), .c(n42804), .o(n42806) );
no02f01 g39015 ( .a(n11670), .b(n11514), .o(n42807) );
no02f01 g39016 ( .a(n42807), .b(n11672), .o(n42808) );
na02f01 g39017 ( .a(n42808), .b(n42806), .o(n42809) );
in01f01 g39018 ( .a(n42806), .o(n42810) );
in01f01 g39019 ( .a(n42808), .o(n42811) );
na02f01 g39020 ( .a(n42811), .b(n42810), .o(n42812) );
na02f01 g39021 ( .a(n42812), .b(n42809), .o(n2068) );
no02f01 g39022 ( .a(n35232), .b(n5978), .o(n42814) );
in01f01 g39023 ( .a(n42814), .o(n42815) );
no02f01 g39024 ( .a(n35233), .b(n34908), .o(n42816) );
no02f01 g39025 ( .a(n35254), .b(n35214), .o(n42817) );
ao12f01 g39026 ( .a(n42816), .b(n42817), .c(n42815), .o(n42818) );
in01f01 g39027 ( .a(n42818), .o(n42819) );
no02f01 g39028 ( .a(n35227), .b(n34908), .o(n42820) );
no02f01 g39029 ( .a(n35226), .b(n5978), .o(n42821) );
no02f01 g39030 ( .a(n42821), .b(n42820), .o(n42822) );
no02f01 g39031 ( .a(n42822), .b(n42819), .o(n42823) );
na02f01 g39032 ( .a(n42822), .b(n42819), .o(n42824) );
in01f01 g39033 ( .a(n42824), .o(n42825) );
no02f01 g39034 ( .a(n42825), .b(n42823), .o(n42826) );
no02f01 g39035 ( .a(n42816), .b(n42814), .o(n42827) );
in01f01 g39036 ( .a(n42827), .o(n42828) );
no03f01 g39037 ( .a(n42828), .b(n35254), .c(n35214), .o(n42829) );
no02f01 g39038 ( .a(n42827), .b(n42817), .o(n42830) );
no02f01 g39039 ( .a(n42830), .b(n42829), .o(n42831) );
ao12f01 g39040 ( .a(n4176), .b(n42831), .c(n42826), .o(n42832) );
in01f01 g39041 ( .a(n42832), .o(n42833) );
no02f01 g39042 ( .a(n35249), .b(n35547), .o(n42834) );
oa12f01 g39043 ( .a(n42834), .b(n35205), .c(n35156), .o(n42835) );
no02f01 g39044 ( .a(n42835), .b(n35252), .o(n42836) );
no02f01 g39045 ( .a(n42836), .b(n35211), .o(n42837) );
in01f01 g39046 ( .a(n42837), .o(n42838) );
no02f01 g39047 ( .a(n35183), .b(n5978), .o(n42839) );
no02f01 g39048 ( .a(n42839), .b(n35185), .o(n42840) );
no02f01 g39049 ( .a(n42840), .b(n42838), .o(n42841) );
na02f01 g39050 ( .a(n42840), .b(n42838), .o(n42842) );
in01f01 g39051 ( .a(n42842), .o(n42843) );
no02f01 g39052 ( .a(n42843), .b(n42841), .o(n42844) );
in01f01 g39053 ( .a(n42844), .o(n42845) );
no02f01 g39054 ( .a(n42845), .b(n35258), .o(n42846) );
in01f01 g39055 ( .a(n35549), .o(n42847) );
oa12f01 g39056 ( .a(n42847), .b(n35550), .c(n35548), .o(n42848) );
no02f01 g39057 ( .a(n35196), .b(n34908), .o(n42849) );
no02f01 g39058 ( .a(n35195), .b(n5978), .o(n42850) );
no02f01 g39059 ( .a(n42850), .b(n42849), .o(n42851) );
in01f01 g39060 ( .a(n42851), .o(n42852) );
no02f01 g39061 ( .a(n42852), .b(n42848), .o(n42853) );
na02f01 g39062 ( .a(n42852), .b(n42848), .o(n42854) );
in01f01 g39063 ( .a(n42854), .o(n42855) );
no03f01 g39064 ( .a(n42855), .b(n42853), .c(n35258), .o(n42856) );
no02f01 g39065 ( .a(n42856), .b(n35557), .o(n42857) );
in01f01 g39066 ( .a(n42857), .o(n42858) );
in01f01 g39067 ( .a(n42835), .o(n42859) );
no02f01 g39068 ( .a(n35252), .b(n35211), .o(n42860) );
no02f01 g39069 ( .a(n42860), .b(n42859), .o(n42861) );
na02f01 g39070 ( .a(n42860), .b(n42859), .o(n42862) );
in01f01 g39071 ( .a(n42862), .o(n42863) );
no02f01 g39072 ( .a(n42863), .b(n42861), .o(n42864) );
in01f01 g39073 ( .a(n42864), .o(n42865) );
no02f01 g39074 ( .a(n42865), .b(n35258), .o(n42866) );
no03f01 g39075 ( .a(n42866), .b(n42858), .c(n42846), .o(n42867) );
in01f01 g39076 ( .a(n42867), .o(n42868) );
ao12f01 g39077 ( .a(n42868), .b(n35543), .c(n35531), .o(n42869) );
no02f01 g39078 ( .a(n42864), .b(n4176), .o(n42870) );
no02f01 g39079 ( .a(n42870), .b(n42845), .o(n42871) );
no02f01 g39080 ( .a(n42855), .b(n42853), .o(n42872) );
ao12f01 g39081 ( .a(n4176), .b(n42872), .c(n35555), .o(n42873) );
in01f01 g39082 ( .a(n42873), .o(n42874) );
oa12f01 g39083 ( .a(n42874), .b(n42871), .c(n4176), .o(n42875) );
no03f01 g39084 ( .a(n42825), .b(n42823), .c(n35258), .o(n42876) );
no03f01 g39085 ( .a(n42830), .b(n42829), .c(n35258), .o(n42877) );
no02f01 g39086 ( .a(n42877), .b(n42876), .o(n42878) );
oa12f01 g39087 ( .a(n42878), .b(n42875), .c(n42869), .o(n42879) );
oa12f01 g39088 ( .a(n35247), .b(n42817), .c(n35234), .o(n42880) );
in01f01 g39089 ( .a(n42880), .o(n42881) );
no02f01 g39090 ( .a(n35245), .b(n5978), .o(n42882) );
no02f01 g39091 ( .a(n42882), .b(n35243), .o(n42883) );
no02f01 g39092 ( .a(n42883), .b(n42881), .o(n42884) );
na02f01 g39093 ( .a(n42883), .b(n42881), .o(n42885) );
in01f01 g39094 ( .a(n42885), .o(n42886) );
no03f01 g39095 ( .a(n42886), .b(n42884), .c(n35258), .o(n42887) );
no02f01 g39096 ( .a(n42886), .b(n42884), .o(n42888) );
no02f01 g39097 ( .a(n42888), .b(n4176), .o(n42889) );
no02f01 g39098 ( .a(n42889), .b(n42887), .o(n42890) );
na03f01 g39099 ( .a(n42890), .b(n42879), .c(n42833), .o(n42891) );
na02f01 g39100 ( .a(n42879), .b(n42833), .o(n42892) );
in01f01 g39101 ( .a(n42890), .o(n42893) );
na02f01 g39102 ( .a(n42893), .b(n42892), .o(n42894) );
na02f01 g39103 ( .a(n42894), .b(n42891), .o(n2077) );
ao12f01 g39104 ( .a(n27060), .b(n27065), .c(n27045), .o(n42896) );
in01f01 g39105 ( .a(n42896), .o(n42897) );
in01f01 g39106 ( .a(n27061), .o(n42898) );
no02f01 g39107 ( .a(n42898), .b(n26869), .o(n42899) );
no02f01 g39108 ( .a(n42899), .b(n42897), .o(n42900) );
in01f01 g39109 ( .a(n42900), .o(n42901) );
na02f01 g39110 ( .a(n42899), .b(n42897), .o(n42902) );
na02f01 g39111 ( .a(n42902), .b(n42901), .o(n2082) );
no02f01 g39112 ( .a(n39861), .b(n39973), .o(n42904) );
no02f01 g39113 ( .a(n39860), .b(n39972), .o(n42905) );
no02f01 g39114 ( .a(n42905), .b(n42904), .o(n42906) );
in01f01 g39115 ( .a(n42906), .o(n42907) );
no02f01 g39116 ( .a(n39861), .b(n39971), .o(n42908) );
in01f01 g39117 ( .a(n42908), .o(n42909) );
in01f01 g39118 ( .a(n39992), .o(n42910) );
no02f01 g39119 ( .a(n39860), .b(n39970), .o(n42911) );
in01f01 g39120 ( .a(n42911), .o(n42912) );
na03f01 g39121 ( .a(n39978), .b(n39969), .c(n39945), .o(n42913) );
na03f01 g39122 ( .a(n42913), .b(n42912), .c(n42910), .o(n42914) );
na03f01 g39123 ( .a(n42914), .b(n42909), .c(n42907), .o(n42915) );
in01f01 g39124 ( .a(n39978), .o(n42916) );
no03f01 g39125 ( .a(n42916), .b(n40048), .c(n40047), .o(n42917) );
no03f01 g39126 ( .a(n42917), .b(n42911), .c(n39992), .o(n42918) );
oa12f01 g39127 ( .a(n42906), .b(n42918), .c(n42908), .o(n42919) );
na03f01 g39128 ( .a(n42919), .b(n42915), .c(n_27923), .o(n42920) );
no03f01 g39129 ( .a(n42918), .b(n42908), .c(n42906), .o(n42921) );
ao12f01 g39130 ( .a(n42907), .b(n42914), .c(n42909), .o(n42922) );
oa12f01 g39131 ( .a(n34420), .b(n42922), .c(n42921), .o(n42923) );
na02f01 g39132 ( .a(n42923), .b(n42920), .o(n2087) );
in01f01 g39133 ( .a(n40447), .o(n42925) );
no02f01 g39134 ( .a(n39260), .b(n29639), .o(n42926) );
no02f01 g39135 ( .a(n36771), .b(n29430), .o(n42927) );
no02f01 g39136 ( .a(n42927), .b(n42926), .o(n42928) );
in01f01 g39137 ( .a(n40448), .o(n42929) );
oa12f01 g39138 ( .a(n42929), .b(n40452), .c(n40451), .o(n42930) );
na03f01 g39139 ( .a(n42930), .b(n42928), .c(n42925), .o(n42931) );
in01f01 g39140 ( .a(n42928), .o(n42932) );
ao12f01 g39141 ( .a(n40448), .b(n36783), .c(n40446), .o(n42933) );
oa12f01 g39142 ( .a(n42932), .b(n42933), .c(n40447), .o(n42934) );
na02f01 g39143 ( .a(n42934), .b(n42931), .o(n2092) );
no02f01 g39144 ( .a(n32433), .b(n42717), .o(n42936) );
in01f01 g39145 ( .a(n42936), .o(n42937) );
na02f01 g39146 ( .a(n42937), .b(n42719), .o(n42938) );
na02f01 g39147 ( .a(n32430), .b(n32427), .o(n42939) );
na03f01 g39148 ( .a(n42936), .b(n42939), .c(n42718), .o(n42940) );
na03f01 g39149 ( .a(n42940), .b(n42938), .c(n3633), .o(n42941) );
na02f01 g39150 ( .a(n42940), .b(n42938), .o(n2672) );
na02f01 g39151 ( .a(n2672), .b(n6203), .o(n42943) );
na02f01 g39152 ( .a(n42943), .b(n42941), .o(n2097) );
no02f01 g39153 ( .a(n35348), .b(n4176), .o(n42945) );
no02f01 g39154 ( .a(n35349), .b(n35258), .o(n42946) );
in01f01 g39155 ( .a(n42946), .o(n42947) );
ao12f01 g39156 ( .a(n42945), .b(n42947), .c(n38979), .o(n42948) );
no02f01 g39157 ( .a(n35359), .b(n35258), .o(n42949) );
no02f01 g39158 ( .a(n35358), .b(n4176), .o(n42950) );
no02f01 g39159 ( .a(n42950), .b(n42949), .o(n42951) );
na02f01 g39160 ( .a(n42951), .b(n42948), .o(n42952) );
in01f01 g39161 ( .a(n42948), .o(n42953) );
in01f01 g39162 ( .a(n42951), .o(n42954) );
na02f01 g39163 ( .a(n42954), .b(n42953), .o(n42955) );
na02f01 g39164 ( .a(n42955), .b(n42952), .o(n2107) );
in01f01 g39165 ( .a(n40182), .o(n42957) );
no02f01 g39166 ( .a(n42957), .b(n40114), .o(n42958) );
in01f01 g39167 ( .a(n42958), .o(n42959) );
no02f01 g39168 ( .a(n42959), .b(n40181), .o(n42960) );
na02f01 g39169 ( .a(n42959), .b(n40181), .o(n42961) );
in01f01 g39170 ( .a(n42961), .o(n42962) );
no02f01 g39171 ( .a(n42962), .b(n42960), .o(n42963) );
na02f01 g39172 ( .a(n42963), .b(n5799), .o(n42964) );
in01f01 g39173 ( .a(n42963), .o(n4241) );
na02f01 g39174 ( .a(n4241), .b(n911), .o(n42966) );
na02f01 g39175 ( .a(n42966), .b(n42964), .o(n2112) );
na02f01 g39176 ( .a(n32732), .b(cos_out_27), .o(n42968) );
no04f01 g39177 ( .a(n41579), .b(n41570), .c(n41547), .d(n39712), .o(n42969) );
no02f01 g39178 ( .a(n42368), .b(n42365), .o(n42970) );
in01f01 g39179 ( .a(n42970), .o(n42971) );
no02f01 g39180 ( .a(n41633), .b(n35944), .o(n42972) );
no02f01 g39181 ( .a(n42972), .b(n41587), .o(n42973) );
in01f01 g39182 ( .a(n42973), .o(n42974) );
no03f01 g39183 ( .a(n42974), .b(n42971), .c(n42969), .o(n42975) );
in01f01 g39184 ( .a(n41579), .o(n42976) );
na04f01 g39185 ( .a(n42976), .b(n41569), .c(n41546), .d(n39691), .o(n42977) );
ao12f01 g39186 ( .a(n42973), .b(n42970), .c(n42977), .o(n42978) );
oa12f01 g39187 ( .a(n32734), .b(n42978), .c(n42975), .o(n42979) );
na02f01 g39188 ( .a(n42979), .b(n42968), .o(n2117) );
no02f01 g39189 ( .a(n30121), .b(n29984), .o(n42981) );
no02f01 g39190 ( .a(n42981), .b(n30120), .o(n42982) );
na02f01 g39191 ( .a(n42981), .b(n30120), .o(n42983) );
in01f01 g39192 ( .a(n42983), .o(n42984) );
no02f01 g39193 ( .a(n42984), .b(n42982), .o(n42985) );
na02f01 g39194 ( .a(n42985), .b(n6037), .o(n42986) );
in01f01 g39195 ( .a(n42985), .o(n5692) );
na02f01 g39196 ( .a(n5692), .b(n5873), .o(n42988) );
na02f01 g39197 ( .a(n42988), .b(n42986), .o(n2121) );
na03f01 g39198 ( .a(n25580), .b(n25552), .c(n6037), .o(n42990) );
no03f01 g39199 ( .a(n25579), .b(n25553), .c(n25025), .o(n42991) );
ao12f01 g39200 ( .a(n25026), .b(n25551), .c(n25047), .o(n42992) );
oa12f01 g39201 ( .a(n5873), .b(n42992), .c(n42991), .o(n42993) );
na02f01 g39202 ( .a(n42993), .b(n42990), .o(n2126) );
no02f01 g39203 ( .a(n27503), .b(n27367), .o(n42995) );
no03f01 g39204 ( .a(n27524), .b(n27505), .c(n27495), .o(n42996) );
no03f01 g39205 ( .a(n42996), .b(n42995), .c(n27625), .o(n42997) );
no02f01 g39206 ( .a(n27535), .b(n27367), .o(n42998) );
no02f01 g39207 ( .a(n42998), .b(n27537), .o(n42999) );
na02f01 g39208 ( .a(n42999), .b(n42997), .o(n43000) );
in01f01 g39209 ( .a(n42997), .o(n43001) );
in01f01 g39210 ( .a(n42999), .o(n43002) );
na02f01 g39211 ( .a(n43002), .b(n43001), .o(n43003) );
na02f01 g39212 ( .a(n43003), .b(n43000), .o(n2136) );
no02f01 g39213 ( .a(n11841), .b(n35569), .o(n43005) );
no02f01 g39214 ( .a(n11843), .b(n11836), .o(n43006) );
oa12f01 g39215 ( .a(n43006), .b(n43005), .c(n11828), .o(n43007) );
no02f01 g39216 ( .a(n43005), .b(n11828), .o(n43008) );
in01f01 g39217 ( .a(n43006), .o(n43009) );
na02f01 g39218 ( .a(n43009), .b(n43008), .o(n43010) );
na02f01 g39219 ( .a(n43010), .b(n43007), .o(n2141) );
na03f01 g39220 ( .a(n16088), .b(n21364), .c(n21350), .o(n43012) );
oa12f01 g39221 ( .a(n16087), .b(n21365), .c(n16056), .o(n43013) );
na02f01 g39222 ( .a(n43013), .b(n43012), .o(n2146) );
na02f01 g39223 ( .a(n32732), .b(cos_out_25), .o(n43015) );
no02f01 g39224 ( .a(n41630), .b(n35944), .o(n43016) );
no02f01 g39225 ( .a(n43016), .b(n41561), .o(n43017) );
in01f01 g39226 ( .a(n43017), .o(n43018) );
in01f01 g39227 ( .a(n41568), .o(n43019) );
na03f01 g39228 ( .a(n43019), .b(n41546), .c(n39691), .o(n43020) );
no02f01 g39229 ( .a(n41566), .b(n35944), .o(n43021) );
no02f01 g39230 ( .a(n43021), .b(n41629), .o(n43022) );
na02f01 g39231 ( .a(n43022), .b(n43020), .o(n43023) );
no02f01 g39232 ( .a(n43023), .b(n43018), .o(n43024) );
ao12f01 g39233 ( .a(n43017), .b(n43022), .c(n43020), .o(n43025) );
oa12f01 g39234 ( .a(n32734), .b(n43025), .c(n43024), .o(n43026) );
na02f01 g39235 ( .a(n43026), .b(n43015), .o(n2151) );
no02f01 g39236 ( .a(n36790), .b(n36737), .o(n43028) );
na03f01 g39237 ( .a(n43028), .b(n36786), .c(n36779), .o(n43029) );
in01f01 g39238 ( .a(n43028), .o(n43030) );
oa12f01 g39239 ( .a(n43030), .b(n36785), .c(n36795), .o(n43031) );
na03f01 g39240 ( .a(n43031), .b(n43029), .c(n_27923), .o(n43032) );
na02f01 g39241 ( .a(n43031), .b(n43029), .o(n2213) );
na02f01 g39242 ( .a(n2213), .b(n34420), .o(n43034) );
na02f01 g39243 ( .a(n43034), .b(n43032), .o(n2155) );
no02f01 g39244 ( .a(n9482), .b(n9225), .o(n43036) );
ao12f01 g39245 ( .a(n43036), .b(n9456), .c(n9436), .o(n43037) );
no02f01 g39246 ( .a(n9485), .b(n9469), .o(n43038) );
na02f01 g39247 ( .a(n43038), .b(n43037), .o(n43039) );
in01f01 g39248 ( .a(n43037), .o(n43040) );
in01f01 g39249 ( .a(n43038), .o(n43041) );
na02f01 g39250 ( .a(n43041), .b(n43040), .o(n43042) );
na02f01 g39251 ( .a(n43042), .b(n43039), .o(n2160) );
na02f01 g39252 ( .a(n32732), .b(cos_out_7), .o(n43044) );
no02f01 g39253 ( .a(n36248), .b(n35944), .o(n43045) );
no03f01 g39254 ( .a(n36266), .b(n43045), .c(n36253), .o(n43046) );
in01f01 g39255 ( .a(n43046), .o(n43047) );
no02f01 g39256 ( .a(n36261), .b(n35944), .o(n43048) );
no02f01 g39257 ( .a(n43048), .b(n36263), .o(n43049) );
in01f01 g39258 ( .a(n43049), .o(n43050) );
no02f01 g39259 ( .a(n43050), .b(n43047), .o(n43051) );
no02f01 g39260 ( .a(n43049), .b(n43046), .o(n43052) );
oa12f01 g39261 ( .a(n32734), .b(n43052), .c(n43051), .o(n43053) );
na02f01 g39262 ( .a(n43053), .b(n43044), .o(n2165) );
no02f01 g39263 ( .a(n42214), .b(n10980), .o(n43055) );
na02f01 g39264 ( .a(n43055), .b(n10976), .o(n43056) );
in01f01 g39265 ( .a(n10976), .o(n43057) );
in01f01 g39266 ( .a(n43055), .o(n43058) );
na02f01 g39267 ( .a(n43058), .b(n43057), .o(n43059) );
na02f01 g39268 ( .a(n43059), .b(n43056), .o(n2169) );
no02f01 g39269 ( .a(n41166), .b(n41010), .o(n43061) );
na03f01 g39270 ( .a(n43061), .b(n41168), .c(n41176), .o(n43062) );
in01f01 g39271 ( .a(n43061), .o(n43063) );
oa12f01 g39272 ( .a(n43063), .b(n41169), .c(n41167), .o(n43064) );
na03f01 g39273 ( .a(n43064), .b(n43062), .c(n3633), .o(n43065) );
na02f01 g39274 ( .a(n43064), .b(n43062), .o(n5578) );
na02f01 g39275 ( .a(n5578), .b(n6203), .o(n43067) );
na02f01 g39276 ( .a(n43067), .b(n43065), .o(n2174) );
na02f01 g39277 ( .a(n8675), .b(n8661), .o(n43069) );
no02f01 g39278 ( .a(n8683), .b(n8471), .o(n43070) );
in01f01 g39279 ( .a(n43070), .o(n43071) );
na02f01 g39280 ( .a(n43071), .b(n43069), .o(n43072) );
no02f01 g39281 ( .a(n8692), .b(n8471), .o(n43073) );
no02f01 g39282 ( .a(n8691), .b(n5973), .o(n43074) );
no02f01 g39283 ( .a(n43074), .b(n43073), .o(n43075) );
na03f01 g39284 ( .a(n43075), .b(n43072), .c(n8752), .o(n43076) );
na02f01 g39285 ( .a(n43072), .b(n8752), .o(n43077) );
in01f01 g39286 ( .a(n43075), .o(n43078) );
na02f01 g39287 ( .a(n43078), .b(n43077), .o(n43079) );
na02f01 g39288 ( .a(n43079), .b(n43076), .o(n2179) );
in01f01 g39289 ( .a(n22571), .o(n43081) );
no02f01 g39290 ( .a(n22591), .b(n22587), .o(n43082) );
na02f01 g39291 ( .a(n43082), .b(n43081), .o(n43083) );
in01f01 g39292 ( .a(n43082), .o(n43084) );
na02f01 g39293 ( .a(n43084), .b(n22571), .o(n43085) );
na02f01 g39294 ( .a(n43085), .b(n43083), .o(n2184) );
no02f01 g39295 ( .a(n11624), .b(n11618), .o(n43087) );
na02f01 g39296 ( .a(n43087), .b(n11621), .o(n43088) );
in01f01 g39297 ( .a(n43087), .o(n43089) );
na02f01 g39298 ( .a(n43089), .b(n11622), .o(n43090) );
na02f01 g39299 ( .a(n43090), .b(n43088), .o(n2189) );
na02f01 g39300 ( .a(n32732), .b(sin_out_15), .o(n43092) );
no02f01 g39301 ( .a(n39575), .b(n34307), .o(n43093) );
in01f01 g39302 ( .a(n43093), .o(n43094) );
na02f01 g39303 ( .a(n43094), .b(n39594), .o(n43095) );
ao12f01 g39304 ( .a(n43095), .b(n39578), .c(n39496), .o(n43096) );
in01f01 g39305 ( .a(n43096), .o(n43097) );
no02f01 g39306 ( .a(n39588), .b(n34307), .o(n43098) );
no02f01 g39307 ( .a(n43098), .b(n39590), .o(n43099) );
in01f01 g39308 ( .a(n43099), .o(n43100) );
no02f01 g39309 ( .a(n43100), .b(n43097), .o(n43101) );
no02f01 g39310 ( .a(n43099), .b(n43096), .o(n43102) );
oa12f01 g39311 ( .a(n32734), .b(n43102), .c(n43101), .o(n43103) );
na02f01 g39312 ( .a(n43103), .b(n43092), .o(n2194) );
no02f01 g39313 ( .a(n40652), .b(n40648), .o(n43105) );
no02f01 g39314 ( .a(n43105), .b(n21270), .o(n43106) );
in01f01 g39315 ( .a(n43106), .o(n43107) );
na02f01 g39316 ( .a(n43105), .b(n21270), .o(n43108) );
na02f01 g39317 ( .a(n43108), .b(n43107), .o(n43109) );
in01f01 g39318 ( .a(n43109), .o(n43110) );
ao12f01 g39319 ( .a(n21305), .b(n40779), .c(n40784), .o(n43111) );
no02f01 g39320 ( .a(n40736), .b(n21305), .o(n43112) );
no02f01 g39321 ( .a(n43112), .b(n43111), .o(n43113) );
na02f01 g39322 ( .a(n43113), .b(n41381), .o(n43114) );
no02f01 g39323 ( .a(n43114), .b(n21264), .o(n43115) );
ao12f01 g39324 ( .a(n21270), .b(n40725), .c(n40744), .o(n43116) );
oa12f01 g39325 ( .a(n21305), .b(n43116), .c(n40736), .o(n43117) );
na02f01 g39326 ( .a(n43117), .b(n41385), .o(n43118) );
no02f01 g39327 ( .a(n43118), .b(n43115), .o(n43119) );
na02f01 g39328 ( .a(n43119), .b(n43110), .o(n43120) );
in01f01 g39329 ( .a(n43118), .o(n43121) );
oa12f01 g39330 ( .a(n43121), .b(n43114), .c(n21264), .o(n43122) );
na02f01 g39331 ( .a(n43122), .b(n43109), .o(n43123) );
na03f01 g39332 ( .a(n43123), .b(n43120), .c(n5799), .o(n43124) );
no02f01 g39333 ( .a(n43122), .b(n43109), .o(n43125) );
no02f01 g39334 ( .a(n43119), .b(n43110), .o(n43126) );
oa12f01 g39335 ( .a(n911), .b(n43126), .c(n43125), .o(n43127) );
na02f01 g39336 ( .a(n43127), .b(n43124), .o(n2198) );
in01f01 g39337 ( .a(n41198), .o(n43129) );
no02f01 g39338 ( .a(n40791), .b(n20431), .o(n43130) );
no02f01 g39339 ( .a(n43130), .b(n43129), .o(n43131) );
in01f01 g39340 ( .a(n43131), .o(n43132) );
no02f01 g39341 ( .a(n40791), .b(n20349), .o(n43133) );
in01f01 g39342 ( .a(n43133), .o(n43134) );
na03f01 g39343 ( .a(n43134), .b(n41196), .c(n41209), .o(n43135) );
na03f01 g39344 ( .a(n43135), .b(n43132), .c(n41199), .o(n43136) );
in01f01 g39345 ( .a(n41199), .o(n43137) );
no03f01 g39346 ( .a(n43133), .b(n41197), .c(n41193), .o(n43138) );
oa12f01 g39347 ( .a(n43131), .b(n43138), .c(n43137), .o(n43139) );
na03f01 g39348 ( .a(n43139), .b(n43136), .c(n5799), .o(n43140) );
no03f01 g39349 ( .a(n43138), .b(n43131), .c(n43137), .o(n43141) );
ao12f01 g39350 ( .a(n43132), .b(n43135), .c(n41199), .o(n43142) );
oa12f01 g39351 ( .a(n911), .b(n43142), .c(n43141), .o(n43143) );
na02f01 g39352 ( .a(n43143), .b(n43140), .o(n2203) );
oa12f01 g39353 ( .a(n39110), .b(n38405), .c(n39089), .o(n43145) );
na03f01 g39354 ( .a(n39111), .b(n38404), .c(n38360), .o(n43146) );
na02f01 g39355 ( .a(n43146), .b(n43145), .o(n2208) );
na03f01 g39356 ( .a(n37147), .b(n37136), .c(n6037), .o(n43148) );
na02f01 g39357 ( .a(n534), .b(n5873), .o(n43149) );
na02f01 g39358 ( .a(n43149), .b(n43148), .o(n2218) );
na02f01 g39359 ( .a(n32732), .b(cos_out_6), .o(n43151) );
no02f01 g39360 ( .a(n35965), .b(n35978), .o(n43152) );
in01f01 g39361 ( .a(n36241), .o(n43153) );
ao12f01 g39362 ( .a(n36266), .b(n43153), .c(n43152), .o(n43154) );
in01f01 g39363 ( .a(n43154), .o(n43155) );
no02f01 g39364 ( .a(n43045), .b(n36250), .o(n43156) );
in01f01 g39365 ( .a(n43156), .o(n43157) );
no02f01 g39366 ( .a(n43157), .b(n43155), .o(n43158) );
no02f01 g39367 ( .a(n43156), .b(n43154), .o(n43159) );
oa12f01 g39368 ( .a(n32734), .b(n43159), .c(n43158), .o(n43160) );
na02f01 g39369 ( .a(n43160), .b(n43151), .o(n2223) );
na02f01 g39370 ( .a(n604), .b(n4116), .o(n43162) );
na02f01 g39371 ( .a(n38183), .b(n2589), .o(n43163) );
na02f01 g39372 ( .a(n43163), .b(n43162), .o(n2227) );
in01f01 g39373 ( .a(n21205), .o(n43165) );
in01f01 g39374 ( .a(n21206), .o(n43166) );
no02f01 g39375 ( .a(n43166), .b(n21093), .o(n43167) );
na02f01 g39376 ( .a(n43167), .b(n43165), .o(n43168) );
oa12f01 g39377 ( .a(n21205), .b(n43166), .c(n21093), .o(n43169) );
na02f01 g39378 ( .a(n43169), .b(n43168), .o(n2232) );
na02f01 g39379 ( .a(n41251), .b(n41242), .o(n2237) );
na03f01 g39380 ( .a(n39449), .b(n40009), .c(n39398), .o(n43172) );
oa12f01 g39381 ( .a(n40026), .b(n39399), .c(n40008), .o(n43173) );
na02f01 g39382 ( .a(n43173), .b(n43172), .o(n2242) );
no02f01 g39383 ( .a(n36094), .b(n36076), .o(n43175) );
oa12f01 g39384 ( .a(n43175), .b(n38779), .c(n36107), .o(n43176) );
in01f01 g39385 ( .a(n43175), .o(n43177) );
na03f01 g39386 ( .a(n36117), .b(n38776), .c(n43177), .o(n43178) );
na02f01 g39387 ( .a(n43178), .b(n43176), .o(n2247) );
in01f01 g39388 ( .a(n41420), .o(n43180) );
ao12f01 g39389 ( .a(n41418), .b(n43180), .c(n41423), .o(n43181) );
in01f01 g39390 ( .a(n36181), .o(n43182) );
no02f01 g39391 ( .a(n43182), .b(n36038), .o(n43183) );
no02f01 g39392 ( .a(n36181), .b(n36122), .o(n43184) );
no02f01 g39393 ( .a(n43184), .b(n43183), .o(n43185) );
na02f01 g39394 ( .a(n43185), .b(n43181), .o(n43186) );
in01f01 g39395 ( .a(n43181), .o(n43187) );
in01f01 g39396 ( .a(n43185), .o(n43188) );
na02f01 g39397 ( .a(n43188), .b(n43187), .o(n43189) );
na02f01 g39398 ( .a(n43189), .b(n43186), .o(n2252) );
no02f01 g39399 ( .a(n10991), .b(n10787), .o(n43191) );
na02f01 g39400 ( .a(n43191), .b(n42173), .o(n43192) );
in01f01 g39401 ( .a(n43191), .o(n43193) );
oa12f01 g39402 ( .a(n43193), .b(n10989), .c(n42172), .o(n43194) );
na02f01 g39403 ( .a(n43194), .b(n43192), .o(n2257) );
ao12f01 g39404 ( .a(n27625), .b(n27525), .c(n27671), .o(n43196) );
no02f01 g39405 ( .a(n42995), .b(n27505), .o(n43197) );
na02f01 g39406 ( .a(n43197), .b(n43196), .o(n43198) );
in01f01 g39407 ( .a(n43196), .o(n43199) );
in01f01 g39408 ( .a(n43197), .o(n43200) );
na02f01 g39409 ( .a(n43200), .b(n43199), .o(n43201) );
na02f01 g39410 ( .a(n43201), .b(n43198), .o(n2262) );
in01f01 g39411 ( .a(n22296), .o(n43203) );
no02f01 g39412 ( .a(n22314), .b(n22302), .o(n43204) );
in01f01 g39413 ( .a(n43204), .o(n43205) );
no02f01 g39414 ( .a(n43205), .b(n43203), .o(n43206) );
no02f01 g39415 ( .a(n43204), .b(n22296), .o(n43207) );
no02f01 g39416 ( .a(n43207), .b(n43206), .o(n43208) );
in01f01 g39417 ( .a(n43208), .o(n2267) );
in01f01 g39418 ( .a(n35279), .o(n43210) );
in01f01 g39419 ( .a(n35280), .o(n43211) );
oa22f01 g39420 ( .a(n35300), .b(n35288), .c(n43211), .d(n43210), .o(n43212) );
no02f01 g39421 ( .a(n35300), .b(n35288), .o(n43213) );
na03f01 g39422 ( .a(n43213), .b(n35280), .c(n35279), .o(n43214) );
na02f01 g39423 ( .a(n43214), .b(n43212), .o(n2272) );
no02f01 g39424 ( .a(n8483), .b(n8471), .o(n43216) );
in01f01 g39425 ( .a(n8483), .o(n43217) );
no02f01 g39426 ( .a(n43217), .b(n5973), .o(n43218) );
no02f01 g39427 ( .a(n43218), .b(n43216), .o(n43219) );
na03f01 g39428 ( .a(n43219), .b(n8476), .c(n8474), .o(n43220) );
in01f01 g39429 ( .a(n8474), .o(n43221) );
in01f01 g39430 ( .a(n43219), .o(n43222) );
oa12f01 g39431 ( .a(n43222), .b(n8475), .c(n43221), .o(n43223) );
na02f01 g39432 ( .a(n43223), .b(n43220), .o(n2277) );
na04f01 g39433 ( .a(n36661), .b(n25487), .c(n25364), .d(n36620), .o(n43225) );
oa22f01 g39434 ( .a(n25491), .b(n25355), .c(n36660), .d(n25363), .o(n43226) );
na02f01 g39435 ( .a(n43226), .b(n43225), .o(n2282) );
in01f01 g39436 ( .a(n39631), .o(n43228) );
ao12f01 g39437 ( .a(n8899), .b(n39629), .c(n9594), .o(n43229) );
in01f01 g39438 ( .a(n43229), .o(n43230) );
no02f01 g39439 ( .a(n43230), .b(n43228), .o(n43231) );
no02f01 g39440 ( .a(n43229), .b(n39631), .o(n43232) );
no02f01 g39441 ( .a(n43232), .b(n43231), .o(n43233) );
in01f01 g39442 ( .a(n43233), .o(n2287) );
no02f01 g39443 ( .a(n11693), .b(n11571), .o(n43235) );
na02f01 g39444 ( .a(n43235), .b(n11691), .o(n43236) );
in01f01 g39445 ( .a(n11691), .o(n43237) );
in01f01 g39446 ( .a(n43235), .o(n43238) );
na02f01 g39447 ( .a(n43238), .b(n43237), .o(n43239) );
na02f01 g39448 ( .a(n43239), .b(n43236), .o(n2292) );
na02f01 g39449 ( .a(n624), .b(n8066), .o(n43241) );
na03f01 g39450 ( .a(n38564), .b(n38559), .c(n1821), .o(n43242) );
na02f01 g39451 ( .a(n43242), .b(n43241), .o(n2297) );
no03f01 g39452 ( .a(n39629), .b(n9595), .c(n8899), .o(n43244) );
no02f01 g39453 ( .a(n3623), .b(n39831), .o(n43245) );
no02f01 g39454 ( .a(n43245), .b(n43244), .o(n43246) );
in01f01 g39455 ( .a(n43246), .o(n2302) );
na03f01 g39456 ( .a(n43246), .b(n9590), .c(n9589), .o(n43248) );
oa12f01 g39457 ( .a(n2302), .b(n9646), .c(n9645), .o(n43249) );
na02f01 g39458 ( .a(n43249), .b(n43248), .o(n2307) );
na02f01 g39459 ( .a(n41984), .b(n41983), .o(n2312) );
no02f01 g39460 ( .a(n32086), .b(n39524), .o(n43252) );
oa12f01 g39461 ( .a(n43252), .b(n32424), .c(n39522), .o(n43253) );
in01f01 g39462 ( .a(n43253), .o(n43254) );
no02f01 g39463 ( .a(n32062), .b(n31607), .o(n43255) );
no02f01 g39464 ( .a(n43255), .b(n32420), .o(n43256) );
na02f01 g39465 ( .a(n43256), .b(n43254), .o(n43257) );
in01f01 g39466 ( .a(n43256), .o(n43258) );
na02f01 g39467 ( .a(n43258), .b(n43253), .o(n43259) );
na02f01 g39468 ( .a(n43259), .b(n43257), .o(n2317) );
na02f01 g39469 ( .a(n41686), .b(n36501), .o(n43261) );
oa12f01 g39470 ( .a(n41698), .b(n41692), .c(n41691), .o(n43262) );
no02f01 g39471 ( .a(n36432), .b(n21959), .o(n43263) );
no02f01 g39472 ( .a(n36447), .b(n21841), .o(n43264) );
no02f01 g39473 ( .a(n43264), .b(n43263), .o(n43265) );
na03f01 g39474 ( .a(n43265), .b(n43262), .c(n43261), .o(n43266) );
no02f01 g39475 ( .a(n41699), .b(n36461), .o(n43267) );
ao12f01 g39476 ( .a(n36448), .b(n41702), .c(n41701), .o(n43268) );
in01f01 g39477 ( .a(n43265), .o(n43269) );
oa12f01 g39478 ( .a(n43269), .b(n43268), .c(n43267), .o(n43270) );
na02f01 g39479 ( .a(n43270), .b(n43266), .o(n3120) );
na02f01 g39480 ( .a(n3120), .b(n4116), .o(n43272) );
na03f01 g39481 ( .a(n43270), .b(n43266), .c(n2589), .o(n43273) );
na02f01 g39482 ( .a(n43273), .b(n43272), .o(n2322) );
no02f01 g39483 ( .a(n40744), .b(n21270), .o(n43275) );
no02f01 g39484 ( .a(n40784), .b(n21305), .o(n43276) );
no02f01 g39485 ( .a(n43276), .b(n43275), .o(n43277) );
no03f01 g39486 ( .a(n41387), .b(n41394), .c(n41393), .o(n43278) );
oa12f01 g39487 ( .a(n43277), .b(n43278), .c(n41386), .o(n43279) );
in01f01 g39488 ( .a(n41386), .o(n43280) );
in01f01 g39489 ( .a(n43277), .o(n43281) );
in01f01 g39490 ( .a(n41387), .o(n43282) );
na03f01 g39491 ( .a(n43282), .b(n41385), .c(n41382), .o(n43283) );
na03f01 g39492 ( .a(n43283), .b(n43281), .c(n43280), .o(n43284) );
na02f01 g39493 ( .a(n43284), .b(n43279), .o(n2327) );
no02f01 g39494 ( .a(n40313), .b(n40265), .o(n43286) );
na03f01 g39495 ( .a(n43286), .b(n41885), .c(n41892), .o(n43287) );
in01f01 g39496 ( .a(n43286), .o(n43288) );
oa12f01 g39497 ( .a(n43288), .b(n41886), .c(n41884), .o(n43289) );
na02f01 g39498 ( .a(n43289), .b(n43287), .o(n2332) );
na04f01 g39499 ( .a(n29712), .b(n29710), .c(n29673), .d(n29672), .o(n43291) );
oa22f01 g39500 ( .a(n29416), .b(n29281), .c(n29412), .d(n29292), .o(n43292) );
na02f01 g39501 ( .a(n43292), .b(n43291), .o(n2337) );
na02f01 g39502 ( .a(n39171), .b(n39167), .o(n43294) );
no02f01 g39503 ( .a(n43294), .b(n39066), .o(n43295) );
no02f01 g39504 ( .a(n39154), .b(n43295), .o(n43296) );
no02f01 g39505 ( .a(n39135), .b(n32240), .o(n43297) );
no02f01 g39506 ( .a(n43297), .b(n39139), .o(n43298) );
na02f01 g39507 ( .a(n43298), .b(n43296), .o(n43299) );
in01f01 g39508 ( .a(n43298), .o(n43300) );
oa12f01 g39509 ( .a(n43300), .b(n39154), .c(n43295), .o(n43301) );
na03f01 g39510 ( .a(n43301), .b(n43299), .c(n3633), .o(n43302) );
na02f01 g39511 ( .a(n43301), .b(n43299), .o(n4275) );
na02f01 g39512 ( .a(n4275), .b(n6203), .o(n43304) );
na02f01 g39513 ( .a(n43304), .b(n43302), .o(n2342) );
no02f01 g39514 ( .a(n29860), .b(n29856), .o(n43306) );
na02f01 g39515 ( .a(n43306), .b(n29858), .o(n43307) );
in01f01 g39516 ( .a(n25663), .o(n43308) );
na02f01 g39517 ( .a(n43308), .b(n25667), .o(n43309) );
in01f01 g39518 ( .a(n43306), .o(n43310) );
na03f01 g39519 ( .a(n43310), .b(n43309), .c(n29857), .o(n43311) );
na02f01 g39520 ( .a(n43311), .b(n43307), .o(n2347) );
no02f01 g39521 ( .a(n39860), .b(n28973), .o(n43313) );
no02f01 g39522 ( .a(n43313), .b(n40564), .o(n43314) );
in01f01 g39523 ( .a(n43314), .o(n43315) );
oa12f01 g39524 ( .a(n43315), .b(n40581), .c(n40591), .o(n43316) );
na03f01 g39525 ( .a(n43314), .b(n40582), .c(n40578), .o(n43317) );
na03f01 g39526 ( .a(n43317), .b(n43316), .c(n_27923), .o(n43318) );
na02f01 g39527 ( .a(n43317), .b(n43316), .o(n4399) );
na02f01 g39528 ( .a(n4399), .b(n34420), .o(n43320) );
na02f01 g39529 ( .a(n43320), .b(n43318), .o(n2352) );
oa12f01 g39530 ( .a(n32332), .b(n32335), .c(n32270), .o(n43322) );
na03f01 g39531 ( .a(n32465), .b(n32464), .c(n32271), .o(n43323) );
na02f01 g39532 ( .a(n43323), .b(n43322), .o(n2357) );
no02f01 g39533 ( .a(n21230), .b(n21227), .o(n43325) );
no02f01 g39534 ( .a(n43325), .b(n42506), .o(n43326) );
na02f01 g39535 ( .a(n43325), .b(n42506), .o(n43327) );
in01f01 g39536 ( .a(n43327), .o(n43328) );
no02f01 g39537 ( .a(n43328), .b(n43326), .o(n43329) );
na02f01 g39538 ( .a(n43329), .b(n5799), .o(n43330) );
in01f01 g39539 ( .a(n43329), .o(n3653) );
na02f01 g39540 ( .a(n3653), .b(n911), .o(n43332) );
na02f01 g39541 ( .a(n43332), .b(n43330), .o(n2362) );
na03f01 g39542 ( .a(n37173), .b(n37031), .c(n37165), .o(n43334) );
oa12f01 g39543 ( .a(n37017), .b(n37039), .c(n37170), .o(n43335) );
na02f01 g39544 ( .a(n43335), .b(n43334), .o(n2367) );
in01f01 g39545 ( .a(n10057), .o(n43337) );
na03f01 g39546 ( .a(n10058), .b(n43337), .c(delay_sub_ln23_0_unr24_stage8_stallmux_q_0_), .o(n43338) );
in01f01 g39547 ( .a(n10058), .o(n43339) );
oa12f01 g39548 ( .a(n9907), .b(n43339), .c(n10057), .o(n43340) );
na02f01 g39549 ( .a(n43340), .b(n43338), .o(n2372) );
no02f01 g39550 ( .a(n43133), .b(n43137), .o(n43342) );
na03f01 g39551 ( .a(n43342), .b(n41196), .c(n41209), .o(n43343) );
oa22f01 g39552 ( .a(n43133), .b(n43137), .c(n41197), .d(n41193), .o(n43344) );
na03f01 g39553 ( .a(n43344), .b(n43343), .c(n5799), .o(n43345) );
na02f01 g39554 ( .a(n43344), .b(n43343), .o(n4126) );
na02f01 g39555 ( .a(n4126), .b(n911), .o(n43347) );
na02f01 g39556 ( .a(n43347), .b(n43345), .o(n2382) );
na03f01 g39557 ( .a(n39837), .b(n9590), .c(n9589), .o(n43349) );
oa12f01 g39558 ( .a(n921), .b(n9646), .c(n9645), .o(n43350) );
na02f01 g39559 ( .a(n43350), .b(n43349), .o(n2387) );
na02f01 g39560 ( .a(n39631), .b(n37390), .o(n43352) );
na02f01 g39561 ( .a(n43228), .b(n39621), .o(n43353) );
na02f01 g39562 ( .a(n43353), .b(n43352), .o(n2392) );
na02f01 g39563 ( .a(n22249), .b(n22247), .o(n43355) );
no02f01 g39564 ( .a(n43355), .b(n22239), .o(n43356) );
na02f01 g39565 ( .a(n43355), .b(n22239), .o(n43357) );
in01f01 g39566 ( .a(n43357), .o(n43358) );
no02f01 g39567 ( .a(n43358), .b(n43356), .o(n43359) );
in01f01 g39568 ( .a(n43359), .o(n4181) );
na02f01 g39569 ( .a(n4181), .b(n4116), .o(n43361) );
na02f01 g39570 ( .a(n43359), .b(n2589), .o(n43362) );
na02f01 g39571 ( .a(n43362), .b(n43361), .o(n2397) );
in01f01 g39572 ( .a(n21207), .o(n43364) );
in01f01 g39573 ( .a(n21080), .o(n43365) );
no02f01 g39574 ( .a(n21208), .b(n43365), .o(n43366) );
in01f01 g39575 ( .a(n43366), .o(n43367) );
no02f01 g39576 ( .a(n43367), .b(n43364), .o(n43368) );
no02f01 g39577 ( .a(n43366), .b(n21207), .o(n43369) );
no02f01 g39578 ( .a(n43369), .b(n43368), .o(n43370) );
in01f01 g39579 ( .a(n43370), .o(n2402) );
no02f01 g39580 ( .a(n42875), .b(n42869), .o(n43372) );
no02f01 g39581 ( .a(n42831), .b(n4176), .o(n43373) );
no02f01 g39582 ( .a(n43373), .b(n42877), .o(n43374) );
na02f01 g39583 ( .a(n43374), .b(n43372), .o(n43375) );
in01f01 g39584 ( .a(n43374), .o(n43376) );
oa12f01 g39585 ( .a(n43376), .b(n42875), .c(n42869), .o(n43377) );
na02f01 g39586 ( .a(n43377), .b(n43375), .o(n2407) );
no02f01 g39587 ( .a(n38004), .b(n38046), .o(n43379) );
ao12f01 g39588 ( .a(n37913), .b(n43379), .c(n37918), .o(n43380) );
no02f01 g39589 ( .a(n37871), .b(n37874), .o(n43381) );
no02f01 g39590 ( .a(n38010), .b(n38027), .o(n43382) );
no02f01 g39591 ( .a(n43382), .b(n43381), .o(n43383) );
no02f01 g39592 ( .a(n43383), .b(n43380), .o(n43384) );
in01f01 g39593 ( .a(n43384), .o(n43385) );
na02f01 g39594 ( .a(n43383), .b(n43380), .o(n43386) );
na03f01 g39595 ( .a(n43386), .b(n43385), .c(n1821), .o(n43387) );
na02f01 g39596 ( .a(n43386), .b(n43385), .o(n5100) );
na02f01 g39597 ( .a(n5100), .b(n8066), .o(n43389) );
na02f01 g39598 ( .a(n43389), .b(n43387), .o(n2412) );
in01f01 g39599 ( .a(mux_while_ln12_psv_q_4_), .o(n43391) );
no03f01 g39600 ( .a(n41416), .b(n43391), .c(n41414), .o(n2417) );
in01f01 g39601 ( .a(n22587), .o(n43393) );
ao12f01 g39602 ( .a(n22591), .b(n43393), .c(n22571), .o(n43394) );
no02f01 g39603 ( .a(n22590), .b(n22579), .o(n43395) );
na02f01 g39604 ( .a(n43395), .b(n43394), .o(n43396) );
in01f01 g39605 ( .a(n43394), .o(n43397) );
in01f01 g39606 ( .a(n43395), .o(n43398) );
na02f01 g39607 ( .a(n43398), .b(n43397), .o(n43399) );
na02f01 g39608 ( .a(n43399), .b(n43396), .o(n2422) );
na02f01 g39609 ( .a(n42725), .b(n42724), .o(n2427) );
in01f01 g39610 ( .a(n10834), .o(n43402) );
oa12f01 g39611 ( .a(n43402), .b(n10854), .c(n10843), .o(n43403) );
no02f01 g39612 ( .a(n10854), .b(n10843), .o(n43404) );
na02f01 g39613 ( .a(n43404), .b(n10834), .o(n43405) );
na02f01 g39614 ( .a(n43405), .b(n43403), .o(n2432) );
in01f01 g39615 ( .a(n22619), .o(n43407) );
ao12f01 g39616 ( .a(n22623), .b(n43407), .c(n22600), .o(n43408) );
no02f01 g39617 ( .a(n22622), .b(n22608), .o(n43409) );
na02f01 g39618 ( .a(n43409), .b(n43408), .o(n43410) );
in01f01 g39619 ( .a(n43408), .o(n43411) );
in01f01 g39620 ( .a(n43409), .o(n43412) );
na02f01 g39621 ( .a(n43412), .b(n43411), .o(n43413) );
na02f01 g39622 ( .a(n43413), .b(n43410), .o(n2437) );
no02f01 g39623 ( .a(n16209), .b(n16155), .o(n43415) );
no02f01 g39624 ( .a(n16208), .b(n16329), .o(n43416) );
in01f01 g39625 ( .a(n43416), .o(n43417) );
no02f01 g39626 ( .a(n16150), .b(n16089), .o(n43418) );
in01f01 g39627 ( .a(n16233), .o(n43419) );
ao12f01 g39628 ( .a(n43419), .b(n21367), .c(n43418), .o(n43420) );
ao12f01 g39629 ( .a(n43415), .b(n43420), .c(n43417), .o(n43421) );
no02f01 g39630 ( .a(n16228), .b(n16155), .o(n43422) );
no02f01 g39631 ( .a(n16227), .b(n16329), .o(n43423) );
no02f01 g39632 ( .a(n43423), .b(n43422), .o(n43424) );
in01f01 g39633 ( .a(n43424), .o(n43425) );
na02f01 g39634 ( .a(n43425), .b(n43421), .o(n43426) );
in01f01 g39635 ( .a(n43421), .o(n43427) );
na02f01 g39636 ( .a(n43424), .b(n43427), .o(n43428) );
na02f01 g39637 ( .a(n43428), .b(n43426), .o(n2442) );
na02f01 g39638 ( .a(n32732), .b(sin_out_22), .o(n43430) );
na02f01 g39639 ( .a(n41315), .b(n41294), .o(n43431) );
no02f01 g39640 ( .a(n41334), .b(n43431), .o(n43432) );
no02f01 g39641 ( .a(n41369), .b(n34307), .o(n43433) );
no02f01 g39642 ( .a(n43433), .b(n41351), .o(n43434) );
in01f01 g39643 ( .a(n43434), .o(n43435) );
no03f01 g39644 ( .a(n43435), .b(n43432), .c(n41367), .o(n43436) );
no02f01 g39645 ( .a(n43432), .b(n41367), .o(n43437) );
no02f01 g39646 ( .a(n43434), .b(n43437), .o(n43438) );
oa12f01 g39647 ( .a(n32734), .b(n43438), .c(n43436), .o(n43439) );
na02f01 g39648 ( .a(n43439), .b(n43430), .o(n2447) );
no02f01 g39649 ( .a(n22623), .b(n22619), .o(n43441) );
in01f01 g39650 ( .a(n43441), .o(n43442) );
na02f01 g39651 ( .a(n43442), .b(n22600), .o(n43443) );
in01f01 g39652 ( .a(n22600), .o(n43444) );
na02f01 g39653 ( .a(n43441), .b(n43444), .o(n43445) );
na02f01 g39654 ( .a(n43445), .b(n43443), .o(n2451) );
na03f01 g39655 ( .a(n41518), .b(n41512), .c(n6037), .o(n43447) );
ao12f01 g39656 ( .a(n41514), .b(n41517), .c(n41513), .o(n43448) );
no03f01 g39657 ( .a(n41511), .b(n41507), .c(n25159), .o(n43449) );
oa12f01 g39658 ( .a(n5873), .b(n43449), .c(n43448), .o(n43450) );
na02f01 g39659 ( .a(n43450), .b(n43447), .o(n2456) );
na03f01 g39660 ( .a(n42126), .b(n42124), .c(n1821), .o(n43452) );
in01f01 g39661 ( .a(n42124), .o(n43453) );
oa12f01 g39662 ( .a(n8066), .b(n42125), .c(n43453), .o(n43454) );
na02f01 g39663 ( .a(n43454), .b(n43452), .o(n2461) );
no02f01 g39664 ( .a(n41801), .b(n41797), .o(n43456) );
na03f01 g39665 ( .a(n43456), .b(n41809), .c(n41808), .o(n43457) );
in01f01 g39666 ( .a(n43456), .o(n43458) );
oa12f01 g39667 ( .a(n43458), .b(n41803), .c(n27121), .o(n43459) );
na03f01 g39668 ( .a(n43459), .b(n43457), .c(n1821), .o(n43460) );
na02f01 g39669 ( .a(n43459), .b(n43457), .o(n5031) );
na02f01 g39670 ( .a(n5031), .b(n8066), .o(n43462) );
na02f01 g39671 ( .a(n43462), .b(n43460), .o(n2466) );
no02f01 g39672 ( .a(n42397), .b(n42393), .o(n43464) );
na02f01 g39673 ( .a(n43464), .b(n41516), .o(n43465) );
in01f01 g39674 ( .a(n43464), .o(n43466) );
na02f01 g39675 ( .a(n43466), .b(n41510), .o(n43467) );
na03f01 g39676 ( .a(n43467), .b(n43465), .c(n6037), .o(n43468) );
na02f01 g39677 ( .a(n43467), .b(n43465), .o(n5844) );
na02f01 g39678 ( .a(n5844), .b(n5873), .o(n43470) );
na02f01 g39679 ( .a(n43470), .b(n43468), .o(n2471) );
in01f01 g39680 ( .a(n10873), .o(n43472) );
no02f01 g39681 ( .a(n43472), .b(n10824), .o(n43473) );
no02f01 g39682 ( .a(n10869), .b(n3521), .o(n43474) );
in01f01 g39683 ( .a(n43474), .o(n43475) );
no02f01 g39684 ( .a(n10806), .b(n3521), .o(n43476) );
no02f01 g39685 ( .a(n43476), .b(n10808), .o(n43477) );
na03f01 g39686 ( .a(n43477), .b(n43475), .c(n43473), .o(n43478) );
na02f01 g39687 ( .a(n43475), .b(n43473), .o(n43479) );
in01f01 g39688 ( .a(n43477), .o(n43480) );
na02f01 g39689 ( .a(n43480), .b(n43479), .o(n43481) );
na02f01 g39690 ( .a(n43481), .b(n43478), .o(n2476) );
ao12f01 g39691 ( .a(n30035), .b(n30028), .c(n30021), .o(n43483) );
no02f01 g39692 ( .a(n30034), .b(n30031), .o(n43484) );
no02f01 g39693 ( .a(n43484), .b(n43483), .o(n43485) );
in01f01 g39694 ( .a(n43485), .o(n43486) );
na02f01 g39695 ( .a(n43484), .b(n43483), .o(n43487) );
na02f01 g39696 ( .a(n43487), .b(n43486), .o(n2481) );
na02f01 g39697 ( .a(n42560), .b(n42558), .o(n2486) );
no02f01 g39698 ( .a(n4201), .b(n8862), .o(n43490) );
no02f01 g39699 ( .a(n9591), .b(n8899), .o(n43491) );
no02f01 g39700 ( .a(n43491), .b(n43490), .o(n43492) );
na03f01 g39701 ( .a(n43492), .b(n9590), .c(n9589), .o(n43493) );
in01f01 g39702 ( .a(n43492), .o(n5345) );
oa12f01 g39703 ( .a(n5345), .b(n9646), .c(n9645), .o(n43495) );
na02f01 g39704 ( .a(n43495), .b(n43493), .o(n2491) );
na02f01 g39705 ( .a(n2013), .b(n4116), .o(n43497) );
na02f01 g39706 ( .a(n42740), .b(n2589), .o(n43498) );
na02f01 g39707 ( .a(n43498), .b(n43497), .o(n2496) );
na03f01 g39708 ( .a(n41178), .b(n41171), .c(n3633), .o(n43500) );
ao12f01 g39709 ( .a(n41173), .b(n41177), .c(n41172), .o(n43501) );
no03f01 g39710 ( .a(n41170), .b(n41165), .c(n41010), .o(n43502) );
oa12f01 g39711 ( .a(n6203), .b(n43502), .c(n43501), .o(n43503) );
na02f01 g39712 ( .a(n43503), .b(n43500), .o(n2501) );
ao12f01 g39713 ( .a(n25474), .b(n25476), .c(n25466), .o(n43505) );
in01f01 g39714 ( .a(n43505), .o(n43506) );
no02f01 g39715 ( .a(n25479), .b(n36628), .o(n43507) );
no02f01 g39716 ( .a(n25483), .b(n25380), .o(n43508) );
no02f01 g39717 ( .a(n43508), .b(n43507), .o(n43509) );
na02f01 g39718 ( .a(n43509), .b(n43506), .o(n43510) );
oa12f01 g39719 ( .a(n43505), .b(n43508), .c(n43507), .o(n43511) );
na02f01 g39720 ( .a(n43511), .b(n43510), .o(n2511) );
in01f01 g39721 ( .a(n39832), .o(n43513) );
no02f01 g39722 ( .a(n40599), .b(n43513), .o(n43514) );
no02f01 g39723 ( .a(n42473), .b(n39832), .o(n43515) );
no02f01 g39724 ( .a(n43515), .b(n43514), .o(n43516) );
in01f01 g39725 ( .a(n43516), .o(n2516) );
na02f01 g39726 ( .a(n32732), .b(sin_out_23), .o(n43518) );
no02f01 g39727 ( .a(n41368), .b(n34307), .o(n43519) );
no02f01 g39728 ( .a(n43519), .b(n41346), .o(n43520) );
in01f01 g39729 ( .a(n43520), .o(n43521) );
in01f01 g39730 ( .a(n41315), .o(n43522) );
no02f01 g39731 ( .a(n43522), .b(n39599), .o(n43523) );
no02f01 g39732 ( .a(n41351), .b(n41334), .o(n43524) );
na02f01 g39733 ( .a(n43524), .b(n43523), .o(n43525) );
no02f01 g39734 ( .a(n43433), .b(n41367), .o(n43526) );
na02f01 g39735 ( .a(n43526), .b(n43525), .o(n43527) );
no02f01 g39736 ( .a(n43527), .b(n43521), .o(n43528) );
ao12f01 g39737 ( .a(n43520), .b(n43526), .c(n43525), .o(n43529) );
oa12f01 g39738 ( .a(n32734), .b(n43529), .c(n43528), .o(n43530) );
na02f01 g39739 ( .a(n43530), .b(n43518), .o(n2521) );
in01f01 g39740 ( .a(n22626), .o(n43532) );
no02f01 g39741 ( .a(n43532), .b(n22518), .o(n43533) );
na03f01 g39742 ( .a(n43533), .b(n22624), .c(n22621), .o(n43534) );
in01f01 g39743 ( .a(n43533), .o(n43535) );
na02f01 g39744 ( .a(n43535), .b(n22625), .o(n43536) );
na02f01 g39745 ( .a(n43536), .b(n43534), .o(n2525) );
na03f01 g39746 ( .a(n42530), .b(n9590), .c(n9589), .o(n43538) );
oa12f01 g39747 ( .a(n1879), .b(n9646), .c(n9645), .o(n43539) );
na02f01 g39748 ( .a(n43539), .b(n43538), .o(n2530) );
na03f01 g39749 ( .a(n21362), .b(n21361), .c(n16076), .o(n43541) );
oa12f01 g39750 ( .a(n16084), .b(n16085), .c(n21358), .o(n43542) );
na02f01 g39751 ( .a(n43542), .b(n43541), .o(n2535) );
na02f01 g39752 ( .a(n22594), .b(n22538), .o(n43544) );
na02f01 g39753 ( .a(n43544), .b(n22593), .o(n43545) );
in01f01 g39754 ( .a(n43544), .o(n43546) );
na03f01 g39755 ( .a(n43546), .b(n22592), .c(n22589), .o(n43547) );
na02f01 g39756 ( .a(n43547), .b(n43545), .o(n2540) );
no02f01 g39757 ( .a(n25295), .b(n25557), .o(n43549) );
ao12f01 g39758 ( .a(n25561), .b(n37145), .c(n25572), .o(n43550) );
in01f01 g39759 ( .a(n43550), .o(n43551) );
na02f01 g39760 ( .a(n43551), .b(n43549), .o(n43552) );
in01f01 g39761 ( .a(n43549), .o(n43553) );
na02f01 g39762 ( .a(n43550), .b(n43553), .o(n43554) );
na03f01 g39763 ( .a(n43554), .b(n43552), .c(n6037), .o(n43555) );
na02f01 g39764 ( .a(n43554), .b(n43552), .o(n5290) );
na02f01 g39765 ( .a(n5290), .b(n5873), .o(n43557) );
na02f01 g39766 ( .a(n43557), .b(n43555), .o(n2545) );
no02f01 g39767 ( .a(n9678), .b(n36536), .o(n43559) );
no02f01 g39768 ( .a(n9694), .b(n5001), .o(n43560) );
in01f01 g39769 ( .a(n43560), .o(n43561) );
na02f01 g39770 ( .a(n9694), .b(n5001), .o(n43562) );
na02f01 g39771 ( .a(n43562), .b(n43561), .o(n43563) );
in01f01 g39772 ( .a(n43563), .o(n43564) );
na02f01 g39773 ( .a(n43564), .b(n43559), .o(n43565) );
in01f01 g39774 ( .a(n43559), .o(n43566) );
na02f01 g39775 ( .a(n43563), .b(n43566), .o(n43567) );
na02f01 g39776 ( .a(n43567), .b(n43565), .o(n2550) );
na02f01 g39777 ( .a(n38854), .b(n38850), .o(n2555) );
no02f01 g39778 ( .a(n8448), .b(n8471), .o(n43570) );
no02f01 g39779 ( .a(n8467), .b(n8471), .o(n43571) );
no02f01 g39780 ( .a(n43571), .b(n8469), .o(n43572) );
in01f01 g39781 ( .a(n43572), .o(n43573) );
oa12f01 g39782 ( .a(n43573), .b(n43570), .c(n8451), .o(n43574) );
in01f01 g39783 ( .a(n8451), .o(n43575) );
in01f01 g39784 ( .a(n43570), .o(n43576) );
na03f01 g39785 ( .a(n43572), .b(n43576), .c(n43575), .o(n43577) );
na02f01 g39786 ( .a(n43577), .b(n43574), .o(n2560) );
in01f01 g39787 ( .a(n38937), .o(n43579) );
no02f01 g39788 ( .a(n38959), .b(n38948), .o(n43580) );
in01f01 g39789 ( .a(n43580), .o(n43581) );
na02f01 g39790 ( .a(n43581), .b(n43579), .o(n43582) );
na02f01 g39791 ( .a(n43580), .b(n38937), .o(n43583) );
na02f01 g39792 ( .a(n43583), .b(n43582), .o(n2565) );
in01f01 g39793 ( .a(n25836), .o(n43585) );
in01f01 g39794 ( .a(n25844), .o(n43586) );
no02f01 g39795 ( .a(n25849), .b(n43586), .o(n43587) );
na02f01 g39796 ( .a(n25849), .b(n43586), .o(n43588) );
in01f01 g39797 ( .a(n43588), .o(n43589) );
oa12f01 g39798 ( .a(n43585), .b(n43589), .c(n43587), .o(n43590) );
in01f01 g39799 ( .a(n43587), .o(n43591) );
na03f01 g39800 ( .a(n43588), .b(n43591), .c(n25836), .o(n43592) );
na02f01 g39801 ( .a(n43592), .b(n43590), .o(n2570) );
na02f01 g39802 ( .a(n32732), .b(sin_out_4), .o(n43594) );
no02f01 g39803 ( .a(n34371), .b(n34369), .o(n43595) );
in01f01 g39804 ( .a(n43595), .o(n43596) );
no02f01 g39805 ( .a(n43596), .b(n36566), .o(n43597) );
no02f01 g39806 ( .a(n43595), .b(n34348), .o(n43598) );
oa12f01 g39807 ( .a(n32734), .b(n43598), .c(n43597), .o(n43599) );
na02f01 g39808 ( .a(n43599), .b(n43594), .o(n2575) );
no02f01 g39809 ( .a(n37303), .b(n37300), .o(n43601) );
na03f01 g39810 ( .a(n5988), .b(n43601), .c(delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(n43602) );
in01f01 g39811 ( .a(n43601), .o(n6222) );
oa12f01 g39812 ( .a(n6222), .b(n37356), .c(n37149), .o(n43604) );
na02f01 g39813 ( .a(n43604), .b(n43602), .o(n2579) );
in01f01 g39814 ( .a(n35302), .o(n43606) );
no02f01 g39815 ( .a(n35311), .b(n43606), .o(n43607) );
no02f01 g39816 ( .a(n35309), .b(n35258), .o(n43608) );
no02f01 g39817 ( .a(n35320), .b(n35258), .o(n43609) );
no02f01 g39818 ( .a(n43609), .b(n35322), .o(n43610) );
in01f01 g39819 ( .a(n43610), .o(n43611) );
oa12f01 g39820 ( .a(n43611), .b(n43608), .c(n43607), .o(n43612) );
no02f01 g39821 ( .a(n43608), .b(n43607), .o(n43613) );
na02f01 g39822 ( .a(n43610), .b(n43613), .o(n43614) );
na02f01 g39823 ( .a(n43614), .b(n43612), .o(n2584) );
in01f01 g39824 ( .a(n32034), .o(n43616) );
no02f01 g39825 ( .a(n36877), .b(n31607), .o(n43617) );
no02f01 g39826 ( .a(n36871), .b(n31606), .o(n43618) );
no02f01 g39827 ( .a(n43618), .b(n43617), .o(n43619) );
in01f01 g39828 ( .a(n32038), .o(n43620) );
oa12f01 g39829 ( .a(n43620), .b(n32496), .c(n32440), .o(n43621) );
na03f01 g39830 ( .a(n43621), .b(n43619), .c(n43616), .o(n43622) );
in01f01 g39831 ( .a(n43619), .o(n43623) );
ao12f01 g39832 ( .a(n32038), .b(n32437), .c(n32130), .o(n43624) );
oa12f01 g39833 ( .a(n43623), .b(n43624), .c(n32034), .o(n43625) );
na03f01 g39834 ( .a(n43625), .b(n43622), .c(n3633), .o(n43626) );
no03f01 g39835 ( .a(n43624), .b(n43623), .c(n32034), .o(n43627) );
ao12f01 g39836 ( .a(n43619), .b(n43621), .c(n43616), .o(n43628) );
oa12f01 g39837 ( .a(n6203), .b(n43628), .c(n43627), .o(n43629) );
na02f01 g39838 ( .a(n43629), .b(n43626), .o(n2594) );
in01f01 g39839 ( .a(n40916), .o(n43631) );
in01f01 g39840 ( .a(n40924), .o(n43632) );
oa12f01 g39841 ( .a(n43632), .b(n40926), .c(n43631), .o(n43633) );
in01f01 g39842 ( .a(n43633), .o(n43634) );
no02f01 g39843 ( .a(n40925), .b(n40897), .o(n43635) );
in01f01 g39844 ( .a(n43635), .o(n43636) );
no02f01 g39845 ( .a(n43636), .b(n43634), .o(n43637) );
no02f01 g39846 ( .a(n43635), .b(n43633), .o(n43638) );
no02f01 g39847 ( .a(n43638), .b(n43637), .o(n43639) );
na02f01 g39848 ( .a(n43639), .b(n5799), .o(n43640) );
in01f01 g39849 ( .a(n43639), .o(n4736) );
na02f01 g39850 ( .a(n4736), .b(n911), .o(n43642) );
na02f01 g39851 ( .a(n43642), .b(n43640), .o(n2599) );
na04f01 g39852 ( .a(n29715), .b(n29714), .c(n29671), .d(n29670), .o(n43644) );
oa22f01 g39853 ( .a(n29424), .b(n29213), .c(n29421), .d(n29267), .o(n43645) );
na02f01 g39854 ( .a(n43645), .b(n43644), .o(n2604) );
no02f01 g39855 ( .a(n39052), .b(n31607), .o(n43647) );
no02f01 g39856 ( .a(n39055), .b(n31606), .o(n43648) );
no02f01 g39857 ( .a(n43648), .b(n43647), .o(n43649) );
no03f01 g39858 ( .a(n39195), .b(n39189), .c(n36874), .o(n43650) );
oa12f01 g39859 ( .a(n43650), .b(n32496), .c(n32440), .o(n43651) );
no02f01 g39860 ( .a(n39192), .b(n38492), .o(n43652) );
oa12f01 g39861 ( .a(n36884), .b(n43652), .c(n31607), .o(n43653) );
in01f01 g39862 ( .a(n43653), .o(n43654) );
na03f01 g39863 ( .a(n43654), .b(n43651), .c(n43649), .o(n43655) );
in01f01 g39864 ( .a(n43649), .o(n43656) );
in01f01 g39865 ( .a(n43650), .o(n43657) );
ao12f01 g39866 ( .a(n43657), .b(n32437), .c(n32130), .o(n43658) );
oa12f01 g39867 ( .a(n43656), .b(n43653), .c(n43658), .o(n43659) );
na03f01 g39868 ( .a(n43659), .b(n43655), .c(n3633), .o(n43660) );
no03f01 g39869 ( .a(n43653), .b(n43658), .c(n43656), .o(n43661) );
ao12f01 g39870 ( .a(n43649), .b(n43654), .c(n43651), .o(n43662) );
oa12f01 g39871 ( .a(n6203), .b(n43662), .c(n43661), .o(n43663) );
na02f01 g39872 ( .a(n43663), .b(n43660), .o(n2609) );
na02f01 g39873 ( .a(n32732), .b(cos_out_18), .o(n43665) );
no02f01 g39874 ( .a(n39664), .b(n36374), .o(n43666) );
no02f01 g39875 ( .a(n39672), .b(n35944), .o(n43667) );
no02f01 g39876 ( .a(n43667), .b(n39674), .o(n43668) );
in01f01 g39877 ( .a(n43668), .o(n43669) );
no03f01 g39878 ( .a(n43669), .b(n43666), .c(n39692), .o(n43670) );
no02f01 g39879 ( .a(n43666), .b(n39692), .o(n43671) );
no02f01 g39880 ( .a(n43668), .b(n43671), .o(n43672) );
oa12f01 g39881 ( .a(n32734), .b(n43672), .c(n43670), .o(n43673) );
na02f01 g39882 ( .a(n43673), .b(n43665), .o(n2614) );
no02f01 g39883 ( .a(n22477), .b(n22392), .o(n43675) );
in01f01 g39884 ( .a(n43675), .o(n43676) );
oa12f01 g39885 ( .a(n43676), .b(n22480), .c(n25639), .o(n43677) );
na03f01 g39886 ( .a(n43675), .b(n22420), .c(n25643), .o(n43678) );
na03f01 g39887 ( .a(n43678), .b(n43677), .c(n2589), .o(n43679) );
na02f01 g39888 ( .a(n43678), .b(n43677), .o(n4667) );
na02f01 g39889 ( .a(n4667), .b(n4116), .o(n43681) );
na02f01 g39890 ( .a(n43681), .b(n43679), .o(n2618) );
no02f01 g39891 ( .a(n8439), .b(n5973), .o(n43683) );
no02f01 g39892 ( .a(n8438), .b(n8471), .o(n43684) );
no02f01 g39893 ( .a(n43684), .b(n43683), .o(n43685) );
in01f01 g39894 ( .a(n43685), .o(n43686) );
na02f01 g39895 ( .a(n43686), .b(n8431), .o(n43687) );
in01f01 g39896 ( .a(n8431), .o(n43688) );
na02f01 g39897 ( .a(n43685), .b(n43688), .o(n43689) );
na02f01 g39898 ( .a(n43689), .b(n43687), .o(n2623) );
no02f01 g39899 ( .a(n10961), .b(n3521), .o(n43691) );
no02f01 g39900 ( .a(n10962), .b(n10735), .o(n43692) );
no02f01 g39901 ( .a(n43692), .b(n43691), .o(n43693) );
na03f01 g39902 ( .a(n43693), .b(n10927), .c(n10924), .o(n43694) );
in01f01 g39903 ( .a(n43693), .o(n43695) );
na02f01 g39904 ( .a(n43695), .b(n10928), .o(n43696) );
na02f01 g39905 ( .a(n43696), .b(n43694), .o(n2628) );
na02f01 g39906 ( .a(n32732), .b(sin_out_2), .o(n43698) );
no02f01 g39907 ( .a(n34345), .b(n34303), .o(n43699) );
in01f01 g39908 ( .a(n43699), .o(n43700) );
no02f01 g39909 ( .a(n43700), .b(n36562), .o(n43701) );
no02f01 g39910 ( .a(n43699), .b(n34327), .o(n43702) );
oa12f01 g39911 ( .a(n32734), .b(n43702), .c(n43701), .o(n43703) );
na02f01 g39912 ( .a(n43703), .b(n43698), .o(n2633) );
no02f01 g39913 ( .a(n9413), .b(n9224), .o(n43705) );
no02f01 g39914 ( .a(n43705), .b(n9415), .o(n43706) );
in01f01 g39915 ( .a(n43706), .o(n43707) );
oa12f01 g39916 ( .a(n43707), .b(n9406), .c(n9329), .o(n43708) );
na03f01 g39917 ( .a(n43706), .b(n9625), .c(n9619), .o(n43709) );
na02f01 g39918 ( .a(n43709), .b(n43708), .o(n2637) );
na04f01 g39919 ( .a(n21180), .b(n21176), .c(n21172), .d(n21153), .o(n43711) );
na02f01 g39920 ( .a(n21180), .b(n21153), .o(n43712) );
na02f01 g39921 ( .a(n43712), .b(n21177), .o(n43713) );
na02f01 g39922 ( .a(n43713), .b(n43711), .o(n2642) );
no02f01 g39923 ( .a(n22598), .b(n22526), .o(n43715) );
na02f01 g39924 ( .a(n43715), .b(n22597), .o(n43716) );
in01f01 g39925 ( .a(n43715), .o(n43717) );
na02f01 g39926 ( .a(n43717), .b(n22596), .o(n43718) );
na02f01 g39927 ( .a(n43718), .b(n43716), .o(n2647) );
in01f01 g39928 ( .a(mux_while_ln12_psv_q_3_), .o(n43720) );
no03f01 g39929 ( .a(n41416), .b(n43720), .c(n41414), .o(n2652) );
ao12f01 g39930 ( .a(n38427), .b(n38432), .c(n38409), .o(n43722) );
in01f01 g39931 ( .a(n43722), .o(n43723) );
no02f01 g39932 ( .a(n38430), .b(n38337), .o(n43724) );
na02f01 g39933 ( .a(n43724), .b(n43723), .o(n43725) );
in01f01 g39934 ( .a(n43724), .o(n43726) );
na02f01 g39935 ( .a(n43726), .b(n43722), .o(n43727) );
na02f01 g39936 ( .a(n43727), .b(n43725), .o(n2657) );
in01f01 g39937 ( .a(n40322), .o(n43729) );
no02f01 g39938 ( .a(n39860), .b(n39984), .o(n43730) );
no02f01 g39939 ( .a(n39861), .b(n28934), .o(n43731) );
no02f01 g39940 ( .a(n43731), .b(n43730), .o(n43732) );
in01f01 g39941 ( .a(n40323), .o(n43733) );
oa12f01 g39942 ( .a(n43733), .b(n40327), .c(n40326), .o(n43734) );
na03f01 g39943 ( .a(n43734), .b(n43732), .c(n43729), .o(n43735) );
in01f01 g39944 ( .a(n43732), .o(n43736) );
ao12f01 g39945 ( .a(n40323), .b(n39994), .c(n40321), .o(n43737) );
oa12f01 g39946 ( .a(n43736), .b(n43737), .c(n40322), .o(n43738) );
na02f01 g39947 ( .a(n43738), .b(n43735), .o(n2662) );
no02f01 g39948 ( .a(n4201), .b(n9232), .o(n43740) );
no02f01 g39949 ( .a(n43740), .b(n42224), .o(n43741) );
na02f01 g39950 ( .a(n43740), .b(n42224), .o(n43742) );
in01f01 g39951 ( .a(n43742), .o(n43743) );
no02f01 g39952 ( .a(n43743), .b(n43741), .o(n43744) );
na03f01 g39953 ( .a(n43744), .b(n9590), .c(n9589), .o(n43745) );
in01f01 g39954 ( .a(n43744), .o(n3663) );
oa12f01 g39955 ( .a(n3663), .b(n9646), .c(n9645), .o(n43747) );
na02f01 g39956 ( .a(n43747), .b(n43745), .o(n2667) );
ao12f01 g39957 ( .a(n30115), .b(n30118), .c(n42796), .o(n43749) );
no02f01 g39958 ( .a(n30009), .b(n29991), .o(n43750) );
in01f01 g39959 ( .a(n43750), .o(n43751) );
no02f01 g39960 ( .a(n43751), .b(n43749), .o(n43752) );
na02f01 g39961 ( .a(n43751), .b(n43749), .o(n43753) );
in01f01 g39962 ( .a(n43753), .o(n43754) );
no02f01 g39963 ( .a(n43754), .b(n43752), .o(n43755) );
na02f01 g39964 ( .a(n43755), .b(n6037), .o(n43756) );
in01f01 g39965 ( .a(n43755), .o(n5735) );
na02f01 g39966 ( .a(n5735), .b(n5873), .o(n43758) );
na02f01 g39967 ( .a(n43758), .b(n43756), .o(n2677) );
no02f01 g39968 ( .a(n9430), .b(n9279), .o(n43760) );
na02f01 g39969 ( .a(n43760), .b(n9428), .o(n43761) );
in01f01 g39970 ( .a(n43760), .o(n43762) );
na02f01 g39971 ( .a(n43762), .b(n9632), .o(n43763) );
na02f01 g39972 ( .a(n43763), .b(n43761), .o(n2682) );
in01f01 g39973 ( .a(n36781), .o(n43765) );
no02f01 g39974 ( .a(n36759), .b(n29639), .o(n43766) );
no02f01 g39975 ( .a(n43766), .b(n36761), .o(n43767) );
na03f01 g39976 ( .a(n36739), .b(n29614), .c(n29721), .o(n43768) );
na03f01 g39977 ( .a(n43768), .b(n43767), .c(n43765), .o(n43769) );
in01f01 g39978 ( .a(n43767), .o(n43770) );
no03f01 g39979 ( .a(n36740), .b(n29615), .c(n29578), .o(n43771) );
oa12f01 g39980 ( .a(n43770), .b(n43771), .c(n36781), .o(n43772) );
na03f01 g39981 ( .a(n43772), .b(n43769), .c(n_27923), .o(n43773) );
na02f01 g39982 ( .a(n43772), .b(n43769), .o(n2791) );
na02f01 g39983 ( .a(n2791), .b(n34420), .o(n43775) );
na02f01 g39984 ( .a(n43775), .b(n43773), .o(n2692) );
no03f01 g39985 ( .a(n42025), .b(n42028), .c(n42009), .o(n43777) );
ao12f01 g39986 ( .a(n10733), .b(n10710), .c(n42016), .o(n43778) );
no02f01 g39987 ( .a(n10731), .b(n4088), .o(n43779) );
no02f01 g39988 ( .a(n43779), .b(n10727), .o(n43780) );
no02f01 g39989 ( .a(n43780), .b(n43778), .o(n43781) );
na02f01 g39990 ( .a(n43780), .b(n43778), .o(n43782) );
in01f01 g39991 ( .a(n43782), .o(n43783) );
no03f01 g39992 ( .a(n43783), .b(n43781), .c(n10735), .o(n43784) );
no02f01 g39993 ( .a(n43783), .b(n43781), .o(n43785) );
no02f01 g39994 ( .a(n43785), .b(n3521), .o(n43786) );
no02f01 g39995 ( .a(n43786), .b(n43784), .o(n43787) );
oa12f01 g39996 ( .a(n43787), .b(n43777), .c(n42023), .o(n43788) );
no02f01 g39997 ( .a(n43777), .b(n42023), .o(n43789) );
in01f01 g39998 ( .a(n43787), .o(n43790) );
na02f01 g39999 ( .a(n43790), .b(n43789), .o(n43791) );
na02f01 g40000 ( .a(n43791), .b(n43788), .o(n2697) );
in01f01 g40001 ( .a(n14142), .o(n43793) );
na03f01 g40002 ( .a(n14151), .b(n14150), .c(n43793), .o(n43794) );
in01f01 g40003 ( .a(n14150), .o(n43795) );
in01f01 g40004 ( .a(n14151), .o(n43796) );
oa12f01 g40005 ( .a(n43795), .b(n43796), .c(n14142), .o(n43797) );
na02f01 g40006 ( .a(n43797), .b(n43794), .o(n2702) );
no02f01 g40007 ( .a(n4201), .b(n9231), .o(n43799) );
no02f01 g40008 ( .a(n40367), .b(n43799), .o(n43800) );
no02f01 g40009 ( .a(n43800), .b(n36403), .o(n43801) );
na02f01 g40010 ( .a(n43800), .b(n36403), .o(n43802) );
in01f01 g40011 ( .a(n43802), .o(n43803) );
no02f01 g40012 ( .a(n43803), .b(n43801), .o(n43804) );
in01f01 g40013 ( .a(n43804), .o(n2707) );
in01f01 g40014 ( .a(n40406), .o(n43806) );
ao12f01 g40015 ( .a(n9707), .b(n40405), .c(n43806), .o(n43807) );
in01f01 g40016 ( .a(n43807), .o(n43808) );
no02f01 g40017 ( .a(n9716), .b(n5001), .o(n43809) );
no02f01 g40018 ( .a(n43809), .b(n9718), .o(n43810) );
na02f01 g40019 ( .a(n43810), .b(n43808), .o(n43811) );
in01f01 g40020 ( .a(n43810), .o(n43812) );
na02f01 g40021 ( .a(n43812), .b(n43807), .o(n43813) );
na02f01 g40022 ( .a(n43813), .b(n43811), .o(n2712) );
no02f01 g40023 ( .a(n41736), .b(n29639), .o(n43815) );
in01f01 g40024 ( .a(n43815), .o(n43816) );
no02f01 g40025 ( .a(n39307), .b(n29639), .o(n43817) );
no02f01 g40026 ( .a(n43817), .b(n41729), .o(n43818) );
oa12f01 g40027 ( .a(n41727), .b(n42382), .c(n42389), .o(n43819) );
na03f01 g40028 ( .a(n43819), .b(n43818), .c(n43816), .o(n43820) );
in01f01 g40029 ( .a(n43818), .o(n43821) );
in01f01 g40030 ( .a(n41727), .o(n43822) );
ao12f01 g40031 ( .a(n43822), .b(n42383), .c(n42380), .o(n43823) );
oa12f01 g40032 ( .a(n43821), .b(n43823), .c(n43815), .o(n43824) );
na02f01 g40033 ( .a(n43824), .b(n43820), .o(n2717) );
na03f01 g40034 ( .a(n36092), .b(n36089), .c(n38767), .o(n43826) );
oa12f01 g40035 ( .a(n36077), .b(n36091), .c(n36088), .o(n43827) );
na02f01 g40036 ( .a(n43827), .b(n43826), .o(n2722) );
na02f01 g40037 ( .a(n32732), .b(cos_out_15), .o(n43829) );
in01f01 g40038 ( .a(n39747), .o(n43830) );
ao12f01 g40039 ( .a(n36362), .b(n39745), .c(n43830), .o(n43831) );
no02f01 g40040 ( .a(n36353), .b(n35944), .o(n43832) );
no02f01 g40041 ( .a(n43832), .b(n36355), .o(n43833) );
in01f01 g40042 ( .a(n43833), .o(n43834) );
no02f01 g40043 ( .a(n43834), .b(n43831), .o(n43835) );
no02f01 g40044 ( .a(n39746), .b(n39747), .o(n43836) );
no03f01 g40045 ( .a(n43833), .b(n43836), .c(n36362), .o(n43837) );
oa12f01 g40046 ( .a(n32734), .b(n43837), .c(n43835), .o(n43838) );
na02f01 g40047 ( .a(n43838), .b(n43829), .o(n2727) );
in01f01 g40048 ( .a(n25035), .o(n43840) );
no02f01 g40049 ( .a(n25044), .b(n25023), .o(n43841) );
no02f01 g40050 ( .a(n43841), .b(n25046), .o(n43842) );
in01f01 g40051 ( .a(n43842), .o(n43843) );
oa12f01 g40052 ( .a(n25545), .b(n25546), .c(n25023), .o(n43844) );
ao12f01 g40053 ( .a(n43844), .b(n25538), .c(n25182), .o(n43845) );
oa12f01 g40054 ( .a(n43845), .b(n25301), .c(n25183), .o(n43846) );
na03f01 g40055 ( .a(n43846), .b(n43843), .c(n43840), .o(n43847) );
in01f01 g40056 ( .a(n43844), .o(n43848) );
na02f01 g40057 ( .a(n43848), .b(n25576), .o(n43849) );
ao12f01 g40058 ( .a(n43849), .b(n25575), .c(n25182), .o(n43850) );
oa12f01 g40059 ( .a(n43842), .b(n43850), .c(n25035), .o(n43851) );
na03f01 g40060 ( .a(n43851), .b(n43847), .c(n6037), .o(n43852) );
no03f01 g40061 ( .a(n43850), .b(n43842), .c(n25035), .o(n43853) );
ao12f01 g40062 ( .a(n43843), .b(n43846), .c(n43840), .o(n43854) );
oa12f01 g40063 ( .a(n5873), .b(n43854), .c(n43853), .o(n43855) );
na02f01 g40064 ( .a(n43855), .b(n43852), .o(n2731) );
no02f01 g40065 ( .a(n42631), .b(n27453), .o(n43857) );
na03f01 g40066 ( .a(n43857), .b(n27490), .c(n42350), .o(n43858) );
in01f01 g40067 ( .a(n43857), .o(n43859) );
oa12f01 g40068 ( .a(n43859), .b(n42354), .c(n42630), .o(n43860) );
na02f01 g40069 ( .a(n43860), .b(n43858), .o(n2736) );
no02f01 g40070 ( .a(n27078), .b(n26440), .o(n43862) );
in01f01 g40071 ( .a(n43862), .o(n43863) );
no02f01 g40072 ( .a(n27073), .b(n26440), .o(n43864) );
in01f01 g40073 ( .a(n27073), .o(n43865) );
no02f01 g40074 ( .a(n43865), .b(n26441), .o(n43866) );
no02f01 g40075 ( .a(n43866), .b(n43864), .o(n43867) );
in01f01 g40076 ( .a(n27078), .o(n43868) );
no02f01 g40077 ( .a(n43868), .b(n26441), .o(n43869) );
in01f01 g40078 ( .a(n43869), .o(n43870) );
no02f01 g40079 ( .a(n27238), .b(n26869), .o(n43871) );
na03f01 g40080 ( .a(n27109), .b(n27098), .c(n43871), .o(n43872) );
na02f01 g40081 ( .a(n43872), .b(n27116), .o(n43873) );
na02f01 g40082 ( .a(n43873), .b(n43870), .o(n43874) );
na03f01 g40083 ( .a(n43874), .b(n43867), .c(n43863), .o(n43875) );
in01f01 g40084 ( .a(n43867), .o(n43876) );
na02f01 g40085 ( .a(n27068), .b(n26870), .o(n43877) );
no03f01 g40086 ( .a(n27243), .b(n27097), .c(n43877), .o(n43878) );
no02f01 g40087 ( .a(n43878), .b(n27246), .o(n43879) );
no02f01 g40088 ( .a(n43879), .b(n43869), .o(n43880) );
oa12f01 g40089 ( .a(n43876), .b(n43880), .c(n43862), .o(n43881) );
na03f01 g40090 ( .a(n43881), .b(n43875), .c(n1821), .o(n43882) );
no03f01 g40091 ( .a(n43880), .b(n43876), .c(n43862), .o(n43883) );
ao12f01 g40092 ( .a(n43867), .b(n43874), .c(n43863), .o(n43884) );
oa12f01 g40093 ( .a(n8066), .b(n43884), .c(n43883), .o(n43885) );
na02f01 g40094 ( .a(n43885), .b(n43882), .o(n2741) );
na03f01 g40095 ( .a(n39187), .b(n39184), .c(n1821), .o(n43887) );
na02f01 g40096 ( .a(n761), .b(n8066), .o(n43888) );
na02f01 g40097 ( .a(n43888), .b(n43887), .o(n2746) );
no02f01 g40098 ( .a(n38042), .b(n37942), .o(n43890) );
oa12f01 g40099 ( .a(n43890), .b(n38001), .c(n37994), .o(n43891) );
in01f01 g40100 ( .a(n43890), .o(n43892) );
na03f01 g40101 ( .a(n38000), .b(n37995), .c(n43892), .o(n43893) );
na02f01 g40102 ( .a(n43893), .b(n43891), .o(n2751) );
no02f01 g40103 ( .a(n9487), .b(n9638), .o(n43895) );
no02f01 g40104 ( .a(n9503), .b(n9224), .o(n43896) );
na02f01 g40105 ( .a(n9503), .b(n9224), .o(n43897) );
in01f01 g40106 ( .a(n43897), .o(n43898) );
no02f01 g40107 ( .a(n43898), .b(n43896), .o(n43899) );
na02f01 g40108 ( .a(n43899), .b(n43895), .o(n43900) );
in01f01 g40109 ( .a(n43895), .o(n43901) );
in01f01 g40110 ( .a(n43899), .o(n43902) );
na02f01 g40111 ( .a(n43902), .b(n43901), .o(n43903) );
na02f01 g40112 ( .a(n43903), .b(n43900), .o(n2756) );
in01f01 g40113 ( .a(n41455), .o(n43905) );
no03f01 g40114 ( .a(n9607), .b(n9605), .c(n9234), .o(n43906) );
ao12f01 g40115 ( .a(n43906), .b(n43905), .c(n9225), .o(n43907) );
in01f01 g40116 ( .a(n43907), .o(n43908) );
oa12f01 g40117 ( .a(n39621), .b(n43908), .c(n37389), .o(n43909) );
in01f01 g40118 ( .a(n43909), .o(n43910) );
no02f01 g40119 ( .a(n43910), .b(n43228), .o(n43911) );
no02f01 g40120 ( .a(n43909), .b(n39631), .o(n43912) );
no02f01 g40121 ( .a(n43912), .b(n43911), .o(n43913) );
na03f01 g40122 ( .a(n43913), .b(n9590), .c(n9589), .o(n43914) );
in01f01 g40123 ( .a(n43913), .o(n4761) );
oa12f01 g40124 ( .a(n4761), .b(n9646), .c(n9645), .o(n43916) );
na02f01 g40125 ( .a(n43916), .b(n43914), .o(n2761) );
no03f01 g40126 ( .a(n41989), .b(n10988), .c(n10976), .o(n43918) );
in01f01 g40127 ( .a(n43918), .o(n43919) );
no02f01 g40128 ( .a(n41998), .b(n3521), .o(n43920) );
no02f01 g40129 ( .a(n41999), .b(n10735), .o(n43921) );
no02f01 g40130 ( .a(n43921), .b(n43920), .o(n43922) );
na03f01 g40131 ( .a(n43922), .b(n42012), .c(n43919), .o(n43923) );
in01f01 g40132 ( .a(n43922), .o(n43924) );
oa12f01 g40133 ( .a(n43924), .b(n42013), .c(n43918), .o(n43925) );
na02f01 g40134 ( .a(n43925), .b(n43923), .o(n2766) );
ao12f01 g40135 ( .a(n38208), .b(n38207), .c(n38196), .o(n43927) );
no03f01 g40136 ( .a(n38204), .b(n38199), .c(n38197), .o(n43928) );
oa12f01 g40137 ( .a(n21621), .b(n43928), .c(n43927), .o(n43929) );
na03f01 g40138 ( .a(n38209), .b(n38205), .c(delay_sub_ln23_0_unr27_stage10_stallmux_z), .o(n43930) );
na02f01 g40139 ( .a(n43930), .b(n43929), .o(n2771) );
na03f01 g40140 ( .a(n40370), .b(n9590), .c(n9589), .o(n43932) );
oa12f01 g40141 ( .a(n1021), .b(n9646), .c(n9645), .o(n43933) );
na02f01 g40142 ( .a(n43933), .b(n43932), .o(n2776) );
na02f01 g40143 ( .a(n43625), .b(n43622), .o(n2786) );
in01f01 g40144 ( .a(n32173), .o(n43936) );
no02f01 g40145 ( .a(n32485), .b(n32192), .o(n43937) );
in01f01 g40146 ( .a(n43937), .o(n43938) );
ao12f01 g40147 ( .a(n32399), .b(n43938), .c(n43936), .o(n43939) );
in01f01 g40148 ( .a(n43939), .o(n43940) );
no02f01 g40149 ( .a(n32163), .b(n32396), .o(n43941) );
na02f01 g40150 ( .a(n43941), .b(n43940), .o(n43942) );
in01f01 g40151 ( .a(n43941), .o(n43943) );
na02f01 g40152 ( .a(n43943), .b(n43939), .o(n43944) );
na02f01 g40153 ( .a(n43944), .b(n43942), .o(n2796) );
no02f01 g40154 ( .a(n21471), .b(n16329), .o(n43946) );
no02f01 g40155 ( .a(n43946), .b(n21473), .o(n43947) );
na03f01 g40156 ( .a(n43947), .b(n21582), .c(n21428), .o(n43948) );
in01f01 g40157 ( .a(n21582), .o(n43949) );
in01f01 g40158 ( .a(n43947), .o(n43950) );
oa12f01 g40159 ( .a(n43950), .b(n43949), .c(n21615), .o(n43951) );
na02f01 g40160 ( .a(n43951), .b(n43948), .o(n2801) );
no02f01 g40161 ( .a(n35461), .b(n4176), .o(n43953) );
no02f01 g40162 ( .a(n43953), .b(n35463), .o(n43954) );
na02f01 g40163 ( .a(n43954), .b(n42338), .o(n43955) );
in01f01 g40164 ( .a(n43954), .o(n43956) );
na02f01 g40165 ( .a(n43956), .b(n35441), .o(n43957) );
na02f01 g40166 ( .a(n43957), .b(n43955), .o(n2806) );
na02f01 g40167 ( .a(n42691), .b(n1821), .o(n43959) );
na02f01 g40168 ( .a(n1983), .b(n8066), .o(n43960) );
na02f01 g40169 ( .a(n43960), .b(n43959), .o(n2811) );
na03f01 g40170 ( .a(n25465), .b(n36642), .c(n36629), .o(n43962) );
oa12f01 g40171 ( .a(n25464), .b(n36646), .c(n25391), .o(n43963) );
na02f01 g40172 ( .a(n43963), .b(n43962), .o(n2816) );
na02f01 g40173 ( .a(n2267), .b(n4116), .o(n43965) );
na02f01 g40174 ( .a(n43208), .b(n2589), .o(n43966) );
na02f01 g40175 ( .a(n43966), .b(n43965), .o(n2821) );
no02f01 g40176 ( .a(n6002), .b(n5983_1), .o(n43968) );
no02f01 g40177 ( .a(n41898), .b(n6005), .o(n43969) );
in01f01 g40178 ( .a(n43969), .o(n43970) );
ao12f01 g40179 ( .a(n43970), .b(n43968), .c(n38635), .o(n43971) );
no02f01 g40180 ( .a(n5991), .b(n5873), .o(n43972) );
no02f01 g40181 ( .a(n43972), .b(n5993_1), .o(n43973) );
na02f01 g40182 ( .a(n43973), .b(n43971), .o(n43974) );
in01f01 g40183 ( .a(n43971), .o(n43975) );
in01f01 g40184 ( .a(n43973), .o(n43976) );
na02f01 g40185 ( .a(n43976), .b(n43975), .o(n43977) );
na02f01 g40186 ( .a(n43977), .b(n43974), .o(n2826) );
no02f01 g40187 ( .a(n20931), .b(n21324), .o(n43979) );
in01f01 g40188 ( .a(n43979), .o(n43980) );
no02f01 g40189 ( .a(n43980), .b(n39214), .o(n43981) );
no02f01 g40190 ( .a(n43979), .b(n39209), .o(n43982) );
no02f01 g40191 ( .a(n43982), .b(n43981), .o(n43983) );
in01f01 g40192 ( .a(n43983), .o(n2831) );
no02f01 g40193 ( .a(n39860), .b(n40571), .o(n43985) );
no02f01 g40194 ( .a(n43985), .b(n40573), .o(n43986) );
no03f01 g40195 ( .a(n39995), .b(n40049), .c(n39863), .o(n43987) );
oa12f01 g40196 ( .a(n43986), .b(n43987), .c(n39862), .o(n43988) );
in01f01 g40197 ( .a(n39862), .o(n43989) );
in01f01 g40198 ( .a(n43986), .o(n43990) );
in01f01 g40199 ( .a(n39863), .o(n43991) );
na03f01 g40200 ( .a(n39996), .b(n39983), .c(n43991), .o(n43992) );
na03f01 g40201 ( .a(n43992), .b(n43990), .c(n43989), .o(n43993) );
na03f01 g40202 ( .a(n43993), .b(n43988), .c(n_27923), .o(n43994) );
ao12f01 g40203 ( .a(n43990), .b(n43992), .c(n43989), .o(n43995) );
no03f01 g40204 ( .a(n43987), .b(n43986), .c(n39862), .o(n43996) );
oa12f01 g40205 ( .a(n34420), .b(n43996), .c(n43995), .o(n43997) );
na02f01 g40206 ( .a(n43997), .b(n43994), .o(n2836) );
no02f01 g40207 ( .a(n27664), .b(n27663), .o(n43999) );
in01f01 g40208 ( .a(n43999), .o(n44000) );
na02f01 g40209 ( .a(n27396), .b(n27395), .o(n44001) );
ao12f01 g40210 ( .a(n27397), .b(n44001), .c(n44000), .o(n44002) );
no02f01 g40211 ( .a(n27388), .b(n27367), .o(n44003) );
no02f01 g40212 ( .a(n44003), .b(n27399), .o(n44004) );
in01f01 g40213 ( .a(n44004), .o(n44005) );
na02f01 g40214 ( .a(n44005), .b(n44002), .o(n44006) );
in01f01 g40215 ( .a(n44002), .o(n44007) );
na02f01 g40216 ( .a(n44004), .b(n44007), .o(n44008) );
na02f01 g40217 ( .a(n44008), .b(n44006), .o(n2841) );
na02f01 g40218 ( .a(n43851), .b(n43847), .o(n2846) );
no02f01 g40219 ( .a(n38111), .b(n6037), .o(n44011) );
in01f01 g40220 ( .a(n44011), .o(n44012) );
in01f01 g40221 ( .a(n38113), .o(n44013) );
in01f01 g40222 ( .a(n41664), .o(n44014) );
na02f01 g40223 ( .a(n44014), .b(n44013), .o(n44015) );
no02f01 g40224 ( .a(n38137), .b(n6037), .o(n44016) );
no02f01 g40225 ( .a(n44016), .b(n38119), .o(n44017) );
na03f01 g40226 ( .a(n44017), .b(n44015), .c(n44012), .o(n44018) );
oa12f01 g40227 ( .a(n44012), .b(n41664), .c(n38113), .o(n44019) );
in01f01 g40228 ( .a(n44017), .o(n44020) );
na02f01 g40229 ( .a(n44020), .b(n44019), .o(n44021) );
na02f01 g40230 ( .a(n44021), .b(n44018), .o(n2851) );
na03f01 g40231 ( .a(n37396), .b(n9590), .c(n9589), .o(n44023) );
oa12f01 g40232 ( .a(n554), .b(n9646), .c(n9645), .o(n44024) );
na02f01 g40233 ( .a(n44024), .b(n44023), .o(n2856) );
na02f01 g40234 ( .a(n40510), .b(n40505), .o(n2866) );
in01f01 g40235 ( .a(n10856), .o(n44027) );
no02f01 g40236 ( .a(n10858), .b(n44027), .o(n44028) );
ao12f01 g40237 ( .a(n10824), .b(n10862), .c(n44028), .o(n44029) );
no02f01 g40238 ( .a(n43474), .b(n10871), .o(n44030) );
na02f01 g40239 ( .a(n44030), .b(n44029), .o(n44031) );
in01f01 g40240 ( .a(n44029), .o(n44032) );
in01f01 g40241 ( .a(n44030), .o(n44033) );
na02f01 g40242 ( .a(n44033), .b(n44032), .o(n44034) );
na02f01 g40243 ( .a(n44034), .b(n44031), .o(n2871) );
in01f01 g40244 ( .a(n29939), .o(n44036) );
no02f01 g40245 ( .a(n29937), .b(n40055), .o(n44037) );
na02f01 g40246 ( .a(n29937), .b(n40055), .o(n44038) );
in01f01 g40247 ( .a(n44038), .o(n44039) );
no02f01 g40248 ( .a(n44039), .b(n44037), .o(n44040) );
in01f01 g40249 ( .a(n44040), .o(n44041) );
in01f01 g40250 ( .a(n29940), .o(n44042) );
na03f01 g40251 ( .a(n30047), .b(n30042), .c(n44042), .o(n44043) );
na03f01 g40252 ( .a(n44043), .b(n44041), .c(n44036), .o(n44044) );
no03f01 g40253 ( .a(n30046), .b(n30134), .c(n29940), .o(n44045) );
oa12f01 g40254 ( .a(n44040), .b(n44045), .c(n29939), .o(n44046) );
na03f01 g40255 ( .a(n44046), .b(n44044), .c(n6037), .o(n44047) );
no03f01 g40256 ( .a(n44045), .b(n44040), .c(n29939), .o(n44048) );
ao12f01 g40257 ( .a(n44041), .b(n44043), .c(n44036), .o(n44049) );
oa12f01 g40258 ( .a(n5873), .b(n44049), .c(n44048), .o(n44050) );
na02f01 g40259 ( .a(n44050), .b(n44047), .o(n2876) );
na02f01 g40260 ( .a(n39491), .b(n2589), .o(n44052) );
na02f01 g40261 ( .a(n785), .b(n4116), .o(n44053) );
na02f01 g40262 ( .a(n44053), .b(n44052), .o(n2881) );
na02f01 g40263 ( .a(n42518), .b(n8765), .o(n44055) );
na02f01 g40264 ( .a(n42517), .b(beta_31), .o(n44056) );
na03f01 g40265 ( .a(n44056), .b(n44055), .c(n42526), .o(n2886) );
in01f01 g40266 ( .a(n35558), .o(n44058) );
in01f01 g40267 ( .a(n35557), .o(n44059) );
na02f01 g40268 ( .a(n44059), .b(n35544), .o(n44060) );
no02f01 g40269 ( .a(n42872), .b(n4176), .o(n44061) );
no02f01 g40270 ( .a(n44061), .b(n42856), .o(n44062) );
na03f01 g40271 ( .a(n44062), .b(n44060), .c(n44058), .o(n44063) );
na02f01 g40272 ( .a(n44060), .b(n44058), .o(n44064) );
in01f01 g40273 ( .a(n44062), .o(n44065) );
na02f01 g40274 ( .a(n44065), .b(n44064), .o(n44066) );
na02f01 g40275 ( .a(n44066), .b(n44063), .o(n2891) );
oa12f01 g40276 ( .a(n9232), .b(n4201), .c(n9228), .o(n44068) );
na03f01 g40277 ( .a(n44068), .b(n9590), .c(n9589), .o(n44069) );
in01f01 g40278 ( .a(n44068), .o(n5774) );
oa12f01 g40279 ( .a(n5774), .b(n9646), .c(n9645), .o(n44071) );
na02f01 g40280 ( .a(n44071), .b(n44069), .o(n2896) );
na03f01 g40281 ( .a(n27355), .b(n27354), .c(n27652), .o(n44073) );
oa12f01 g40282 ( .a(n27655), .b(n27656), .c(n27345), .o(n44074) );
na02f01 g40283 ( .a(n44074), .b(n44073), .o(n2901) );
in01f01 g40284 ( .a(n40885), .o(n44076) );
oa12f01 g40285 ( .a(n44076), .b(n42059), .c(n42060), .o(n44077) );
na02f01 g40286 ( .a(n40857), .b(n40854), .o(n44078) );
na02f01 g40287 ( .a(n44078), .b(n44077), .o(n44079) );
no02f01 g40288 ( .a(n44078), .b(n44077), .o(n44080) );
in01f01 g40289 ( .a(n44080), .o(n44081) );
na02f01 g40290 ( .a(n44081), .b(n44079), .o(n2906) );
no02f01 g40291 ( .a(n29815), .b(n29756), .o(n44083) );
na02f01 g40292 ( .a(n44083), .b(n29813), .o(n44084) );
in01f01 g40293 ( .a(n29813), .o(n44085) );
oa12f01 g40294 ( .a(n44085), .b(n29815), .c(n29756), .o(n44086) );
na02f01 g40295 ( .a(n44086), .b(n44084), .o(n2911) );
no02f01 g40296 ( .a(n38637), .b(n6015), .o(n44088) );
na03f01 g40297 ( .a(n44088), .b(n6007_1), .c(n38636), .o(n44089) );
in01f01 g40298 ( .a(n44088), .o(n44090) );
na02f01 g40299 ( .a(n44090), .b(n6008), .o(n44091) );
na02f01 g40300 ( .a(n44091), .b(n44089), .o(n2916) );
na03f01 g40301 ( .a(n27228), .b(n27030), .c(n26969), .o(n44093) );
oa12f01 g40302 ( .a(n27227), .b(n27031), .c(n27202), .o(n44094) );
na02f01 g40303 ( .a(n44094), .b(n44093), .o(n2921) );
no02f01 g40304 ( .a(n39860), .b(n29010), .o(n44096) );
no02f01 g40305 ( .a(n39861), .b(n29019), .o(n44097) );
no02f01 g40306 ( .a(n44097), .b(n44096), .o(n44098) );
no03f01 g40307 ( .a(n40585), .b(n40576), .c(n40590), .o(n44099) );
oa12f01 g40308 ( .a(n44099), .b(n40327), .c(n40326), .o(n44100) );
ao12f01 g40309 ( .a(n39860), .b(n40568), .c(n28833), .o(n44101) );
no03f01 g40310 ( .a(n44101), .b(n40579), .c(n39985), .o(n44102) );
na03f01 g40311 ( .a(n44102), .b(n44100), .c(n44098), .o(n44103) );
in01f01 g40312 ( .a(n44098), .o(n44104) );
in01f01 g40313 ( .a(n44099), .o(n44105) );
ao12f01 g40314 ( .a(n44105), .b(n39994), .c(n40321), .o(n44106) );
in01f01 g40315 ( .a(n44102), .o(n44107) );
oa12f01 g40316 ( .a(n44104), .b(n44107), .c(n44106), .o(n44108) );
na03f01 g40317 ( .a(n44108), .b(n44103), .c(n_27923), .o(n44109) );
no03f01 g40318 ( .a(n44107), .b(n44106), .c(n44104), .o(n44110) );
ao12f01 g40319 ( .a(n44098), .b(n44102), .c(n44100), .o(n44111) );
oa12f01 g40320 ( .a(n34420), .b(n44111), .c(n44110), .o(n44112) );
na02f01 g40321 ( .a(n44112), .b(n44109), .o(n2926) );
no02f01 g40322 ( .a(n40522), .b(n6934), .o(n44114) );
no02f01 g40323 ( .a(n9659), .b(n5001), .o(n44115) );
no02f01 g40324 ( .a(n44115), .b(n44114), .o(n44116) );
na03f01 g40325 ( .a(n44116), .b(n9899), .c(n40523), .o(n44117) );
in01f01 g40326 ( .a(n44116), .o(n44118) );
oa12f01 g40327 ( .a(n44118), .b(n9900), .c(n9894), .o(n44119) );
na02f01 g40328 ( .a(n44119), .b(n44117), .o(n2931) );
no03f01 g40329 ( .a(n21174), .b(n21173), .c(n21170), .o(n44121) );
no02f01 g40330 ( .a(n21175), .b(n21171), .o(n44122) );
oa12f01 g40331 ( .a(n21163), .b(n44122), .c(n44121), .o(n44123) );
in01f01 g40332 ( .a(n21163), .o(n44124) );
no02f01 g40333 ( .a(n44122), .b(n44121), .o(n44125) );
na02f01 g40334 ( .a(n44125), .b(n44124), .o(n44126) );
na02f01 g40335 ( .a(n44126), .b(n44123), .o(n2936) );
in01f01 g40336 ( .a(n21243), .o(n44128) );
ao12f01 g40337 ( .a(n21254), .b(n21257), .c(n44128), .o(n44129) );
in01f01 g40338 ( .a(n21256), .o(n44130) );
no02f01 g40339 ( .a(n44130), .b(n21026), .o(n44131) );
in01f01 g40340 ( .a(n44131), .o(n44132) );
no02f01 g40341 ( .a(n44132), .b(n44129), .o(n44133) );
na02f01 g40342 ( .a(n44132), .b(n44129), .o(n44134) );
in01f01 g40343 ( .a(n44134), .o(n44135) );
no02f01 g40344 ( .a(n44135), .b(n44133), .o(n44136) );
in01f01 g40345 ( .a(n44136), .o(n2941) );
in01f01 g40346 ( .a(n27640), .o(n44138) );
na02f01 g40347 ( .a(n44138), .b(n27676), .o(n44139) );
no02f01 g40348 ( .a(n27639), .b(n27677), .o(n44140) );
no02f01 g40349 ( .a(n27367), .b(n38193), .o(n44141) );
no02f01 g40350 ( .a(n44141), .b(n38195), .o(n44142) );
na03f01 g40351 ( .a(n44142), .b(n44140), .c(n44139), .o(n44143) );
no02f01 g40352 ( .a(n27640), .b(n27624), .o(n44144) );
in01f01 g40353 ( .a(n44140), .o(n44145) );
in01f01 g40354 ( .a(n44142), .o(n44146) );
oa12f01 g40355 ( .a(n44146), .b(n44145), .c(n44144), .o(n44147) );
na03f01 g40356 ( .a(n44147), .b(n44143), .c(delay_sub_ln23_0_unr27_stage10_stallmux_z), .o(n44148) );
no03f01 g40357 ( .a(n44146), .b(n44145), .c(n44144), .o(n44149) );
ao12f01 g40358 ( .a(n44142), .b(n44140), .c(n44139), .o(n44150) );
oa12f01 g40359 ( .a(n21621), .b(n44150), .c(n44149), .o(n44151) );
na02f01 g40360 ( .a(n44151), .b(n44148), .o(n2946) );
no02f01 g40361 ( .a(n29425), .b(n29213), .o(n44153) );
in01f01 g40362 ( .a(n29532), .o(n44154) );
ao12f01 g40363 ( .a(n44154), .b(n29717), .c(n44153), .o(n44155) );
no02f01 g40364 ( .a(n29507), .b(n29430), .o(n44156) );
no02f01 g40365 ( .a(n29506), .b(n29639), .o(n44157) );
no02f01 g40366 ( .a(n44157), .b(n44156), .o(n44158) );
na02f01 g40367 ( .a(n44158), .b(n44155), .o(n44159) );
in01f01 g40368 ( .a(n44155), .o(n44160) );
in01f01 g40369 ( .a(n44158), .o(n44161) );
na02f01 g40370 ( .a(n44161), .b(n44160), .o(n44162) );
na02f01 g40371 ( .a(n44162), .b(n44159), .o(n2951) );
no02f01 g40372 ( .a(n21608), .b(n21576), .o(n44164) );
in01f01 g40373 ( .a(n44164), .o(n44165) );
no02f01 g40374 ( .a(n27300), .b(n16155), .o(n44166) );
no02f01 g40375 ( .a(n44166), .b(n44165), .o(n44167) );
in01f01 g40376 ( .a(n44167), .o(n44168) );
no04f01 g40377 ( .a(n44168), .b(n21559), .c(n21475), .d(n21428), .o(n44169) );
ao12f01 g40378 ( .a(n16329), .b(n21606), .c(n21595), .o(n44170) );
in01f01 g40379 ( .a(n44170), .o(n44171) );
ao12f01 g40380 ( .a(n16329), .b(n44171), .c(n27291), .o(n44172) );
in01f01 g40381 ( .a(n44172), .o(n44173) );
na02f01 g40382 ( .a(n44173), .b(n21593), .o(n44174) );
no02f01 g40383 ( .a(n27275), .b(n16329), .o(n44175) );
in01f01 g40384 ( .a(n27275), .o(n44176) );
no02f01 g40385 ( .a(n44176), .b(n16155), .o(n44177) );
no02f01 g40386 ( .a(n44177), .b(n44175), .o(n44178) );
in01f01 g40387 ( .a(n44178), .o(n44179) );
oa12f01 g40388 ( .a(n44179), .b(n44174), .c(n44169), .o(n44180) );
na04f01 g40389 ( .a(n44167), .b(n21558), .c(n21474), .d(n21615), .o(n44181) );
in01f01 g40390 ( .a(n44174), .o(n44182) );
na03f01 g40391 ( .a(n44178), .b(n44182), .c(n44181), .o(n44183) );
na03f01 g40392 ( .a(n44183), .b(n44180), .c(delay_sub_ln23_0_unr27_stage10_stallmux_z), .o(n44184) );
ao12f01 g40393 ( .a(n44178), .b(n44182), .c(n44181), .o(n44185) );
no03f01 g40394 ( .a(n44179), .b(n44174), .c(n44169), .o(n44186) );
oa12f01 g40395 ( .a(n21621), .b(n44186), .c(n44185), .o(n44187) );
na02f01 g40396 ( .a(n44187), .b(n44184), .o(n2956) );
in01f01 g40397 ( .a(n34412), .o(n44189) );
na02f01 g40398 ( .a(n34413), .b(n6050), .o(n44190) );
no02f01 g40399 ( .a(n5895), .b(n5873), .o(n44191) );
no02f01 g40400 ( .a(n44191), .b(n38088), .o(n44192) );
na03f01 g40401 ( .a(n44192), .b(n44190), .c(n44189), .o(n44193) );
na02f01 g40402 ( .a(n44190), .b(n44189), .o(n44194) );
in01f01 g40403 ( .a(n44192), .o(n44195) );
na02f01 g40404 ( .a(n44195), .b(n44194), .o(n44196) );
na02f01 g40405 ( .a(n44196), .b(n44193), .o(n2961) );
in01f01 g40406 ( .a(n9234), .o(n44198) );
ao12f01 g40407 ( .a(n9233), .b(n39834), .c(n44198), .o(n44199) );
no02f01 g40408 ( .a(n44199), .b(n40599), .o(n44200) );
na02f01 g40409 ( .a(n44199), .b(n40599), .o(n44201) );
in01f01 g40410 ( .a(n44201), .o(n44202) );
no02f01 g40411 ( .a(n44202), .b(n44200), .o(n44203) );
na03f01 g40412 ( .a(n44203), .b(n9590), .c(n9589), .o(n44204) );
in01f01 g40413 ( .a(n44203), .o(n3466) );
oa12f01 g40414 ( .a(n3466), .b(n9646), .c(n9645), .o(n44206) );
na02f01 g40415 ( .a(n44206), .b(n44204), .o(n2966) );
na03f01 g40416 ( .a(n38407), .b(n39112), .c(n38350), .o(n44208) );
oa12f01 g40417 ( .a(n38406), .b(n38408), .c(n38349), .o(n44209) );
na02f01 g40418 ( .a(n44209), .b(n44208), .o(n2971) );
no02f01 g40419 ( .a(n39137), .b(n39075), .o(n44211) );
no02f01 g40420 ( .a(n39064), .b(n39135), .o(n44212) );
no02f01 g40421 ( .a(n39065), .b(n39059), .o(n44213) );
no02f01 g40422 ( .a(n44213), .b(n44212), .o(n44214) );
in01f01 g40423 ( .a(n44214), .o(n44215) );
na02f01 g40424 ( .a(n44215), .b(n44211), .o(n44216) );
na02f01 g40425 ( .a(n44214), .b(n43294), .o(n44217) );
na02f01 g40426 ( .a(n44217), .b(n44216), .o(n2976) );
in01f01 g40427 ( .a(n21211), .o(n44219) );
no02f01 g40428 ( .a(n21212), .b(n21049), .o(n44220) );
in01f01 g40429 ( .a(n44220), .o(n44221) );
no02f01 g40430 ( .a(n44221), .b(n44219), .o(n44222) );
no02f01 g40431 ( .a(n44220), .b(n21211), .o(n44223) );
no02f01 g40432 ( .a(n44223), .b(n44222), .o(n44224) );
na02f01 g40433 ( .a(n44224), .b(n5799), .o(n44225) );
in01f01 g40434 ( .a(n44224), .o(n5420) );
na02f01 g40435 ( .a(n5420), .b(n911), .o(n44227) );
na02f01 g40436 ( .a(n44227), .b(n44225), .o(n2981) );
na02f01 g40437 ( .a(n42297), .b(n42296), .o(n2986) );
oa12f01 g40438 ( .a(n38166), .b(n43513), .c(n9596), .o(n44230) );
in01f01 g40439 ( .a(n44230), .o(n44231) );
no02f01 g40440 ( .a(n44231), .b(n41456), .o(n44232) );
no02f01 g40441 ( .a(n44230), .b(n41457), .o(n44233) );
no02f01 g40442 ( .a(n44233), .b(n44232), .o(n44234) );
na03f01 g40443 ( .a(n44234), .b(n9590), .c(n9589), .o(n44235) );
in01f01 g40444 ( .a(n44234), .o(n5628) );
oa12f01 g40445 ( .a(n5628), .b(n9646), .c(n9645), .o(n44237) );
na02f01 g40446 ( .a(n44237), .b(n44235), .o(n2991) );
in01f01 g40447 ( .a(n41195), .o(n44239) );
no02f01 g40448 ( .a(n40791), .b(n20334), .o(n44240) );
no02f01 g40449 ( .a(n44240), .b(n41206), .o(n44241) );
na02f01 g40450 ( .a(n41189), .b(n40950), .o(n44242) );
na03f01 g40451 ( .a(n44242), .b(n44241), .c(n44239), .o(n44243) );
in01f01 g40452 ( .a(n44241), .o(n44244) );
oa12f01 g40453 ( .a(n44239), .b(n41205), .c(n40936), .o(n44245) );
na02f01 g40454 ( .a(n44245), .b(n44244), .o(n44246) );
na02f01 g40455 ( .a(n44246), .b(n44243), .o(n2996) );
na02f01 g40456 ( .a(n32732), .b(cos_out_11), .o(n44248) );
no02f01 g40457 ( .a(n36292), .b(n36269), .o(n44249) );
in01f01 g40458 ( .a(n44249), .o(n44250) );
no02f01 g40459 ( .a(n44250), .b(n36313), .o(n44251) );
no02f01 g40460 ( .a(n36311), .b(n35944), .o(n44252) );
in01f01 g40461 ( .a(n44252), .o(n44253) );
in01f01 g40462 ( .a(n36367), .o(n44254) );
na02f01 g40463 ( .a(n44254), .b(n44253), .o(n44255) );
no02f01 g40464 ( .a(n36302), .b(n35944), .o(n44256) );
no02f01 g40465 ( .a(n44256), .b(n36304), .o(n44257) );
in01f01 g40466 ( .a(n44257), .o(n44258) );
no03f01 g40467 ( .a(n44258), .b(n44255), .c(n44251), .o(n44259) );
no02f01 g40468 ( .a(n44255), .b(n44251), .o(n44260) );
no02f01 g40469 ( .a(n44257), .b(n44260), .o(n44261) );
oa12f01 g40470 ( .a(n32734), .b(n44261), .c(n44259), .o(n44262) );
na02f01 g40471 ( .a(n44262), .b(n44248), .o(n3001) );
na02f01 g40472 ( .a(n43983), .b(n5799), .o(n44264) );
na02f01 g40473 ( .a(n2831), .b(n911), .o(n44265) );
na02f01 g40474 ( .a(n44265), .b(n44264), .o(n3005) );
no02f01 g40475 ( .a(n21319), .b(n20904), .o(n44267) );
no02f01 g40476 ( .a(n39210), .b(n21324), .o(n44268) );
na02f01 g40477 ( .a(n44268), .b(n44267), .o(n44269) );
in01f01 g40478 ( .a(n44267), .o(n44270) );
oa12f01 g40479 ( .a(n44270), .b(n39210), .c(n21324), .o(n44271) );
na02f01 g40480 ( .a(n44271), .b(n44269), .o(n3010) );
na03f01 g40481 ( .a(n38871), .b(n38869), .c(n1821), .o(n44273) );
na02f01 g40482 ( .a(n688), .b(n8066), .o(n44274) );
na02f01 g40483 ( .a(n44274), .b(n44273), .o(n3015) );
na03f01 g40484 ( .a(n4991), .b(n4947_1), .c(n4981), .o(n44276) );
oa12f01 g40485 ( .a(n4968), .b(n4982_1), .c(n4946), .o(n44277) );
na02f01 g40486 ( .a(n44277), .b(n44276), .o(n3025) );
no02f01 g40487 ( .a(n11758), .b(n11734), .o(n44279) );
na02f01 g40488 ( .a(n44279), .b(n38076), .o(n44280) );
in01f01 g40489 ( .a(n44279), .o(n44281) );
na03f01 g40490 ( .a(n44281), .b(n11717), .c(n11716), .o(n44282) );
na02f01 g40491 ( .a(n44282), .b(n44280), .o(n3030) );
no02f01 g40492 ( .a(n38167), .b(n9598), .o(n44284) );
no02f01 g40493 ( .a(n44284), .b(n41456), .o(n44285) );
na02f01 g40494 ( .a(n44284), .b(n41456), .o(n44286) );
in01f01 g40495 ( .a(n44286), .o(n44287) );
no02f01 g40496 ( .a(n44287), .b(n44285), .o(n44288) );
na03f01 g40497 ( .a(n44288), .b(n9590), .c(n9589), .o(n44289) );
in01f01 g40498 ( .a(n44288), .o(n3456) );
oa12f01 g40499 ( .a(n3456), .b(n9646), .c(n9645), .o(n44291) );
na02f01 g40500 ( .a(n44291), .b(n44289), .o(n3035) );
no03f01 g40501 ( .a(n42887), .b(n42877), .c(n42876), .o(n44293) );
ao12f01 g40502 ( .a(n4176), .b(n42888), .c(n42833), .o(n44294) );
no02f01 g40503 ( .a(n44294), .b(n42875), .o(n44295) );
in01f01 g40504 ( .a(n44295), .o(n44296) );
ao12f01 g40505 ( .a(n44296), .b(n44293), .c(n42869), .o(n3040) );
na02f01 g40506 ( .a(n39540), .b(n5799), .o(n44298) );
na02f01 g40507 ( .a(n799), .b(n911), .o(n44299) );
na02f01 g40508 ( .a(n44299), .b(n44298), .o(n3045) );
no02f01 g40509 ( .a(n22267), .b(n22266), .o(n44301) );
no02f01 g40510 ( .a(n22270), .b(n22142), .o(n44302) );
in01f01 g40511 ( .a(n44302), .o(n44303) );
no02f01 g40512 ( .a(n44303), .b(n44301), .o(n44304) );
na02f01 g40513 ( .a(n44303), .b(n44301), .o(n44305) );
in01f01 g40514 ( .a(n44305), .o(n44306) );
no02f01 g40515 ( .a(n44306), .b(n44304), .o(n44307) );
in01f01 g40516 ( .a(n44307), .o(n3050) );
na03f01 g40517 ( .a(n29406), .b(n29404), .c(n29701), .o(n44309) );
oa12f01 g40518 ( .a(n29390), .b(n29706), .c(n29403), .o(n44310) );
na02f01 g40519 ( .a(n44310), .b(n44309), .o(n3060) );
na02f01 g40520 ( .a(n21376), .b(n16489), .o(n44312) );
in01f01 g40521 ( .a(n44312), .o(n44313) );
in01f01 g40522 ( .a(n21403), .o(n44314) );
na02f01 g40523 ( .a(n44314), .b(n44313), .o(n44315) );
no02f01 g40524 ( .a(n21401), .b(n16329), .o(n44316) );
no02f01 g40525 ( .a(n44316), .b(n21580), .o(n44317) );
no02f01 g40526 ( .a(n21424), .b(n16329), .o(n44318) );
no02f01 g40527 ( .a(n44318), .b(n21426), .o(n44319) );
na03f01 g40528 ( .a(n44319), .b(n44317), .c(n44315), .o(n44320) );
na02f01 g40529 ( .a(n44317), .b(n44315), .o(n44321) );
in01f01 g40530 ( .a(n44319), .o(n44322) );
na02f01 g40531 ( .a(n44322), .b(n44321), .o(n44323) );
na02f01 g40532 ( .a(n44323), .b(n44320), .o(n3070) );
no02f01 g40533 ( .a(n29379), .b(n29364), .o(n44325) );
no02f01 g40534 ( .a(n29380), .b(n29688), .o(n44326) );
oa12f01 g40535 ( .a(n29372), .b(n44326), .c(n44325), .o(n44327) );
in01f01 g40536 ( .a(n29372), .o(n44328) );
no02f01 g40537 ( .a(n44326), .b(n44325), .o(n44329) );
na02f01 g40538 ( .a(n44329), .b(n44328), .o(n44330) );
na02f01 g40539 ( .a(n44330), .b(n44327), .o(n3075) );
in01f01 g40540 ( .a(n29806), .o(n44332) );
na02f01 g40541 ( .a(n44332), .b(n29802), .o(n44333) );
na03f01 g40542 ( .a(n29806), .b(n29801), .c(n29799), .o(n44334) );
na02f01 g40543 ( .a(n44334), .b(n44333), .o(n3080) );
no02f01 g40544 ( .a(n39135), .b(n31401), .o(n44336) );
no02f01 g40545 ( .a(n44336), .b(n39145), .o(n44337) );
in01f01 g40546 ( .a(n39156), .o(n44338) );
no02f01 g40547 ( .a(n44338), .b(n39142), .o(n44339) );
na02f01 g40548 ( .a(n44339), .b(n44337), .o(n44340) );
in01f01 g40549 ( .a(n44337), .o(n44341) );
oa12f01 g40550 ( .a(n44341), .b(n44338), .c(n39142), .o(n44342) );
na03f01 g40551 ( .a(n44342), .b(n44340), .c(n3633), .o(n44343) );
na02f01 g40552 ( .a(n44342), .b(n44340), .o(n6017) );
na02f01 g40553 ( .a(n6017), .b(n6203), .o(n44345) );
na02f01 g40554 ( .a(n44345), .b(n44343), .o(n3085) );
no02f01 g40555 ( .a(n10823), .b(n3521), .o(n44347) );
no02f01 g40556 ( .a(n44347), .b(n10858), .o(n44348) );
in01f01 g40557 ( .a(n44348), .o(n44349) );
na02f01 g40558 ( .a(n44349), .b(n10856), .o(n44350) );
na02f01 g40559 ( .a(n44348), .b(n44027), .o(n44351) );
na02f01 g40560 ( .a(n44351), .b(n44350), .o(n3090) );
na03f01 g40561 ( .a(n40050), .b(n39997), .c(n_27923), .o(n44353) );
na02f01 g40562 ( .a(n926), .b(n34420), .o(n44354) );
na02f01 g40563 ( .a(n44354), .b(n44353), .o(n3095) );
no02f01 g40564 ( .a(n42805), .b(n11662), .o(n44356) );
na02f01 g40565 ( .a(n44356), .b(n42803), .o(n44357) );
in01f01 g40566 ( .a(n44356), .o(n44358) );
na02f01 g40567 ( .a(n44358), .b(n42804), .o(n44359) );
na02f01 g40568 ( .a(n44359), .b(n44357), .o(n3100) );
in01f01 g40569 ( .a(n40792), .o(n44361) );
in01f01 g40570 ( .a(n40795), .o(n44362) );
na02f01 g40571 ( .a(n40950), .b(n44362), .o(n44363) );
no02f01 g40572 ( .a(n40791), .b(n20424), .o(n44364) );
no02f01 g40573 ( .a(n40794), .b(n20337), .o(n44365) );
no02f01 g40574 ( .a(n44365), .b(n44364), .o(n44366) );
na03f01 g40575 ( .a(n44366), .b(n44363), .c(n44361), .o(n44367) );
oa12f01 g40576 ( .a(n44361), .b(n40936), .c(n40795), .o(n44368) );
in01f01 g40577 ( .a(n44366), .o(n44369) );
na02f01 g40578 ( .a(n44369), .b(n44368), .o(n44370) );
na03f01 g40579 ( .a(n44370), .b(n44367), .c(n5799), .o(n44371) );
na02f01 g40580 ( .a(n44370), .b(n44367), .o(n3673) );
na02f01 g40581 ( .a(n3673), .b(n911), .o(n44373) );
na02f01 g40582 ( .a(n44373), .b(n44371), .o(n3105) );
ao12f01 g40583 ( .a(n9233), .b(n39624), .c(n44198), .o(n44375) );
in01f01 g40584 ( .a(n44375), .o(n44376) );
no02f01 g40585 ( .a(n44376), .b(n9228), .o(n44377) );
no02f01 g40586 ( .a(n44375), .b(n936), .o(n44378) );
no02f01 g40587 ( .a(n44378), .b(n44377), .o(n44379) );
na03f01 g40588 ( .a(n44379), .b(n9590), .c(n9589), .o(n44380) );
in01f01 g40589 ( .a(n44379), .o(n3855) );
oa12f01 g40590 ( .a(n3855), .b(n9646), .c(n9645), .o(n44382) );
na02f01 g40591 ( .a(n44382), .b(n44380), .o(n3110) );
no02f01 g40592 ( .a(n29481), .b(n29639), .o(n44384) );
no02f01 g40593 ( .a(n29482), .b(n29430), .o(n44385) );
in01f01 g40594 ( .a(n44385), .o(n44386) );
ao12f01 g40595 ( .a(n44384), .b(n44386), .c(n44153), .o(n44387) );
no02f01 g40596 ( .a(n29476), .b(n29430), .o(n44388) );
no02f01 g40597 ( .a(n29475), .b(n29639), .o(n44389) );
no02f01 g40598 ( .a(n44389), .b(n44388), .o(n44390) );
na02f01 g40599 ( .a(n44390), .b(n44387), .o(n44391) );
in01f01 g40600 ( .a(n44387), .o(n44392) );
in01f01 g40601 ( .a(n44390), .o(n44393) );
na02f01 g40602 ( .a(n44393), .b(n44392), .o(n44394) );
na02f01 g40603 ( .a(n44394), .b(n44391), .o(n3115) );
no02f01 g40604 ( .a(n44316), .b(n21403), .o(n44396) );
na03f01 g40605 ( .a(n44396), .b(n21579), .c(n44312), .o(n44397) );
in01f01 g40606 ( .a(n44396), .o(n44398) );
oa12f01 g40607 ( .a(n44398), .b(n21580), .c(n44313), .o(n44399) );
na02f01 g40608 ( .a(n44399), .b(n44397), .o(n3125) );
na02f01 g40609 ( .a(n5988), .b(n37149), .o(n44401) );
na02f01 g40610 ( .a(n44401), .b(n37312), .o(n3130) );
na03f01 g40611 ( .a(n29389), .b(n29388), .c(n29676), .o(n44403) );
oa12f01 g40612 ( .a(n29699), .b(n29700), .c(n29337), .o(n44404) );
na02f01 g40613 ( .a(n44404), .b(n44403), .o(n3135) );
na03f01 g40614 ( .a(n39811), .b(n39807), .c(delay_sub_ln23_0_unr27_stage10_stallmux_z), .o(n44406) );
no03f01 g40615 ( .a(n39810), .b(n39809), .c(n39808), .o(n44407) );
ao12f01 g40616 ( .a(n39802), .b(n39806), .c(n39804), .o(n44408) );
oa12f01 g40617 ( .a(n21621), .b(n44408), .c(n44407), .o(n44409) );
na02f01 g40618 ( .a(n44409), .b(n44406), .o(n3140) );
no02f01 g40619 ( .a(n42908), .b(n42911), .o(n44411) );
na03f01 g40620 ( .a(n44411), .b(n42913), .c(n42910), .o(n44412) );
in01f01 g40621 ( .a(n44411), .o(n44413) );
oa12f01 g40622 ( .a(n44413), .b(n42917), .c(n39992), .o(n44414) );
na03f01 g40623 ( .a(n44414), .b(n44412), .c(n_27923), .o(n44415) );
na02f01 g40624 ( .a(n44414), .b(n44412), .o(n3841) );
na02f01 g40625 ( .a(n3841), .b(n34420), .o(n44417) );
na02f01 g40626 ( .a(n44417), .b(n44415), .o(n3145) );
no03f01 g40627 ( .a(n30125), .b(n30016), .c(n29961), .o(n44419) );
ao12f01 g40628 ( .a(n30124), .b(n30018), .c(n29960), .o(n44420) );
no02f01 g40629 ( .a(n44420), .b(n44419), .o(n44421) );
in01f01 g40630 ( .a(n44421), .o(n3150) );
no02f01 g40631 ( .a(n22251), .b(n22155), .o(n44423) );
no02f01 g40632 ( .a(n22253), .b(n22148), .o(n44424) );
in01f01 g40633 ( .a(n44424), .o(n44425) );
no02f01 g40634 ( .a(n44425), .b(n44423), .o(n44426) );
na02f01 g40635 ( .a(n44425), .b(n44423), .o(n44427) );
in01f01 g40636 ( .a(n44427), .o(n44428) );
no02f01 g40637 ( .a(n44428), .b(n44426), .o(n44429) );
na02f01 g40638 ( .a(n44429), .b(n2589), .o(n44430) );
in01f01 g40639 ( .a(n44429), .o(n3277) );
na02f01 g40640 ( .a(n3277), .b(n4116), .o(n44432) );
na02f01 g40641 ( .a(n44432), .b(n44430), .o(n3155) );
in01f01 g40642 ( .a(n32416), .o(n44434) );
no02f01 g40643 ( .a(n44434), .b(n32414), .o(n44435) );
na02f01 g40644 ( .a(n44435), .b(n32489), .o(n44436) );
oa12f01 g40645 ( .a(n32402), .b(n44434), .c(n32414), .o(n44437) );
na02f01 g40646 ( .a(n44437), .b(n44436), .o(n3160) );
in01f01 g40647 ( .a(n22222), .o(n44439) );
na03f01 g40648 ( .a(n22231), .b(n22230), .c(n44439), .o(n44440) );
in01f01 g40649 ( .a(n22230), .o(n44441) );
in01f01 g40650 ( .a(n22231), .o(n44442) );
oa12f01 g40651 ( .a(n44441), .b(n44442), .c(n22222), .o(n44443) );
na02f01 g40652 ( .a(n44443), .b(n44440), .o(n3165) );
no02f01 g40653 ( .a(n36124), .b(n36057), .o(n44445) );
in01f01 g40654 ( .a(n44445), .o(n44446) );
no02f01 g40655 ( .a(n36132), .b(n36122), .o(n44447) );
no02f01 g40656 ( .a(n36133), .b(n36038), .o(n44448) );
no02f01 g40657 ( .a(n44448), .b(n44447), .o(n44449) );
na02f01 g40658 ( .a(n44449), .b(n44446), .o(n44450) );
in01f01 g40659 ( .a(n44449), .o(n44451) );
na02f01 g40660 ( .a(n44451), .b(n44445), .o(n44452) );
na02f01 g40661 ( .a(n44452), .b(n44450), .o(n3170) );
na02f01 g40662 ( .a(n37333), .b(n37331), .o(n3175) );
no02f01 g40663 ( .a(n9230), .b(n9229), .o(n44455) );
in01f01 g40664 ( .a(n44455), .o(n3180) );
no02f01 g40665 ( .a(n6946), .b(n6934), .o(n44457) );
no02f01 g40666 ( .a(n44457), .b(n6948), .o(n44458) );
na02f01 g40667 ( .a(n44458), .b(n6938), .o(n44459) );
in01f01 g40668 ( .a(n44458), .o(n44460) );
na02f01 g40669 ( .a(n44460), .b(n36532), .o(n44461) );
na02f01 g40670 ( .a(n44461), .b(n44459), .o(n3185) );
na02f01 g40671 ( .a(n32732), .b(sin_out_0), .o(n44463) );
ao12f01 g40672 ( .a(n34324), .b(n36558), .c(n36557), .o(n44464) );
no03f01 g40673 ( .a(n36559), .b(n34319), .c(n34318), .o(n44465) );
oa12f01 g40674 ( .a(n32734), .b(n44465), .c(n44464), .o(n44466) );
na02f01 g40675 ( .a(n44466), .b(n44463), .o(n3190) );
no02f01 g40676 ( .a(n22273), .b(n22133), .o(n44468) );
in01f01 g40677 ( .a(n44468), .o(n44469) );
no03f01 g40678 ( .a(n44469), .b(n22271), .c(n22142), .o(n44470) );
no02f01 g40679 ( .a(n22271), .b(n22142), .o(n44471) );
no02f01 g40680 ( .a(n44468), .b(n44471), .o(n44472) );
no02f01 g40681 ( .a(n44472), .b(n44470), .o(n44473) );
in01f01 g40682 ( .a(n44473), .o(n4727) );
na02f01 g40683 ( .a(n4727), .b(n4116), .o(n44475) );
na02f01 g40684 ( .a(n44473), .b(n2589), .o(n44476) );
na02f01 g40685 ( .a(n44476), .b(n44475), .o(n3194) );
no02f01 g40686 ( .a(n43608), .b(n35311), .o(n44478) );
in01f01 g40687 ( .a(n44478), .o(n44479) );
na02f01 g40688 ( .a(n44479), .b(n35302), .o(n44480) );
na02f01 g40689 ( .a(n44478), .b(n43606), .o(n44481) );
na02f01 g40690 ( .a(n44481), .b(n44480), .o(n3204) );
na02f01 g40691 ( .a(n43139), .b(n43136), .o(n3209) );
in01f01 g40692 ( .a(n41221), .o(n44484) );
no02f01 g40693 ( .a(n37871), .b(n26272), .o(n44485) );
no02f01 g40694 ( .a(n44485), .b(n41222), .o(n44486) );
in01f01 g40695 ( .a(n44486), .o(n44487) );
in01f01 g40696 ( .a(n41237), .o(n44488) );
no02f01 g40697 ( .a(n37871), .b(n26407), .o(n44489) );
in01f01 g40698 ( .a(n44489), .o(n44490) );
in01f01 g40699 ( .a(n41225), .o(n44491) );
oa12f01 g40700 ( .a(n44491), .b(n41247), .c(n41246), .o(n44492) );
na03f01 g40701 ( .a(n44492), .b(n44490), .c(n44488), .o(n44493) );
na03f01 g40702 ( .a(n44493), .b(n44487), .c(n44484), .o(n44494) );
ao12f01 g40703 ( .a(n41225), .b(n40990), .c(n40988), .o(n44495) );
no03f01 g40704 ( .a(n44495), .b(n44489), .c(n41237), .o(n44496) );
oa12f01 g40705 ( .a(n44486), .b(n44496), .c(n41221), .o(n44497) );
na03f01 g40706 ( .a(n44497), .b(n44494), .c(n1821), .o(n44498) );
no03f01 g40707 ( .a(n44496), .b(n44486), .c(n41221), .o(n44499) );
ao12f01 g40708 ( .a(n44487), .b(n44493), .c(n44484), .o(n44500) );
oa12f01 g40709 ( .a(n8066), .b(n44500), .c(n44499), .o(n44501) );
na02f01 g40710 ( .a(n44501), .b(n44498), .o(n3214) );
no02f01 g40711 ( .a(n36432), .b(n41680), .o(n44503) );
no02f01 g40712 ( .a(n44503), .b(n41682), .o(n44504) );
in01f01 g40713 ( .a(n44504), .o(n44505) );
in01f01 g40714 ( .a(n41684), .o(n44506) );
na03f01 g40715 ( .a(n43262), .b(n43261), .c(n44506), .o(n44507) );
ao12f01 g40716 ( .a(n44505), .b(n44507), .c(n41689), .o(n44508) );
no03f01 g40717 ( .a(n43268), .b(n43267), .c(n41684), .o(n44509) );
no03f01 g40718 ( .a(n44509), .b(n44504), .c(n41688), .o(n44510) );
oa12f01 g40719 ( .a(n4116), .b(n44510), .c(n44508), .o(n44511) );
oa12f01 g40720 ( .a(n44504), .b(n44509), .c(n41688), .o(n44512) );
na03f01 g40721 ( .a(n44507), .b(n44505), .c(n41689), .o(n44513) );
na03f01 g40722 ( .a(n44513), .b(n44512), .c(n2589), .o(n44514) );
na02f01 g40723 ( .a(n44514), .b(n44511), .o(n3219) );
na02f01 g40724 ( .a(n32732), .b(cos_out_23), .o(n44516) );
na03f01 g40725 ( .a(n41493), .b(n41498), .c(n39691), .o(n44517) );
no02f01 g40726 ( .a(n41492), .b(n41480), .o(n44518) );
na02f01 g40727 ( .a(n44518), .b(n44517), .o(n44519) );
no02f01 g40728 ( .a(n41626), .b(n35944), .o(n44520) );
no02f01 g40729 ( .a(n44520), .b(n41545), .o(n44521) );
in01f01 g40730 ( .a(n44521), .o(n44522) );
no02f01 g40731 ( .a(n44522), .b(n44519), .o(n44523) );
ao12f01 g40732 ( .a(n44521), .b(n44518), .c(n44517), .o(n44524) );
oa12f01 g40733 ( .a(n32734), .b(n44524), .c(n44523), .o(n44525) );
na02f01 g40734 ( .a(n44525), .b(n44516), .o(n3224) );
no02f01 g40735 ( .a(n25282), .b(n25250), .o(n44527) );
no02f01 g40736 ( .a(n44527), .b(n39017), .o(n44528) );
in01f01 g40737 ( .a(n44528), .o(n44529) );
na02f01 g40738 ( .a(n44527), .b(n39017), .o(n44530) );
na03f01 g40739 ( .a(n44530), .b(n44529), .c(n6037), .o(n44531) );
na02f01 g40740 ( .a(n44530), .b(n44529), .o(n5834) );
na02f01 g40741 ( .a(n5834), .b(n5873), .o(n44533) );
na02f01 g40742 ( .a(n44533), .b(n44531), .o(n3238) );
na02f01 g40743 ( .a(n38808), .b(n38803), .o(n3243) );
na02f01 g40744 ( .a(n32732), .b(sin_out_27), .o(n44536) );
no02f01 g40745 ( .a(n35886), .b(n35818), .o(n44537) );
oa12f01 g40746 ( .a(n44537), .b(n35847), .c(n35906), .o(n44538) );
ao12f01 g40747 ( .a(n35884), .b(n44538), .c(n35829), .o(n44539) );
no02f01 g40748 ( .a(n35887), .b(n35858), .o(n44540) );
no02f01 g40749 ( .a(n44540), .b(n44539), .o(n44541) );
na02f01 g40750 ( .a(n44540), .b(n44539), .o(n44542) );
in01f01 g40751 ( .a(n44542), .o(n44543) );
no03f01 g40752 ( .a(n44543), .b(n44541), .c(n34267), .o(n44544) );
no02f01 g40753 ( .a(n44543), .b(n44541), .o(n44545) );
no02f01 g40754 ( .a(n44545), .b(n34307), .o(n44546) );
no02f01 g40755 ( .a(n44546), .b(n44544), .o(n44547) );
no02f01 g40756 ( .a(n35884), .b(n35828), .o(n44548) );
in01f01 g40757 ( .a(n44548), .o(n44549) );
no02f01 g40758 ( .a(n44549), .b(n44538), .o(n44550) );
na02f01 g40759 ( .a(n44549), .b(n44538), .o(n44551) );
in01f01 g40760 ( .a(n44551), .o(n44552) );
no03f01 g40761 ( .a(n44552), .b(n44550), .c(n34267), .o(n44553) );
in01f01 g40762 ( .a(n41352), .o(n44554) );
no02f01 g40763 ( .a(n41291), .b(n41280), .o(n44555) );
in01f01 g40764 ( .a(n44555), .o(n44556) );
no04f01 g40765 ( .a(n44556), .b(n44554), .c(n43522), .d(n39599), .o(n44557) );
ao12f01 g40766 ( .a(n34307), .b(n41356), .c(n41281), .o(n44558) );
in01f01 g40767 ( .a(n44550), .o(n44559) );
ao12f01 g40768 ( .a(n34307), .b(n44551), .c(n44559), .o(n44560) );
no02f01 g40769 ( .a(n44560), .b(n44558), .o(n44561) );
na02f01 g40770 ( .a(n44561), .b(n41371), .o(n44562) );
no02f01 g40771 ( .a(n44562), .b(n44557), .o(n44563) );
no03f01 g40772 ( .a(n44563), .b(n44553), .c(n44547), .o(n44564) );
in01f01 g40773 ( .a(n44547), .o(n44565) );
na04f01 g40774 ( .a(n44555), .b(n41352), .c(n41315), .d(n41294), .o(n44566) );
in01f01 g40775 ( .a(n44562), .o(n44567) );
ao12f01 g40776 ( .a(n44553), .b(n44567), .c(n44566), .o(n44568) );
no02f01 g40777 ( .a(n44568), .b(n44565), .o(n44569) );
oa12f01 g40778 ( .a(n32734), .b(n44569), .c(n44564), .o(n44570) );
na02f01 g40779 ( .a(n44570), .b(n44536), .o(n3248) );
na03f01 g40780 ( .a(n43824), .b(n43820), .c(n_27923), .o(n44572) );
no03f01 g40781 ( .a(n43823), .b(n43821), .c(n43815), .o(n44573) );
ao12f01 g40782 ( .a(n43818), .b(n43819), .c(n43816), .o(n44574) );
oa12f01 g40783 ( .a(n34420), .b(n44574), .c(n44573), .o(n44575) );
na02f01 g40784 ( .a(n44575), .b(n44572), .o(n3252) );
na02f01 g40785 ( .a(n1796), .b(n37149), .o(n44577) );
na03f01 g40786 ( .a(n44577), .b(n38834), .c(n42787), .o(n44578) );
na02f01 g40787 ( .a(n44577), .b(n38834), .o(n44579) );
na02f01 g40788 ( .a(n44579), .b(n42788), .o(n44580) );
na02f01 g40789 ( .a(n44580), .b(n44578), .o(n3257) );
na02f01 g40790 ( .a(n27672), .b(n42461), .o(n44582) );
no02f01 g40791 ( .a(n27572), .b(n27367), .o(n44583) );
no02f01 g40792 ( .a(n44583), .b(n27574), .o(n44584) );
na03f01 g40793 ( .a(n44584), .b(n27630), .c(n44582), .o(n44585) );
na02f01 g40794 ( .a(n27630), .b(n44582), .o(n44586) );
in01f01 g40795 ( .a(n44584), .o(n44587) );
na02f01 g40796 ( .a(n44587), .b(n44586), .o(n44588) );
na02f01 g40797 ( .a(n44588), .b(n44585), .o(n3262) );
in01f01 g40798 ( .a(n22566), .o(n44590) );
in01f01 g40799 ( .a(n22567), .o(n44591) );
no02f01 g40800 ( .a(n44591), .b(n22551), .o(n44592) );
na02f01 g40801 ( .a(n44592), .b(n44590), .o(n44593) );
oa12f01 g40802 ( .a(n22566), .b(n44591), .c(n22551), .o(n44594) );
na02f01 g40803 ( .a(n44594), .b(n44593), .o(n3267) );
oa12f01 g40804 ( .a(n29386), .b(n29698), .c(n29345), .o(n44596) );
na03f01 g40805 ( .a(n29387), .b(n29694), .c(n29677), .o(n44597) );
na02f01 g40806 ( .a(n44597), .b(n44596), .o(n3272) );
no03f01 g40807 ( .a(n37230), .b(n37208), .c(n37182), .o(n44599) );
in01f01 g40808 ( .a(n37239), .o(n44600) );
no02f01 g40809 ( .a(n37237), .b(n36963), .o(n44601) );
in01f01 g40810 ( .a(n44601), .o(n44602) );
na02f01 g40811 ( .a(n44602), .b(n37255), .o(n44603) );
ao12f01 g40812 ( .a(n44603), .b(n44600), .c(n44599), .o(n44604) );
no02f01 g40813 ( .a(n36963), .b(n7373), .o(n44605) );
no02f01 g40814 ( .a(n44605), .b(n37231), .o(n44606) );
na02f01 g40815 ( .a(n44606), .b(n44604), .o(n44607) );
in01f01 g40816 ( .a(n44604), .o(n44608) );
in01f01 g40817 ( .a(n44606), .o(n44609) );
na02f01 g40818 ( .a(n44609), .b(n44608), .o(n44610) );
na02f01 g40819 ( .a(n44610), .b(n44607), .o(n3282) );
ao12f01 g40820 ( .a(n37039), .b(n37031), .c(n37017), .o(n44612) );
no02f01 g40821 ( .a(n37040), .b(n37171), .o(n44613) );
na02f01 g40822 ( .a(n44613), .b(n44612), .o(n44614) );
in01f01 g40823 ( .a(n44612), .o(n44615) );
in01f01 g40824 ( .a(n44613), .o(n44616) );
na02f01 g40825 ( .a(n44616), .b(n44615), .o(n44617) );
na02f01 g40826 ( .a(n44617), .b(n44614), .o(n3292) );
no02f01 g40827 ( .a(n22292), .b(n22281), .o(n44619) );
no02f01 g40828 ( .a(n44619), .b(n42312), .o(n44620) );
na02f01 g40829 ( .a(n44619), .b(n42312), .o(n44621) );
in01f01 g40830 ( .a(n44621), .o(n44622) );
no02f01 g40831 ( .a(n44622), .b(n44620), .o(n44623) );
in01f01 g40832 ( .a(n44623), .o(n3297) );
ao12f01 g40833 ( .a(n13962), .b(n41155), .c(n13966), .o(n44625) );
in01f01 g40834 ( .a(n44625), .o(n44626) );
ao12f01 g40835 ( .a(n13926), .b(n44626), .c(n13963), .o(n44627) );
na02f01 g40836 ( .a(n13910), .b(n13909), .o(n44628) );
in01f01 g40837 ( .a(n44628), .o(n44629) );
no02f01 g40838 ( .a(n44629), .b(n44627), .o(n44630) );
na02f01 g40839 ( .a(n44629), .b(n44627), .o(n44631) );
in01f01 g40840 ( .a(n44631), .o(n44632) );
no02f01 g40841 ( .a(n44632), .b(n44630), .o(n44633) );
in01f01 g40842 ( .a(n44633), .o(n6061) );
na02f01 g40843 ( .a(n6061), .b(n4116), .o(n44635) );
na02f01 g40844 ( .a(n44633), .b(n2589), .o(n44636) );
na02f01 g40845 ( .a(n44636), .b(n44635), .o(n3302) );
na02f01 g40846 ( .a(n41162), .b(n2589), .o(n44638) );
na02f01 g40847 ( .a(n1290), .b(n4116), .o(n44639) );
na02f01 g40848 ( .a(n44639), .b(n44638), .o(n3307) );
ao12f01 g40849 ( .a(delay_sub_ln23_0_unr23_stage8_stallmux_q), .b(n38753), .c(n38751), .o(n44641) );
ao12f01 g40850 ( .a(n37149), .b(n38753), .c(n38751), .o(n44642) );
no02f01 g40851 ( .a(n44642), .b(n44641), .o(n44643) );
oa12f01 g40852 ( .a(n44643), .b(n38855), .c(n38845), .o(n44644) );
in01f01 g40853 ( .a(n38855), .o(n44645) );
in01f01 g40854 ( .a(n38751), .o(n44646) );
oa12f01 g40855 ( .a(n37149), .b(n38752), .c(n44646), .o(n44647) );
oa12f01 g40856 ( .a(delay_sub_ln23_0_unr23_stage8_stallmux_q), .b(n38752), .c(n44646), .o(n44648) );
na02f01 g40857 ( .a(n44648), .b(n44647), .o(n44649) );
na03f01 g40858 ( .a(n44649), .b(n44645), .c(n42455), .o(n44650) );
na02f01 g40859 ( .a(n44650), .b(n44644), .o(n3312) );
no02f01 g40860 ( .a(n36752), .b(n29639), .o(n44652) );
no02f01 g40861 ( .a(n44652), .b(n36754), .o(n44653) );
no03f01 g40862 ( .a(n43771), .b(n43766), .c(n36781), .o(n44654) );
oa12f01 g40863 ( .a(n44653), .b(n44654), .c(n36761), .o(n44655) );
in01f01 g40864 ( .a(n36761), .o(n44656) );
in01f01 g40865 ( .a(n44653), .o(n44657) );
in01f01 g40866 ( .a(n43766), .o(n44658) );
na03f01 g40867 ( .a(n43768), .b(n44658), .c(n43765), .o(n44659) );
na03f01 g40868 ( .a(n44659), .b(n44657), .c(n44656), .o(n44660) );
na02f01 g40869 ( .a(n44660), .b(n44655), .o(n3317) );
no02f01 g40870 ( .a(n40791), .b(n20159), .o(n44662) );
no02f01 g40871 ( .a(n44662), .b(n41207), .o(n44663) );
in01f01 g40872 ( .a(n44663), .o(n44664) );
na02f01 g40873 ( .a(n41190), .b(n41189), .o(n44665) );
no02f01 g40874 ( .a(n41195), .b(n44240), .o(n44666) );
oa12f01 g40875 ( .a(n44666), .b(n44665), .c(n40936), .o(n44667) );
no02f01 g40876 ( .a(n44667), .b(n44664), .o(n44668) );
in01f01 g40877 ( .a(n44668), .o(n44669) );
na02f01 g40878 ( .a(n44667), .b(n44664), .o(n44670) );
na03f01 g40879 ( .a(n44670), .b(n44669), .c(n5799), .o(n44671) );
in01f01 g40880 ( .a(n44670), .o(n44672) );
oa12f01 g40881 ( .a(n911), .b(n44672), .c(n44668), .o(n44673) );
na02f01 g40882 ( .a(n44673), .b(n44671), .o(n3322) );
no02f01 g40883 ( .a(n37871), .b(n26250), .o(n44675) );
in01f01 g40884 ( .a(n26250), .o(n44676) );
no02f01 g40885 ( .a(n38010), .b(n44676), .o(n44677) );
no02f01 g40886 ( .a(n44677), .b(n44675), .o(n44678) );
no03f01 g40887 ( .a(n41240), .b(n42671), .c(n41228), .o(n44679) );
oa12f01 g40888 ( .a(n44678), .b(n44679), .c(n42673), .o(n44680) );
in01f01 g40889 ( .a(n42673), .o(n44681) );
in01f01 g40890 ( .a(n44678), .o(n44682) );
in01f01 g40891 ( .a(n42671), .o(n44683) );
na03f01 g40892 ( .a(n41239), .b(n44683), .c(n41248), .o(n44684) );
na03f01 g40893 ( .a(n44684), .b(n44682), .c(n44681), .o(n44685) );
na03f01 g40894 ( .a(n44685), .b(n44680), .c(n1821), .o(n44686) );
ao12f01 g40895 ( .a(n44682), .b(n44684), .c(n44681), .o(n44687) );
no03f01 g40896 ( .a(n44679), .b(n44678), .c(n42673), .o(n44688) );
oa12f01 g40897 ( .a(n8066), .b(n44688), .c(n44687), .o(n44689) );
na02f01 g40898 ( .a(n44689), .b(n44686), .o(n3327) );
no02f01 g40899 ( .a(n42539), .b(n42538), .o(n44691) );
oa12f01 g40900 ( .a(n44691), .b(n32428), .c(n32493), .o(n44692) );
in01f01 g40901 ( .a(n44692), .o(n44693) );
no02f01 g40902 ( .a(n38228), .b(n31607), .o(n44694) );
no02f01 g40903 ( .a(n44694), .b(n32429), .o(n44695) );
na02f01 g40904 ( .a(n44695), .b(n44693), .o(n44696) );
in01f01 g40905 ( .a(n44695), .o(n44697) );
na02f01 g40906 ( .a(n44697), .b(n44692), .o(n44698) );
na02f01 g40907 ( .a(n44698), .b(n44696), .o(n3337) );
no02f01 g40908 ( .a(n37856), .b(n26440), .o(n44700) );
no02f01 g40909 ( .a(n37857), .b(n26441), .o(n44701) );
no02f01 g40910 ( .a(n44701), .b(n44700), .o(n44702) );
no02f01 g40911 ( .a(n27194), .b(n26740), .o(n44703) );
na02f01 g40912 ( .a(n44703), .b(n27166), .o(n44704) );
ao12f01 g40913 ( .a(n26440), .b(n27250), .c(n26738), .o(n44705) );
no02f01 g40914 ( .a(n44705), .b(n27172), .o(n44706) );
na03f01 g40915 ( .a(n44706), .b(n44704), .c(n44702), .o(n44707) );
in01f01 g40916 ( .a(n44702), .o(n44708) );
no03f01 g40917 ( .a(n27194), .b(n27249), .c(n26740), .o(n44709) );
in01f01 g40918 ( .a(n44706), .o(n44710) );
oa12f01 g40919 ( .a(n44708), .b(n44710), .c(n44709), .o(n44711) );
na02f01 g40920 ( .a(n44711), .b(n44707), .o(n3342) );
in01f01 g40921 ( .a(n40132), .o(n44713) );
no02f01 g40922 ( .a(n40177), .b(n44713), .o(n44714) );
in01f01 g40923 ( .a(n44714), .o(n44715) );
no02f01 g40924 ( .a(n44715), .b(n40176), .o(n44716) );
na02f01 g40925 ( .a(n44715), .b(n40176), .o(n44717) );
in01f01 g40926 ( .a(n44717), .o(n44718) );
no02f01 g40927 ( .a(n44718), .b(n44716), .o(n44719) );
na02f01 g40928 ( .a(n44719), .b(n5799), .o(n44720) );
in01f01 g40929 ( .a(n44719), .o(n4573) );
na02f01 g40930 ( .a(n4573), .b(n911), .o(n44722) );
na02f01 g40931 ( .a(n44722), .b(n44720), .o(n3347) );
na02f01 g40932 ( .a(n353), .b(n34420), .o(n44724) );
na03f01 g40933 ( .a(n29725), .b(n29669), .c(n_27923), .o(n44725) );
na02f01 g40934 ( .a(n44725), .b(n44724), .o(n3352) );
na02f01 g40935 ( .a(n42452), .b(n42451), .o(n3357) );
na02f01 g40936 ( .a(n22229), .b(n22225), .o(n44728) );
na02f01 g40937 ( .a(n44728), .b(n44441), .o(n3362) );
in01f01 g40938 ( .a(n39146), .o(n44730) );
no02f01 g40939 ( .a(n39157), .b(n44338), .o(n44731) );
oa12f01 g40940 ( .a(n44731), .b(n44730), .c(n39172), .o(n44732) );
in01f01 g40941 ( .a(n44732), .o(n44733) );
no02f01 g40942 ( .a(n39135), .b(n31502), .o(n44734) );
no02f01 g40943 ( .a(n44734), .b(n39148), .o(n44735) );
na02f01 g40944 ( .a(n44735), .b(n44733), .o(n44736) );
in01f01 g40945 ( .a(n44735), .o(n44737) );
na02f01 g40946 ( .a(n44737), .b(n44732), .o(n44738) );
na02f01 g40947 ( .a(n44738), .b(n44736), .o(n3367) );
na03f01 g40948 ( .a(n4967_1), .b(n4966), .c(n4985), .o(n44740) );
oa12f01 g40949 ( .a(n4989), .b(n4990), .c(n4959), .o(n44741) );
na02f01 g40950 ( .a(n44741), .b(n44740), .o(n3372) );
in01f01 g40951 ( .a(n40140), .o(n44743) );
no02f01 g40952 ( .a(n40175), .b(n44743), .o(n44744) );
na02f01 g40953 ( .a(n44744), .b(n40174), .o(n44745) );
in01f01 g40954 ( .a(n40174), .o(n44746) );
oa12f01 g40955 ( .a(n44746), .b(n40175), .c(n44743), .o(n44747) );
na02f01 g40956 ( .a(n44747), .b(n44745), .o(n3377) );
na02f01 g40957 ( .a(n42747), .b(n27412), .o(n44749) );
in01f01 g40958 ( .a(n44749), .o(n44750) );
na03f01 g40959 ( .a(n44750), .b(n42743), .c(n42745), .o(n44751) );
oa12f01 g40960 ( .a(n44749), .b(n42744), .c(n27488), .o(n44752) );
na02f01 g40961 ( .a(n44752), .b(n44751), .o(n3382) );
no02f01 g40962 ( .a(n29641), .b(n29430), .o(n44754) );
no02f01 g40963 ( .a(n29568), .b(n29639), .o(n44755) );
no02f01 g40964 ( .a(n44755), .b(n44754), .o(n44756) );
na02f01 g40965 ( .a(n29720), .b(n29719), .o(n44757) );
no02f01 g40966 ( .a(n29574), .b(n29639), .o(n44758) );
no02f01 g40967 ( .a(n29642), .b(n29430), .o(n44759) );
in01f01 g40968 ( .a(n44759), .o(n44760) );
ao12f01 g40969 ( .a(n44758), .b(n44760), .c(n44757), .o(n44761) );
na02f01 g40970 ( .a(n44761), .b(n44756), .o(n44762) );
in01f01 g40971 ( .a(n44756), .o(n44763) );
in01f01 g40972 ( .a(n44761), .o(n44764) );
na02f01 g40973 ( .a(n44764), .b(n44763), .o(n44765) );
na02f01 g40974 ( .a(n44765), .b(n44762), .o(n3387) );
no02f01 g40975 ( .a(n5912), .b(n5911), .o(n44767) );
no02f01 g40976 ( .a(n5920), .b(n6037), .o(n44768) );
no02f01 g40977 ( .a(n5919), .b(n5873), .o(n44769) );
no02f01 g40978 ( .a(n44769), .b(n44768), .o(n44770) );
na02f01 g40979 ( .a(n44770), .b(n44767), .o(n44771) );
oa22f01 g40980 ( .a(n44769), .b(n44768), .c(n5912), .d(n5911), .o(n44772) );
na02f01 g40981 ( .a(n44772), .b(n44771), .o(n3392) );
na03f01 g40982 ( .a(n42902), .b(n42901), .c(n1821), .o(n44774) );
na02f01 g40983 ( .a(n2082), .b(n8066), .o(n44775) );
na02f01 g40984 ( .a(n44775), .b(n44774), .o(n3397) );
na03f01 g40985 ( .a(n37362), .b(n37361), .c(n37358), .o(n44777) );
na02f01 g40986 ( .a(n1595), .b(n37149), .o(n44778) );
na03f01 g40987 ( .a(n44778), .b(n37365), .c(n44777), .o(n44779) );
na02f01 g40988 ( .a(n37361), .b(n37358), .o(n44780) );
in01f01 g40989 ( .a(n44780), .o(n44781) );
na02f01 g40990 ( .a(n44778), .b(n37365), .o(n44782) );
na03f01 g40991 ( .a(n44782), .b(n37362), .c(n44781), .o(n44783) );
na02f01 g40992 ( .a(n44783), .b(n44779), .o(n3402) );
na02f01 g40993 ( .a(n32732), .b(sin_out_29), .o(n44785) );
no02f01 g40994 ( .a(n35860), .b(n41267), .o(n44786) );
no02f01 g40995 ( .a(n44786), .b(n35889), .o(n44787) );
no02f01 g40996 ( .a(n35877), .b(n34336), .o(n44788) );
no02f01 g40997 ( .a(n35876), .b(n34287), .o(n44789) );
no02f01 g40998 ( .a(n44789), .b(n44788), .o(n44790) );
no02f01 g40999 ( .a(n44790), .b(n44787), .o(n44791) );
na02f01 g41000 ( .a(n44790), .b(n44787), .o(n44792) );
in01f01 g41001 ( .a(n44792), .o(n44793) );
no02f01 g41002 ( .a(n44793), .b(n44791), .o(n44794) );
in01f01 g41003 ( .a(n44794), .o(n44795) );
no02f01 g41004 ( .a(n44795), .b(n34267), .o(n44796) );
no03f01 g41005 ( .a(n44556), .b(n44553), .c(n44544), .o(n44797) );
in01f01 g41006 ( .a(n44797), .o(n44798) );
no04f01 g41007 ( .a(n44798), .b(n44554), .c(n43522), .d(n39599), .o(n44799) );
na02f01 g41008 ( .a(n44561), .b(n44545), .o(n44800) );
na02f01 g41009 ( .a(n44800), .b(n34267), .o(n44801) );
na02f01 g41010 ( .a(n44801), .b(n41371), .o(n44802) );
no02f01 g41011 ( .a(n44794), .b(n34307), .o(n44803) );
no03f01 g41012 ( .a(n44803), .b(n44802), .c(n44799), .o(n44804) );
no02f01 g41013 ( .a(n44788), .b(n44787), .o(n44805) );
no02f01 g41014 ( .a(n44805), .b(n44789), .o(n44806) );
no02f01 g41015 ( .a(n35870), .b(n34287), .o(n44807) );
no02f01 g41016 ( .a(n35871), .b(n34336), .o(n44808) );
no02f01 g41017 ( .a(n44808), .b(n44807), .o(n44809) );
no02f01 g41018 ( .a(n44809), .b(n44806), .o(n44810) );
na02f01 g41019 ( .a(n44809), .b(n44806), .o(n44811) );
in01f01 g41020 ( .a(n44811), .o(n44812) );
no03f01 g41021 ( .a(n44812), .b(n44810), .c(n34267), .o(n44813) );
no02f01 g41022 ( .a(n44812), .b(n44810), .o(n44814) );
no02f01 g41023 ( .a(n44814), .b(n34307), .o(n44815) );
no02f01 g41024 ( .a(n44815), .b(n44813), .o(n44816) );
no03f01 g41025 ( .a(n44816), .b(n44804), .c(n44796), .o(n44817) );
in01f01 g41026 ( .a(n44796), .o(n44818) );
na04f01 g41027 ( .a(n44797), .b(n41352), .c(n41315), .d(n41294), .o(n44819) );
in01f01 g41028 ( .a(n44802), .o(n44820) );
in01f01 g41029 ( .a(n44803), .o(n44821) );
na03f01 g41030 ( .a(n44821), .b(n44820), .c(n44819), .o(n44822) );
in01f01 g41031 ( .a(n44816), .o(n44823) );
ao12f01 g41032 ( .a(n44823), .b(n44822), .c(n44818), .o(n44824) );
oa12f01 g41033 ( .a(n32734), .b(n44824), .c(n44817), .o(n44825) );
na02f01 g41034 ( .a(n44825), .b(n44785), .o(n3407) );
no02f01 g41035 ( .a(n38907), .b(n38896), .o(n44827) );
in01f01 g41036 ( .a(n44827), .o(n44828) );
na03f01 g41037 ( .a(n44828), .b(n38888), .c(n38886), .o(n44829) );
na02f01 g41038 ( .a(n38888), .b(n38886), .o(n44830) );
na02f01 g41039 ( .a(n44827), .b(n44830), .o(n44831) );
na02f01 g41040 ( .a(n44831), .b(n44829), .o(n3411) );
na03f01 g41041 ( .a(n32471), .b(n32355), .c(n32336), .o(n44833) );
oa12f01 g41042 ( .a(n32466), .b(n32376), .c(n32356), .o(n44834) );
na02f01 g41043 ( .a(n44834), .b(n44833), .o(n3416) );
in01f01 g41044 ( .a(n22178), .o(n44836) );
oa12f01 g41045 ( .a(n22236), .b(n44836), .c(n22177), .o(n44837) );
in01f01 g41046 ( .a(n22236), .o(n44838) );
no02f01 g41047 ( .a(n44836), .b(n22177), .o(n44839) );
na02f01 g41048 ( .a(n44839), .b(n44838), .o(n44840) );
na02f01 g41049 ( .a(n44840), .b(n44837), .o(n3421) );
no02f01 g41050 ( .a(n42445), .b(n42444), .o(n44842) );
in01f01 g41051 ( .a(n44842), .o(n3426) );
na03f01 g41052 ( .a(n38173), .b(n9590), .c(n9589), .o(n44844) );
oa12f01 g41053 ( .a(n599), .b(n9646), .c(n9645), .o(n44845) );
na02f01 g41054 ( .a(n44845), .b(n44844), .o(n3431) );
no02f01 g41055 ( .a(n10852), .b(n10735), .o(n44847) );
no02f01 g41056 ( .a(n10851), .b(n3521), .o(n44848) );
oa22f01 g41057 ( .a(n44848), .b(n44847), .c(n10854), .d(n10844), .o(n44849) );
no02f01 g41058 ( .a(n10854), .b(n10844), .o(n44850) );
no02f01 g41059 ( .a(n44848), .b(n44847), .o(n44851) );
na02f01 g41060 ( .a(n44851), .b(n44850), .o(n44852) );
na02f01 g41061 ( .a(n44852), .b(n44849), .o(n3436) );
na02f01 g41062 ( .a(n1075), .b(n34420), .o(n44854) );
na03f01 g41063 ( .a(n40454), .b(n40450), .c(n_27923), .o(n44855) );
na02f01 g41064 ( .a(n44855), .b(n44854), .o(n3441) );
no02f01 g41065 ( .a(n9829), .b(n5001), .o(n44857) );
in01f01 g41066 ( .a(n44857), .o(n44858) );
no02f01 g41067 ( .a(n9842), .b(n5001), .o(n44859) );
no02f01 g41068 ( .a(n44859), .b(n9844), .o(n44860) );
na03f01 g41069 ( .a(n44860), .b(n44858), .c(n39647), .o(n44861) );
in01f01 g41070 ( .a(n44860), .o(n44862) );
oa12f01 g41071 ( .a(n44862), .b(n44857), .c(n9832), .o(n44863) );
na02f01 g41072 ( .a(n44863), .b(n44861), .o(n3446) );
no02f01 g41073 ( .a(n9425), .b(n9295), .o(n44865) );
na02f01 g41074 ( .a(n44865), .b(n9423), .o(n44866) );
in01f01 g41075 ( .a(n44865), .o(n44867) );
na02f01 g41076 ( .a(n44867), .b(n9629), .o(n44868) );
na02f01 g41077 ( .a(n44868), .b(n44866), .o(n3451) );
oa12f01 g41078 ( .a(n21161), .b(n21156), .c(n21155), .o(n44870) );
na02f01 g41079 ( .a(n44870), .b(n21163), .o(n3461) );
ao12f01 g41080 ( .a(n36088), .b(n36092), .c(n38767), .o(n44872) );
in01f01 g41081 ( .a(n44872), .o(n44873) );
no02f01 g41082 ( .a(n38770), .b(n36076), .o(n44874) );
na02f01 g41083 ( .a(n44874), .b(n44873), .o(n44875) );
in01f01 g41084 ( .a(n44874), .o(n44876) );
na02f01 g41085 ( .a(n44876), .b(n44872), .o(n44877) );
na02f01 g41086 ( .a(n44877), .b(n44875), .o(n3471) );
oa12f01 g41087 ( .a(n29692), .b(n29385), .c(n29680), .o(n44879) );
na03f01 g41088 ( .a(n29693), .b(n29384), .c(n29352), .o(n44880) );
na02f01 g41089 ( .a(n44880), .b(n44879), .o(n3476) );
no02f01 g41090 ( .a(n9797), .b(n40341), .o(n44882) );
no02f01 g41091 ( .a(n44882), .b(n9819), .o(n44883) );
in01f01 g41092 ( .a(n9815), .o(n44884) );
na02f01 g41093 ( .a(n9821), .b(n44884), .o(n44885) );
in01f01 g41094 ( .a(n44885), .o(n44886) );
na02f01 g41095 ( .a(n44886), .b(n44883), .o(n44887) );
oa12f01 g41096 ( .a(n44885), .b(n44882), .c(n9819), .o(n44888) );
na02f01 g41097 ( .a(n44888), .b(n44887), .o(n3481) );
na02f01 g41098 ( .a(n42919), .b(n42915), .o(n3486) );
na03f01 g41099 ( .a(n25476), .b(n36650), .c(n25466), .o(n44891) );
oa12f01 g41100 ( .a(n36647), .b(n25482), .c(n25474), .o(n44892) );
na02f01 g41101 ( .a(n44892), .b(n44891), .o(n3491) );
ao12f01 g41102 ( .a(n32356), .b(n32471), .c(n32336), .o(n44894) );
in01f01 g41103 ( .a(n44894), .o(n44895) );
no02f01 g41104 ( .a(n32382), .b(n32375), .o(n44896) );
na02f01 g41105 ( .a(n44896), .b(n44895), .o(n44897) );
in01f01 g41106 ( .a(n44896), .o(n44898) );
na02f01 g41107 ( .a(n44898), .b(n44894), .o(n44899) );
na02f01 g41108 ( .a(n44899), .b(n44897), .o(n3496) );
no02f01 g41109 ( .a(n25600), .b(n36454), .o(n44901) );
no02f01 g41110 ( .a(n44901), .b(n25608), .o(n44902) );
na02f01 g41111 ( .a(n44901), .b(n25608), .o(n44903) );
in01f01 g41112 ( .a(n44903), .o(n44904) );
no02f01 g41113 ( .a(n44904), .b(n44902), .o(n44905) );
in01f01 g41114 ( .a(n44905), .o(n4613) );
na02f01 g41115 ( .a(n4613), .b(n4116), .o(n44907) );
na02f01 g41116 ( .a(n44905), .b(n2589), .o(n44908) );
na02f01 g41117 ( .a(n44908), .b(n44907), .o(n3501) );
in01f01 g41118 ( .a(n40178), .o(n44910) );
no02f01 g41119 ( .a(n40180), .b(n40123), .o(n44911) );
in01f01 g41120 ( .a(n44911), .o(n44912) );
no02f01 g41121 ( .a(n44912), .b(n44910), .o(n44913) );
no02f01 g41122 ( .a(n44911), .b(n40178), .o(n44914) );
no02f01 g41123 ( .a(n44914), .b(n44913), .o(n44915) );
na02f01 g41124 ( .a(n44915), .b(n5799), .o(n44916) );
in01f01 g41125 ( .a(n44915), .o(n4349) );
na02f01 g41126 ( .a(n4349), .b(n911), .o(n44918) );
na02f01 g41127 ( .a(n44918), .b(n44916), .o(n3506) );
in01f01 g41128 ( .a(n8473), .o(n44920) );
oa12f01 g41129 ( .a(n44920), .b(n8469), .c(n43575), .o(n44921) );
no02f01 g41130 ( .a(n8475), .b(n8460), .o(n44922) );
in01f01 g41131 ( .a(n44922), .o(n44923) );
na02f01 g41132 ( .a(n44923), .b(n44921), .o(n44924) );
in01f01 g41133 ( .a(n44921), .o(n44925) );
na02f01 g41134 ( .a(n44922), .b(n44925), .o(n44926) );
na02f01 g41135 ( .a(n44926), .b(n44924), .o(n3511) );
ao12f01 g41136 ( .a(n22467), .b(n42735), .c(n22463), .o(n44928) );
no02f01 g41137 ( .a(n22459), .b(n22069), .o(n44929) );
in01f01 g41138 ( .a(n44929), .o(n44930) );
no02f01 g41139 ( .a(n44930), .b(n44928), .o(n44931) );
na02f01 g41140 ( .a(n44930), .b(n44928), .o(n44932) );
in01f01 g41141 ( .a(n44932), .o(n44933) );
no02f01 g41142 ( .a(n44933), .b(n44931), .o(n44934) );
in01f01 g41143 ( .a(n44934), .o(n5440) );
na02f01 g41144 ( .a(n5440), .b(n4116), .o(n44936) );
na02f01 g41145 ( .a(n44934), .b(n2589), .o(n44937) );
na02f01 g41146 ( .a(n44937), .b(n44936), .o(n3516) );
in01f01 g41147 ( .a(n22360), .o(n44939) );
no02f01 g41148 ( .a(n22361), .b(n22465), .o(n44940) );
no02f01 g41149 ( .a(n44940), .b(n44939), .o(n44941) );
na02f01 g41150 ( .a(n44940), .b(n44939), .o(n44942) );
in01f01 g41151 ( .a(n44942), .o(n44943) );
no02f01 g41152 ( .a(n44943), .b(n44941), .o(n44944) );
in01f01 g41153 ( .a(n44944), .o(n3526) );
na02f01 g41154 ( .a(n32732), .b(sin_out_14), .o(n44946) );
ao12f01 g41155 ( .a(n39595), .b(n39565), .c(n39496), .o(n44947) );
in01f01 g41156 ( .a(n44947), .o(n44948) );
no02f01 g41157 ( .a(n43093), .b(n39577), .o(n44949) );
in01f01 g41158 ( .a(n44949), .o(n44950) );
no02f01 g41159 ( .a(n44950), .b(n44948), .o(n44951) );
no02f01 g41160 ( .a(n44949), .b(n44947), .o(n44952) );
oa12f01 g41161 ( .a(n32734), .b(n44952), .c(n44951), .o(n44953) );
na02f01 g41162 ( .a(n44953), .b(n44946), .o(n3531) );
in01f01 g41163 ( .a(n43920), .o(n44955) );
in01f01 g41164 ( .a(n43921), .o(n44956) );
oa12f01 g41165 ( .a(n44956), .b(n42013), .c(n43918), .o(n44957) );
no02f01 g41166 ( .a(n42007), .b(n10735), .o(n44958) );
no02f01 g41167 ( .a(n42006), .b(n3521), .o(n44959) );
no02f01 g41168 ( .a(n44959), .b(n44958), .o(n44960) );
na03f01 g41169 ( .a(n44960), .b(n44957), .c(n44955), .o(n44961) );
na02f01 g41170 ( .a(n44957), .b(n44955), .o(n44962) );
in01f01 g41171 ( .a(n44960), .o(n44963) );
na02f01 g41172 ( .a(n44963), .b(n44962), .o(n44964) );
na02f01 g41173 ( .a(n44964), .b(n44961), .o(n3535) );
no02f01 g41174 ( .a(n37375), .b(n8420), .o(n44966) );
na02f01 g41175 ( .a(n44966), .b(cordic_combinational_sub_ln23_0_unr16_z_0_), .o(n44967) );
oa12f01 g41176 ( .a(n7703), .b(n37375), .c(n8420), .o(n44968) );
na02f01 g41177 ( .a(n44968), .b(n44967), .o(n3540) );
no02f01 g41178 ( .a(n38004), .b(n38024), .o(n44970) );
no02f01 g41179 ( .a(n44970), .b(n38046), .o(n44971) );
na02f01 g41180 ( .a(n44970), .b(n38046), .o(n44972) );
in01f01 g41181 ( .a(n44972), .o(n44973) );
no02f01 g41182 ( .a(n44973), .b(n44971), .o(n44974) );
in01f01 g41183 ( .a(n44974), .o(n3545) );
in01f01 g41184 ( .a(n10972), .o(n44976) );
oa12f01 g41185 ( .a(n10927), .b(n10970), .c(n10924), .o(n44977) );
in01f01 g41186 ( .a(n44977), .o(n44978) );
no02f01 g41187 ( .a(n10944), .b(n3521), .o(n44979) );
no02f01 g41188 ( .a(n44979), .b(n10946), .o(n44980) );
na03f01 g41189 ( .a(n44980), .b(n44978), .c(n44976), .o(n44981) );
in01f01 g41190 ( .a(n44980), .o(n44982) );
oa12f01 g41191 ( .a(n44982), .b(n44977), .c(n10972), .o(n44983) );
na02f01 g41192 ( .a(n44983), .b(n44981), .o(n3550) );
ao12f01 g41193 ( .a(n22465), .b(n22362), .c(n22360), .o(n44985) );
no02f01 g41194 ( .a(n22116), .b(n22464), .o(n44986) );
no02f01 g41195 ( .a(n44986), .b(n44985), .o(n44987) );
na02f01 g41196 ( .a(n44986), .b(n44985), .o(n44988) );
in01f01 g41197 ( .a(n44988), .o(n44989) );
no02f01 g41198 ( .a(n44989), .b(n44987), .o(n44990) );
in01f01 g41199 ( .a(n44990), .o(n4389) );
na02f01 g41200 ( .a(n4389), .b(n4116), .o(n44992) );
na02f01 g41201 ( .a(n44990), .b(n2589), .o(n44993) );
na02f01 g41202 ( .a(n44993), .b(n44992), .o(n3555) );
na02f01 g41203 ( .a(n44014), .b(n38120), .o(n44995) );
no02f01 g41204 ( .a(n38135), .b(n38127), .o(n44996) );
na03f01 g41205 ( .a(n44996), .b(n44995), .c(n38139), .o(n44997) );
oa12f01 g41206 ( .a(n38139), .b(n41664), .c(n38121), .o(n44998) );
in01f01 g41207 ( .a(n44996), .o(n44999) );
na02f01 g41208 ( .a(n44999), .b(n44998), .o(n45000) );
na02f01 g41209 ( .a(n45000), .b(n44997), .o(n3560) );
no02f01 g41210 ( .a(n29416), .b(n29413), .o(n45002) );
oa12f01 g41211 ( .a(n45002), .b(n29420), .c(n29267), .o(n45003) );
in01f01 g41212 ( .a(n45002), .o(n45004) );
na03f01 g41213 ( .a(n29713), .b(n45004), .c(n29671), .o(n45005) );
na02f01 g41214 ( .a(n45005), .b(n45003), .o(n3565) );
no02f01 g41215 ( .a(n42384), .b(n41724), .o(n45007) );
na03f01 g41216 ( .a(n45007), .b(n42383), .c(n42380), .o(n45008) );
in01f01 g41217 ( .a(n45007), .o(n45009) );
oa12f01 g41218 ( .a(n45009), .b(n42382), .c(n42389), .o(n45010) );
na02f01 g41219 ( .a(n45010), .b(n45008), .o(n3570) );
na03f01 g41220 ( .a(n44738), .b(n44736), .c(n3633), .o(n45012) );
na02f01 g41221 ( .a(n3367), .b(n6203), .o(n45013) );
na02f01 g41222 ( .a(n45013), .b(n45012), .o(n3575) );
ao12f01 g41223 ( .a(n9634), .b(n9633), .c(n9615), .o(n45015) );
no02f01 g41224 ( .a(n9435), .b(n9260), .o(n45016) );
in01f01 g41225 ( .a(n45016), .o(n45017) );
na02f01 g41226 ( .a(n45017), .b(n45015), .o(n45018) );
in01f01 g41227 ( .a(n45015), .o(n45019) );
na02f01 g41228 ( .a(n45016), .b(n45019), .o(n45020) );
na02f01 g41229 ( .a(n45020), .b(n45018), .o(n3580) );
no02f01 g41230 ( .a(n9528), .b(n9506), .o(n45022) );
no02f01 g41231 ( .a(n9530), .b(n9515), .o(n45023) );
na02f01 g41232 ( .a(n45023), .b(n45022), .o(n45024) );
in01f01 g41233 ( .a(n45022), .o(n45025) );
in01f01 g41234 ( .a(n45023), .o(n45026) );
na02f01 g41235 ( .a(n45026), .b(n45025), .o(n45027) );
na02f01 g41236 ( .a(n45027), .b(n45024), .o(n3585) );
na02f01 g41237 ( .a(n42417), .b(n6037), .o(n45029) );
na02f01 g41238 ( .a(n1816), .b(n5873), .o(n45030) );
na02f01 g41239 ( .a(n45030), .b(n45029), .o(n3590) );
na03f01 g41240 ( .a(n17957), .b(n17956), .c(n17916), .o(n45032) );
oa12f01 g41241 ( .a(n17937), .b(n17938), .c(n17946), .o(n45033) );
na02f01 g41242 ( .a(n45033), .b(n45032), .o(n3595) );
na02f01 g41243 ( .a(n32732), .b(cos_out_21), .o(n45035) );
na02f01 g41244 ( .a(n39707), .b(n39691), .o(n45036) );
no02f01 g41245 ( .a(n39706), .b(n39695), .o(n45037) );
na02f01 g41246 ( .a(n45037), .b(n45036), .o(n45038) );
in01f01 g41247 ( .a(n41481), .o(n45039) );
no02f01 g41248 ( .a(n41477), .b(n35944), .o(n45040) );
no02f01 g41249 ( .a(n45040), .b(n45039), .o(n45041) );
in01f01 g41250 ( .a(n45041), .o(n45042) );
no02f01 g41251 ( .a(n45042), .b(n45038), .o(n45043) );
ao12f01 g41252 ( .a(n45041), .b(n45037), .c(n45036), .o(n45044) );
oa12f01 g41253 ( .a(n32734), .b(n45044), .c(n45043), .o(n45045) );
na02f01 g41254 ( .a(n45045), .b(n45035), .o(n3600) );
in01f01 g41255 ( .a(n37080), .o(n45047) );
ao12f01 g41256 ( .a(n37105), .b(n45047), .c(n37180), .o(n45048) );
no02f01 g41257 ( .a(n37100), .b(n36963), .o(n45049) );
no02f01 g41258 ( .a(n45049), .b(n37102), .o(n45050) );
na02f01 g41259 ( .a(n45050), .b(n45048), .o(n45051) );
in01f01 g41260 ( .a(n45048), .o(n45052) );
in01f01 g41261 ( .a(n45050), .o(n45053) );
na02f01 g41262 ( .a(n45053), .b(n45052), .o(n45054) );
na02f01 g41263 ( .a(n45054), .b(n45051), .o(n3604) );
oa12f01 g41264 ( .a(n8738), .b(n8758), .c(n8716), .o(n45056) );
no02f01 g41265 ( .a(n8745), .b(n5973), .o(n45057) );
no02f01 g41266 ( .a(n45057), .b(n8747), .o(n45058) );
na03f01 g41267 ( .a(n45058), .b(n45056), .c(n8760), .o(n45059) );
na02f01 g41268 ( .a(n45056), .b(n8760), .o(n45060) );
in01f01 g41269 ( .a(n45058), .o(n45061) );
na02f01 g41270 ( .a(n45061), .b(n45060), .o(n45062) );
na02f01 g41271 ( .a(n45062), .b(n45059), .o(n3609) );
na03f01 g41272 ( .a(n32457), .b(n32456), .c(n32314), .o(n45064) );
oa12f01 g41273 ( .a(n32321), .b(n32322), .c(n32453), .o(n45065) );
na02f01 g41274 ( .a(n45065), .b(n45064), .o(n3614) );
na02f01 g41275 ( .a(n32732), .b(sin_out_19), .o(n45067) );
na02f01 g41276 ( .a(n41295), .b(n41294), .o(n45068) );
no02f01 g41277 ( .a(n45068), .b(n41314), .o(n45069) );
no02f01 g41278 ( .a(n41358), .b(n34307), .o(n45070) );
in01f01 g41279 ( .a(n45070), .o(n45071) );
in01f01 g41280 ( .a(n41360), .o(n45072) );
na02f01 g41281 ( .a(n45072), .b(n45071), .o(n45073) );
no02f01 g41282 ( .a(n41357), .b(n34307), .o(n45074) );
no02f01 g41283 ( .a(n45074), .b(n41308), .o(n45075) );
in01f01 g41284 ( .a(n45075), .o(n45076) );
no03f01 g41285 ( .a(n45076), .b(n45073), .c(n45069), .o(n45077) );
no02f01 g41286 ( .a(n45073), .b(n45069), .o(n45078) );
no02f01 g41287 ( .a(n45075), .b(n45078), .o(n45079) );
oa12f01 g41288 ( .a(n32734), .b(n45079), .c(n45077), .o(n45080) );
na02f01 g41289 ( .a(n45080), .b(n45067), .o(n3619) );
in01f01 g41290 ( .a(n42866), .o(n45082) );
in01f01 g41291 ( .a(n42870), .o(n45083) );
no02f01 g41292 ( .a(n42858), .b(n35531), .o(n45084) );
no02f01 g41293 ( .a(n42873), .b(n35542), .o(n45085) );
in01f01 g41294 ( .a(n45085), .o(n45086) );
no02f01 g41295 ( .a(n45086), .b(n45084), .o(n45087) );
na02f01 g41296 ( .a(n45087), .b(n45083), .o(n45088) );
na02f01 g41297 ( .a(n45088), .b(n45082), .o(n45089) );
no02f01 g41298 ( .a(n42844), .b(n4176), .o(n45090) );
no02f01 g41299 ( .a(n45090), .b(n42846), .o(n45091) );
na02f01 g41300 ( .a(n45091), .b(n45089), .o(n45092) );
in01f01 g41301 ( .a(n45091), .o(n45093) );
na03f01 g41302 ( .a(n45093), .b(n45088), .c(n45082), .o(n45094) );
na02f01 g41303 ( .a(n45094), .b(n45092), .o(n3628) );
in01f01 g41304 ( .a(n35529), .o(n45096) );
no02f01 g41305 ( .a(n35527), .b(n4176), .o(n45097) );
in01f01 g41306 ( .a(n45097), .o(n45098) );
na02f01 g41307 ( .a(n35486), .b(n35441), .o(n45099) );
in01f01 g41308 ( .a(n35536), .o(n45100) );
no02f01 g41309 ( .a(n35538), .b(n45100), .o(n45101) );
oa12f01 g41310 ( .a(n45101), .b(n35509), .c(n45099), .o(n45102) );
in01f01 g41311 ( .a(n45102), .o(n45103) );
na02f01 g41312 ( .a(n45103), .b(n45098), .o(n45104) );
na02f01 g41313 ( .a(n45104), .b(n45096), .o(n45105) );
no02f01 g41314 ( .a(n35539), .b(n4176), .o(n45106) );
no02f01 g41315 ( .a(n45106), .b(n35520), .o(n45107) );
na02f01 g41316 ( .a(n45107), .b(n45105), .o(n45108) );
in01f01 g41317 ( .a(n45107), .o(n45109) );
na03f01 g41318 ( .a(n45109), .b(n45104), .c(n45096), .o(n45110) );
na02f01 g41319 ( .a(n45110), .b(n45108), .o(n3638) );
in01f01 g41320 ( .a(n27397), .o(n45112) );
na02f01 g41321 ( .a(n45112), .b(n44001), .o(n45113) );
in01f01 g41322 ( .a(n45113), .o(n45114) );
na02f01 g41323 ( .a(n45114), .b(n44000), .o(n45115) );
na02f01 g41324 ( .a(n45113), .b(n43999), .o(n45116) );
na02f01 g41325 ( .a(n45116), .b(n45115), .o(n3643) );
no02f01 g41326 ( .a(n25916), .b(n25780), .o(n45118) );
no02f01 g41327 ( .a(n25917), .b(n30065), .o(n45119) );
no02f01 g41328 ( .a(n45119), .b(n45118), .o(n45120) );
na03f01 g41329 ( .a(n45120), .b(n30103), .c(n30102), .o(n45121) );
oa22f01 g41330 ( .a(n45119), .b(n45118), .c(n25911), .d(n25908), .o(n45122) );
na02f01 g41331 ( .a(n45122), .b(n45121), .o(n3648) );
na02f01 g41332 ( .a(n41706), .b(n41696), .o(n3658) );
na02f01 g41333 ( .a(n44147), .b(n44143), .o(n3668) );
na02f01 g41334 ( .a(n609), .b(n4116), .o(n45126) );
na02f01 g41335 ( .a(n38191), .b(n2589), .o(n45127) );
na02f01 g41336 ( .a(n45127), .b(n45126), .o(n3678) );
no02f01 g41337 ( .a(n41080), .b(n41077), .o(n45129) );
in01f01 g41338 ( .a(n45129), .o(n45130) );
no03f01 g41339 ( .a(n45130), .b(n30131), .c(n30129), .o(n45131) );
no02f01 g41340 ( .a(n45129), .b(n41079), .o(n45132) );
no02f01 g41341 ( .a(n45132), .b(n45131), .o(n45133) );
na02f01 g41342 ( .a(n45133), .b(n6037), .o(n45134) );
in01f01 g41343 ( .a(n45133), .o(n5903) );
na02f01 g41344 ( .a(n5903), .b(n5873), .o(n45136) );
na02f01 g41345 ( .a(n45136), .b(n45134), .o(n3683) );
no02f01 g41346 ( .a(n27522), .b(n27367), .o(n45138) );
na02f01 g41347 ( .a(n27522), .b(n27367), .o(n45139) );
in01f01 g41348 ( .a(n45139), .o(n45140) );
no02f01 g41349 ( .a(n45140), .b(n45138), .o(n45141) );
na02f01 g41350 ( .a(n45141), .b(n27495), .o(n45142) );
in01f01 g41351 ( .a(n45141), .o(n45143) );
na02f01 g41352 ( .a(n45143), .b(n27671), .o(n45144) );
na02f01 g41353 ( .a(n45144), .b(n45142), .o(n3688) );
na02f01 g41354 ( .a(n42801), .b(n6037), .o(n45146) );
na02f01 g41355 ( .a(n2058), .b(n5873), .o(n45147) );
na02f01 g41356 ( .a(n45147), .b(n45146), .o(n3693) );
in01f01 g41357 ( .a(n43692), .o(n45149) );
ao12f01 g41358 ( .a(n43691), .b(n45149), .c(n10928), .o(n45150) );
no02f01 g41359 ( .a(n10969), .b(n10735), .o(n45151) );
no02f01 g41360 ( .a(n10968), .b(n3521), .o(n45152) );
no02f01 g41361 ( .a(n45152), .b(n45151), .o(n45153) );
na02f01 g41362 ( .a(n45153), .b(n45150), .o(n45154) );
in01f01 g41363 ( .a(n45150), .o(n45155) );
in01f01 g41364 ( .a(n45153), .o(n45156) );
na02f01 g41365 ( .a(n45156), .b(n45155), .o(n45157) );
na02f01 g41366 ( .a(n45157), .b(n45154), .o(n3698) );
na02f01 g41367 ( .a(n32732), .b(cos_out_13), .o(n45159) );
no02f01 g41368 ( .a(n36339), .b(n39048), .o(n45160) );
no02f01 g41369 ( .a(n36329), .b(n35944), .o(n45161) );
no02f01 g41370 ( .a(n45161), .b(n36331), .o(n45162) );
in01f01 g41371 ( .a(n45162), .o(n45163) );
no04f01 g41372 ( .a(n45163), .b(n45160), .c(n39044), .d(n36369), .o(n45164) );
no03f01 g41373 ( .a(n45160), .b(n39044), .c(n36369), .o(n45165) );
no02f01 g41374 ( .a(n45162), .b(n45165), .o(n45166) );
oa12f01 g41375 ( .a(n32734), .b(n45166), .c(n45164), .o(n45167) );
na02f01 g41376 ( .a(n45167), .b(n45159), .o(n3703) );
na03f01 g41377 ( .a(n44246), .b(n44243), .c(n5799), .o(n45169) );
na02f01 g41378 ( .a(n2996), .b(n911), .o(n45170) );
na02f01 g41379 ( .a(n45170), .b(n45169), .o(n3712) );
na03f01 g41380 ( .a(n25862), .b(n30085), .c(n25852), .o(n45172) );
oa12f01 g41381 ( .a(n30082), .b(n30086), .c(n25861), .o(n45173) );
na02f01 g41382 ( .a(n45173), .b(n45172), .o(n3717) );
no02f01 g41383 ( .a(n40046), .b(n40045), .o(n45175) );
in01f01 g41384 ( .a(n45175), .o(n45176) );
no02f01 g41385 ( .a(n39872), .b(n39860), .o(n45177) );
no02f01 g41386 ( .a(n39873), .b(n39861), .o(n45178) );
in01f01 g41387 ( .a(n45178), .o(n45179) );
ao12f01 g41388 ( .a(n45177), .b(n45179), .c(n45176), .o(n45180) );
no02f01 g41389 ( .a(n39882), .b(n39860), .o(n45181) );
no02f01 g41390 ( .a(n39883), .b(n39861), .o(n45182) );
no02f01 g41391 ( .a(n45182), .b(n45181), .o(n45183) );
na02f01 g41392 ( .a(n45183), .b(n45180), .o(n45184) );
in01f01 g41393 ( .a(n45180), .o(n45185) );
in01f01 g41394 ( .a(n45183), .o(n45186) );
na02f01 g41395 ( .a(n45186), .b(n45185), .o(n45187) );
na02f01 g41396 ( .a(n45187), .b(n45184), .o(n3722) );
no02f01 g41397 ( .a(n40771), .b(n21305), .o(n45189) );
no02f01 g41398 ( .a(n40715), .b(n21270), .o(n45190) );
no02f01 g41399 ( .a(n45190), .b(n45189), .o(n45191) );
in01f01 g41400 ( .a(n21309), .o(n45192) );
oa12f01 g41401 ( .a(n45192), .b(n21302), .c(n21335), .o(n45193) );
na02f01 g41402 ( .a(n45193), .b(n45191), .o(n45194) );
no02f01 g41403 ( .a(n45193), .b(n45191), .o(n45195) );
in01f01 g41404 ( .a(n45195), .o(n45196) );
na03f01 g41405 ( .a(n45196), .b(n45194), .c(n5799), .o(n45197) );
in01f01 g41406 ( .a(n45194), .o(n45198) );
oa12f01 g41407 ( .a(n911), .b(n45195), .c(n45198), .o(n45199) );
na02f01 g41408 ( .a(n45199), .b(n45197), .o(n3727) );
no02f01 g41409 ( .a(n8561), .b(n8557), .o(n45201) );
no02f01 g41410 ( .a(n8576), .b(n5973), .o(n45202) );
no02f01 g41411 ( .a(n8582), .b(n45202), .o(n45203) );
na02f01 g41412 ( .a(n45203), .b(n45201), .o(n45204) );
in01f01 g41413 ( .a(n45201), .o(n45205) );
in01f01 g41414 ( .a(n45203), .o(n45206) );
na02f01 g41415 ( .a(n45206), .b(n45205), .o(n45207) );
na02f01 g41416 ( .a(n45207), .b(n45204), .o(n3732) );
ao12f01 g41417 ( .a(n38323), .b(n38436), .c(n39827), .o(n45209) );
no02f01 g41418 ( .a(n38309), .b(n39081), .o(n45210) );
na02f01 g41419 ( .a(n45210), .b(n45209), .o(n45211) );
in01f01 g41420 ( .a(n45209), .o(n45212) );
in01f01 g41421 ( .a(n45210), .o(n45213) );
na02f01 g41422 ( .a(n45213), .b(n45212), .o(n45214) );
na02f01 g41423 ( .a(n45214), .b(n45211), .o(n3737) );
in01f01 g41424 ( .a(n44448), .o(n45216) );
ao12f01 g41425 ( .a(n44447), .b(n45216), .c(n44445), .o(n45217) );
no02f01 g41426 ( .a(n36141), .b(n36038), .o(n45218) );
no02f01 g41427 ( .a(n36140), .b(n36122), .o(n45219) );
no02f01 g41428 ( .a(n45219), .b(n45218), .o(n45220) );
na02f01 g41429 ( .a(n45220), .b(n45217), .o(n45221) );
in01f01 g41430 ( .a(n45217), .o(n45222) );
in01f01 g41431 ( .a(n45220), .o(n45223) );
na02f01 g41432 ( .a(n45223), .b(n45222), .o(n45224) );
na02f01 g41433 ( .a(n45224), .b(n45221), .o(n3742) );
na03f01 g41434 ( .a(n38432), .b(n38426), .c(n38409), .o(n45226) );
oa12f01 g41435 ( .a(n39113), .b(n38433), .c(n38427), .o(n45227) );
na02f01 g41436 ( .a(n45227), .b(n45226), .o(n3752) );
no02f01 g41437 ( .a(n39135), .b(n31485), .o(n45229) );
no02f01 g41438 ( .a(n45229), .b(n39138), .o(n45230) );
in01f01 g41439 ( .a(n39139), .o(n45231) );
na02f01 g41440 ( .a(n45231), .b(n43295), .o(n45232) );
no02f01 g41441 ( .a(n43297), .b(n39154), .o(n45233) );
na03f01 g41442 ( .a(n45233), .b(n45232), .c(n45230), .o(n45234) );
in01f01 g41443 ( .a(n45230), .o(n45235) );
na02f01 g41444 ( .a(n44211), .b(n39166), .o(n45236) );
oa12f01 g41445 ( .a(n45233), .b(n39139), .c(n45236), .o(n45237) );
na02f01 g41446 ( .a(n45237), .b(n45235), .o(n45238) );
na03f01 g41447 ( .a(n45238), .b(n45234), .c(n3633), .o(n45239) );
na02f01 g41448 ( .a(n45238), .b(n45234), .o(n4141) );
na02f01 g41449 ( .a(n4141), .b(n6203), .o(n45241) );
na02f01 g41450 ( .a(n45241), .b(n45239), .o(n3757) );
no02f01 g41451 ( .a(n27115), .b(n27243), .o(n45243) );
ao12f01 g41452 ( .a(n27114), .b(n27098), .c(n43871), .o(n45244) );
na02f01 g41453 ( .a(n45244), .b(n45243), .o(n45245) );
in01f01 g41454 ( .a(n45243), .o(n45246) );
in01f01 g41455 ( .a(n45244), .o(n45247) );
na02f01 g41456 ( .a(n45247), .b(n45246), .o(n45248) );
na02f01 g41457 ( .a(n45248), .b(n45245), .o(n3762) );
no02f01 g41458 ( .a(n41443), .b(n41442), .o(n45250) );
na02f01 g41459 ( .a(n45250), .b(n16236), .o(n45251) );
in01f01 g41460 ( .a(n45250), .o(n45252) );
na02f01 g41461 ( .a(n45252), .b(n21371), .o(n45253) );
na02f01 g41462 ( .a(n45253), .b(n45251), .o(n3767) );
no04f01 g41463 ( .a(n44165), .b(n21559), .c(n21475), .d(n21428), .o(n45255) );
na02f01 g41464 ( .a(n44171), .b(n21593), .o(n45256) );
no02f01 g41465 ( .a(n27291), .b(n16329), .o(n45257) );
no02f01 g41466 ( .a(n45257), .b(n44166), .o(n45258) );
in01f01 g41467 ( .a(n45258), .o(n45259) );
oa12f01 g41468 ( .a(n45259), .b(n45256), .c(n45255), .o(n45260) );
na04f01 g41469 ( .a(n44164), .b(n21558), .c(n21474), .d(n21615), .o(n45261) );
in01f01 g41470 ( .a(n45256), .o(n45262) );
na03f01 g41471 ( .a(n45258), .b(n45262), .c(n45261), .o(n45263) );
na03f01 g41472 ( .a(n45263), .b(n45260), .c(delay_sub_ln23_0_unr27_stage10_stallmux_z), .o(n45264) );
ao12f01 g41473 ( .a(n45258), .b(n45262), .c(n45261), .o(n45265) );
no03f01 g41474 ( .a(n45259), .b(n45256), .c(n45255), .o(n45266) );
oa12f01 g41475 ( .a(n21621), .b(n45266), .c(n45265), .o(n45267) );
na02f01 g41476 ( .a(n45267), .b(n45264), .o(n3772) );
no03f01 g41477 ( .a(n43737), .b(n43736), .c(n40322), .o(n45269) );
ao12f01 g41478 ( .a(n43732), .b(n43734), .c(n43729), .o(n45270) );
oa12f01 g41479 ( .a(n34420), .b(n45270), .c(n45269), .o(n45271) );
na03f01 g41480 ( .a(n43738), .b(n43735), .c(n_27923), .o(n45272) );
na02f01 g41481 ( .a(n45272), .b(n45271), .o(n3777) );
in01f01 g41482 ( .a(n29807), .o(n45274) );
in01f01 g41483 ( .a(n29808), .o(n45275) );
na03f01 g41484 ( .a(n45275), .b(n45274), .c(n29798), .o(n45276) );
in01f01 g41485 ( .a(n29798), .o(n45277) );
oa12f01 g41486 ( .a(n29807), .b(n29808), .c(n45277), .o(n45278) );
na02f01 g41487 ( .a(n45278), .b(n45276), .o(n3787) );
no02f01 g41488 ( .a(n11638), .b(n11590), .o(n45280) );
na02f01 g41489 ( .a(n45280), .b(n11636), .o(n45281) );
in01f01 g41490 ( .a(n45280), .o(n45282) );
na03f01 g41491 ( .a(n45282), .b(n11635), .c(n11599), .o(n45283) );
na02f01 g41492 ( .a(n45283), .b(n45281), .o(n3792) );
no02f01 g41493 ( .a(n25442), .b(n25434), .o(n45285) );
no03f01 g41494 ( .a(n25441), .b(n25440), .c(n25433), .o(n45286) );
oa12f01 g41495 ( .a(n25426), .b(n45286), .c(n45285), .o(n45287) );
in01f01 g41496 ( .a(n25426), .o(n45288) );
no02f01 g41497 ( .a(n45286), .b(n45285), .o(n45289) );
na02f01 g41498 ( .a(n45289), .b(n45288), .o(n45290) );
na02f01 g41499 ( .a(n45290), .b(n45287), .o(n3797) );
na02f01 g41500 ( .a(n32732), .b(cos_out_5), .o(n45292) );
no02f01 g41501 ( .a(n36239), .b(n35944), .o(n45293) );
no02f01 g41502 ( .a(n45293), .b(n36241), .o(n45294) );
in01f01 g41503 ( .a(n45294), .o(n45295) );
no03f01 g41504 ( .a(n45295), .b(n43152), .c(n35966), .o(n45296) );
no02f01 g41505 ( .a(n43152), .b(n35966), .o(n45297) );
no02f01 g41506 ( .a(n45294), .b(n45297), .o(n45298) );
oa12f01 g41507 ( .a(n32734), .b(n45298), .c(n45296), .o(n45299) );
na02f01 g41508 ( .a(n45299), .b(n45292), .o(n3802) );
no02f01 g41509 ( .a(n30035), .b(n30027), .o(n45301) );
no02f01 g41510 ( .a(n45301), .b(n30128), .o(n45302) );
na02f01 g41511 ( .a(n45301), .b(n30128), .o(n45303) );
in01f01 g41512 ( .a(n45303), .o(n45304) );
no02f01 g41513 ( .a(n45304), .b(n45302), .o(n45305) );
na02f01 g41514 ( .a(n45305), .b(n6037), .o(n45306) );
in01f01 g41515 ( .a(n45305), .o(n4558) );
na02f01 g41516 ( .a(n4558), .b(n5873), .o(n45308) );
na02f01 g41517 ( .a(n45308), .b(n45306), .o(n3806) );
no02f01 g41518 ( .a(n42442), .b(n42441), .o(n45310) );
na03f01 g41519 ( .a(n3426), .b(n45310), .c(delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(n45311) );
in01f01 g41520 ( .a(n45310), .o(n4883) );
oa12f01 g41521 ( .a(n4883), .b(n44842), .c(n37149), .o(n45313) );
na02f01 g41522 ( .a(n45313), .b(n45311), .o(n3811) );
no02f01 g41523 ( .a(n39016), .b(n25277), .o(n45315) );
no02f01 g41524 ( .a(n25264), .b(n25261), .o(n45316) );
na02f01 g41525 ( .a(n45316), .b(n45315), .o(n45317) );
no02f01 g41526 ( .a(n45316), .b(n45315), .o(n45318) );
in01f01 g41527 ( .a(n45318), .o(n45319) );
na03f01 g41528 ( .a(n45319), .b(n45317), .c(n6037), .o(n45320) );
na02f01 g41529 ( .a(n45319), .b(n45317), .o(n4196) );
na02f01 g41530 ( .a(n4196), .b(n5873), .o(n45322) );
na02f01 g41531 ( .a(n45322), .b(n45320), .o(n3816) );
in01f01 g41532 ( .a(n41042), .o(n45324) );
no02f01 g41533 ( .a(n41044), .b(n38708), .o(n45325) );
na03f01 g41534 ( .a(n45325), .b(n38717), .c(n45324), .o(n45326) );
in01f01 g41535 ( .a(n38717), .o(n45327) );
in01f01 g41536 ( .a(n45325), .o(n45328) );
oa12f01 g41537 ( .a(n45328), .b(n45327), .c(n41042), .o(n45329) );
na02f01 g41538 ( .a(n45329), .b(n45326), .o(n3821) );
na02f01 g41539 ( .a(n36512), .b(n36510), .o(n45331) );
in01f01 g41540 ( .a(n45331), .o(n45332) );
na02f01 g41541 ( .a(n45332), .b(n36509), .o(n45333) );
na02f01 g41542 ( .a(n45331), .b(n36485), .o(n45334) );
na02f01 g41543 ( .a(n45334), .b(n45333), .o(n3826) );
in01f01 g41544 ( .a(n44213), .o(n45336) );
ao12f01 g41545 ( .a(n44212), .b(n45336), .c(n44211), .o(n45337) );
no02f01 g41546 ( .a(n39135), .b(n32243), .o(n45338) );
no02f01 g41547 ( .a(n39059), .b(n31474), .o(n45339) );
no02f01 g41548 ( .a(n45339), .b(n45338), .o(n45340) );
na02f01 g41549 ( .a(n45340), .b(n45337), .o(n45341) );
in01f01 g41550 ( .a(n45337), .o(n45342) );
in01f01 g41551 ( .a(n45340), .o(n45343) );
na02f01 g41552 ( .a(n45343), .b(n45342), .o(n45344) );
na02f01 g41553 ( .a(n45344), .b(n45341), .o(n3831) );
in01f01 g41554 ( .a(n35589), .o(n45346) );
ao12f01 g41555 ( .a(n35588), .b(n45346), .c(n9436), .o(n45347) );
no02f01 g41556 ( .a(n9447), .b(n9225), .o(n45348) );
no02f01 g41557 ( .a(n9448), .b(n9224), .o(n45349) );
no02f01 g41558 ( .a(n45349), .b(n45348), .o(n45350) );
na02f01 g41559 ( .a(n45350), .b(n45347), .o(n45351) );
in01f01 g41560 ( .a(n45347), .o(n45352) );
in01f01 g41561 ( .a(n45350), .o(n45353) );
na02f01 g41562 ( .a(n45353), .b(n45352), .o(n45354) );
na02f01 g41563 ( .a(n45354), .b(n45351), .o(n3836) );
na02f01 g41564 ( .a(n32732), .b(cos_out_0), .o(n45356) );
ao12f01 g41565 ( .a(n35973), .b(n35972), .c(n35971), .o(n45357) );
oa12f01 g41566 ( .a(n32734), .b(n45357), .c(n35930), .o(n45358) );
na02f01 g41567 ( .a(n45358), .b(n45356), .o(n3846) );
no02f01 g41568 ( .a(n40034), .b(n39372), .o(n45360) );
oa12f01 g41569 ( .a(n45360), .b(n40038), .c(n39354), .o(n45361) );
in01f01 g41570 ( .a(n45360), .o(n45362) );
na03f01 g41571 ( .a(n39476), .b(n45362), .c(n39355), .o(n45363) );
na02f01 g41572 ( .a(n45363), .b(n45361), .o(n3850) );
no02f01 g41573 ( .a(n21259), .b(n21026), .o(n45365) );
in01f01 g41574 ( .a(n45365), .o(n45366) );
in01f01 g41575 ( .a(n21003), .o(n45367) );
no02f01 g41576 ( .a(n21260), .b(n45367), .o(n45368) );
no02f01 g41577 ( .a(n45368), .b(n45366), .o(n45369) );
na02f01 g41578 ( .a(n45368), .b(n45366), .o(n45370) );
in01f01 g41579 ( .a(n45370), .o(n45371) );
no02f01 g41580 ( .a(n45371), .b(n45369), .o(n45372) );
na02f01 g41581 ( .a(n45372), .b(n5799), .o(n45373) );
in01f01 g41582 ( .a(n45372), .o(n6081) );
na02f01 g41583 ( .a(n6081), .b(n911), .o(n45375) );
na02f01 g41584 ( .a(n45375), .b(n45373), .o(n3860) );
no02f01 g41585 ( .a(n29650), .b(n29636), .o(n45377) );
na03f01 g41586 ( .a(n45377), .b(n29645), .c(n29722), .o(n45378) );
in01f01 g41587 ( .a(n45377), .o(n45379) );
oa12f01 g41588 ( .a(n45379), .b(n29646), .c(n29616), .o(n45380) );
na02f01 g41589 ( .a(n45380), .b(n45378), .o(n3870) );
no02f01 g41590 ( .a(n36882), .b(n31607), .o(n45382) );
no02f01 g41591 ( .a(n45382), .b(n36862), .o(n45383) );
in01f01 g41592 ( .a(n45383), .o(n45384) );
na03f01 g41593 ( .a(n41651), .b(n41650), .c(n41652), .o(n45385) );
na03f01 g41594 ( .a(n45385), .b(n45384), .c(n36852), .o(n45386) );
no03f01 g41595 ( .a(n41657), .b(n41656), .c(n41653), .o(n45387) );
oa12f01 g41596 ( .a(n45383), .b(n45387), .c(n36851), .o(n45388) );
na03f01 g41597 ( .a(n45388), .b(n45386), .c(n3633), .o(n45389) );
no03f01 g41598 ( .a(n45387), .b(n45383), .c(n36851), .o(n45390) );
ao12f01 g41599 ( .a(n45384), .b(n45385), .c(n36852), .o(n45391) );
oa12f01 g41600 ( .a(n6203), .b(n45391), .c(n45390), .o(n45392) );
na02f01 g41601 ( .a(n45392), .b(n45389), .o(n3875) );
no02f01 g41602 ( .a(n35297), .b(n35258), .o(n45394) );
no02f01 g41603 ( .a(n35298), .b(n4176), .o(n45395) );
oa22f01 g41604 ( .a(n45395), .b(n45394), .c(n35300), .d(n35289), .o(n45396) );
no02f01 g41605 ( .a(n35300), .b(n35289), .o(n45397) );
no02f01 g41606 ( .a(n45395), .b(n45394), .o(n45398) );
na02f01 g41607 ( .a(n45398), .b(n45397), .o(n45399) );
na02f01 g41608 ( .a(n45399), .b(n45396), .o(n3880) );
no02f01 g41609 ( .a(n8544), .b(n42037), .o(n45401) );
no02f01 g41610 ( .a(n45401), .b(n8558), .o(n45402) );
no02f01 g41611 ( .a(n8559), .b(n8554), .o(n45403) );
na02f01 g41612 ( .a(n45403), .b(n45402), .o(n45404) );
in01f01 g41613 ( .a(n45403), .o(n45405) );
oa12f01 g41614 ( .a(n45405), .b(n45401), .c(n8558), .o(n45406) );
na02f01 g41615 ( .a(n45406), .b(n45404), .o(n3885) );
na03f01 g41616 ( .a(n43284), .b(n43279), .c(n5799), .o(n45408) );
ao12f01 g41617 ( .a(n43281), .b(n43283), .c(n43280), .o(n45409) );
no03f01 g41618 ( .a(n43278), .b(n43277), .c(n41386), .o(n45410) );
oa12f01 g41619 ( .a(n911), .b(n45410), .c(n45409), .o(n45411) );
na02f01 g41620 ( .a(n45411), .b(n45408), .o(n3890) );
ao12f01 g41621 ( .a(n43560), .b(n43562), .c(n43566), .o(n45413) );
in01f01 g41622 ( .a(n45413), .o(n45414) );
in01f01 g41623 ( .a(n9688), .o(n45415) );
no02f01 g41624 ( .a(n45415), .b(n6934), .o(n45416) );
no02f01 g41625 ( .a(n9688), .b(n5001), .o(n45417) );
no02f01 g41626 ( .a(n45417), .b(n45416), .o(n45418) );
in01f01 g41627 ( .a(n45418), .o(n45419) );
na02f01 g41628 ( .a(n45419), .b(n45414), .o(n45420) );
na02f01 g41629 ( .a(n45418), .b(n45413), .o(n45421) );
na02f01 g41630 ( .a(n45421), .b(n45420), .o(n3895) );
no02f01 g41631 ( .a(n40791), .b(n21265), .o(n45423) );
na02f01 g41632 ( .a(n40791), .b(n21265), .o(n45424) );
in01f01 g41633 ( .a(n45424), .o(n45425) );
no02f01 g41634 ( .a(n45425), .b(n45423), .o(n45426) );
no02f01 g41635 ( .a(n41200), .b(n41180), .o(n45427) );
na02f01 g41636 ( .a(n45427), .b(n41193), .o(n45428) );
oa12f01 g41637 ( .a(n40794), .b(n41183), .c(n20360), .o(n45429) );
na02f01 g41638 ( .a(n45429), .b(n41196), .o(n45430) );
in01f01 g41639 ( .a(n45430), .o(n45431) );
na03f01 g41640 ( .a(n45431), .b(n45428), .c(n45426), .o(n45432) );
in01f01 g41641 ( .a(n45426), .o(n45433) );
no03f01 g41642 ( .a(n41200), .b(n41209), .c(n41180), .o(n45434) );
oa12f01 g41643 ( .a(n45433), .b(n45430), .c(n45434), .o(n45435) );
na02f01 g41644 ( .a(n45435), .b(n45432), .o(n3900) );
in01f01 g41645 ( .a(n43264), .o(n45437) );
no02f01 g41646 ( .a(n36432), .b(n21835), .o(n45438) );
no02f01 g41647 ( .a(n36447), .b(n22376), .o(n45439) );
no02f01 g41648 ( .a(n45439), .b(n45438), .o(n45440) );
in01f01 g41649 ( .a(n45440), .o(n45441) );
in01f01 g41650 ( .a(n43263), .o(n45442) );
na03f01 g41651 ( .a(n43262), .b(n43261), .c(n45442), .o(n45443) );
ao12f01 g41652 ( .a(n45441), .b(n45443), .c(n45437), .o(n45444) );
no03f01 g41653 ( .a(n43268), .b(n43267), .c(n43263), .o(n45445) );
no03f01 g41654 ( .a(n45445), .b(n45440), .c(n43264), .o(n45446) );
oa12f01 g41655 ( .a(n4116), .b(n45446), .c(n45444), .o(n45447) );
oa12f01 g41656 ( .a(n45440), .b(n45445), .c(n43264), .o(n45448) );
na03f01 g41657 ( .a(n45443), .b(n45441), .c(n45437), .o(n45449) );
na03f01 g41658 ( .a(n45449), .b(n45448), .c(n2589), .o(n45450) );
na02f01 g41659 ( .a(n45450), .b(n45447), .o(n3905) );
no02f01 g41660 ( .a(n9600), .b(n9599), .o(n45452) );
no03f01 g41661 ( .a(n41455), .b(n45452), .c(n9591), .o(n45453) );
no02f01 g41662 ( .a(n41455), .b(n45452), .o(n45454) );
no02f01 g41663 ( .a(n45454), .b(n4201), .o(n45455) );
no02f01 g41664 ( .a(n45455), .b(n45453), .o(n45456) );
in01f01 g41665 ( .a(n45456), .o(n3910) );
no02f01 g41666 ( .a(n42696), .b(n41379), .o(n45458) );
na03f01 g41667 ( .a(n45458), .b(n42703), .c(n42702), .o(n45459) );
in01f01 g41668 ( .a(n45458), .o(n45460) );
oa12f01 g41669 ( .a(n45460), .b(n42697), .c(n41384), .o(n45461) );
na03f01 g41670 ( .a(n45461), .b(n45459), .c(n5799), .o(n45462) );
na02f01 g41671 ( .a(n45461), .b(n45459), .o(n4424) );
na02f01 g41672 ( .a(n4424), .b(n911), .o(n45464) );
na02f01 g41673 ( .a(n45464), .b(n45462), .o(n3915) );
in01f01 g41674 ( .a(n8440), .o(n45466) );
no02f01 g41675 ( .a(n43570), .b(n8450), .o(n45467) );
in01f01 g41676 ( .a(n45467), .o(n45468) );
oa12f01 g41677 ( .a(n45468), .b(n8441), .c(n45466), .o(n45469) );
na03f01 g41678 ( .a(n45467), .b(n8442), .c(n8440), .o(n45470) );
na02f01 g41679 ( .a(n45470), .b(n45469), .o(n3920) );
na04f01 g41680 ( .a(n32386), .b(n32385), .c(n32235), .d(n32224), .o(n45472) );
oa22f01 g41681 ( .a(n32479), .b(n32223), .c(n32477), .d(n32234), .o(n45473) );
na02f01 g41682 ( .a(n45473), .b(n45472), .o(n3925) );
na02f01 g41683 ( .a(n742), .b(n4116), .o(n45475) );
na02f01 g41684 ( .a(n39037), .b(n2589), .o(n45476) );
na02f01 g41685 ( .a(n45476), .b(n45475), .o(n3930) );
no02f01 g41686 ( .a(n14235), .b(n13960), .o(n45478) );
in01f01 g41687 ( .a(n45478), .o(n45479) );
no02f01 g41688 ( .a(n45479), .b(n14232), .o(n45480) );
no02f01 g41689 ( .a(n45478), .b(n41154), .o(n45481) );
no02f01 g41690 ( .a(n45481), .b(n45480), .o(n45482) );
in01f01 g41691 ( .a(n45482), .o(n5080) );
na02f01 g41692 ( .a(n5080), .b(n4116), .o(n45484) );
na02f01 g41693 ( .a(n45482), .b(n2589), .o(n45485) );
na02f01 g41694 ( .a(n45485), .b(n45484), .o(n3940) );
na03f01 g41695 ( .a(n40329), .b(n40325), .c(n_27923), .o(n45487) );
na02f01 g41696 ( .a(n996), .b(n34420), .o(n45488) );
na02f01 g41697 ( .a(n45488), .b(n45487), .o(n3945) );
na03f01 g41698 ( .a(n41107), .b(n9590), .c(n9589), .o(n45490) );
oa12f01 g41699 ( .a(n1255), .b(n9646), .c(n9645), .o(n45491) );
na02f01 g41700 ( .a(n45491), .b(n45490), .o(n3950) );
in01f01 g41701 ( .a(n16284), .o(n45493) );
no02f01 g41702 ( .a(n16302), .b(n16236), .o(n45494) );
na02f01 g41703 ( .a(n16283), .b(n16155), .o(n45495) );
na02f01 g41704 ( .a(n45495), .b(n16433), .o(n45496) );
ao12f01 g41705 ( .a(n45496), .b(n45494), .c(n45493), .o(n45497) );
no02f01 g41706 ( .a(n16322), .b(n16329), .o(n45498) );
no02f01 g41707 ( .a(n45498), .b(n16324), .o(n45499) );
na02f01 g41708 ( .a(n45499), .b(n45497), .o(n45500) );
in01f01 g41709 ( .a(n45497), .o(n45501) );
in01f01 g41710 ( .a(n45499), .o(n45502) );
na02f01 g41711 ( .a(n45502), .b(n45501), .o(n45503) );
na02f01 g41712 ( .a(n45503), .b(n45500), .o(n3955) );
in01f01 g41713 ( .a(n21339), .o(n45505) );
no02f01 g41714 ( .a(n16356), .b(n45505), .o(n45506) );
no03f01 g41715 ( .a(n45506), .b(n21341), .c(n16435), .o(n45507) );
no02f01 g41716 ( .a(n16377), .b(n16329), .o(n45508) );
no02f01 g41717 ( .a(n45508), .b(n16379), .o(n45509) );
na02f01 g41718 ( .a(n45509), .b(n45507), .o(n45510) );
in01f01 g41719 ( .a(n45507), .o(n45511) );
in01f01 g41720 ( .a(n45509), .o(n45512) );
na02f01 g41721 ( .a(n45512), .b(n45511), .o(n45513) );
na02f01 g41722 ( .a(n45513), .b(n45510), .o(n3960) );
no02f01 g41723 ( .a(n42583), .b(n39976), .o(n45515) );
na03f01 g41724 ( .a(n45515), .b(n39989), .c(n42588), .o(n45516) );
in01f01 g41725 ( .a(n45515), .o(n45517) );
oa12f01 g41726 ( .a(n45517), .b(n42582), .c(n42579), .o(n45518) );
na02f01 g41727 ( .a(n45518), .b(n45516), .o(n3965) );
na03f01 g41728 ( .a(n25850), .b(n25827), .c(n30080), .o(n45520) );
oa12f01 g41729 ( .a(n25851), .b(n30081), .c(n25826), .o(n45521) );
na02f01 g41730 ( .a(n45521), .b(n45520), .o(n3970) );
na02f01 g41731 ( .a(n41878), .b(n41874), .o(n3975) );
no02f01 g41732 ( .a(n9623), .b(n9336), .o(n45524) );
in01f01 g41733 ( .a(n45524), .o(n45525) );
oa12f01 g41734 ( .a(n45525), .b(n9401), .c(n9397), .o(n45526) );
na03f01 g41735 ( .a(n45524), .b(n9400), .c(n9622), .o(n45527) );
na02f01 g41736 ( .a(n45527), .b(n45526), .o(n3980) );
na03f01 g41737 ( .a(n32678), .b(n32720), .c(n32694), .o(n45529) );
oa12f01 g41738 ( .a(n32677), .b(n32724), .c(n32598), .o(n45530) );
na02f01 g41739 ( .a(n45530), .b(n45529), .o(n3985) );
no02f01 g41740 ( .a(n36887), .b(n36840), .o(n45532) );
na03f01 g41741 ( .a(n45532), .b(n36886), .c(n36876), .o(n45533) );
in01f01 g41742 ( .a(n45532), .o(n45534) );
oa12f01 g41743 ( .a(n45534), .b(n36885), .c(n36891), .o(n45535) );
na02f01 g41744 ( .a(n45535), .b(n45533), .o(n3990) );
in01f01 g41745 ( .a(n39435), .o(n45537) );
in01f01 g41746 ( .a(n39436), .o(n45538) );
oa12f01 g41747 ( .a(n39440), .b(n45538), .c(n45537), .o(n45539) );
na03f01 g41748 ( .a(n39439), .b(n39436), .c(n39435), .o(n45540) );
na02f01 g41749 ( .a(n45540), .b(n45539), .o(n3999) );
no02f01 g41750 ( .a(n16515), .b(n16489), .o(n45542) );
no02f01 g41751 ( .a(n16516), .b(n16512), .o(n45543) );
na02f01 g41752 ( .a(n45543), .b(n45542), .o(n45544) );
in01f01 g41753 ( .a(n45543), .o(n45545) );
oa12f01 g41754 ( .a(n45545), .b(n16515), .c(n16489), .o(n45546) );
na02f01 g41755 ( .a(n45546), .b(n45544), .o(n4004) );
na02f01 g41756 ( .a(n971), .b(n37149), .o(n45548) );
na03f01 g41757 ( .a(n45548), .b(n37361), .c(n37313), .o(n45549) );
na02f01 g41758 ( .a(n45548), .b(n37361), .o(n45550) );
na02f01 g41759 ( .a(n45550), .b(n37358), .o(n45551) );
na02f01 g41760 ( .a(n45551), .b(n45549), .o(n4009) );
no02f01 g41761 ( .a(n29937), .b(n24273), .o(n45553) );
in01f01 g41762 ( .a(n24273), .o(n45554) );
no02f01 g41763 ( .a(n29938), .b(n45554), .o(n45555) );
no02f01 g41764 ( .a(n45555), .b(n45553), .o(n45556) );
no02f01 g41765 ( .a(n40059), .b(n40052), .o(n45557) );
na02f01 g41766 ( .a(n45557), .b(n30134), .o(n45558) );
ao12f01 g41767 ( .a(n29937), .b(n40057), .c(n24608), .o(n45559) );
no02f01 g41768 ( .a(n45559), .b(n30046), .o(n45560) );
na03f01 g41769 ( .a(n45560), .b(n45558), .c(n45556), .o(n45561) );
in01f01 g41770 ( .a(n45556), .o(n45562) );
no03f01 g41771 ( .a(n40059), .b(n40052), .c(n30042), .o(n45563) );
in01f01 g41772 ( .a(n45560), .o(n45564) );
oa12f01 g41773 ( .a(n45562), .b(n45564), .c(n45563), .o(n45565) );
na02f01 g41774 ( .a(n45565), .b(n45561), .o(n4014) );
na03f01 g41775 ( .a(n43259), .b(n43257), .c(n3633), .o(n45567) );
na02f01 g41776 ( .a(n2317), .b(n6203), .o(n45568) );
na02f01 g41777 ( .a(n45568), .b(n45567), .o(n4019) );
na02f01 g41778 ( .a(n32732), .b(cos_out_10), .o(n45570) );
no02f01 g41779 ( .a(n44252), .b(n36313), .o(n45571) );
in01f01 g41780 ( .a(n45571), .o(n45572) );
no03f01 g41781 ( .a(n45572), .b(n44249), .c(n36367), .o(n45573) );
ao12f01 g41782 ( .a(n45571), .b(n44250), .c(n44254), .o(n45574) );
oa12f01 g41783 ( .a(n32734), .b(n45574), .c(n45573), .o(n45575) );
na02f01 g41784 ( .a(n45575), .b(n45570), .o(n4024) );
no02f01 g41785 ( .a(n38020), .b(n37902), .o(n45577) );
in01f01 g41786 ( .a(n45577), .o(n45578) );
no03f01 g41787 ( .a(n45578), .b(n43379), .c(n38024), .o(n45579) );
no02f01 g41788 ( .a(n43379), .b(n38024), .o(n45580) );
no02f01 g41789 ( .a(n45577), .b(n45580), .o(n45581) );
no02f01 g41790 ( .a(n45581), .b(n45579), .o(n45582) );
in01f01 g41791 ( .a(n45582), .o(n4028) );
na03f01 g41792 ( .a(n36526), .b(n36524), .c(n6037), .o(n45584) );
in01f01 g41793 ( .a(n36524), .o(n45585) );
oa12f01 g41794 ( .a(n5873), .b(n36525), .c(n45585), .o(n45586) );
na02f01 g41795 ( .a(n45586), .b(n45584), .o(n4033) );
in01f01 g41796 ( .a(n40958), .o(n45588) );
no02f01 g41797 ( .a(n40956), .b(n6044), .o(n45589) );
in01f01 g41798 ( .a(n45589), .o(n45590) );
na02f01 g41799 ( .a(n45590), .b(n45588), .o(n45591) );
na02f01 g41800 ( .a(n45589), .b(n40958), .o(n45592) );
na02f01 g41801 ( .a(n45592), .b(n45591), .o(n4038) );
no02f01 g41802 ( .a(n41416), .b(n41414), .o(n4048) );
ao12f01 g41803 ( .a(n9602), .b(n45452), .c(n44198), .o(n45595) );
no02f01 g41804 ( .a(n45595), .b(n9226), .o(n45596) );
no03f01 g41805 ( .a(n45596), .b(n9591), .c(n9227), .o(n45597) );
no02f01 g41806 ( .a(n45596), .b(n9227), .o(n45598) );
no02f01 g41807 ( .a(n45598), .b(n4201), .o(n45599) );
no02f01 g41808 ( .a(n45599), .b(n45597), .o(n45600) );
in01f01 g41809 ( .a(n45600), .o(n4053) );
na02f01 g41810 ( .a(n44944), .b(n2589), .o(n45602) );
na02f01 g41811 ( .a(n3526), .b(n4116), .o(n45603) );
na02f01 g41812 ( .a(n45603), .b(n45602), .o(n4058) );
oa12f01 g41813 ( .a(n27233), .b(n27042), .c(n26917), .o(n45605) );
na03f01 g41814 ( .a(n27041), .b(n27040), .c(n26918), .o(n45606) );
na02f01 g41815 ( .a(n45606), .b(n45605), .o(n4063) );
ao12f01 g41816 ( .a(n38541), .b(n39133), .c(n38511), .o(n45608) );
no02f01 g41817 ( .a(n39073), .b(n39135), .o(n45609) );
no02f01 g41818 ( .a(n45609), .b(n39075), .o(n45610) );
in01f01 g41819 ( .a(n45610), .o(n45611) );
na02f01 g41820 ( .a(n45611), .b(n45608), .o(n45612) );
in01f01 g41821 ( .a(n45608), .o(n45613) );
na02f01 g41822 ( .a(n45610), .b(n45613), .o(n45614) );
na02f01 g41823 ( .a(n45614), .b(n45612), .o(n4068) );
in01f01 g41824 ( .a(n10913), .o(n45616) );
no02f01 g41825 ( .a(n45616), .b(n25629), .o(n45617) );
no03f01 g41826 ( .a(n10926), .b(n25632), .c(n45617), .o(n45618) );
no02f01 g41827 ( .a(n10920), .b(n3521), .o(n45619) );
no02f01 g41828 ( .a(n45619), .b(n10922), .o(n45620) );
na02f01 g41829 ( .a(n45620), .b(n45618), .o(n45621) );
in01f01 g41830 ( .a(n45618), .o(n45622) );
in01f01 g41831 ( .a(n45620), .o(n45623) );
na02f01 g41832 ( .a(n45623), .b(n45622), .o(n45624) );
na02f01 g41833 ( .a(n45624), .b(n45621), .o(n4073) );
no02f01 g41834 ( .a(n38189), .b(n22347), .o(n45626) );
no02f01 g41835 ( .a(n45626), .b(n22356), .o(n45627) );
na02f01 g41836 ( .a(n22350), .b(n22340), .o(n45628) );
in01f01 g41837 ( .a(n45628), .o(n45629) );
no02f01 g41838 ( .a(n45629), .b(n45627), .o(n45630) );
na02f01 g41839 ( .a(n45629), .b(n45627), .o(n45631) );
in01f01 g41840 ( .a(n45631), .o(n45632) );
no02f01 g41841 ( .a(n45632), .b(n45630), .o(n45633) );
in01f01 g41842 ( .a(n45633), .o(n5648) );
na02f01 g41843 ( .a(n5648), .b(n4116), .o(n45635) );
na02f01 g41844 ( .a(n45633), .b(n2589), .o(n45636) );
na02f01 g41845 ( .a(n45636), .b(n45635), .o(n4078) );
in01f01 g41846 ( .a(n11631), .o(n45638) );
no02f01 g41847 ( .a(n45638), .b(n11606), .o(n45639) );
na02f01 g41848 ( .a(n45639), .b(n11629), .o(n45640) );
in01f01 g41849 ( .a(n45639), .o(n45641) );
na02f01 g41850 ( .a(n45641), .b(n11630), .o(n45642) );
na02f01 g41851 ( .a(n45642), .b(n45640), .o(n4083) );
ao12f01 g41852 ( .a(n37994), .b(n38000), .c(n43892), .o(n45644) );
no02f01 g41853 ( .a(n37999), .b(n37925), .o(n45645) );
in01f01 g41854 ( .a(n45645), .o(n45646) );
no02f01 g41855 ( .a(n45646), .b(n45644), .o(n45647) );
na02f01 g41856 ( .a(n45646), .b(n45644), .o(n45648) );
in01f01 g41857 ( .a(n45648), .o(n45649) );
no02f01 g41858 ( .a(n45649), .b(n45647), .o(n45650) );
na02f01 g41859 ( .a(n45650), .b(n1821), .o(n45651) );
in01f01 g41860 ( .a(n45650), .o(n5603) );
na02f01 g41861 ( .a(n5603), .b(n8066), .o(n45653) );
na02f01 g41862 ( .a(n45653), .b(n45651), .o(n4093) );
na02f01 g41863 ( .a(n32732), .b(sin_out_13), .o(n45655) );
no02f01 g41864 ( .a(n39512), .b(n39499), .o(n45656) );
oa12f01 g41865 ( .a(n45656), .b(n39511), .c(n39516), .o(n45657) );
no02f01 g41866 ( .a(n39592), .b(n34307), .o(n45658) );
no02f01 g41867 ( .a(n45658), .b(n39564), .o(n45659) );
in01f01 g41868 ( .a(n45659), .o(n45660) );
no02f01 g41869 ( .a(n45660), .b(n45657), .o(n45661) );
in01f01 g41870 ( .a(n45657), .o(n45662) );
no02f01 g41871 ( .a(n45659), .b(n45662), .o(n45663) );
oa12f01 g41872 ( .a(n32734), .b(n45663), .c(n45661), .o(n45664) );
na02f01 g41873 ( .a(n45664), .b(n45655), .o(n4103) );
na02f01 g41874 ( .a(n11651), .b(n11649), .o(n45666) );
oa12f01 g41875 ( .a(n45666), .b(n11639), .c(n11590), .o(n45667) );
in01f01 g41876 ( .a(n45666), .o(n45668) );
na02f01 g41877 ( .a(n45668), .b(n11640), .o(n45669) );
na02f01 g41878 ( .a(n45669), .b(n45667), .o(n4107) );
na02f01 g41879 ( .a(n32732), .b(cos_out_3), .o(n45671) );
in01f01 g41880 ( .a(n35953), .o(n45672) );
no02f01 g41881 ( .a(n35952), .b(n35944), .o(n45673) );
no02f01 g41882 ( .a(n45673), .b(n45672), .o(n45674) );
in01f01 g41883 ( .a(n45674), .o(n45675) );
no03f01 g41884 ( .a(n45675), .b(n41428), .c(n35977), .o(n45676) );
no02f01 g41885 ( .a(n41428), .b(n35977), .o(n45677) );
no02f01 g41886 ( .a(n45674), .b(n45677), .o(n45678) );
oa12f01 g41887 ( .a(n32734), .b(n45678), .c(n45676), .o(n45679) );
na02f01 g41888 ( .a(n45679), .b(n45671), .o(n4112) );
no02f01 g41889 ( .a(n42045), .b(n37194), .o(n45681) );
no03f01 g41890 ( .a(n45681), .b(n42046), .c(n37250), .o(n45682) );
no02f01 g41891 ( .a(n37204), .b(n36963), .o(n45683) );
no02f01 g41892 ( .a(n45683), .b(n37206), .o(n45684) );
na02f01 g41893 ( .a(n45684), .b(n45682), .o(n45685) );
in01f01 g41894 ( .a(n45682), .o(n45686) );
in01f01 g41895 ( .a(n45684), .o(n45687) );
na02f01 g41896 ( .a(n45687), .b(n45686), .o(n45688) );
na02f01 g41897 ( .a(n45688), .b(n45685), .o(n4121) );
in01f01 g41898 ( .a(n9768), .o(n45690) );
in01f01 g41899 ( .a(n42269), .o(n45691) );
na02f01 g41900 ( .a(n42268), .b(n45691), .o(n45692) );
ao12f01 g41901 ( .a(n45692), .b(n45690), .c(n42266), .o(n45693) );
no02f01 g41902 ( .a(n9757), .b(n5001), .o(n45694) );
no02f01 g41903 ( .a(n45694), .b(n9759), .o(n45695) );
na02f01 g41904 ( .a(n45695), .b(n45693), .o(n45696) );
in01f01 g41905 ( .a(n45693), .o(n45697) );
in01f01 g41906 ( .a(n45695), .o(n45698) );
na02f01 g41907 ( .a(n45698), .b(n45697), .o(n45699) );
na02f01 g41908 ( .a(n45699), .b(n45696), .o(n4131) );
na02f01 g41909 ( .a(n42571), .b(n5799), .o(n45701) );
na02f01 g41910 ( .a(n1914), .b(n911), .o(n45702) );
na02f01 g41911 ( .a(n45702), .b(n45701), .o(n4136) );
na03f01 g41912 ( .a(n40416), .b(n9590), .c(n9589), .o(n45704) );
oa12f01 g41913 ( .a(n1050), .b(n9646), .c(n9645), .o(n45705) );
na02f01 g41914 ( .a(n45705), .b(n45704), .o(n4146) );
oa12f01 g41915 ( .a(n32681), .b(n32728), .c(n32577), .o(n45707) );
na03f01 g41916 ( .a(n32682), .b(n32727), .c(n32690), .o(n45708) );
na02f01 g41917 ( .a(n45708), .b(n45707), .o(n4151) );
na02f01 g41918 ( .a(n1090), .b(n4116), .o(n45710) );
na03f01 g41919 ( .a(n40474), .b(n40473), .c(n2589), .o(n45711) );
na02f01 g41920 ( .a(n45711), .b(n45710), .o(n4161) );
na03f01 g41921 ( .a(n45456), .b(n9590), .c(n9589), .o(n45713) );
oa12f01 g41922 ( .a(n3910), .b(n9646), .c(n9645), .o(n45714) );
na02f01 g41923 ( .a(n45714), .b(n45713), .o(n4166) );
no02f01 g41924 ( .a(n14237), .b(n13926), .o(n45716) );
in01f01 g41925 ( .a(n45716), .o(n45717) );
no02f01 g41926 ( .a(n45717), .b(n44626), .o(n45718) );
no02f01 g41927 ( .a(n45716), .b(n44625), .o(n45719) );
no02f01 g41928 ( .a(n45719), .b(n45718), .o(n45720) );
in01f01 g41929 ( .a(n45720), .o(n4171) );
na02f01 g41930 ( .a(n44046), .b(n44044), .o(n4186) );
na02f01 g41931 ( .a(n42705), .b(n42699), .o(n4191) );
na03f01 g41932 ( .a(n45010), .b(n45008), .c(n_27923), .o(n45724) );
na02f01 g41933 ( .a(n3570), .b(n34420), .o(n45725) );
na02f01 g41934 ( .a(n45725), .b(n45724), .o(n4206) );
in01f01 g41935 ( .a(mux_while_ln12_psv_q_5_), .o(n45727) );
in01f01 g41936 ( .a(n4048), .o(n45728) );
no02f01 g41937 ( .a(n45728), .b(n45727), .o(n4211) );
na03f01 g41938 ( .a(n43804), .b(n9590), .c(n9589), .o(n45730) );
oa12f01 g41939 ( .a(n2707), .b(n9646), .c(n9645), .o(n45731) );
na02f01 g41940 ( .a(n45731), .b(n45730), .o(n4216) );
na02f01 g41941 ( .a(n44421), .b(n6037), .o(n45733) );
na02f01 g41942 ( .a(n3150), .b(n5873), .o(n45734) );
na02f01 g41943 ( .a(n45734), .b(n45733), .o(n4221) );
in01f01 g41944 ( .a(n5949), .o(n45736) );
no02f01 g41945 ( .a(n5950), .b(n45736), .o(n45737) );
na02f01 g41946 ( .a(n5962), .b(n45737), .o(n45738) );
in01f01 g41947 ( .a(n5959), .o(n45739) );
no02f01 g41948 ( .a(n45739), .b(n6037), .o(n45740) );
no02f01 g41949 ( .a(n5959), .b(n5873), .o(n45741) );
no02f01 g41950 ( .a(n45741), .b(n45740), .o(n45742) );
in01f01 g41951 ( .a(n45742), .o(n45743) );
na02f01 g41952 ( .a(n45743), .b(n45738), .o(n45744) );
na03f01 g41953 ( .a(n45742), .b(n5962), .c(n45737), .o(n45745) );
na02f01 g41954 ( .a(n45745), .b(n45744), .o(n4226) );
no02f01 g41955 ( .a(n8726), .b(n8471), .o(n45747) );
no02f01 g41956 ( .a(n8725), .b(n5973), .o(n45748) );
no03f01 g41957 ( .a(n45748), .b(n8758), .c(n8716), .o(n45749) );
no02f01 g41958 ( .a(n45749), .b(n45747), .o(n45750) );
no02f01 g41959 ( .a(n8736), .b(n8471), .o(n45751) );
no02f01 g41960 ( .a(n8735), .b(n5973), .o(n45752) );
no02f01 g41961 ( .a(n45752), .b(n45751), .o(n45753) );
in01f01 g41962 ( .a(n45753), .o(n45754) );
na02f01 g41963 ( .a(n45754), .b(n45750), .o(n45755) );
oa12f01 g41964 ( .a(n45753), .b(n45749), .c(n45747), .o(n45756) );
na02f01 g41965 ( .a(n45756), .b(n45755), .o(n4231) );
na03f01 g41966 ( .a(n25921), .b(n30106), .c(n30063), .o(n45758) );
oa12f01 g41967 ( .a(n25920), .b(n30107), .c(n25772), .o(n45759) );
na02f01 g41968 ( .a(n45759), .b(n45758), .o(n4236) );
no02f01 g41969 ( .a(n5930), .b(n42263), .o(n45761) );
ao12f01 g41970 ( .a(n5961), .b(n5938_1), .c(n45761), .o(n45762) );
in01f01 g41971 ( .a(n45762), .o(n45763) );
na02f01 g41972 ( .a(n5951), .b(n5946), .o(n45764) );
na02f01 g41973 ( .a(n45764), .b(n45763), .o(n45765) );
in01f01 g41974 ( .a(n45764), .o(n45766) );
na02f01 g41975 ( .a(n45766), .b(n45762), .o(n45767) );
na02f01 g41976 ( .a(n45767), .b(n45765), .o(n4246) );
in01f01 g41977 ( .a(n485), .o(n4251) );
na02f01 g41978 ( .a(n43659), .b(n43655), .o(n4261) );
in01f01 g41979 ( .a(n37132), .o(n45771) );
in01f01 g41980 ( .a(n37131), .o(n45772) );
na03f01 g41981 ( .a(n37135), .b(n45772), .c(n25297), .o(n45773) );
no02f01 g41982 ( .a(n25212), .b(n25023), .o(n45774) );
no02f01 g41983 ( .a(n25290), .b(n24613), .o(n45775) );
no02f01 g41984 ( .a(n45775), .b(n45774), .o(n45776) );
in01f01 g41985 ( .a(n45776), .o(n45777) );
na03f01 g41986 ( .a(n45777), .b(n45773), .c(n45771), .o(n45778) );
no03f01 g41987 ( .a(n37146), .b(n37131), .c(n25573), .o(n45779) );
oa12f01 g41988 ( .a(n45776), .b(n45779), .c(n37132), .o(n45780) );
na02f01 g41989 ( .a(n45780), .b(n45778), .o(n4266) );
na02f01 g41990 ( .a(n32732), .b(sin_out_20), .o(n45782) );
no02f01 g41991 ( .a(n41363), .b(n34307), .o(n45783) );
no02f01 g41992 ( .a(n45783), .b(n41324), .o(n45784) );
in01f01 g41993 ( .a(n45784), .o(n45785) );
no03f01 g41994 ( .a(n45785), .b(n41362), .c(n43523), .o(n45786) );
ao12f01 g41995 ( .a(n45784), .b(n41361), .c(n43431), .o(n45787) );
oa12f01 g41996 ( .a(n32734), .b(n45787), .c(n45786), .o(n45788) );
na02f01 g41997 ( .a(n45788), .b(n45782), .o(n4271) );
na03f01 g41998 ( .a(n32664), .b(n32703), .c(n32629), .o(n45790) );
oa12f01 g41999 ( .a(n32713), .b(n32630), .c(n32702), .o(n45791) );
na02f01 g42000 ( .a(n45791), .b(n45790), .o(n4280) );
in01f01 g42001 ( .a(n10775), .o(n45793) );
oa12f01 g42002 ( .a(n45793), .b(n10982), .c(n10976), .o(n45794) );
in01f01 g42003 ( .a(n45794), .o(n45795) );
no02f01 g42004 ( .a(n10748), .b(n3521), .o(n45796) );
no02f01 g42005 ( .a(n10986), .b(n45796), .o(n45797) );
na02f01 g42006 ( .a(n45797), .b(n45795), .o(n45798) );
in01f01 g42007 ( .a(n45797), .o(n45799) );
na02f01 g42008 ( .a(n45799), .b(n45794), .o(n45800) );
na02f01 g42009 ( .a(n45800), .b(n45798), .o(n4285) );
na03f01 g42010 ( .a(n39718), .b(n9590), .c(n9589), .o(n45802) );
oa12f01 g42011 ( .a(n847), .b(n9646), .c(n9645), .o(n45803) );
na02f01 g42012 ( .a(n45803), .b(n45802), .o(n4290) );
oa12f01 g42013 ( .a(n32325), .b(n32326), .c(n32446), .o(n45805) );
na03f01 g42014 ( .a(n32461), .b(n32460), .c(n32294), .o(n45806) );
na02f01 g42015 ( .a(n45806), .b(n45805), .o(n4295) );
no02f01 g42016 ( .a(n40486), .b(n22484), .o(n45808) );
no02f01 g42017 ( .a(n22446), .b(n22050), .o(n45809) );
no02f01 g42018 ( .a(n22452), .b(n21993), .o(n45810) );
no02f01 g42019 ( .a(n45810), .b(n45809), .o(n45811) );
oa12f01 g42020 ( .a(n45811), .b(n45808), .c(n40487), .o(n45812) );
in01f01 g42021 ( .a(n40487), .o(n45813) );
oa12f01 g42022 ( .a(n22426), .b(n22436), .c(n22050), .o(n45814) );
in01f01 g42023 ( .a(n45811), .o(n45815) );
na03f01 g42024 ( .a(n45815), .b(n45814), .c(n45813), .o(n45816) );
na03f01 g42025 ( .a(n45816), .b(n45812), .c(n2589), .o(n45817) );
ao12f01 g42026 ( .a(n45815), .b(n45814), .c(n45813), .o(n45818) );
no03f01 g42027 ( .a(n45811), .b(n45808), .c(n40487), .o(n45819) );
oa12f01 g42028 ( .a(n4116), .b(n45819), .c(n45818), .o(n45820) );
na02f01 g42029 ( .a(n45820), .b(n45817), .o(n4300) );
na02f01 g42030 ( .a(n45816), .b(n45812), .o(n4305) );
na04f01 g42031 ( .a(n32391), .b(n32389), .c(n32208), .d(n32193), .o(n45823) );
oa22f01 g42032 ( .a(n32390), .b(n32192), .c(n32484), .d(n32207), .o(n45824) );
na02f01 g42033 ( .a(n45824), .b(n45823), .o(n4310) );
na02f01 g42034 ( .a(n41811), .b(n41805), .o(n4315) );
no02f01 g42035 ( .a(n6948), .b(n6938), .o(n45827) );
in01f01 g42036 ( .a(n6969), .o(n45828) );
ao12f01 g42037 ( .a(n6985), .b(n45828), .c(n45827), .o(n45829) );
no02f01 g42038 ( .a(n6955), .b(n6934), .o(n45830) );
no02f01 g42039 ( .a(n45830), .b(n6957), .o(n45831) );
na02f01 g42040 ( .a(n45831), .b(n45829), .o(n45832) );
in01f01 g42041 ( .a(n45829), .o(n45833) );
in01f01 g42042 ( .a(n45831), .o(n45834) );
na02f01 g42043 ( .a(n45834), .b(n45833), .o(n45835) );
na02f01 g42044 ( .a(n45835), .b(n45832), .o(n4320) );
na02f01 g42045 ( .a(n44670), .b(n44669), .o(n4325) );
na02f01 g42046 ( .a(n32732), .b(cos_out_28), .o(n45838) );
na03f01 g42047 ( .a(n41588), .b(n41546), .c(n39691), .o(n45839) );
in01f01 g42048 ( .a(n45839), .o(n45840) );
no02f01 g42049 ( .a(n41609), .b(n35944), .o(n45841) );
no02f01 g42050 ( .a(n45841), .b(n41611), .o(n45842) );
in01f01 g42051 ( .a(n45842), .o(n45843) );
no03f01 g42052 ( .a(n45843), .b(n41636), .c(n45840), .o(n45844) );
in01f01 g42053 ( .a(n41636), .o(n45845) );
ao12f01 g42054 ( .a(n45842), .b(n45845), .c(n45839), .o(n45846) );
oa12f01 g42055 ( .a(n32734), .b(n45846), .c(n45844), .o(n45847) );
na02f01 g42056 ( .a(n45847), .b(n45838), .o(n4330) );
na02f01 g42057 ( .a(n45196), .b(n45194), .o(n4334) );
na03f01 g42058 ( .a(n44271), .b(n44269), .c(n5799), .o(n45850) );
na02f01 g42059 ( .a(n3010), .b(n911), .o(n45851) );
na02f01 g42060 ( .a(n45851), .b(n45850), .o(n4339) );
oa12f01 g42061 ( .a(n40266), .b(n41886), .c(n41884), .o(n45853) );
no02f01 g42062 ( .a(n40311), .b(n6037), .o(n45854) );
no02f01 g42063 ( .a(n45854), .b(n40274), .o(n45855) );
na03f01 g42064 ( .a(n45855), .b(n45853), .c(n40316), .o(n45856) );
ao12f01 g42065 ( .a(n40267), .b(n41885), .c(n41892), .o(n45857) );
in01f01 g42066 ( .a(n45855), .o(n45858) );
oa12f01 g42067 ( .a(n45858), .b(n45857), .c(n40315), .o(n45859) );
na02f01 g42068 ( .a(n45859), .b(n45856), .o(n4344) );
in01f01 g42069 ( .a(n37048), .o(n45861) );
no02f01 g42070 ( .a(n45861), .b(n36972), .o(n45862) );
no02f01 g42071 ( .a(n45862), .b(n37049), .o(n45863) );
na02f01 g42072 ( .a(n45863), .b(n37176), .o(n45864) );
in01f01 g42073 ( .a(n45863), .o(n45865) );
na02f01 g42074 ( .a(n45865), .b(n37042), .o(n45866) );
na02f01 g42075 ( .a(n45866), .b(n45864), .o(n4354) );
no02f01 g42076 ( .a(n9343), .b(n9225), .o(n45868) );
no02f01 g42077 ( .a(n9344), .b(n9224), .o(n45869) );
oa12f01 g42078 ( .a(n9350), .b(n45869), .c(n45868), .o(n45870) );
no02f01 g42079 ( .a(n45869), .b(n45868), .o(n45871) );
na02f01 g42080 ( .a(n45871), .b(n452), .o(n45872) );
na02f01 g42081 ( .a(n45872), .b(n45870), .o(n4359) );
na02f01 g42082 ( .a(n45263), .b(n45260), .o(n4364) );
na04f01 g42083 ( .a(n39121), .b(n39120), .c(n39077), .d(n39076), .o(n45875) );
oa22f01 g42084 ( .a(n38445), .b(n38282), .c(n38442), .d(n38296), .o(n45876) );
na02f01 g42085 ( .a(n45876), .b(n45875), .o(n4369) );
na02f01 g42086 ( .a(n41743), .b(n41739), .o(n4374) );
na02f01 g42087 ( .a(n44513), .b(n44512), .o(n4379) );
no02f01 g42088 ( .a(n11734), .b(n38076), .o(n45880) );
no02f01 g42089 ( .a(n11759), .b(n11725), .o(n45881) );
in01f01 g42090 ( .a(n45881), .o(n45882) );
oa12f01 g42091 ( .a(n45882), .b(n45880), .c(n11758), .o(n45883) );
no02f01 g42092 ( .a(n45880), .b(n11758), .o(n45884) );
na02f01 g42093 ( .a(n45881), .b(n45884), .o(n45885) );
na02f01 g42094 ( .a(n45885), .b(n45883), .o(n4384) );
na03f01 g42095 ( .a(n9225), .b(n8862), .c(n8765), .o(n45887) );
na02f01 g42096 ( .a(n45887), .b(n42526), .o(n4394) );
in01f01 g42097 ( .a(n44157), .o(n45889) );
ao12f01 g42098 ( .a(n44156), .b(n44155), .c(n45889), .o(n45890) );
no02f01 g42099 ( .a(n29528), .b(n29430), .o(n45891) );
no02f01 g42100 ( .a(n29527), .b(n29639), .o(n45892) );
no02f01 g42101 ( .a(n45892), .b(n45891), .o(n45893) );
in01f01 g42102 ( .a(n45893), .o(n45894) );
na02f01 g42103 ( .a(n45894), .b(n45890), .o(n45895) );
in01f01 g42104 ( .a(n45890), .o(n45896) );
na02f01 g42105 ( .a(n45893), .b(n45896), .o(n45897) );
na02f01 g42106 ( .a(n45897), .b(n45895), .o(n4404) );
in01f01 g42107 ( .a(n22164), .o(n45899) );
na03f01 g42108 ( .a(n22238), .b(n22237), .c(n45899), .o(n45900) );
in01f01 g42109 ( .a(n22237), .o(n45901) );
in01f01 g42110 ( .a(n22238), .o(n45902) );
oa12f01 g42111 ( .a(n45901), .b(n45902), .c(n22164), .o(n45903) );
na02f01 g42112 ( .a(n45903), .b(n45900), .o(n4409) );
oa12f01 g42113 ( .a(n22354), .b(n22332), .c(n22760), .o(n45905) );
in01f01 g42114 ( .a(n45905), .o(n45906) );
in01f01 g42115 ( .a(n22351), .o(n45907) );
no02f01 g42116 ( .a(n45907), .b(n22326), .o(n45908) );
no02f01 g42117 ( .a(n45908), .b(n45906), .o(n45909) );
na02f01 g42118 ( .a(n45908), .b(n45906), .o(n45910) );
in01f01 g42119 ( .a(n45910), .o(n45911) );
no02f01 g42120 ( .a(n45911), .b(n45909), .o(n45912) );
in01f01 g42121 ( .a(n45912), .o(n5849) );
na02f01 g42122 ( .a(n5849), .b(n4116), .o(n45914) );
na02f01 g42123 ( .a(n45912), .b(n2589), .o(n45915) );
na02f01 g42124 ( .a(n45915), .b(n45914), .o(n4414) );
na03f01 g42125 ( .a(n39447), .b(n40018), .c(n39427), .o(n45917) );
oa12f01 g42126 ( .a(n40024), .b(n39428), .c(n40017), .o(n45918) );
na02f01 g42127 ( .a(n45918), .b(n45917), .o(n4419) );
in01f01 g42128 ( .a(n42357), .o(n45920) );
na02f01 g42129 ( .a(n42355), .b(n45920), .o(n45921) );
ao12f01 g42130 ( .a(n45921), .b(n42352), .c(n27485), .o(n45922) );
in01f01 g42131 ( .a(n27479), .o(n45923) );
no02f01 g42132 ( .a(n27478), .b(n27367), .o(n45924) );
no02f01 g42133 ( .a(n45924), .b(n45923), .o(n45925) );
na02f01 g42134 ( .a(n45925), .b(n45922), .o(n45926) );
in01f01 g42135 ( .a(n45922), .o(n45927) );
in01f01 g42136 ( .a(n45925), .o(n45928) );
na02f01 g42137 ( .a(n45928), .b(n45927), .o(n45929) );
na02f01 g42138 ( .a(n45929), .b(n45926), .o(n4429) );
in01f01 g42139 ( .a(n37049), .o(n45931) );
oa12f01 g42140 ( .a(n45931), .b(n45862), .c(n37176), .o(n45932) );
in01f01 g42141 ( .a(n45932), .o(n45933) );
no02f01 g42142 ( .a(n37057), .b(n36963), .o(n45934) );
no02f01 g42143 ( .a(n37058), .b(n36972), .o(n45935) );
no02f01 g42144 ( .a(n45935), .b(n45934), .o(n45936) );
na02f01 g42145 ( .a(n45936), .b(n45933), .o(n45937) );
in01f01 g42146 ( .a(n45936), .o(n45938) );
na02f01 g42147 ( .a(n45938), .b(n45932), .o(n45939) );
na02f01 g42148 ( .a(n45939), .b(n45937), .o(n4434) );
oa12f01 g42149 ( .a(n30089), .b(n25810), .c(n30071), .o(n45941) );
na03f01 g42150 ( .a(n25865), .b(n30072), .c(n25809), .o(n45942) );
na02f01 g42151 ( .a(n45942), .b(n45941), .o(n4439) );
in01f01 g42152 ( .a(n43116), .o(n45944) );
no02f01 g42153 ( .a(n40748), .b(n21270), .o(n45945) );
no02f01 g42154 ( .a(n45945), .b(n43112), .o(n45946) );
in01f01 g42155 ( .a(n43111), .o(n45947) );
oa12f01 g42156 ( .a(n45947), .b(n41394), .c(n41393), .o(n45948) );
na03f01 g42157 ( .a(n45948), .b(n45946), .c(n45944), .o(n45949) );
in01f01 g42158 ( .a(n45946), .o(n45950) );
ao12f01 g42159 ( .a(n43111), .b(n41385), .c(n41382), .o(n45951) );
oa12f01 g42160 ( .a(n45950), .b(n45951), .c(n43116), .o(n45952) );
na03f01 g42161 ( .a(n45952), .b(n45949), .c(n5799), .o(n45953) );
no03f01 g42162 ( .a(n45951), .b(n45950), .c(n43116), .o(n45954) );
ao12f01 g42163 ( .a(n45946), .b(n45948), .c(n45944), .o(n45955) );
oa12f01 g42164 ( .a(n911), .b(n45955), .c(n45954), .o(n45956) );
na02f01 g42165 ( .a(n45956), .b(n45953), .o(n4453) );
in01f01 g42166 ( .a(n9515), .o(n45958) );
in01f01 g42167 ( .a(n9530), .o(n45959) );
na02f01 g42168 ( .a(n45022), .b(n45959), .o(n45960) );
no02f01 g42169 ( .a(n9531), .b(n9525), .o(n45961) );
in01f01 g42170 ( .a(n45961), .o(n45962) );
na03f01 g42171 ( .a(n45962), .b(n45960), .c(n45958), .o(n45963) );
na02f01 g42172 ( .a(n45960), .b(n45958), .o(n45964) );
na02f01 g42173 ( .a(n45961), .b(n45964), .o(n45965) );
na02f01 g42174 ( .a(n45965), .b(n45963), .o(n4458) );
no02f01 g42175 ( .a(n44385), .b(n44384), .o(n45967) );
oa12f01 g42176 ( .a(n45967), .b(n29425), .c(n29213), .o(n45968) );
oa12f01 g42177 ( .a(n44153), .b(n44385), .c(n44384), .o(n45969) );
na02f01 g42178 ( .a(n45969), .b(n45968), .o(n4463) );
na02f01 g42179 ( .a(n25640), .b(n22424), .o(n45971) );
no02f01 g42180 ( .a(n22474), .b(n22402), .o(n45972) );
in01f01 g42181 ( .a(n45972), .o(n45973) );
na03f01 g42182 ( .a(n45973), .b(n45971), .c(n22418), .o(n45974) );
oa12f01 g42183 ( .a(n22418), .b(n25644), .c(n22423), .o(n45975) );
na02f01 g42184 ( .a(n45972), .b(n45975), .o(n45976) );
na02f01 g42185 ( .a(n45976), .b(n45974), .o(n4468) );
no02f01 g42186 ( .a(n32480), .b(n32223), .o(n45978) );
oa12f01 g42187 ( .a(n45978), .b(n32483), .c(n32207), .o(n45979) );
in01f01 g42188 ( .a(n45978), .o(n45980) );
na03f01 g42189 ( .a(n32388), .b(n45980), .c(n32208), .o(n45981) );
na02f01 g42190 ( .a(n45981), .b(n45979), .o(n4473) );
no02f01 g42191 ( .a(n37366), .b(n37278), .o(n45983) );
na03f01 g42192 ( .a(n41103), .b(n41102), .c(delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(n45984) );
na02f01 g42193 ( .a(n1250), .b(n37149), .o(n45985) );
ao22f01 g42194 ( .a(n45985), .b(n45984), .c(n45983), .d(delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(n4478) );
ao12f01 g42195 ( .a(n38779), .b(n38776), .c(n43175), .o(n45987) );
no02f01 g42196 ( .a(n38780), .b(n36115), .o(n45988) );
na02f01 g42197 ( .a(n45988), .b(n45987), .o(n45989) );
in01f01 g42198 ( .a(n45987), .o(n45990) );
in01f01 g42199 ( .a(n45988), .o(n45991) );
na02f01 g42200 ( .a(n45991), .b(n45990), .o(n45992) );
na02f01 g42201 ( .a(n45992), .b(n45989), .o(n4483) );
in01f01 g42202 ( .a(n35463), .o(n45994) );
ao12f01 g42203 ( .a(n43953), .b(n45994), .c(n35441), .o(n45995) );
no02f01 g42204 ( .a(n35453), .b(n4176), .o(n45996) );
no02f01 g42205 ( .a(n45996), .b(n35455), .o(n45997) );
na02f01 g42206 ( .a(n45997), .b(n45995), .o(n45998) );
in01f01 g42207 ( .a(n45995), .o(n45999) );
in01f01 g42208 ( .a(n45997), .o(n46000) );
na02f01 g42209 ( .a(n46000), .b(n45999), .o(n46001) );
na02f01 g42210 ( .a(n46001), .b(n45998), .o(n4493) );
na03f01 g42211 ( .a(n45780), .b(n45778), .c(n6037), .o(n46003) );
no03f01 g42212 ( .a(n45776), .b(n45779), .c(n37132), .o(n46004) );
ao12f01 g42213 ( .a(n45777), .b(n45773), .c(n45771), .o(n46005) );
oa12f01 g42214 ( .a(n5873), .b(n46005), .c(n46004), .o(n46006) );
na02f01 g42215 ( .a(n46006), .b(n46003), .o(n4503) );
na02f01 g42216 ( .a(n21525), .b(n42236), .o(n46008) );
no02f01 g42217 ( .a(n21586), .b(n21585), .o(n46009) );
no02f01 g42218 ( .a(n21555), .b(n16329), .o(n46010) );
no02f01 g42219 ( .a(n46010), .b(n21557), .o(n46011) );
na03f01 g42220 ( .a(n46011), .b(n46009), .c(n46008), .o(n46012) );
oa12f01 g42221 ( .a(n46009), .b(n21526), .c(n42235), .o(n46013) );
in01f01 g42222 ( .a(n46011), .o(n46014) );
na02f01 g42223 ( .a(n46014), .b(n46013), .o(n46015) );
na02f01 g42224 ( .a(n46015), .b(n46012), .o(n4508) );
no02f01 g42225 ( .a(n43416), .b(n43415), .o(n46017) );
na02f01 g42226 ( .a(n46017), .b(n43420), .o(n46018) );
in01f01 g42227 ( .a(n43420), .o(n46019) );
in01f01 g42228 ( .a(n46017), .o(n46020) );
na02f01 g42229 ( .a(n46020), .b(n46019), .o(n46021) );
na02f01 g42230 ( .a(n46021), .b(n46018), .o(n4513) );
na03f01 g42231 ( .a(n9590), .b(n9589), .c(n9243), .o(n46023) );
oa12f01 g42232 ( .a(n233), .b(n9646), .c(n9645), .o(n46024) );
na02f01 g42233 ( .a(n46024), .b(n46023), .o(n4518) );
oa12f01 g42234 ( .a(n27028), .b(n27029), .c(n27206), .o(n46026) );
na03f01 g42235 ( .a(n27226), .b(n27225), .c(n26982), .o(n46027) );
na02f01 g42236 ( .a(n46027), .b(n46026), .o(n4523) );
no02f01 g42237 ( .a(n10898), .b(n25629), .o(n46029) );
no02f01 g42238 ( .a(n46029), .b(n40539), .o(n46030) );
no02f01 g42239 ( .a(n10886), .b(n3521), .o(n46031) );
no02f01 g42240 ( .a(n46031), .b(n10888), .o(n46032) );
na02f01 g42241 ( .a(n46032), .b(n46030), .o(n46033) );
in01f01 g42242 ( .a(n46032), .o(n46034) );
oa12f01 g42243 ( .a(n46034), .b(n46029), .c(n40539), .o(n46035) );
na02f01 g42244 ( .a(n46035), .b(n46033), .o(n4528) );
in01f01 g42245 ( .a(n14205), .o(n46037) );
no02f01 g42246 ( .a(n46037), .b(n14048), .o(n46038) );
no02f01 g42247 ( .a(n14206), .b(n14035), .o(n46039) );
no02f01 g42248 ( .a(n46039), .b(n46038), .o(n46040) );
na02f01 g42249 ( .a(n46039), .b(n46038), .o(n46041) );
in01f01 g42250 ( .a(n46041), .o(n46042) );
no02f01 g42251 ( .a(n46042), .b(n46040), .o(n46043) );
in01f01 g42252 ( .a(n46043), .o(n5220) );
na02f01 g42253 ( .a(n5220), .b(n4116), .o(n46045) );
na02f01 g42254 ( .a(n46043), .b(n2589), .o(n46046) );
na02f01 g42255 ( .a(n46046), .b(n46045), .o(n4533) );
in01f01 g42256 ( .a(n42764), .o(n46048) );
ao12f01 g42257 ( .a(n42765), .b(n46048), .c(n39521), .o(n46049) );
no02f01 g42258 ( .a(n32078), .b(n31606), .o(n46050) );
no02f01 g42259 ( .a(n38250), .b(n31607), .o(n46051) );
no02f01 g42260 ( .a(n46051), .b(n46050), .o(n46052) );
na02f01 g42261 ( .a(n46052), .b(n46049), .o(n46053) );
in01f01 g42262 ( .a(n46049), .o(n46054) );
in01f01 g42263 ( .a(n46052), .o(n46055) );
na02f01 g42264 ( .a(n46055), .b(n46054), .o(n46056) );
na02f01 g42265 ( .a(n46056), .b(n46053), .o(n4538) );
na03f01 g42266 ( .a(n42543), .b(n42542), .c(n3633), .o(n46058) );
na02f01 g42267 ( .a(n1894), .b(n6203), .o(n46059) );
na02f01 g42268 ( .a(n46059), .b(n46058), .o(n4543) );
no02f01 g42269 ( .a(n11695), .b(n11559), .o(n46061) );
in01f01 g42270 ( .a(n46061), .o(n46062) );
na02f01 g42271 ( .a(n46062), .b(n11694), .o(n46063) );
in01f01 g42272 ( .a(n11694), .o(n46064) );
na02f01 g42273 ( .a(n46061), .b(n46064), .o(n46065) );
na02f01 g42274 ( .a(n46065), .b(n46063), .o(n4548) );
na02f01 g42275 ( .a(n37277), .b(n37274), .o(n4553) );
no02f01 g42276 ( .a(n42946), .b(n42945), .o(n46068) );
na02f01 g42277 ( .a(n46068), .b(n38980), .o(n46069) );
in01f01 g42278 ( .a(n46068), .o(n46070) );
na02f01 g42279 ( .a(n46070), .b(n38979), .o(n46071) );
na02f01 g42280 ( .a(n46071), .b(n46069), .o(n4563) );
in01f01 g42281 ( .a(n43418), .o(n46073) );
no02f01 g42282 ( .a(n16231), .b(n16184), .o(n46074) );
na03f01 g42283 ( .a(n46074), .b(n39733), .c(n46073), .o(n46075) );
oa22f01 g42284 ( .a(n16232), .b(n43418), .c(n16231), .d(n16184), .o(n46076) );
na02f01 g42285 ( .a(n46076), .b(n46075), .o(n4578) );
no03f01 g42286 ( .a(n9815), .b(n9797), .c(n40341), .o(n46078) );
in01f01 g42287 ( .a(n9819), .o(n46079) );
na02f01 g42288 ( .a(n9821), .b(n46079), .o(n46080) );
no02f01 g42289 ( .a(n46080), .b(n46078), .o(n46081) );
no02f01 g42290 ( .a(n9820), .b(n5001), .o(n46082) );
no02f01 g42291 ( .a(n46082), .b(n9808), .o(n46083) );
na02f01 g42292 ( .a(n46083), .b(n46081), .o(n46084) );
in01f01 g42293 ( .a(n46083), .o(n46085) );
oa12f01 g42294 ( .a(n46085), .b(n46080), .c(n46078), .o(n46086) );
na02f01 g42295 ( .a(n46086), .b(n46084), .o(n4583) );
no03f01 g42296 ( .a(n4201), .b(n9231), .c(n9228), .o(n46088) );
no02f01 g42297 ( .a(n9232), .b(n936), .o(n46089) );
no02f01 g42298 ( .a(n46089), .b(n46088), .o(n46090) );
na03f01 g42299 ( .a(n46090), .b(n9590), .c(n9589), .o(n46091) );
in01f01 g42300 ( .a(n46090), .o(n5210) );
oa12f01 g42301 ( .a(n5210), .b(n9646), .c(n9645), .o(n46093) );
na02f01 g42302 ( .a(n46093), .b(n46091), .o(n4588) );
in01f01 g42303 ( .a(n22233), .o(n46095) );
oa12f01 g42304 ( .a(n22232), .b(n46095), .c(n22209), .o(n46096) );
in01f01 g42305 ( .a(n22209), .o(n46097) );
in01f01 g42306 ( .a(n22232), .o(n46098) );
na03f01 g42307 ( .a(n22233), .b(n46098), .c(n46097), .o(n46099) );
na02f01 g42308 ( .a(n46099), .b(n46096), .o(n4593) );
na02f01 g42309 ( .a(n45388), .b(n45386), .o(n4598) );
in01f01 g42310 ( .a(n44284), .o(n46102) );
oa12f01 g42311 ( .a(n39830), .b(n46102), .c(n41455), .o(n46103) );
no02f01 g42312 ( .a(n46103), .b(n4201), .o(n46104) );
na02f01 g42313 ( .a(n46103), .b(n4201), .o(n46105) );
in01f01 g42314 ( .a(n46105), .o(n46106) );
no02f01 g42315 ( .a(n46106), .b(n46104), .o(n46107) );
in01f01 g42316 ( .a(n46107), .o(n4603) );
in01f01 g42317 ( .a(n14199), .o(n46109) );
in01f01 g42318 ( .a(n14200), .o(n46110) );
no02f01 g42319 ( .a(n46110), .b(n14060), .o(n46111) );
in01f01 g42320 ( .a(n46111), .o(n46112) );
no03f01 g42321 ( .a(n46112), .b(n46109), .c(n14071), .o(n46113) );
ao12f01 g42322 ( .a(n46111), .b(n14199), .c(n14072), .o(n46114) );
no02f01 g42323 ( .a(n46114), .b(n46113), .o(n46115) );
in01f01 g42324 ( .a(n46115), .o(n4608) );
na03f01 g42325 ( .a(n45565), .b(n45561), .c(n6037), .o(n46117) );
no03f01 g42326 ( .a(n45564), .b(n45563), .c(n45562), .o(n46118) );
ao12f01 g42327 ( .a(n45556), .b(n45560), .c(n45558), .o(n46119) );
oa12f01 g42328 ( .a(n5873), .b(n46119), .c(n46118), .o(n46120) );
na02f01 g42329 ( .a(n46120), .b(n46117), .o(n4618) );
in01f01 g42330 ( .a(n27574), .o(n46122) );
na03f01 g42331 ( .a(n46122), .b(n27672), .c(n42461), .o(n46123) );
no02f01 g42332 ( .a(n44583), .b(n27631), .o(n46124) );
no02f01 g42333 ( .a(n27583), .b(n27367), .o(n46125) );
no02f01 g42334 ( .a(n46125), .b(n27585), .o(n46126) );
na03f01 g42335 ( .a(n46126), .b(n46124), .c(n46123), .o(n46127) );
na02f01 g42336 ( .a(n46124), .b(n46123), .o(n46128) );
in01f01 g42337 ( .a(n46126), .o(n46129) );
na02f01 g42338 ( .a(n46129), .b(n46128), .o(n46130) );
na02f01 g42339 ( .a(n46130), .b(n46127), .o(n4623) );
na02f01 g42340 ( .a(n41036), .b(n41031), .o(n4628) );
ao12f01 g42341 ( .a(n45138), .b(n45139), .c(n27671), .o(n46133) );
in01f01 g42342 ( .a(n27517), .o(n46134) );
no02f01 g42343 ( .a(n46134), .b(n27395), .o(n46135) );
no02f01 g42344 ( .a(n27517), .b(n27367), .o(n46136) );
no02f01 g42345 ( .a(n46136), .b(n46135), .o(n46137) );
na02f01 g42346 ( .a(n46137), .b(n46133), .o(n46138) );
in01f01 g42347 ( .a(n46133), .o(n46139) );
in01f01 g42348 ( .a(n46137), .o(n46140) );
na02f01 g42349 ( .a(n46140), .b(n46139), .o(n46141) );
na02f01 g42350 ( .a(n46141), .b(n46138), .o(n4633) );
no02f01 g42351 ( .a(n6967), .b(n6934), .o(n46143) );
no02f01 g42352 ( .a(n46143), .b(n6969), .o(n46144) );
in01f01 g42353 ( .a(n46144), .o(n46145) );
oa12f01 g42354 ( .a(n46145), .b(n44457), .c(n45827), .o(n46146) );
in01f01 g42355 ( .a(n45827), .o(n46147) );
in01f01 g42356 ( .a(n44457), .o(n46148) );
na03f01 g42357 ( .a(n46144), .b(n46148), .c(n46147), .o(n46149) );
na02f01 g42358 ( .a(n46149), .b(n46146), .o(n4638) );
no02f01 g42359 ( .a(n41919), .b(n41915), .o(n46151) );
na03f01 g42360 ( .a(n46151), .b(n27171), .c(n27249), .o(n46152) );
in01f01 g42361 ( .a(n46151), .o(n46153) );
oa12f01 g42362 ( .a(n46153), .b(n27172), .c(n27166), .o(n46154) );
na02f01 g42363 ( .a(n46154), .b(n46152), .o(n4643) );
na02f01 g42364 ( .a(n32732), .b(sin_out_8), .o(n46156) );
no02f01 g42365 ( .a(n36597), .b(n36553), .o(n46157) );
in01f01 g42366 ( .a(n46157), .o(n46158) );
no02f01 g42367 ( .a(n46158), .b(n36595), .o(n46159) );
no02f01 g42368 ( .a(n46157), .b(n38595), .o(n46160) );
oa12f01 g42369 ( .a(n32734), .b(n46160), .c(n46159), .o(n46161) );
na02f01 g42370 ( .a(n46161), .b(n46156), .o(n4648) );
oa12f01 g42371 ( .a(n17949), .b(n17918), .c(n17917), .o(n46163) );
na03f01 g42372 ( .a(n17922), .b(n17948), .c(n17947), .o(n46164) );
na02f01 g42373 ( .a(n46164), .b(n46163), .o(n4652) );
na02f01 g42374 ( .a(n42212), .b(n6037), .o(n46166) );
na02f01 g42375 ( .a(n1689), .b(n5873), .o(n46167) );
na02f01 g42376 ( .a(n46167), .b(n46166), .o(n4657) );
no02f01 g42377 ( .a(n16381), .b(n45505), .o(n46169) );
in01f01 g42378 ( .a(n16403), .o(n46170) );
na02f01 g42379 ( .a(n16402), .b(n16155), .o(n46171) );
na02f01 g42380 ( .a(n46171), .b(n16437), .o(n46172) );
ao12f01 g42381 ( .a(n46172), .b(n46170), .c(n46169), .o(n46173) );
no02f01 g42382 ( .a(n16423), .b(n16329), .o(n46174) );
no02f01 g42383 ( .a(n46174), .b(n16425), .o(n46175) );
na02f01 g42384 ( .a(n46175), .b(n46173), .o(n46176) );
in01f01 g42385 ( .a(n46173), .o(n46177) );
in01f01 g42386 ( .a(n46175), .o(n46178) );
na02f01 g42387 ( .a(n46178), .b(n46177), .o(n46179) );
na02f01 g42388 ( .a(n46179), .b(n46176), .o(n4662) );
no03f01 g42389 ( .a(n5716), .b(n9646), .c(n9645), .o(n46181) );
ao12f01 g42390 ( .a(n3707), .b(n9590), .c(n9589), .o(n46182) );
no02f01 g42391 ( .a(n46182), .b(n46181), .o(n4672) );
no02f01 g42392 ( .a(n9398), .b(n9381), .o(n46184) );
na02f01 g42393 ( .a(n46184), .b(n35575), .o(n46185) );
in01f01 g42394 ( .a(n46184), .o(n46186) );
na02f01 g42395 ( .a(n46186), .b(n35576), .o(n46187) );
na02f01 g42396 ( .a(n46187), .b(n46185), .o(n4677) );
na02f01 g42397 ( .a(n3297), .b(n4116), .o(n46189) );
na02f01 g42398 ( .a(n44623), .b(n2589), .o(n46190) );
na02f01 g42399 ( .a(n46190), .b(n46189), .o(n4682) );
na02f01 g42400 ( .a(n1739), .b(n4116), .o(n46192) );
na02f01 g42401 ( .a(n42281), .b(n2589), .o(n46193) );
na02f01 g42402 ( .a(n46193), .b(n46192), .o(n4687) );
no03f01 g42403 ( .a(n42933), .b(n42932), .c(n40447), .o(n46195) );
ao12f01 g42404 ( .a(n42928), .b(n42930), .c(n42925), .o(n46196) );
oa12f01 g42405 ( .a(n34420), .b(n46196), .c(n46195), .o(n46197) );
na03f01 g42406 ( .a(n42934), .b(n42931), .c(n_27923), .o(n46198) );
na02f01 g42407 ( .a(n46198), .b(n46197), .o(n4692) );
no02f01 g42408 ( .a(n7013), .b(n6989), .o(n46200) );
no02f01 g42409 ( .a(n46200), .b(n37369), .o(n46201) );
no02f01 g42410 ( .a(n7004), .b(n6934), .o(n46202) );
no02f01 g42411 ( .a(n46202), .b(n7006), .o(n46203) );
na02f01 g42412 ( .a(n46203), .b(n46201), .o(n46204) );
in01f01 g42413 ( .a(n46203), .o(n46205) );
oa12f01 g42414 ( .a(n46205), .b(n46200), .c(n37369), .o(n46206) );
na02f01 g42415 ( .a(n46206), .b(n46204), .o(n4697) );
no02f01 g42416 ( .a(n45178), .b(n45177), .o(n46208) );
na02f01 g42417 ( .a(n46208), .b(n45175), .o(n46209) );
in01f01 g42418 ( .a(n46208), .o(n46210) );
na02f01 g42419 ( .a(n46210), .b(n45176), .o(n46211) );
na02f01 g42420 ( .a(n46211), .b(n46209), .o(n4702) );
no02f01 g42421 ( .a(n41764), .b(n41763), .o(n46213) );
in01f01 g42422 ( .a(n46213), .o(n46214) );
na02f01 g42423 ( .a(n46214), .b(n41762), .o(n46215) );
na02f01 g42424 ( .a(n46213), .b(n41761), .o(n46216) );
na02f01 g42425 ( .a(n46216), .b(n46215), .o(n4707) );
no02f01 g42426 ( .a(n36625), .b(n36624), .o(n46218) );
in01f01 g42427 ( .a(n46218), .o(n46219) );
na04f01 g42428 ( .a(n46219), .b(n25484), .c(n25481), .d(n36621), .o(n46220) );
oa22f01 g42429 ( .a(n46218), .b(n25377), .c(n36654), .d(n36653), .o(n46221) );
na02f01 g42430 ( .a(n46221), .b(n46220), .o(n4712) );
in01f01 g42431 ( .a(n41832), .o(n46223) );
no02f01 g42432 ( .a(n39135), .b(n31586), .o(n46224) );
na02f01 g42433 ( .a(n39135), .b(n31586), .o(n46225) );
in01f01 g42434 ( .a(n46225), .o(n46226) );
no02f01 g42435 ( .a(n46226), .b(n46224), .o(n46227) );
in01f01 g42436 ( .a(n46227), .o(n46228) );
in01f01 g42437 ( .a(n41830), .o(n46229) );
na03f01 g42438 ( .a(n41829), .b(n41828), .c(n46229), .o(n46230) );
na03f01 g42439 ( .a(n46230), .b(n46228), .c(n46223), .o(n46231) );
no03f01 g42440 ( .a(n41836), .b(n41835), .c(n41830), .o(n46232) );
oa12f01 g42441 ( .a(n46227), .b(n46232), .c(n41832), .o(n46233) );
na02f01 g42442 ( .a(n46233), .b(n46231), .o(n4717) );
no03f01 g42443 ( .a(n4201), .b(n9231), .c(n9228), .o(n46235) );
ao12f01 g42444 ( .a(n9591), .b(n9231), .c(n936), .o(n46236) );
no02f01 g42445 ( .a(n46236), .b(n46235), .o(n46237) );
in01f01 g42446 ( .a(n46237), .o(n4722) );
na02f01 g42447 ( .a(n32732), .b(cos_out_19), .o(n46239) );
no02f01 g42448 ( .a(n39676), .b(n36374), .o(n46240) );
no02f01 g42449 ( .a(n39686), .b(n35944), .o(n46241) );
no02f01 g42450 ( .a(n46241), .b(n39688), .o(n46242) );
in01f01 g42451 ( .a(n46242), .o(n46243) );
no04f01 g42452 ( .a(n46243), .b(n46240), .c(n43667), .d(n39692), .o(n46244) );
no03f01 g42453 ( .a(n46240), .b(n43667), .c(n39692), .o(n46245) );
no02f01 g42454 ( .a(n46242), .b(n46245), .o(n46246) );
oa12f01 g42455 ( .a(n32734), .b(n46246), .c(n46244), .o(n46247) );
na02f01 g42456 ( .a(n46247), .b(n46239), .o(n4732) );
na02f01 g42457 ( .a(n20974), .b(n20969), .o(n46249) );
in01f01 g42458 ( .a(n46249), .o(n46250) );
no02f01 g42459 ( .a(n46250), .b(n38879), .o(n46251) );
no02f01 g42460 ( .a(n46249), .b(n38880), .o(n46252) );
no02f01 g42461 ( .a(n46252), .b(n46251), .o(n46253) );
na02f01 g42462 ( .a(n46253), .b(n5799), .o(n46254) );
in01f01 g42463 ( .a(n46253), .o(n4907) );
na02f01 g42464 ( .a(n4907), .b(n911), .o(n46256) );
na02f01 g42465 ( .a(n46256), .b(n46254), .o(n4741) );
oa12f01 g42466 ( .a(n7514), .b(n7544), .c(n7477), .o(n46258) );
na03f01 g42467 ( .a(n7515), .b(n7540), .c(n7525), .o(n46259) );
na02f01 g42468 ( .a(n46259), .b(n46258), .o(n4746) );
no02f01 g42469 ( .a(n35278), .b(n4176), .o(n46261) );
in01f01 g42470 ( .a(n46261), .o(n46262) );
na03f01 g42471 ( .a(n46262), .b(n35279), .c(n_186), .o(n46263) );
oa12f01 g42472 ( .a(n34438), .b(n46261), .c(n43210), .o(n46264) );
na02f01 g42473 ( .a(n46264), .b(n46263), .o(n4751) );
no02f01 g42474 ( .a(n40528), .b(n27600), .o(n46266) );
na03f01 g42475 ( .a(n46266), .b(n27633), .c(n27673), .o(n46267) );
in01f01 g42476 ( .a(n27633), .o(n46268) );
in01f01 g42477 ( .a(n46266), .o(n46269) );
oa12f01 g42478 ( .a(n46269), .b(n46268), .c(n27588), .o(n46270) );
na02f01 g42479 ( .a(n46270), .b(n46267), .o(n4756) );
na02f01 g42480 ( .a(n21257), .b(n21255), .o(n46272) );
in01f01 g42481 ( .a(n46272), .o(n46273) );
no02f01 g42482 ( .a(n46273), .b(n44128), .o(n46274) );
no02f01 g42483 ( .a(n46272), .b(n21243), .o(n46275) );
no02f01 g42484 ( .a(n46275), .b(n46274), .o(n46276) );
in01f01 g42485 ( .a(n46276), .o(n4766) );
na03f01 g42486 ( .a(n45535), .b(n45533), .c(n3633), .o(n46278) );
na02f01 g42487 ( .a(n3990), .b(n6203), .o(n46279) );
na02f01 g42488 ( .a(n46279), .b(n46278), .o(n4771) );
in01f01 g42489 ( .a(mux_while_ln12_psv_q_2_), .o(n46281) );
no02f01 g42490 ( .a(n45728), .b(n46281), .o(n4776) );
na02f01 g42491 ( .a(n44183), .b(n44180), .o(n4781) );
no02f01 g42492 ( .a(n9371), .b(n9224), .o(n46284) );
no02f01 g42493 ( .a(n9367), .b(n9225), .o(n46285) );
no02f01 g42494 ( .a(n38973), .b(n38972), .o(n46286) );
oa22f01 g42495 ( .a(n46286), .b(n38974), .c(n46285), .d(n46284), .o(n46287) );
no02f01 g42496 ( .a(n46286), .b(n38974), .o(n46288) );
no02f01 g42497 ( .a(n46285), .b(n46284), .o(n46289) );
na02f01 g42498 ( .a(n46289), .b(n46288), .o(n46290) );
na02f01 g42499 ( .a(n46290), .b(n46287), .o(n4791) );
na02f01 g42500 ( .a(n39201), .b(n39198), .o(n4796) );
no02f01 g42501 ( .a(n43037), .b(n9469), .o(n46293) );
no02f01 g42502 ( .a(n46293), .b(n9485), .o(n46294) );
no02f01 g42503 ( .a(n9484), .b(n9479), .o(n46295) );
na02f01 g42504 ( .a(n46295), .b(n46294), .o(n46296) );
in01f01 g42505 ( .a(n46295), .o(n46297) );
oa12f01 g42506 ( .a(n46297), .b(n46293), .c(n9485), .o(n46298) );
na02f01 g42507 ( .a(n46298), .b(n46296), .o(n4801) );
na02f01 g42508 ( .a(n32732), .b(sin_out_30), .o(n46300) );
no02f01 g42509 ( .a(n35882), .b(n34287), .o(n46301) );
no02f01 g42510 ( .a(n44787), .b(n35878), .o(n46302) );
no02f01 g42511 ( .a(n46302), .b(n46301), .o(n46303) );
no02f01 g42512 ( .a(n34287), .b(n33506), .o(n46304) );
no02f01 g42513 ( .a(n46304), .b(n35879), .o(n46305) );
no02f01 g42514 ( .a(n46305), .b(n46303), .o(n46306) );
na02f01 g42515 ( .a(n46305), .b(n46303), .o(n46307) );
in01f01 g42516 ( .a(n46307), .o(n46308) );
no03f01 g42517 ( .a(n46308), .b(n46306), .c(n34267), .o(n46309) );
no02f01 g42518 ( .a(n46308), .b(n46306), .o(n46310) );
no02f01 g42519 ( .a(n46310), .b(n34307), .o(n46311) );
no02f01 g42520 ( .a(n46311), .b(n46309), .o(n46312) );
in01f01 g42521 ( .a(n46312), .o(n46313) );
no02f01 g42522 ( .a(n44813), .b(n44796), .o(n46314) );
ao12f01 g42523 ( .a(n34307), .b(n44814), .c(n44794), .o(n46315) );
in01f01 g42524 ( .a(n46315), .o(n46316) );
na03f01 g42525 ( .a(n46316), .b(n44820), .c(n44819), .o(n46317) );
ao12f01 g42526 ( .a(n46313), .b(n46317), .c(n46314), .o(n46318) );
in01f01 g42527 ( .a(n46314), .o(n46319) );
no03f01 g42528 ( .a(n46315), .b(n44802), .c(n44799), .o(n46320) );
no03f01 g42529 ( .a(n46320), .b(n46319), .c(n46312), .o(n46321) );
oa12f01 g42530 ( .a(n32734), .b(n46321), .c(n46318), .o(n46322) );
na02f01 g42531 ( .a(n46322), .b(n46300), .o(n4806) );
in01f01 g42532 ( .a(n10826), .o(n46324) );
na03f01 g42533 ( .a(n5618), .b(n10827), .c(n46324), .o(n46325) );
in01f01 g42534 ( .a(n10827), .o(n46326) );
oa12f01 g42535 ( .a(n10833), .b(n46326), .c(n10826), .o(n46327) );
na02f01 g42536 ( .a(n46327), .b(n46325), .o(n4810) );
oa12f01 g42537 ( .a(n39448), .b(n40014), .c(n39411), .o(n46329) );
na03f01 g42538 ( .a(n40025), .b(n39412), .c(n40013), .o(n46330) );
na02f01 g42539 ( .a(n46330), .b(n46329), .o(n4815) );
na02f01 g42540 ( .a(n46276), .b(n5799), .o(n46332) );
na02f01 g42541 ( .a(n4766), .b(n911), .o(n46333) );
na02f01 g42542 ( .a(n46333), .b(n46332), .o(n4820) );
na02f01 g42543 ( .a(n32732), .b(sin_out_24), .o(n46335) );
no03f01 g42544 ( .a(n44554), .b(n43522), .c(n39599), .o(n46336) );
in01f01 g42545 ( .a(n41371), .o(n46337) );
no02f01 g42546 ( .a(n41355), .b(n41291), .o(n46338) );
in01f01 g42547 ( .a(n46338), .o(n46339) );
no03f01 g42548 ( .a(n46339), .b(n46337), .c(n46336), .o(n46340) );
ao12f01 g42549 ( .a(n46338), .b(n41371), .c(n41353), .o(n46341) );
oa12f01 g42550 ( .a(n32734), .b(n46341), .c(n46340), .o(n46342) );
na02f01 g42551 ( .a(n46342), .b(n46335), .o(n4825) );
in01f01 g42552 ( .a(n11619), .o(n46344) );
oa12f01 g42553 ( .a(delay_sub_ln23_0_unr1_stage2_stallmux_q_0_), .b(n11620), .c(n46344), .o(n46345) );
in01f01 g42554 ( .a(delay_sub_ln23_0_unr1_stage2_stallmux_q_0_), .o(n5255) );
in01f01 g42555 ( .a(n11620), .o(n46347) );
na03f01 g42556 ( .a(n46347), .b(n11619), .c(n5255), .o(n46348) );
na02f01 g42557 ( .a(n46348), .b(n46345), .o(n4829) );
no02f01 g42558 ( .a(n7025), .b(n7016), .o(n46350) );
no02f01 g42559 ( .a(n9670), .b(n6934), .o(n46351) );
no02f01 g42560 ( .a(n9669), .b(n5001), .o(n46352) );
no02f01 g42561 ( .a(n46352), .b(n46351), .o(n46353) );
in01f01 g42562 ( .a(n46353), .o(n46354) );
oa12f01 g42563 ( .a(n46354), .b(n46350), .c(n7026), .o(n46355) );
no02f01 g42564 ( .a(n46350), .b(n7026), .o(n46356) );
na02f01 g42565 ( .a(n46353), .b(n46356), .o(n46357) );
na02f01 g42566 ( .a(n46357), .b(n46355), .o(n4834) );
no02f01 g42567 ( .a(n11802), .b(n11775), .o(n46359) );
in01f01 g42568 ( .a(n46359), .o(n46360) );
na02f01 g42569 ( .a(n46360), .b(n11765), .o(n46361) );
na02f01 g42570 ( .a(n46359), .b(n41856), .o(n46362) );
na02f01 g42571 ( .a(n46362), .b(n46361), .o(n4839) );
no02f01 g42572 ( .a(n43070), .b(n8751), .o(n46364) );
na03f01 g42573 ( .a(n46364), .b(n8675), .c(n8661), .o(n46365) );
in01f01 g42574 ( .a(n46364), .o(n46366) );
na02f01 g42575 ( .a(n46366), .b(n43069), .o(n46367) );
na02f01 g42576 ( .a(n46367), .b(n46365), .o(n4848) );
oa12f01 g42577 ( .a(n16082), .b(n21360), .c(n21359), .o(n46369) );
na02f01 g42578 ( .a(n46369), .b(n16084), .o(n4853) );
na03f01 g42579 ( .a(n45600), .b(n9590), .c(n9589), .o(n46371) );
oa12f01 g42580 ( .a(n4053), .b(n9646), .c(n9645), .o(n46372) );
na02f01 g42581 ( .a(n46372), .b(n46371), .o(n4858) );
na03f01 g42582 ( .a(n27679), .b(n27642), .c(delay_sub_ln23_0_unr27_stage10_stallmux_z), .o(n46374) );
na02f01 g42583 ( .a(n348), .b(n21621), .o(n46375) );
na02f01 g42584 ( .a(n46375), .b(n46374), .o(n4863) );
na02f01 g42585 ( .a(n40230), .b(n6037), .o(n46377) );
na02f01 g42586 ( .a(n976), .b(n5873), .o(n46378) );
na02f01 g42587 ( .a(n46378), .b(n46377), .o(n4868) );
no02f01 g42588 ( .a(n38896), .b(n44830), .o(n46380) );
no02f01 g42589 ( .a(n46380), .b(n38907), .o(n46381) );
no02f01 g42590 ( .a(n38909), .b(n38903), .o(n46382) );
na02f01 g42591 ( .a(n46382), .b(n46381), .o(n46383) );
in01f01 g42592 ( .a(n46382), .o(n46384) );
oa12f01 g42593 ( .a(n46384), .b(n46380), .c(n38907), .o(n46385) );
na02f01 g42594 ( .a(n46385), .b(n46383), .o(n4873) );
na02f01 g42595 ( .a(n43123), .b(n43120), .o(n4878) );
na03f01 g42596 ( .a(n44711), .b(n44707), .c(n1821), .o(n46388) );
no03f01 g42597 ( .a(n44710), .b(n44709), .c(n44708), .o(n46389) );
ao12f01 g42598 ( .a(n44702), .b(n44706), .c(n44704), .o(n46390) );
oa12f01 g42599 ( .a(n8066), .b(n46390), .c(n46389), .o(n46391) );
na02f01 g42600 ( .a(n46391), .b(n46388), .o(n4888) );
na02f01 g42601 ( .a(n32732), .b(sin_out_7), .o(n46393) );
no03f01 g42602 ( .a(n36593), .b(n38999), .c(n38592), .o(n46394) );
in01f01 g42603 ( .a(n46394), .o(n46395) );
no02f01 g42604 ( .a(n36589), .b(n34307), .o(n46396) );
no02f01 g42605 ( .a(n46396), .b(n36591), .o(n46397) );
in01f01 g42606 ( .a(n46397), .o(n46398) );
no02f01 g42607 ( .a(n46398), .b(n46395), .o(n46399) );
no02f01 g42608 ( .a(n46397), .b(n46394), .o(n46400) );
oa12f01 g42609 ( .a(n32734), .b(n46400), .c(n46399), .o(n46401) );
na02f01 g42610 ( .a(n46401), .b(n46393), .o(n4893) );
na02f01 g42611 ( .a(n44108), .b(n44103), .o(n4897) );
na02f01 g42612 ( .a(n4171), .b(n4116), .o(n46404) );
na02f01 g42613 ( .a(n45720), .b(n2589), .o(n46405) );
na02f01 g42614 ( .a(n46405), .b(n46404), .o(n4902) );
in01f01 g42615 ( .a(n44979), .o(n46407) );
in01f01 g42616 ( .a(n10946), .o(n46408) );
na02f01 g42617 ( .a(n44977), .b(n46408), .o(n46409) );
no02f01 g42618 ( .a(n10951), .b(n3521), .o(n46410) );
no02f01 g42619 ( .a(n46410), .b(n10953), .o(n46411) );
na04f01 g42620 ( .a(n46411), .b(n46409), .c(n46407), .d(n44976), .o(n46412) );
na03f01 g42621 ( .a(n46409), .b(n46407), .c(n44976), .o(n46413) );
in01f01 g42622 ( .a(n46411), .o(n46414) );
na02f01 g42623 ( .a(n46414), .b(n46413), .o(n46415) );
na02f01 g42624 ( .a(n46415), .b(n46412), .o(n4912) );
oa12f01 g42625 ( .a(n11804), .b(n11785), .c(n41858), .o(n46417) );
no02f01 g42626 ( .a(n11809), .b(n11794), .o(n46418) );
in01f01 g42627 ( .a(n46418), .o(n46419) );
na02f01 g42628 ( .a(n46419), .b(n46417), .o(n46420) );
in01f01 g42629 ( .a(n46417), .o(n46421) );
na02f01 g42630 ( .a(n46418), .b(n46421), .o(n46422) );
na02f01 g42631 ( .a(n46422), .b(n46420), .o(n4917) );
no02f01 g42632 ( .a(n46417), .b(n11809), .o(n46424) );
no02f01 g42633 ( .a(n46424), .b(n11794), .o(n46425) );
no02f01 g42634 ( .a(n11807), .b(n11799), .o(n46426) );
in01f01 g42635 ( .a(n46426), .o(n46427) );
na02f01 g42636 ( .a(n46427), .b(n46425), .o(n46428) );
oa12f01 g42637 ( .a(n46426), .b(n46424), .c(n11794), .o(n46429) );
na02f01 g42638 ( .a(n46429), .b(n46428), .o(n4922) );
no02f01 g42639 ( .a(n42339), .b(n35535), .o(n46431) );
no02f01 g42640 ( .a(n42341), .b(n35485), .o(n46432) );
na02f01 g42641 ( .a(n46432), .b(n46431), .o(n46433) );
in01f01 g42642 ( .a(n46432), .o(n46434) );
oa12f01 g42643 ( .a(n46434), .b(n42339), .c(n35535), .o(n46435) );
na02f01 g42644 ( .a(n46435), .b(n46433), .o(n4927) );
na02f01 g42645 ( .a(n42320), .b(n2589), .o(n46437) );
na02f01 g42646 ( .a(n1754), .b(n4116), .o(n46438) );
na02f01 g42647 ( .a(n46438), .b(n46437), .o(n4937) );
na02f01 g42648 ( .a(n298), .b(n4116), .o(n46440) );
na02f01 g42649 ( .a(n22765), .b(n2589), .o(n46441) );
na02f01 g42650 ( .a(n46441), .b(n46440), .o(n4942) );
na03f01 g42651 ( .a(n42391), .b(n42387), .c(n_27923), .o(n46443) );
no03f01 g42652 ( .a(n42390), .b(n42378), .c(n41724), .o(n46444) );
ao12f01 g42653 ( .a(n42379), .b(n42386), .c(n42376), .o(n46445) );
oa12f01 g42654 ( .a(n34420), .b(n46445), .c(n46444), .o(n46446) );
na02f01 g42655 ( .a(n46446), .b(n46443), .o(n4947) );
in01f01 g42656 ( .a(n3040), .o(n4952) );
no02f01 g42657 ( .a(n6911), .b(cordic_combinational_sub_ln23_0_unr20_z_0_), .o(n46449) );
no02f01 g42658 ( .a(n6910), .b(n6079), .o(n46450) );
no02f01 g42659 ( .a(n46450), .b(n46449), .o(n46451) );
in01f01 g42660 ( .a(n46451), .o(n46452) );
no02f01 g42661 ( .a(n5001), .b(n46452), .o(n46453) );
no02f01 g42662 ( .a(n6934), .b(n46451), .o(n46454) );
no02f01 g42663 ( .a(n46454), .b(n46453), .o(n46455) );
na02f01 g42664 ( .a(n46455), .b(cordic_combinational_sub_ln23_0_unr20_z_0_), .o(n46456) );
oa12f01 g42665 ( .a(n6079), .b(n46454), .c(n46453), .o(n46457) );
na02f01 g42666 ( .a(n46457), .b(n46456), .o(n4957) );
na02f01 g42667 ( .a(n44974), .b(n1821), .o(n46459) );
na02f01 g42668 ( .a(n3545), .b(n8066), .o(n46460) );
na02f01 g42669 ( .a(n46460), .b(n46459), .o(n4962) );
no03f01 g42670 ( .a(n4251), .b(n9646), .c(n9645), .o(n46462) );
ao12f01 g42671 ( .a(n485), .b(n9590), .c(n9589), .o(n46463) );
no02f01 g42672 ( .a(n46463), .b(n46462), .o(n4967) );
no02f01 g42673 ( .a(n9795), .b(n39642), .o(n46465) );
no03f01 g42674 ( .a(n46465), .b(n40342), .c(n9775), .o(n46466) );
no02f01 g42675 ( .a(n9818), .b(n5001), .o(n46467) );
no02f01 g42676 ( .a(n46467), .b(n9787), .o(n46468) );
na02f01 g42677 ( .a(n46468), .b(n46466), .o(n46469) );
in01f01 g42678 ( .a(n46466), .o(n46470) );
in01f01 g42679 ( .a(n46468), .o(n46471) );
na02f01 g42680 ( .a(n46471), .b(n46470), .o(n46472) );
na02f01 g42681 ( .a(n46472), .b(n46469), .o(n4972) );
in01f01 g42682 ( .a(n11674), .o(n46474) );
no02f01 g42683 ( .a(n11675), .b(n46474), .o(n46475) );
no02f01 g42684 ( .a(n11688), .b(n11685), .o(n46476) );
na02f01 g42685 ( .a(n46476), .b(n46475), .o(n46477) );
in01f01 g42686 ( .a(n46476), .o(n46478) );
oa12f01 g42687 ( .a(n46478), .b(n11675), .c(n46474), .o(n46479) );
na02f01 g42688 ( .a(n46479), .b(n46477), .o(n4977) );
na02f01 g42689 ( .a(n3175), .b(n37149), .o(n46481) );
na03f01 g42690 ( .a(n46481), .b(n37362), .c(n44780), .o(n46482) );
na02f01 g42691 ( .a(n46481), .b(n37362), .o(n46483) );
na02f01 g42692 ( .a(n46483), .b(n44781), .o(n46484) );
na02f01 g42693 ( .a(n46484), .b(n46482), .o(n4982) );
oa22f01 g42694 ( .a(n30099), .b(n25793), .c(n25891), .d(n25886), .o(n46486) );
na04f01 g42695 ( .a(n25892), .b(n30095), .c(n30094), .d(n25794), .o(n46487) );
na02f01 g42696 ( .a(n46487), .b(n46486), .o(n4987) );
no02f01 g42697 ( .a(n43907), .b(n37391), .o(n46489) );
no02f01 g42698 ( .a(n43908), .b(n3623), .o(n46490) );
no02f01 g42699 ( .a(n46490), .b(n46489), .o(n46491) );
in01f01 g42700 ( .a(n46491), .o(n4992) );
na02f01 g42701 ( .a(n32732), .b(cos_out_29), .o(n46493) );
no04f01 g42702 ( .a(n41611), .b(n41589), .c(n41547), .d(n39712), .o(n46494) );
no02f01 g42703 ( .a(n45841), .b(n41636), .o(n46495) );
in01f01 g42704 ( .a(n46495), .o(n46496) );
no02f01 g42705 ( .a(n41638), .b(n35944), .o(n46497) );
no02f01 g42706 ( .a(n46497), .b(n41603), .o(n46498) );
in01f01 g42707 ( .a(n46498), .o(n46499) );
no03f01 g42708 ( .a(n46499), .b(n46496), .c(n46494), .o(n46500) );
in01f01 g42709 ( .a(n41611), .o(n46501) );
na04f01 g42710 ( .a(n46501), .b(n41588), .c(n41546), .d(n39691), .o(n46502) );
ao12f01 g42711 ( .a(n46498), .b(n46495), .c(n46502), .o(n46503) );
oa12f01 g42712 ( .a(n32734), .b(n46503), .c(n46500), .o(n46504) );
na02f01 g42713 ( .a(n46504), .b(n46493), .o(n4997) );
no02f01 g42714 ( .a(n40820), .b(n40817), .o(n46506) );
in01f01 g42715 ( .a(n46506), .o(n46507) );
no03f01 g42716 ( .a(n46507), .b(n42481), .c(n40827), .o(n46508) );
in01f01 g42717 ( .a(n46508), .o(n46509) );
oa12f01 g42718 ( .a(n46507), .b(n42481), .c(n40827), .o(n46510) );
na03f01 g42719 ( .a(n46510), .b(n46509), .c(n5799), .o(n46511) );
na02f01 g42720 ( .a(n46510), .b(n46509), .o(n5913) );
na02f01 g42721 ( .a(n5913), .b(n911), .o(n46513) );
na02f01 g42722 ( .a(n46513), .b(n46511), .o(n5006) );
no02f01 g42723 ( .a(n44857), .b(n9831), .o(n46515) );
na03f01 g42724 ( .a(n46515), .b(n9823), .c(n9817), .o(n46516) );
in01f01 g42725 ( .a(n46515), .o(n46517) );
oa12f01 g42726 ( .a(n46517), .b(n39645), .c(n39644), .o(n46518) );
na02f01 g42727 ( .a(n46518), .b(n46516), .o(n5011) );
no03f01 g42728 ( .a(n43373), .b(n42875), .c(n42869), .o(n46520) );
no02f01 g42729 ( .a(n42826), .b(n4176), .o(n46521) );
no02f01 g42730 ( .a(n46521), .b(n42876), .o(n46522) );
oa12f01 g42731 ( .a(n46522), .b(n46520), .c(n42877), .o(n46523) );
no02f01 g42732 ( .a(n46520), .b(n42877), .o(n46524) );
in01f01 g42733 ( .a(n46522), .o(n46525) );
na02f01 g42734 ( .a(n46525), .b(n46524), .o(n46526) );
na02f01 g42735 ( .a(n46526), .b(n46523), .o(n5016) );
no02f01 g42736 ( .a(n22735), .b(n22718), .o(n46528) );
in01f01 g42737 ( .a(n46528), .o(n46529) );
oa12f01 g42738 ( .a(n46529), .b(n22734), .c(n22706), .o(n46530) );
in01f01 g42739 ( .a(n22706), .o(n46531) );
na03f01 g42740 ( .a(n46528), .b(n22733), .c(n46531), .o(n46532) );
na02f01 g42741 ( .a(n46532), .b(n46530), .o(n5021) );
no02f01 g42742 ( .a(n40931), .b(n40929), .o(n46534) );
no02f01 g42743 ( .a(n46534), .b(n40882), .o(n46535) );
in01f01 g42744 ( .a(n40875), .o(n46536) );
na02f01 g42745 ( .a(n40876), .b(n46536), .o(n46537) );
in01f01 g42746 ( .a(n46537), .o(n46538) );
no02f01 g42747 ( .a(n46538), .b(n46535), .o(n46539) );
na02f01 g42748 ( .a(n46538), .b(n46535), .o(n46540) );
in01f01 g42749 ( .a(n46540), .o(n46541) );
no02f01 g42750 ( .a(n46541), .b(n46539), .o(n46542) );
in01f01 g42751 ( .a(n46542), .o(n5041) );
in01f01 g42752 ( .a(mux_while_ln12_psv_q_1_), .o(n46544) );
no02f01 g42753 ( .a(n45728), .b(n46544), .o(n5046) );
no02f01 g42754 ( .a(n32399), .b(n32173), .o(n46546) );
in01f01 g42755 ( .a(n46546), .o(n46547) );
na02f01 g42756 ( .a(n46547), .b(n43937), .o(n46548) );
na02f01 g42757 ( .a(n46546), .b(n43938), .o(n46549) );
na02f01 g42758 ( .a(n46549), .b(n46548), .o(n5056) );
na02f01 g42759 ( .a(n42515), .b(n5799), .o(n46551) );
na02f01 g42760 ( .a(n1874), .b(n911), .o(n46552) );
na02f01 g42761 ( .a(n46552), .b(n46551), .o(n5061) );
na03f01 g42762 ( .a(n27038), .b(n27232), .c(n26935), .o(n46554) );
oa12f01 g42763 ( .a(n27037), .b(n27039), .c(n26934), .o(n46555) );
na02f01 g42764 ( .a(n46555), .b(n46554), .o(n5066) );
in01f01 g42765 ( .a(n14155), .o(n46557) );
in01f01 g42766 ( .a(n14156), .o(n46558) );
no02f01 g42767 ( .a(n46558), .b(n14100), .o(n46559) );
na02f01 g42768 ( .a(n46559), .b(n46557), .o(n46560) );
oa12f01 g42769 ( .a(n14155), .b(n46558), .c(n14100), .o(n46561) );
na02f01 g42770 ( .a(n46561), .b(n46560), .o(n5075) );
no02f01 g42771 ( .a(n37871), .b(n37873), .o(n46563) );
no02f01 g42772 ( .a(n38010), .b(n38026), .o(n46564) );
no02f01 g42773 ( .a(n46564), .b(n46563), .o(n46565) );
no02f01 g42774 ( .a(n43382), .b(n43380), .o(n46566) );
no02f01 g42775 ( .a(n46566), .b(n43381), .o(n46567) );
na02f01 g42776 ( .a(n46567), .b(n46565), .o(n46568) );
in01f01 g42777 ( .a(n46565), .o(n46569) );
oa12f01 g42778 ( .a(n46569), .b(n46566), .c(n43381), .o(n46570) );
na03f01 g42779 ( .a(n46570), .b(n46568), .c(n1821), .o(n46571) );
na02f01 g42780 ( .a(n46570), .b(n46568), .o(n5760) );
na02f01 g42781 ( .a(n5760), .b(n8066), .o(n46573) );
na02f01 g42782 ( .a(n46573), .b(n46571), .o(n5085) );
na03f01 g42783 ( .a(n40969), .b(n9590), .c(n9589), .o(n46575) );
oa12f01 g42784 ( .a(n1195), .b(n9646), .c(n9645), .o(n46576) );
na02f01 g42785 ( .a(n46576), .b(n46575), .o(n5090) );
in01f01 g42786 ( .a(n45595), .o(n46578) );
no02f01 g42787 ( .a(n46578), .b(n936), .o(n46579) );
no02f01 g42788 ( .a(n45595), .b(n9228), .o(n46580) );
no02f01 g42789 ( .a(n46580), .b(n46579), .o(n46581) );
na03f01 g42790 ( .a(n46581), .b(n9590), .c(n9589), .o(n46582) );
in01f01 g42791 ( .a(n46581), .o(n5250) );
oa12f01 g42792 ( .a(n5250), .b(n9646), .c(n9645), .o(n46584) );
na02f01 g42793 ( .a(n46584), .b(n46582), .o(n5095) );
na03f01 g42794 ( .a(n42403), .b(n42399), .c(n6037), .o(n46586) );
ao12f01 g42795 ( .a(n42400), .b(n42402), .c(n25146), .o(n46587) );
no03f01 g42796 ( .a(n42398), .b(n42396), .c(n42393), .o(n46588) );
oa12f01 g42797 ( .a(n5873), .b(n46588), .c(n46587), .o(n46589) );
na02f01 g42798 ( .a(n46589), .b(n46586), .o(n5105) );
na02f01 g42799 ( .a(n42065), .b(n5799), .o(n46591) );
na02f01 g42800 ( .a(n1580), .b(n911), .o(n46592) );
na02f01 g42801 ( .a(n46592), .b(n46591), .o(n5110) );
no02f01 g42802 ( .a(n22657), .b(n22653), .o(n46594) );
in01f01 g42803 ( .a(n22681), .o(n46595) );
ao12f01 g42804 ( .a(n22669), .b(n46595), .c(n46594), .o(n46596) );
in01f01 g42805 ( .a(n46596), .o(n46597) );
no02f01 g42806 ( .a(n22682), .b(n22678), .o(n46598) );
na02f01 g42807 ( .a(n46598), .b(n46597), .o(n46599) );
in01f01 g42808 ( .a(n46598), .o(n46600) );
na02f01 g42809 ( .a(n46600), .b(n46596), .o(n46601) );
na02f01 g42810 ( .a(n46601), .b(n46599), .o(n5115) );
na04f01 g42811 ( .a(n39899), .b(n39898), .c(n39897), .d(n39327), .o(n46603) );
oa22f01 g42812 ( .a(n40043), .b(n39896), .c(n40041), .d(n39326), .o(n46604) );
na02f01 g42813 ( .a(n46604), .b(n46603), .o(n5120) );
no02f01 g42814 ( .a(n5981), .b(n5964), .o(n46606) );
no02f01 g42815 ( .a(n46606), .b(n41712), .o(n46607) );
no02f01 g42816 ( .a(n5971), .b(n5873), .o(n46608) );
no02f01 g42817 ( .a(n46608), .b(n5973_1), .o(n46609) );
na02f01 g42818 ( .a(n46609), .b(n46607), .o(n46610) );
in01f01 g42819 ( .a(n46609), .o(n46611) );
oa12f01 g42820 ( .a(n46611), .b(n46606), .c(n41712), .o(n46612) );
na02f01 g42821 ( .a(n46612), .b(n46610), .o(n5125) );
na02f01 g42822 ( .a(n3826), .b(n4116), .o(n46614) );
na03f01 g42823 ( .a(n45334), .b(n45333), .c(n2589), .o(n46615) );
na02f01 g42824 ( .a(n46615), .b(n46614), .o(n5130) );
no02f01 g42825 ( .a(n36142), .b(n44446), .o(n46617) );
no02f01 g42826 ( .a(n36161), .b(n36122), .o(n46618) );
no03f01 g42827 ( .a(n46618), .b(n36167), .c(n46617), .o(n46619) );
no02f01 g42828 ( .a(n46619), .b(n36163), .o(n46620) );
no02f01 g42829 ( .a(n36154), .b(n36122), .o(n46621) );
no02f01 g42830 ( .a(n46621), .b(n36156), .o(n46622) );
in01f01 g42831 ( .a(n46622), .o(n46623) );
na02f01 g42832 ( .a(n46623), .b(n46620), .o(n46624) );
oa12f01 g42833 ( .a(n46622), .b(n46619), .c(n36163), .o(n46625) );
na02f01 g42834 ( .a(n46625), .b(n46624), .o(n5135) );
no02f01 g42835 ( .a(n44336), .b(n44338), .o(n46627) );
oa12f01 g42836 ( .a(n46627), .b(n39145), .c(n39172), .o(n46628) );
in01f01 g42837 ( .a(n46628), .o(n46629) );
no02f01 g42838 ( .a(n39135), .b(n31515), .o(n46630) );
no02f01 g42839 ( .a(n46630), .b(n39144), .o(n46631) );
na02f01 g42840 ( .a(n46631), .b(n46629), .o(n46632) );
in01f01 g42841 ( .a(n46631), .o(n46633) );
na02f01 g42842 ( .a(n46633), .b(n46628), .o(n46634) );
na02f01 g42843 ( .a(n46634), .b(n46632), .o(n5140) );
na04f01 g42844 ( .a(n39477), .b(n39355), .c(n40001), .d(n40000), .o(n46636) );
oa22f01 g42845 ( .a(n40039), .b(n39354), .c(n39342), .d(n39338), .o(n46637) );
na02f01 g42846 ( .a(n46637), .b(n46636), .o(n5145) );
na03f01 g42847 ( .a(n46107), .b(n9590), .c(n9589), .o(n46639) );
oa12f01 g42848 ( .a(n4603), .b(n9646), .c(n9645), .o(n46640) );
na02f01 g42849 ( .a(n46640), .b(n46639), .o(n5150) );
no02f01 g42850 ( .a(n44489), .b(n41221), .o(n46642) );
na03f01 g42851 ( .a(n46642), .b(n44492), .c(n44488), .o(n46643) );
in01f01 g42852 ( .a(n46642), .o(n46644) );
oa12f01 g42853 ( .a(n46644), .b(n44495), .c(n41237), .o(n46645) );
na03f01 g42854 ( .a(n46645), .b(n46643), .c(n1821), .o(n46646) );
na02f01 g42855 ( .a(n46645), .b(n46643), .o(n5908) );
na02f01 g42856 ( .a(n5908), .b(n8066), .o(n46648) );
na02f01 g42857 ( .a(n46648), .b(n46646), .o(n5155) );
na02f01 g42858 ( .a(n46115), .b(n2589), .o(n46650) );
na02f01 g42859 ( .a(n4608), .b(n4116), .o(n46651) );
na02f01 g42860 ( .a(n46651), .b(n46650), .o(n5165) );
na03f01 g42861 ( .a(n42439), .b(n42435), .c(delay_sub_ln23_0_unr27_stage10_stallmux_z), .o(n46653) );
no03f01 g42862 ( .a(n42438), .b(n42437), .c(n42436), .o(n46654) );
ao12f01 g42863 ( .a(n42434), .b(n21593), .c(n42433), .o(n46655) );
oa12f01 g42864 ( .a(n21621), .b(n46655), .c(n46654), .o(n46656) );
na02f01 g42865 ( .a(n46656), .b(n46653), .o(n5170) );
no02f01 g42866 ( .a(n27114), .b(n27097), .o(n46658) );
no02f01 g42867 ( .a(n46658), .b(n43877), .o(n46659) );
in01f01 g42868 ( .a(n46659), .o(n46660) );
na02f01 g42869 ( .a(n46658), .b(n43877), .o(n46661) );
na02f01 g42870 ( .a(n46661), .b(n46660), .o(n5175) );
no02f01 g42871 ( .a(n42870), .b(n42866), .o(n46663) );
na02f01 g42872 ( .a(n46663), .b(n45087), .o(n46664) );
in01f01 g42873 ( .a(n46663), .o(n46665) );
oa12f01 g42874 ( .a(n46665), .b(n45086), .c(n45084), .o(n46666) );
na02f01 g42875 ( .a(n46666), .b(n46664), .o(n5180) );
no02f01 g42876 ( .a(n37871), .b(n26438), .o(n46668) );
no02f01 g42877 ( .a(n46668), .b(n41229), .o(n46669) );
in01f01 g42878 ( .a(n41231), .o(n46670) );
oa12f01 g42879 ( .a(n46670), .b(n41240), .c(n41228), .o(n46671) );
na03f01 g42880 ( .a(n46671), .b(n46669), .c(n41235), .o(n46672) );
in01f01 g42881 ( .a(n46669), .o(n46673) );
ao12f01 g42882 ( .a(n41231), .b(n41239), .c(n41248), .o(n46674) );
oa12f01 g42883 ( .a(n46673), .b(n46674), .c(n41234), .o(n46675) );
na03f01 g42884 ( .a(n46675), .b(n46672), .c(n1821), .o(n46676) );
no03f01 g42885 ( .a(n46674), .b(n46673), .c(n41234), .o(n46677) );
ao12f01 g42886 ( .a(n46669), .b(n46671), .c(n41235), .o(n46678) );
oa12f01 g42887 ( .a(n8066), .b(n46678), .c(n46677), .o(n46679) );
na02f01 g42888 ( .a(n46679), .b(n46676), .o(n5185) );
na02f01 g42889 ( .a(n46542), .b(n5799), .o(n46681) );
na02f01 g42890 ( .a(n5041), .b(n911), .o(n46682) );
na02f01 g42891 ( .a(n46682), .b(n46681), .o(n5190) );
no03f01 g42892 ( .a(n43313), .b(n40581), .c(n40591), .o(n46684) );
no02f01 g42893 ( .a(n39860), .b(n28982), .o(n46685) );
no02f01 g42894 ( .a(n46685), .b(n40566), .o(n46686) );
oa12f01 g42895 ( .a(n46686), .b(n46684), .c(n40564), .o(n46687) );
in01f01 g42896 ( .a(n40564), .o(n46688) );
in01f01 g42897 ( .a(n43313), .o(n46689) );
na03f01 g42898 ( .a(n46689), .b(n40582), .c(n40578), .o(n46690) );
in01f01 g42899 ( .a(n46686), .o(n46691) );
na03f01 g42900 ( .a(n46691), .b(n46690), .c(n46688), .o(n46692) );
na03f01 g42901 ( .a(n46692), .b(n46687), .c(n_27923), .o(n46693) );
ao12f01 g42902 ( .a(n46691), .b(n46690), .c(n46688), .o(n46694) );
no03f01 g42903 ( .a(n46686), .b(n46684), .c(n40564), .o(n46695) );
oa12f01 g42904 ( .a(n34420), .b(n46695), .c(n46694), .o(n46696) );
na02f01 g42905 ( .a(n46696), .b(n46693), .o(n5200) );
no02f01 g42906 ( .a(n22735), .b(n22734), .o(n46698) );
oa12f01 g42907 ( .a(n46698), .b(n22718), .c(n46531), .o(n46699) );
no02f01 g42908 ( .a(n22736), .b(n22729), .o(n46700) );
in01f01 g42909 ( .a(n46700), .o(n46701) );
na02f01 g42910 ( .a(n46701), .b(n46699), .o(n46702) );
in01f01 g42911 ( .a(n46699), .o(n46703) );
na02f01 g42912 ( .a(n46700), .b(n46703), .o(n46704) );
na02f01 g42913 ( .a(n46704), .b(n46702), .o(n5205) );
no02f01 g42914 ( .a(n37357), .b(n37353), .o(n46706) );
ao12f01 g42915 ( .a(delay_sub_ln23_0_unr23_stage8_stallmux_q), .b(n37349), .c(n37348), .o(n46707) );
oa12f01 g42916 ( .a(n46706), .b(n46707), .c(n37350), .o(n46708) );
no02f01 g42917 ( .a(n46707), .b(n37350), .o(n46709) );
oa12f01 g42918 ( .a(n46709), .b(n37357), .c(n37353), .o(n46710) );
na02f01 g42919 ( .a(n46710), .b(n46708), .o(n5225) );
na03f01 g42920 ( .a(n4993), .b(n4969), .c(n4924), .o(n46712) );
oa12f01 g42921 ( .a(n4992_1), .b(n4970), .c(n4977_1), .o(n46713) );
na02f01 g42922 ( .a(n46713), .b(n46712), .o(n5230) );
na03f01 g42923 ( .a(n43516), .b(n9590), .c(n9589), .o(n46715) );
oa12f01 g42924 ( .a(n2516), .b(n9646), .c(n9645), .o(n46716) );
na02f01 g42925 ( .a(n46716), .b(n46715), .o(n5235) );
in01f01 g42926 ( .a(n32655), .o(n46718) );
in01f01 g42927 ( .a(n32650), .o(n46719) );
no02f01 g42928 ( .a(n32711), .b(n46719), .o(n46720) );
no02f01 g42929 ( .a(n32662), .b(n32650), .o(n46721) );
oa12f01 g42930 ( .a(n46718), .b(n46721), .c(n46720), .o(n46722) );
no02f01 g42931 ( .a(n46721), .b(n46720), .o(n46723) );
na02f01 g42932 ( .a(n46723), .b(n32655), .o(n46724) );
na02f01 g42933 ( .a(n46724), .b(n46722), .o(n5240) );
no02f01 g42934 ( .a(n41405), .b(n8506), .o(n46726) );
in01f01 g42935 ( .a(n46726), .o(n46727) );
na02f01 g42936 ( .a(n46727), .b(n37800), .o(n46728) );
na02f01 g42937 ( .a(n46726), .b(n37801), .o(n46729) );
na02f01 g42938 ( .a(n46729), .b(n46728), .o(n5245) );
no02f01 g42939 ( .a(n22693), .b(n38574), .o(n46731) );
no02f01 g42940 ( .a(n46731), .b(n22731), .o(n46732) );
no02f01 g42941 ( .a(n22732), .b(n22703), .o(n46733) );
na02f01 g42942 ( .a(n46733), .b(n46732), .o(n46734) );
in01f01 g42943 ( .a(n46733), .o(n46735) );
oa12f01 g42944 ( .a(n46735), .b(n46731), .c(n22731), .o(n46736) );
na02f01 g42945 ( .a(n46736), .b(n46734), .o(n5260) );
na03f01 g42946 ( .a(n27363), .b(n27661), .c(n27311), .o(n46738) );
oa12f01 g42947 ( .a(n27360), .b(n27362), .c(n27310), .o(n46739) );
na02f01 g42948 ( .a(n46739), .b(n46738), .o(n5265) );
oa12f01 g42949 ( .a(n32319), .b(n32455), .c(n32454), .o(n46741) );
na02f01 g42950 ( .a(n46741), .b(n32321), .o(n5270) );
oa12f01 g42951 ( .a(n38784), .b(n36167), .c(n44445), .o(n46743) );
no02f01 g42952 ( .a(n46618), .b(n36163), .o(n46744) );
na02f01 g42953 ( .a(n46744), .b(n46743), .o(n46745) );
in01f01 g42954 ( .a(n46743), .o(n46746) );
in01f01 g42955 ( .a(n46744), .o(n46747) );
na02f01 g42956 ( .a(n46747), .b(n46746), .o(n46748) );
na02f01 g42957 ( .a(n46748), .b(n46745), .o(n5275) );
na03f01 g42958 ( .a(n44455), .b(n9590), .c(n9589), .o(n46750) );
oa12f01 g42959 ( .a(n3180), .b(n9646), .c(n9645), .o(n46751) );
na02f01 g42960 ( .a(n46751), .b(n46750), .o(n5280) );
ao12f01 g42961 ( .a(n37983), .b(n37988), .c(n37973), .o(n46753) );
in01f01 g42962 ( .a(n46753), .o(n46754) );
no02f01 g42963 ( .a(n37986), .b(n37942), .o(n46755) );
na02f01 g42964 ( .a(n46755), .b(n46754), .o(n46756) );
in01f01 g42965 ( .a(n46755), .o(n46757) );
na02f01 g42966 ( .a(n46757), .b(n46753), .o(n46758) );
na02f01 g42967 ( .a(n46758), .b(n46756), .o(n5285) );
na03f01 g42968 ( .a(n37972), .b(n38037), .c(n38034), .o(n46760) );
oa12f01 g42969 ( .a(n37971), .b(n38038), .c(n37956), .o(n46761) );
na02f01 g42970 ( .a(n46761), .b(n46760), .o(n5295) );
na02f01 g42971 ( .a(n1105), .b(n4116), .o(n46763) );
na03f01 g42972 ( .a(n40491), .b(n40489), .c(n2589), .o(n46764) );
na02f01 g42973 ( .a(n46764), .b(n46763), .o(n5300) );
no02f01 g42974 ( .a(n39988), .b(n40419), .o(n46766) );
oa12f01 g42975 ( .a(n46766), .b(n39968), .c(n40047), .o(n46767) );
in01f01 g42976 ( .a(n46767), .o(n46768) );
no02f01 g42977 ( .a(n39958), .b(n39860), .o(n46769) );
no02f01 g42978 ( .a(n46769), .b(n39960), .o(n46770) );
na02f01 g42979 ( .a(n46770), .b(n46768), .o(n46771) );
in01f01 g42980 ( .a(n46770), .o(n46772) );
na02f01 g42981 ( .a(n46772), .b(n46767), .o(n46773) );
na02f01 g42982 ( .a(n46773), .b(n46771), .o(n5305) );
na03f01 g42983 ( .a(n37400), .b(n9590), .c(n9589), .o(n46775) );
oa12f01 g42984 ( .a(n559), .b(n9646), .c(n9645), .o(n46776) );
na02f01 g42985 ( .a(n46776), .b(n46775), .o(n5310) );
no02f01 g42986 ( .a(n9225), .b(n8765), .o(n46778) );
no02f01 g42987 ( .a(n9224), .b(n8765), .o(n46779) );
no02f01 g42988 ( .a(n46779), .b(n46778), .o(n46780) );
na03f01 g42989 ( .a(n46780), .b(n9590), .c(n9589), .o(n46781) );
in01f01 g42990 ( .a(n46780), .o(n5888) );
oa12f01 g42991 ( .a(n5888), .b(n9646), .c(n9645), .o(n46783) );
na02f01 g42992 ( .a(n46783), .b(n46781), .o(n5315) );
na02f01 g42993 ( .a(n490), .b(n4116), .o(n46785) );
na03f01 g42994 ( .a(n36513), .b(n36495), .c(n2589), .o(n46786) );
na02f01 g42995 ( .a(n46786), .b(n46785), .o(n5320) );
oa12f01 g42996 ( .a(n40029), .b(n39473), .c(n39466), .o(n46788) );
na03f01 g42997 ( .a(n40032), .b(n40030), .c(n39452), .o(n46789) );
na02f01 g42998 ( .a(n46789), .b(n46788), .o(n5325) );
in01f01 g42999 ( .a(n38153), .o(n46791) );
in01f01 g43000 ( .a(n38152), .o(n46792) );
na02f01 g43001 ( .a(n46792), .b(n38162), .o(n46793) );
no02f01 g43002 ( .a(n40306), .b(n6037), .o(n46794) );
no02f01 g43003 ( .a(n46794), .b(n40299), .o(n46795) );
na03f01 g43004 ( .a(n46795), .b(n46793), .c(n46791), .o(n46796) );
oa12f01 g43005 ( .a(n46791), .b(n38152), .c(n38143), .o(n46797) );
in01f01 g43006 ( .a(n46795), .o(n46798) );
na02f01 g43007 ( .a(n46798), .b(n46797), .o(n46799) );
na02f01 g43008 ( .a(n46799), .b(n46796), .o(n5335) );
na02f01 g43009 ( .a(n37349), .b(n37348), .o(n5340) );
na03f01 g43010 ( .a(n46237), .b(n9590), .c(n9589), .o(n46802) );
oa12f01 g43011 ( .a(n4722), .b(n9646), .c(n9645), .o(n46803) );
na02f01 g43012 ( .a(n46803), .b(n46802), .o(n5350) );
in01f01 g43013 ( .a(n46169), .o(n46805) );
na02f01 g43014 ( .a(n46171), .b(n46170), .o(n46806) );
in01f01 g43015 ( .a(n46806), .o(n46807) );
na03f01 g43016 ( .a(n46807), .b(n16437), .c(n46805), .o(n46808) );
in01f01 g43017 ( .a(n16437), .o(n46809) );
oa12f01 g43018 ( .a(n46806), .b(n46809), .c(n46169), .o(n46810) );
na02f01 g43019 ( .a(n46810), .b(n46808), .o(n5355) );
ao12f01 g43020 ( .a(n44657), .b(n44659), .c(n44656), .o(n46812) );
no03f01 g43021 ( .a(n44654), .b(n44653), .c(n36761), .o(n46813) );
oa12f01 g43022 ( .a(n34420), .b(n46813), .c(n46812), .o(n46814) );
na03f01 g43023 ( .a(n44660), .b(n44655), .c(n_27923), .o(n46815) );
na02f01 g43024 ( .a(n46815), .b(n46814), .o(n5360) );
no03f01 g43025 ( .a(n42406), .b(n9581), .c(n9579), .o(n46817) );
no02f01 g43026 ( .a(n9583), .b(n9565), .o(n46818) );
oa12f01 g43027 ( .a(n46818), .b(n46817), .c(n9573), .o(n46819) );
no02f01 g43028 ( .a(n46817), .b(n9573), .o(n46820) );
in01f01 g43029 ( .a(n46818), .o(n46821) );
na02f01 g43030 ( .a(n46821), .b(n46820), .o(n46822) );
na02f01 g43031 ( .a(n46822), .b(n46819), .o(n5365) );
no02f01 g43032 ( .a(n29937), .b(n24598), .o(n46824) );
no02f01 g43033 ( .a(n46824), .b(n30038), .o(n46825) );
in01f01 g43034 ( .a(n30039), .o(n46826) );
in01f01 g43035 ( .a(n30045), .o(n46827) );
ao12f01 g43036 ( .a(n46827), .b(n46826), .c(n36520), .o(n46828) );
oa12f01 g43037 ( .a(n46825), .b(n46828), .c(n30040), .o(n46829) );
in01f01 g43038 ( .a(n30040), .o(n46830) );
in01f01 g43039 ( .a(n46825), .o(n46831) );
oa12f01 g43040 ( .a(n30045), .b(n30039), .c(n40213), .o(n46832) );
na03f01 g43041 ( .a(n46832), .b(n46831), .c(n46830), .o(n46833) );
na03f01 g43042 ( .a(n46833), .b(n46829), .c(n6037), .o(n46834) );
ao12f01 g43043 ( .a(n46831), .b(n46832), .c(n46830), .o(n46835) );
no03f01 g43044 ( .a(n46828), .b(n46825), .c(n30040), .o(n46836) );
oa12f01 g43045 ( .a(n5873), .b(n46836), .c(n46835), .o(n46837) );
na02f01 g43046 ( .a(n46837), .b(n46834), .o(n5370) );
na03f01 g43047 ( .a(n485), .b(n9590), .c(n9589), .o(n46839) );
oa12f01 g43048 ( .a(n4251), .b(n9646), .c(n9645), .o(n46840) );
na02f01 g43049 ( .a(n46840), .b(n46839), .o(n5375) );
no02f01 g43050 ( .a(n25296), .b(n25561), .o(n46842) );
in01f01 g43051 ( .a(n46842), .o(n46843) );
no02f01 g43052 ( .a(n46843), .b(n37134), .o(n46844) );
in01f01 g43053 ( .a(n46844), .o(n46845) );
na02f01 g43054 ( .a(n46843), .b(n37134), .o(n46846) );
na02f01 g43055 ( .a(n46846), .b(n46845), .o(n5390) );
na02f01 g43056 ( .a(n41211), .b(n41203), .o(n5395) );
in01f01 g43057 ( .a(n21260), .o(n46849) );
ao12f01 g43058 ( .a(n45367), .b(n46849), .c(n45365), .o(n46850) );
na02f01 g43059 ( .a(n20993), .b(n20988), .o(n46851) );
in01f01 g43060 ( .a(n46851), .o(n46852) );
no02f01 g43061 ( .a(n46852), .b(n46850), .o(n46853) );
na02f01 g43062 ( .a(n46852), .b(n46850), .o(n46854) );
in01f01 g43063 ( .a(n46854), .o(n46855) );
no02f01 g43064 ( .a(n46855), .b(n46853), .o(n46856) );
in01f01 g43065 ( .a(n46856), .o(n5400) );
na02f01 g43066 ( .a(n46833), .b(n46829), .o(n5405) );
no02f01 g43067 ( .a(n9231), .b(n936), .o(n46859) );
no02f01 g43068 ( .a(n9232), .b(n9228), .o(n46860) );
no02f01 g43069 ( .a(n46860), .b(n46859), .o(n46861) );
in01f01 g43070 ( .a(n46861), .o(n5410) );
no02f01 g43071 ( .a(n41123), .b(n41121), .o(n46863) );
in01f01 g43072 ( .a(n46863), .o(n46864) );
na02f01 g43073 ( .a(n46864), .b(n41120), .o(n46865) );
oa12f01 g43074 ( .a(n46863), .b(n27401), .c(n27394), .o(n46866) );
na02f01 g43075 ( .a(n46866), .b(n46865), .o(n5415) );
na03f01 g43076 ( .a(n27660), .b(n27358), .c(n27324), .o(n46868) );
oa12f01 g43077 ( .a(n27659), .b(n27359), .c(n27645), .o(n46869) );
na02f01 g43078 ( .a(n46869), .b(n46868), .o(n5435) );
na03f01 g43079 ( .a(n44698), .b(n44696), .c(n3633), .o(n46871) );
na02f01 g43080 ( .a(n3337), .b(n6203), .o(n46872) );
na02f01 g43081 ( .a(n46872), .b(n46871), .o(n5445) );
no02f01 g43082 ( .a(n22681), .b(n22669), .o(n46874) );
na02f01 g43083 ( .a(n46874), .b(n46594), .o(n46875) );
in01f01 g43084 ( .a(n46874), .o(n46876) );
oa12f01 g43085 ( .a(n46876), .b(n22657), .c(n22653), .o(n46877) );
na02f01 g43086 ( .a(n46877), .b(n46875), .o(n5450) );
na02f01 g43087 ( .a(n32732), .b(cos_out_24), .o(n46879) );
na02f01 g43088 ( .a(n41546), .b(n39691), .o(n46880) );
in01f01 g43089 ( .a(n41629), .o(n46881) );
na02f01 g43090 ( .a(n46881), .b(n46880), .o(n46882) );
no02f01 g43091 ( .a(n43021), .b(n41568), .o(n46883) );
in01f01 g43092 ( .a(n46883), .o(n46884) );
no02f01 g43093 ( .a(n46884), .b(n46882), .o(n46885) );
ao12f01 g43094 ( .a(n46883), .b(n46881), .c(n46880), .o(n46886) );
oa12f01 g43095 ( .a(n32734), .b(n46886), .c(n46885), .o(n46887) );
na02f01 g43096 ( .a(n46887), .b(n46879), .o(n5455) );
no02f01 g43097 ( .a(n21589), .b(n16329), .o(n46889) );
no02f01 g43098 ( .a(n46889), .b(n21549), .o(n46890) );
no03f01 g43099 ( .a(n21557), .b(n21526), .c(n42235), .o(n46891) );
no03f01 g43100 ( .a(n46010), .b(n21586), .c(n21585), .o(n46892) );
in01f01 g43101 ( .a(n46892), .o(n46893) );
no02f01 g43102 ( .a(n46893), .b(n46891), .o(n46894) );
na02f01 g43103 ( .a(n46894), .b(n46890), .o(n46895) );
in01f01 g43104 ( .a(n46890), .o(n46896) );
oa12f01 g43105 ( .a(n46896), .b(n46893), .c(n46891), .o(n46897) );
na02f01 g43106 ( .a(n46897), .b(n46895), .o(n5459) );
in01f01 g43107 ( .a(n8758), .o(n46899) );
no02f01 g43108 ( .a(n45747), .b(n45748), .o(n46900) );
na03f01 g43109 ( .a(n46900), .b(n46899), .c(n8717), .o(n46901) );
in01f01 g43110 ( .a(n46900), .o(n46902) );
oa12f01 g43111 ( .a(n46902), .b(n8758), .c(n8716), .o(n46903) );
na02f01 g43112 ( .a(n46903), .b(n46901), .o(n5464) );
na02f01 g43113 ( .a(n44685), .b(n44680), .o(n5469) );
na02f01 g43114 ( .a(n32732), .b(sin_out_21), .o(n46906) );
no02f01 g43115 ( .a(n41364), .b(n34307), .o(n46907) );
no02f01 g43116 ( .a(n46907), .b(n41332), .o(n46908) );
in01f01 g43117 ( .a(n46908), .o(n46909) );
no02f01 g43118 ( .a(n41324), .b(n43431), .o(n46910) );
in01f01 g43119 ( .a(n45783), .o(n46911) );
na02f01 g43120 ( .a(n46911), .b(n41361), .o(n46912) );
no03f01 g43121 ( .a(n46912), .b(n46910), .c(n46909), .o(n46913) );
no02f01 g43122 ( .a(n46912), .b(n46910), .o(n46914) );
no02f01 g43123 ( .a(n46914), .b(n46908), .o(n46915) );
oa12f01 g43124 ( .a(n32734), .b(n46915), .c(n46913), .o(n46916) );
na02f01 g43125 ( .a(n46916), .b(n46906), .o(n5479) );
no02f01 g43126 ( .a(n5897), .b(cordic_combinational_sub_ln23_0_unr12_z_0_), .o(n46918) );
na02f01 g43127 ( .a(n5897), .b(cordic_combinational_sub_ln23_0_unr12_z_0_), .o(n46919) );
in01f01 g43128 ( .a(n46919), .o(n46920) );
no02f01 g43129 ( .a(n46920), .b(n46918), .o(n46921) );
in01f01 g43130 ( .a(n46921), .o(n46922) );
no02f01 g43131 ( .a(n46922), .b(n6037), .o(n46923) );
no02f01 g43132 ( .a(n46921), .b(n5873), .o(n46924) );
no02f01 g43133 ( .a(n46924), .b(n46923), .o(n46925) );
na02f01 g43134 ( .a(n46925), .b(cordic_combinational_sub_ln23_0_unr12_z_0_), .o(n46926) );
oa12f01 g43135 ( .a(n5151), .b(n46924), .c(n46923), .o(n46927) );
na02f01 g43136 ( .a(n46927), .b(n46926), .o(n5483) );
in01f01 g43137 ( .a(n11707), .o(n46929) );
ao12f01 g43138 ( .a(n11706), .b(n46929), .c(n11696), .o(n46930) );
in01f01 g43139 ( .a(n11717), .o(n46931) );
no02f01 g43140 ( .a(n46931), .b(n11714), .o(n46932) );
in01f01 g43141 ( .a(n46932), .o(n46933) );
na02f01 g43142 ( .a(n46933), .b(n46930), .o(n46934) );
in01f01 g43143 ( .a(n46930), .o(n46935) );
na02f01 g43144 ( .a(n46932), .b(n46935), .o(n46936) );
na02f01 g43145 ( .a(n46936), .b(n46934), .o(n5488) );
na02f01 g43146 ( .a(n39823), .b(n6037), .o(n46938) );
na02f01 g43147 ( .a(n906), .b(n5873), .o(n46939) );
na02f01 g43148 ( .a(n46939), .b(n46938), .o(n5498) );
no02f01 g43149 ( .a(n39008), .b(n39010), .o(n46941) );
no02f01 g43150 ( .a(n8672), .b(n5973), .o(n46942) );
no02f01 g43151 ( .a(n46942), .b(n8636), .o(n46943) );
oa12f01 g43152 ( .a(n46943), .b(n46941), .c(n8659), .o(n46944) );
no02f01 g43153 ( .a(n46941), .b(n8659), .o(n46945) );
in01f01 g43154 ( .a(n46943), .o(n46946) );
na02f01 g43155 ( .a(n46946), .b(n46945), .o(n46947) );
na02f01 g43156 ( .a(n46947), .b(n46944), .o(n5503) );
na03f01 g43157 ( .a(n45435), .b(n45432), .c(n5799), .o(n46949) );
no03f01 g43158 ( .a(n45430), .b(n45434), .c(n45433), .o(n46950) );
ao12f01 g43159 ( .a(n45426), .b(n45431), .c(n45428), .o(n46951) );
oa12f01 g43160 ( .a(n911), .b(n46951), .c(n46950), .o(n46952) );
na02f01 g43161 ( .a(n46952), .b(n46949), .o(n5508) );
ao12f01 g43162 ( .a(n45494), .b(n16432), .c(n16155), .o(n46954) );
na02f01 g43163 ( .a(n45495), .b(n45493), .o(n46955) );
in01f01 g43164 ( .a(n46955), .o(n46956) );
na02f01 g43165 ( .a(n46956), .b(n46954), .o(n46957) );
in01f01 g43166 ( .a(n46954), .o(n46958) );
na02f01 g43167 ( .a(n46955), .b(n46958), .o(n46959) );
na02f01 g43168 ( .a(n46959), .b(n46957), .o(n5513) );
no02f01 g43169 ( .a(n40074), .b(n40073), .o(n46961) );
na02f01 g43170 ( .a(n46961), .b(n40202), .o(n46962) );
in01f01 g43171 ( .a(n46961), .o(n46963) );
na02f01 g43172 ( .a(n46963), .b(n40072), .o(n46964) );
na02f01 g43173 ( .a(n46964), .b(n46962), .o(n5518) );
na03f01 g43174 ( .a(n42104), .b(n42102), .c(n1821), .o(n46966) );
na02f01 g43175 ( .a(n1610), .b(n8066), .o(n46967) );
na02f01 g43176 ( .a(n46967), .b(n46966), .o(n5523) );
no02f01 g43177 ( .a(n43784), .b(n42023), .o(n46969) );
na02f01 g43178 ( .a(n46969), .b(n42009), .o(n46970) );
ao12f01 g43179 ( .a(n3521), .b(n43785), .c(n42024), .o(n46971) );
no02f01 g43180 ( .a(n46971), .b(n42028), .o(n46972) );
in01f01 g43181 ( .a(n43779), .o(n46973) );
ao12f01 g43182 ( .a(n10727), .b(n43778), .c(n46973), .o(n46974) );
no02f01 g43183 ( .a(n10730), .b(n4088), .o(n46975) );
no02f01 g43184 ( .a(n46975), .b(n10718), .o(n46976) );
in01f01 g43185 ( .a(n46976), .o(n46977) );
no02f01 g43186 ( .a(n46977), .b(n46974), .o(n46978) );
na02f01 g43187 ( .a(n46977), .b(n46974), .o(n46979) );
in01f01 g43188 ( .a(n46979), .o(n46980) );
no02f01 g43189 ( .a(n46980), .b(n46978), .o(n46981) );
no02f01 g43190 ( .a(n46981), .b(n3521), .o(n46982) );
in01f01 g43191 ( .a(n46981), .o(n46983) );
no02f01 g43192 ( .a(n46983), .b(n10735), .o(n46984) );
no02f01 g43193 ( .a(n46984), .b(n46982), .o(n46985) );
na03f01 g43194 ( .a(n46985), .b(n46972), .c(n46970), .o(n46986) );
na02f01 g43195 ( .a(n46972), .b(n46970), .o(n46987) );
in01f01 g43196 ( .a(n46985), .o(n46988) );
na02f01 g43197 ( .a(n46988), .b(n46987), .o(n46989) );
na02f01 g43198 ( .a(n46989), .b(n46986), .o(n5528) );
in01f01 g43199 ( .a(n40293), .o(n46991) );
na03f01 g43200 ( .a(n40300), .b(n46991), .c(n38162), .o(n46992) );
no02f01 g43201 ( .a(n40291), .b(n6037), .o(n46993) );
no02f01 g43202 ( .a(n46993), .b(n40307), .o(n46994) );
no02f01 g43203 ( .a(n40283), .b(n6037), .o(n46995) );
no02f01 g43204 ( .a(n46995), .b(n40285), .o(n46996) );
na03f01 g43205 ( .a(n46996), .b(n46994), .c(n46992), .o(n46997) );
no03f01 g43206 ( .a(n40301), .b(n40293), .c(n38143), .o(n46998) );
in01f01 g43207 ( .a(n46994), .o(n46999) );
in01f01 g43208 ( .a(n46996), .o(n47000) );
oa12f01 g43209 ( .a(n47000), .b(n46999), .c(n46998), .o(n47001) );
na02f01 g43210 ( .a(n47001), .b(n46997), .o(n5533) );
oa12f01 g43211 ( .a(n38378), .b(n39095), .c(n39094), .o(n47003) );
na03f01 g43212 ( .a(n38377), .b(n38373), .c(n38372), .o(n47004) );
na02f01 g43213 ( .a(n47004), .b(n47003), .o(n5538) );
oa12f01 g43214 ( .a(n42662), .b(n39129), .c(n38468), .o(n47006) );
na03f01 g43215 ( .a(n38505), .b(n39126), .c(n42663), .o(n47007) );
na02f01 g43216 ( .a(n47007), .b(n47006), .o(n5543) );
na03f01 g43217 ( .a(n42257), .b(n42255), .c(n6037), .o(n47009) );
in01f01 g43218 ( .a(n42255), .o(n47010) );
oa12f01 g43219 ( .a(n5873), .b(n42256), .c(n47010), .o(n47011) );
na02f01 g43220 ( .a(n47011), .b(n47009), .o(n5553) );
na03f01 g43221 ( .a(n32463), .b(n32327), .c(n32280), .o(n47013) );
oa12f01 g43222 ( .a(n32462), .b(n32331), .c(n32279), .o(n47014) );
na02f01 g43223 ( .a(n47014), .b(n47013), .o(n5558) );
no02f01 g43224 ( .a(n45097), .b(n35529), .o(n47016) );
na02f01 g43225 ( .a(n47016), .b(n45103), .o(n47017) );
in01f01 g43226 ( .a(n47016), .o(n47018) );
na02f01 g43227 ( .a(n47018), .b(n45102), .o(n47019) );
na02f01 g43228 ( .a(n47019), .b(n47017), .o(n5563) );
ao12f01 g43229 ( .a(n32724), .b(n32720), .c(n32694), .o(n47021) );
in01f01 g43230 ( .a(n47021), .o(n47022) );
na03f01 g43231 ( .a(n47022), .b(n32726), .c(n32590), .o(n47023) );
oa12f01 g43232 ( .a(n47021), .b(n32680), .c(n32693), .o(n47024) );
na02f01 g43233 ( .a(n47024), .b(n47023), .o(n5568) );
in01f01 g43234 ( .a(n21182), .o(n47026) );
oa12f01 g43235 ( .a(n21181), .b(n47026), .c(n21141), .o(n47027) );
na04f01 g43236 ( .a(n21182), .b(n21180), .c(n21178), .d(n21142), .o(n47028) );
na02f01 g43237 ( .a(n47028), .b(n47027), .o(n5573) );
na02f01 g43238 ( .a(n45449), .b(n45448), .o(n5583) );
ao12f01 g43239 ( .a(delay_sub_ln23_0_unr23_stage8_stallmux_q), .b(n42452), .c(n42451), .o(n47031) );
oa12f01 g43240 ( .a(n38810), .b(n47031), .c(n42453), .o(n47032) );
no02f01 g43241 ( .a(n47031), .b(n42453), .o(n47033) );
na02f01 g43242 ( .a(n47033), .b(n42450), .o(n47034) );
na02f01 g43243 ( .a(n47034), .b(n47032), .o(n5588) );
na04f01 g43244 ( .a(n21185), .b(n21183), .c(n21142), .d(n21131), .o(n47036) );
na02f01 g43245 ( .a(n21185), .b(n21131), .o(n47037) );
na02f01 g43246 ( .a(n47037), .b(n21184), .o(n47038) );
na02f01 g43247 ( .a(n47038), .b(n47036), .o(n5593) );
na03f01 g43248 ( .a(n39218), .b(n39213), .c(n5799), .o(n47040) );
no02f01 g43249 ( .a(n39217), .b(n39207), .o(n47041) );
no02f01 g43250 ( .a(n39212), .b(n39208), .o(n47042) );
oa12f01 g43251 ( .a(n911), .b(n47042), .c(n47041), .o(n47043) );
na02f01 g43252 ( .a(n47043), .b(n47040), .o(n5598) );
na02f01 g43253 ( .a(n45582), .b(n1821), .o(n47045) );
na02f01 g43254 ( .a(n4028), .b(n8066), .o(n47046) );
na02f01 g43255 ( .a(n47046), .b(n47045), .o(n5608) );
na03f01 g43256 ( .a(n7513), .b(n7529), .c(n7490), .o(n47048) );
oa12f01 g43257 ( .a(n7539), .b(n7491), .c(n7528), .o(n47049) );
na02f01 g43258 ( .a(n47049), .b(n47048), .o(n5613) );
no02f01 g43259 ( .a(n38798), .b(n38791), .o(n47051) );
ao12f01 g43260 ( .a(delay_sub_ln23_0_unr23_stage8_stallmux_q), .b(n38808), .c(n38803), .o(n47052) );
oa12f01 g43261 ( .a(n47051), .b(n47052), .c(n38809), .o(n47053) );
no02f01 g43262 ( .a(n47052), .b(n38809), .o(n47054) );
oa12f01 g43263 ( .a(n47054), .b(n38798), .c(n38791), .o(n47055) );
na02f01 g43264 ( .a(n47055), .b(n47053), .o(n5623) );
na02f01 g43265 ( .a(n32732), .b(cos_out_1), .o(n47057) );
no03f01 g43266 ( .a(n35932), .b(n35974), .c(n35970), .o(n47058) );
ao12f01 g43267 ( .a(n35930), .b(n35975), .c(n35920), .o(n47059) );
oa12f01 g43268 ( .a(n32734), .b(n47059), .c(n47058), .o(n47060) );
na02f01 g43269 ( .a(n47060), .b(n47057), .o(n5653) );
na03f01 g43270 ( .a(n46154), .b(n46152), .c(n1821), .o(n47062) );
na02f01 g43271 ( .a(n4643), .b(n8066), .o(n47063) );
na02f01 g43272 ( .a(n47063), .b(n47062), .o(n5657) );
in01f01 g43273 ( .a(n42070), .o(n47065) );
no02f01 g43274 ( .a(n42072), .b(n37228), .o(n47066) );
na03f01 g43275 ( .a(n47066), .b(n37252), .c(n47065), .o(n47067) );
in01f01 g43276 ( .a(n47066), .o(n47068) );
oa12f01 g43277 ( .a(n47068), .b(n37253), .c(n42070), .o(n47069) );
na02f01 g43278 ( .a(n47069), .b(n47067), .o(n5662) );
in01f01 g43279 ( .a(n21585), .o(n47071) );
no02f01 g43280 ( .a(n42239), .b(n21502), .o(n47072) );
na03f01 g43281 ( .a(n47072), .b(n47071), .c(n42235), .o(n47073) );
in01f01 g43282 ( .a(n47072), .o(n47074) );
oa12f01 g43283 ( .a(n47074), .b(n21585), .c(n42236), .o(n47075) );
na02f01 g43284 ( .a(n47075), .b(n47073), .o(n5667) );
in01f01 g43285 ( .a(n25448), .o(n47077) );
no02f01 g43286 ( .a(n25458), .b(n47077), .o(n47078) );
na02f01 g43287 ( .a(n25458), .b(n47077), .o(n47079) );
in01f01 g43288 ( .a(n47079), .o(n47080) );
oa22f01 g43289 ( .a(n47080), .b(n47078), .c(n25444), .d(n25436), .o(n47081) );
in01f01 g43290 ( .a(n47078), .o(n47082) );
na03f01 g43291 ( .a(n47079), .b(n47082), .c(n25445), .o(n47083) );
na02f01 g43292 ( .a(n47083), .b(n47081), .o(n5672) );
na03f01 g43293 ( .a(n43233), .b(n9590), .c(n9589), .o(n47085) );
oa12f01 g43294 ( .a(n2287), .b(n9646), .c(n9645), .o(n47086) );
na02f01 g43295 ( .a(n47086), .b(n47085), .o(n5677) );
ao12f01 g43296 ( .a(n32414), .b(n32416), .c(n32489), .o(n47088) );
in01f01 g43297 ( .a(n47088), .o(n47089) );
no02f01 g43298 ( .a(n32137), .b(n31607), .o(n47090) );
no02f01 g43299 ( .a(n47090), .b(n32139), .o(n47091) );
na02f01 g43300 ( .a(n47091), .b(n47089), .o(n47092) );
in01f01 g43301 ( .a(n47091), .o(n47093) );
na02f01 g43302 ( .a(n47093), .b(n47088), .o(n47094) );
na02f01 g43303 ( .a(n47094), .b(n47092), .o(n5682) );
in01f01 g43304 ( .a(n21473), .o(n47096) );
na02f01 g43305 ( .a(n47096), .b(n21615), .o(n47097) );
no02f01 g43306 ( .a(n43946), .b(n43949), .o(n47098) );
no02f01 g43307 ( .a(n21463), .b(n16329), .o(n47099) );
no02f01 g43308 ( .a(n47099), .b(n21465), .o(n47100) );
na03f01 g43309 ( .a(n47100), .b(n47098), .c(n47097), .o(n47101) );
na02f01 g43310 ( .a(n47098), .b(n47097), .o(n47102) );
in01f01 g43311 ( .a(n47100), .o(n47103) );
na02f01 g43312 ( .a(n47103), .b(n47102), .o(n47104) );
na02f01 g43313 ( .a(n47104), .b(n47101), .o(n5687) );
na02f01 g43314 ( .a(n32732), .b(sin_out_16), .o(n47106) );
no02f01 g43315 ( .a(n39601), .b(n39554), .o(n47107) );
in01f01 g43316 ( .a(n47107), .o(n47108) );
no02f01 g43317 ( .a(n47108), .b(n41294), .o(n47109) );
no02f01 g43318 ( .a(n47107), .b(n39599), .o(n47110) );
oa12f01 g43319 ( .a(n32734), .b(n47110), .c(n47109), .o(n47111) );
na02f01 g43320 ( .a(n47111), .b(n47106), .o(n5697) );
in01f01 g43321 ( .a(n38948), .o(n47113) );
in01f01 g43322 ( .a(n38959), .o(n47114) );
na02f01 g43323 ( .a(n47114), .b(n38937), .o(n47115) );
no02f01 g43324 ( .a(n38961), .b(n38956), .o(n47116) );
in01f01 g43325 ( .a(n47116), .o(n47117) );
na03f01 g43326 ( .a(n47117), .b(n47115), .c(n47113), .o(n47118) );
na02f01 g43327 ( .a(n47115), .b(n47113), .o(n47119) );
na02f01 g43328 ( .a(n47116), .b(n47119), .o(n47120) );
na02f01 g43329 ( .a(n47120), .b(n47118), .o(n5701) );
na03f01 g43330 ( .a(n37160), .b(n37010), .c(n37009), .o(n47122) );
oa12f01 g43331 ( .a(n37158), .b(n37011), .c(n37157), .o(n47123) );
na02f01 g43332 ( .a(n47123), .b(n47122), .o(n5706) );
na03f01 g43333 ( .a(n46861), .b(n9590), .c(n9589), .o(n47125) );
oa12f01 g43334 ( .a(n5410), .b(n9646), .c(n9645), .o(n47126) );
na02f01 g43335 ( .a(n47126), .b(n47125), .o(n5711) );
na03f01 g43336 ( .a(n44081), .b(n44079), .c(n5799), .o(n47128) );
na02f01 g43337 ( .a(n2906), .b(n911), .o(n47129) );
na02f01 g43338 ( .a(n47129), .b(n47128), .o(n5721) );
na02f01 g43339 ( .a(n32732), .b(sin_out_28), .o(n47131) );
no02f01 g43340 ( .a(n44803), .b(n44796), .o(n47132) );
in01f01 g43341 ( .a(n47132), .o(n47133) );
no03f01 g43342 ( .a(n47133), .b(n44802), .c(n44799), .o(n47134) );
ao12f01 g43343 ( .a(n47132), .b(n44820), .c(n44819), .o(n47135) );
oa12f01 g43344 ( .a(n32734), .b(n47135), .c(n47134), .o(n47136) );
na02f01 g43345 ( .a(n47136), .b(n47131), .o(n5726) );
na02f01 g43346 ( .a(n3050), .b(n4116), .o(n47138) );
na02f01 g43347 ( .a(n44307), .b(n2589), .o(n47139) );
na02f01 g43348 ( .a(n47139), .b(n47138), .o(n5740) );
na02f01 g43349 ( .a(n45952), .b(n45949), .o(n5745) );
na03f01 g43350 ( .a(n46491), .b(n9590), .c(n9589), .o(n47142) );
oa12f01 g43351 ( .a(n4992), .b(n9646), .c(n9645), .o(n47143) );
na02f01 g43352 ( .a(n47143), .b(n47142), .o(n5750) );
no02f01 g43353 ( .a(n6971), .b(n46147), .o(n47145) );
no03f01 g43354 ( .a(n45830), .b(n6985), .c(n47145), .o(n47146) );
no02f01 g43355 ( .a(n6981), .b(n6934), .o(n47147) );
no02f01 g43356 ( .a(n47147), .b(n6983), .o(n47148) );
na02f01 g43357 ( .a(n47148), .b(n47146), .o(n47149) );
in01f01 g43358 ( .a(n47146), .o(n47150) );
in01f01 g43359 ( .a(n47148), .o(n47151) );
na02f01 g43360 ( .a(n47151), .b(n47150), .o(n47152) );
na02f01 g43361 ( .a(n47152), .b(n47149), .o(n5755) );
na02f01 g43362 ( .a(n32732), .b(sin_out_18), .o(n47154) );
na02f01 g43363 ( .a(n45068), .b(n45072), .o(n47155) );
no02f01 g43364 ( .a(n45070), .b(n41314), .o(n47156) );
in01f01 g43365 ( .a(n47156), .o(n47157) );
no02f01 g43366 ( .a(n47157), .b(n47155), .o(n47158) );
ao12f01 g43367 ( .a(n47156), .b(n45068), .c(n45072), .o(n47159) );
oa12f01 g43368 ( .a(n32734), .b(n47159), .c(n47158), .o(n47160) );
na02f01 g43369 ( .a(n47160), .b(n47154), .o(n5765) );
oa22f01 g43370 ( .a(n21203), .b(n41939), .c(n21190), .d(n21119), .o(n47162) );
na03f01 g43371 ( .a(n41940), .b(n21199), .c(n41938), .o(n47163) );
na02f01 g43372 ( .a(n47163), .b(n47162), .o(n5769) );
na03f01 g43373 ( .a(n36637), .b(n36636), .c(n25415), .o(n47165) );
oa12f01 g43374 ( .a(n25460), .b(n25461), .c(n36634), .o(n47166) );
na02f01 g43375 ( .a(n47166), .b(n47165), .o(n5779) );
na03f01 g43376 ( .a(n45976), .b(n45974), .c(n2589), .o(n47168) );
na02f01 g43377 ( .a(n4468), .b(n4116), .o(n47169) );
na02f01 g43378 ( .a(n47169), .b(n47168), .o(n5784) );
na02f01 g43379 ( .a(n21619), .b(n21612), .o(n5789) );
no02f01 g43380 ( .a(n42147), .b(n35412), .o(n47172) );
na02f01 g43381 ( .a(n47172), .b(n42144), .o(n47173) );
in01f01 g43382 ( .a(n47172), .o(n47174) );
na02f01 g43383 ( .a(n47174), .b(n42145), .o(n47175) );
na02f01 g43384 ( .a(n47175), .b(n47173), .o(n5794) );
in01f01 g43385 ( .a(n39148), .o(n47177) );
na02f01 g43386 ( .a(n47177), .b(n39146), .o(n47178) );
no03f01 g43387 ( .a(n44734), .b(n39157), .c(n44338), .o(n47179) );
oa12f01 g43388 ( .a(n47179), .b(n47178), .c(n39172), .o(n47180) );
in01f01 g43389 ( .a(n47180), .o(n47181) );
no02f01 g43390 ( .a(n39135), .b(n32344), .o(n47182) );
no02f01 g43391 ( .a(n47182), .b(n39149), .o(n47183) );
na02f01 g43392 ( .a(n47183), .b(n47181), .o(n47184) );
in01f01 g43393 ( .a(n47183), .o(n47185) );
na02f01 g43394 ( .a(n47185), .b(n47180), .o(n47186) );
na03f01 g43395 ( .a(n47186), .b(n47184), .c(n3633), .o(n47187) );
na02f01 g43396 ( .a(n47186), .b(n47184), .o(n6106) );
na02f01 g43397 ( .a(n6106), .b(n6203), .o(n47189) );
na02f01 g43398 ( .a(n47189), .b(n47187), .o(n5804) );
no02f01 g43399 ( .a(n29408), .b(n29327), .o(n47191) );
oa12f01 g43400 ( .a(n47191), .b(n29411), .c(n29292), .o(n47192) );
in01f01 g43401 ( .a(n47191), .o(n47193) );
na03f01 g43402 ( .a(n29709), .b(n47193), .c(n29673), .o(n47194) );
na02f01 g43403 ( .a(n47194), .b(n47192), .o(n5809) );
no02f01 g43404 ( .a(n9315), .b(n9225), .o(n47196) );
no02f01 g43405 ( .a(n47196), .b(n9317), .o(n47197) );
in01f01 g43406 ( .a(n47197), .o(n47198) );
oa12f01 g43407 ( .a(n47198), .b(n43705), .c(n9626), .o(n47199) );
in01f01 g43408 ( .a(n43705), .o(n47200) );
na03f01 g43409 ( .a(n47197), .b(n47200), .c(n9417), .o(n47201) );
na02f01 g43410 ( .a(n47201), .b(n47199), .o(n5814) );
no02f01 g43411 ( .a(n22631), .b(n22501), .o(n47203) );
in01f01 g43412 ( .a(n47203), .o(n47204) );
na02f01 g43413 ( .a(n47204), .b(n22630), .o(n47205) );
na02f01 g43414 ( .a(n47203), .b(n22629), .o(n47206) );
na02f01 g43415 ( .a(n47206), .b(n47205), .o(n5819) );
na03f01 g43416 ( .a(n39792), .b(n39789), .c(n3633), .o(n47208) );
no03f01 g43417 ( .a(n39791), .b(n39790), .c(n39162), .o(n47209) );
ao12f01 g43418 ( .a(n39786), .b(n39788), .c(n39782), .o(n47210) );
oa12f01 g43419 ( .a(n6203), .b(n47210), .c(n47209), .o(n47211) );
na02f01 g43420 ( .a(n47211), .b(n47208), .o(n5824) );
na03f01 g43421 ( .a(n36893), .b(n36890), .c(n3633), .o(n47213) );
no03f01 g43422 ( .a(n36892), .b(n36840), .c(n36831), .o(n47214) );
ao12f01 g43423 ( .a(n36832), .b(n36889), .c(n36841), .o(n47215) );
oa12f01 g43424 ( .a(n6203), .b(n47215), .c(n47214), .o(n47216) );
na02f01 g43425 ( .a(n47216), .b(n47213), .o(n5829) );
na02f01 g43426 ( .a(n43370), .b(n5799), .o(n47218) );
na02f01 g43427 ( .a(n2402), .b(n911), .o(n47219) );
na02f01 g43428 ( .a(n47219), .b(n47218), .o(n5839) );
no02f01 g43429 ( .a(n42771), .b(n35336), .o(n47221) );
in01f01 g43430 ( .a(n47221), .o(n47222) );
na02f01 g43431 ( .a(n47222), .b(n35327), .o(n47223) );
na03f01 g43432 ( .a(n47221), .b(n35326), .c(n35324), .o(n47224) );
na02f01 g43433 ( .a(n47224), .b(n47223), .o(n5854) );
no02f01 g43434 ( .a(n27235), .b(n26904), .o(n47226) );
na02f01 g43435 ( .a(n47226), .b(n27234), .o(n47227) );
in01f01 g43436 ( .a(n47226), .o(n47228) );
na02f01 g43437 ( .a(n47228), .b(n27043), .o(n47229) );
na02f01 g43438 ( .a(n47229), .b(n47227), .o(n5859) );
na02f01 g43439 ( .a(n46675), .b(n46672), .o(n5864) );
no02f01 g43440 ( .a(n11688), .b(n11686), .o(n47232) );
no02f01 g43441 ( .a(n11687), .b(n11579), .o(n47233) );
na02f01 g43442 ( .a(n47233), .b(n47232), .o(n47234) );
in01f01 g43443 ( .a(n47233), .o(n47235) );
oa12f01 g43444 ( .a(n47235), .b(n11688), .c(n11686), .o(n47236) );
na02f01 g43445 ( .a(n47236), .b(n47234), .o(n5869) );
na02f01 g43446 ( .a(n32732), .b(cos_out_8), .o(n47238) );
no02f01 g43447 ( .a(n36277), .b(n35944), .o(n47239) );
no02f01 g43448 ( .a(n47239), .b(n36279), .o(n47240) );
in01f01 g43449 ( .a(n47240), .o(n47241) );
no02f01 g43450 ( .a(n47241), .b(n39661), .o(n47242) );
no02f01 g43451 ( .a(n47240), .b(n36269), .o(n47243) );
oa12f01 g43452 ( .a(n32734), .b(n47243), .c(n47242), .o(n47244) );
na02f01 g43453 ( .a(n47244), .b(n47238), .o(n5874) );
no02f01 g43454 ( .a(n42259), .b(n45761), .o(n47246) );
in01f01 g43455 ( .a(n5938_1), .o(n47247) );
no02f01 g43456 ( .a(n5937), .b(n5873), .o(n47248) );
no02f01 g43457 ( .a(n47248), .b(n47247), .o(n47249) );
na02f01 g43458 ( .a(n47249), .b(n47246), .o(n47250) );
in01f01 g43459 ( .a(n47249), .o(n47251) );
oa12f01 g43460 ( .a(n47251), .b(n42259), .c(n45761), .o(n47252) );
na02f01 g43461 ( .a(n47252), .b(n47250), .o(n5878) );
na02f01 g43462 ( .a(n46692), .b(n46687), .o(n5883) );
na02f01 g43463 ( .a(n44497), .b(n44494), .o(n5893) );
na03f01 g43464 ( .a(n38401), .b(n39106), .c(n38391), .o(n47256) );
oa12f01 g43465 ( .a(n39103), .b(n39107), .c(n38400), .o(n47257) );
na02f01 g43466 ( .a(n47257), .b(n47256), .o(n5898) );
no02f01 g43467 ( .a(n9405), .b(n9329), .o(n47259) );
na03f01 g43468 ( .a(n47259), .b(n9403), .c(n9337), .o(n47260) );
in01f01 g43469 ( .a(n47259), .o(n47261) );
oa12f01 g43470 ( .a(n47261), .b(n9624), .c(n9336), .o(n47262) );
na02f01 g43471 ( .a(n47262), .b(n47260), .o(n5918) );
no02f01 g43472 ( .a(n35505), .b(n4176), .o(n47264) );
in01f01 g43473 ( .a(n47264), .o(n47265) );
in01f01 g43474 ( .a(n35507), .o(n47266) );
na02f01 g43475 ( .a(n35536), .b(n45099), .o(n47267) );
na02f01 g43476 ( .a(n47267), .b(n47266), .o(n47268) );
no02f01 g43477 ( .a(n35537), .b(n4176), .o(n47269) );
no02f01 g43478 ( .a(n47269), .b(n35499), .o(n47270) );
na03f01 g43479 ( .a(n47270), .b(n47268), .c(n47265), .o(n47271) );
na02f01 g43480 ( .a(n47268), .b(n47265), .o(n47272) );
in01f01 g43481 ( .a(n47270), .o(n47273) );
na02f01 g43482 ( .a(n47273), .b(n47272), .o(n47274) );
na02f01 g43483 ( .a(n47274), .b(n47271), .o(n5923) );
ao12f01 g43484 ( .a(n43896), .b(n43897), .c(n43901), .o(n47276) );
in01f01 g43485 ( .a(n9497), .o(n47277) );
no02f01 g43486 ( .a(n47277), .b(n9224), .o(n47278) );
no02f01 g43487 ( .a(n9497), .b(n9225), .o(n47279) );
no02f01 g43488 ( .a(n47279), .b(n47278), .o(n47280) );
na02f01 g43489 ( .a(n47280), .b(n47276), .o(n47281) );
in01f01 g43490 ( .a(n47276), .o(n47282) );
in01f01 g43491 ( .a(n47280), .o(n47283) );
na02f01 g43492 ( .a(n47283), .b(n47282), .o(n47284) );
na02f01 g43493 ( .a(n47284), .b(n47281), .o(n5928) );
no02f01 g43494 ( .a(n27674), .b(n27673), .o(n47286) );
in01f01 g43495 ( .a(n27621), .o(n47287) );
na02f01 g43496 ( .a(n47287), .b(n47286), .o(n47288) );
no02f01 g43497 ( .a(n27619), .b(n27367), .o(n47289) );
no02f01 g43498 ( .a(n47289), .b(n27636), .o(n47290) );
no02f01 g43499 ( .a(n27367), .b(n15984), .o(n47291) );
no02f01 g43500 ( .a(n47291), .b(n27622), .o(n47292) );
na03f01 g43501 ( .a(n47292), .b(n47290), .c(n47288), .o(n47293) );
na02f01 g43502 ( .a(n47290), .b(n47288), .o(n47294) );
in01f01 g43503 ( .a(n47292), .o(n47295) );
na02f01 g43504 ( .a(n47295), .b(n47294), .o(n47296) );
na02f01 g43505 ( .a(n47296), .b(n47293), .o(n5933) );
ao12f01 g43506 ( .a(n46981), .b(n46970), .c(n42012), .o(n47298) );
oa22f01 g43507 ( .a(n47298), .b(n10735), .c(n46983), .d(n46987), .o(n5938) );
na02f01 g43508 ( .a(n683), .b(n4116), .o(n47300) );
na02f01 g43509 ( .a(n38866), .b(n2589), .o(n47301) );
na02f01 g43510 ( .a(n47301), .b(n47300), .o(n5943) );
no02f01 g43511 ( .a(n44011), .b(n38113), .o(n47303) );
na02f01 g43512 ( .a(n47303), .b(n41664), .o(n47304) );
in01f01 g43513 ( .a(n47303), .o(n47305) );
na02f01 g43514 ( .a(n47305), .b(n44014), .o(n47306) );
na02f01 g43515 ( .a(n47306), .b(n47304), .o(n5948) );
na03f01 g43516 ( .a(n27224), .b(n27026), .c(n26994), .o(n47308) );
oa12f01 g43517 ( .a(n27223), .b(n27027), .c(n27209), .o(n47309) );
na02f01 g43518 ( .a(n47309), .b(n47308), .o(n5953) );
na03f01 g43519 ( .a(n46661), .b(n46660), .c(n1821), .o(n47311) );
na02f01 g43520 ( .a(n5175), .b(n8066), .o(n47312) );
na02f01 g43521 ( .a(n47312), .b(n47311), .o(n5958) );
na02f01 g43522 ( .a(n46856), .b(n5799), .o(n47314) );
na02f01 g43523 ( .a(n5400), .b(n911), .o(n47315) );
na02f01 g43524 ( .a(n47315), .b(n47314), .o(n5963) );
na03f01 g43525 ( .a(n32714), .b(n32609), .c(n32698), .o(n47317) );
oa12f01 g43526 ( .a(n32665), .b(n32699), .c(n32608), .o(n47318) );
na02f01 g43527 ( .a(n47318), .b(n47317), .o(n5968) );
na03f01 g43528 ( .a(n46634), .b(n46632), .c(n3633), .o(n47320) );
na02f01 g43529 ( .a(n5140), .b(n6203), .o(n47321) );
na02f01 g43530 ( .a(n47321), .b(n47320), .o(n5983) );
na02f01 g43531 ( .a(n32654), .b(n27063), .o(n47323) );
na02f01 g43532 ( .a(n47323), .b(n46718), .o(n5993) );
na03f01 g43533 ( .a(n46233), .b(n46231), .c(n3633), .o(n47325) );
no03f01 g43534 ( .a(n46232), .b(n46227), .c(n41832), .o(n47326) );
ao12f01 g43535 ( .a(n46228), .b(n46230), .c(n46223), .o(n47327) );
oa12f01 g43536 ( .a(n6203), .b(n47327), .c(n47326), .o(n47328) );
na02f01 g43537 ( .a(n47328), .b(n47325), .o(n5998) );
na02f01 g43538 ( .a(n32732), .b(cos_out_16), .o(n47330) );
no02f01 g43539 ( .a(n36376), .b(n36231), .o(n47331) );
in01f01 g43540 ( .a(n47331), .o(n47332) );
no03f01 g43541 ( .a(n47332), .b(n36373), .c(n36365), .o(n47333) );
no02f01 g43542 ( .a(n47331), .b(n36374), .o(n47334) );
oa12f01 g43543 ( .a(n32734), .b(n47334), .c(n47333), .o(n47335) );
na02f01 g43544 ( .a(n47335), .b(n47330), .o(n6003) );
na03f01 g43545 ( .a(n39175), .b(n39165), .c(n3633), .o(n47337) );
na02f01 g43546 ( .a(n756), .b(n6203), .o(n47338) );
na02f01 g43547 ( .a(n47338), .b(n47337), .o(n6007) );
no02f01 g43548 ( .a(n47264), .b(n35507), .o(n47340) );
na03f01 g43549 ( .a(n47340), .b(n35536), .c(n45099), .o(n47341) );
in01f01 g43550 ( .a(n47340), .o(n47342) );
na02f01 g43551 ( .a(n47342), .b(n47267), .o(n47343) );
na02f01 g43552 ( .a(n47343), .b(n47341), .o(n6012) );
in01f01 g43553 ( .a(n44599), .o(n47345) );
no02f01 g43554 ( .a(n44601), .b(n37239), .o(n47346) );
na03f01 g43555 ( .a(n47346), .b(n37255), .c(n47345), .o(n47347) );
in01f01 g43556 ( .a(n47346), .o(n47348) );
oa12f01 g43557 ( .a(n47348), .b(n37256), .c(n44599), .o(n47349) );
na02f01 g43558 ( .a(n47349), .b(n47347), .o(n6022) );
na03f01 g43559 ( .a(n32719), .b(n32675), .c(n32666), .o(n47351) );
oa12f01 g43560 ( .a(n32715), .b(n32676), .c(n32718), .o(n47352) );
na02f01 g43561 ( .a(n47352), .b(n47351), .o(n6027) );
na03f01 g43562 ( .a(n46846), .b(n46845), .c(n6037), .o(n47354) );
na02f01 g43563 ( .a(n5390), .b(n5873), .o(n47355) );
na02f01 g43564 ( .a(n47355), .b(n47354), .o(n6032) );
in01f01 g43565 ( .a(n40158), .o(n47357) );
no02f01 g43566 ( .a(n40171), .b(n40168), .o(n47358) );
in01f01 g43567 ( .a(n47358), .o(n47359) );
na02f01 g43568 ( .a(n47359), .b(n47357), .o(n47360) );
na02f01 g43569 ( .a(n47358), .b(n40158), .o(n47361) );
na02f01 g43570 ( .a(n47361), .b(n47360), .o(n6042) );
in01f01 g43571 ( .a(n9745), .o(n47363) );
ao12f01 g43572 ( .a(n36528), .b(n47363), .c(n36539), .o(n47364) );
no02f01 g43573 ( .a(n9736), .b(n5001), .o(n47365) );
no02f01 g43574 ( .a(n47365), .b(n9738), .o(n47366) );
na02f01 g43575 ( .a(n47366), .b(n47364), .o(n47367) );
in01f01 g43576 ( .a(n47364), .o(n47368) );
in01f01 g43577 ( .a(n47366), .o(n47369) );
na02f01 g43578 ( .a(n47369), .b(n47368), .o(n47370) );
na02f01 g43579 ( .a(n47370), .b(n47367), .o(n6056) );
no02f01 g43580 ( .a(n44591), .b(n44590), .o(n47372) );
no02f01 g43581 ( .a(n22570), .b(n22544), .o(n47373) );
in01f01 g43582 ( .a(n47373), .o(n47374) );
oa12f01 g43583 ( .a(n47374), .b(n47372), .c(n22551), .o(n47375) );
na02f01 g43584 ( .a(n47373), .b(n22568), .o(n47376) );
na02f01 g43585 ( .a(n47376), .b(n47375), .o(n6066) );
no02f01 g43586 ( .a(n43869), .b(n43862), .o(n47378) );
na02f01 g43587 ( .a(n47378), .b(n43879), .o(n47379) );
in01f01 g43588 ( .a(n47378), .o(n47380) );
na02f01 g43589 ( .a(n47380), .b(n43873), .o(n47381) );
na03f01 g43590 ( .a(n47381), .b(n47379), .c(n1821), .o(n47382) );
na02f01 g43591 ( .a(n47381), .b(n47379), .o(n6125) );
na02f01 g43592 ( .a(n6125), .b(n8066), .o(n47384) );
na02f01 g43593 ( .a(n47384), .b(n47382), .o(n6071) );
in01f01 g43594 ( .a(n29644), .o(n47386) );
na02f01 g43595 ( .a(n29599), .b(n29430), .o(n47387) );
na02f01 g43596 ( .a(n47387), .b(n42136), .o(n47388) );
in01f01 g43597 ( .a(n47388), .o(n47389) );
na03f01 g43598 ( .a(n47389), .b(n47386), .c(n29578), .o(n47390) );
oa12f01 g43599 ( .a(n47388), .b(n29644), .c(n29721), .o(n47391) );
na02f01 g43600 ( .a(n47391), .b(n47390), .o(n6076) );
na03f01 g43601 ( .a(n43487), .b(n43486), .c(n6037), .o(n47393) );
na02f01 g43602 ( .a(n2481), .b(n5873), .o(n47394) );
na02f01 g43603 ( .a(n47394), .b(n47393), .o(n6086) );
na03f01 g43604 ( .a(n42608), .b(n42606), .c(n5799), .o(n47396) );
in01f01 g43605 ( .a(n42606), .o(n47397) );
oa12f01 g43606 ( .a(n911), .b(n42607), .c(n47397), .o(n47398) );
na02f01 g43607 ( .a(n47398), .b(n47396), .o(n6091) );
in01f01 g43608 ( .a(n45049), .o(n47400) );
ao12f01 g43609 ( .a(n37102), .b(n45048), .c(n47400), .o(n47401) );
in01f01 g43610 ( .a(n47401), .o(n47402) );
no02f01 g43611 ( .a(n37091), .b(n36963), .o(n47403) );
no02f01 g43612 ( .a(n47403), .b(n37093), .o(n47404) );
na02f01 g43613 ( .a(n47404), .b(n47402), .o(n47405) );
in01f01 g43614 ( .a(n47404), .o(n47406) );
na02f01 g43615 ( .a(n47406), .b(n47401), .o(n47407) );
na02f01 g43616 ( .a(n47407), .b(n47405), .o(n6096) );
oa12f01 g43617 ( .a(n8581), .b(n45202), .c(n45205), .o(n47409) );
no02f01 g43618 ( .a(n8570), .b(n5973), .o(n47410) );
no02f01 g43619 ( .a(n47410), .b(n8580), .o(n47411) );
na02f01 g43620 ( .a(n47411), .b(n47409), .o(n47412) );
in01f01 g43621 ( .a(n47409), .o(n47413) );
in01f01 g43622 ( .a(n47411), .o(n47414) );
na02f01 g43623 ( .a(n47414), .b(n47413), .o(n47415) );
na02f01 g43624 ( .a(n47415), .b(n47412), .o(n6101) );
na04f01 g43625 ( .a(n30103), .b(n30101), .c(n25893), .d(n25794), .o(n47417) );
oa22f01 g43626 ( .a(n25911), .b(n25907), .c(n30100), .d(n25793), .o(n47418) );
na02f01 g43627 ( .a(n47418), .b(n47417), .o(n6111) );
na02f01 g43628 ( .a(n43881), .b(n43875), .o(n6116) );
na02f01 g43629 ( .a(n32732), .b(sin_out_26), .o(n47421) );
no02f01 g43630 ( .a(n44558), .b(n46337), .o(n47422) );
in01f01 g43631 ( .a(n47422), .o(n47423) );
no02f01 g43632 ( .a(n44560), .b(n44553), .o(n47424) );
in01f01 g43633 ( .a(n47424), .o(n47425) );
no03f01 g43634 ( .a(n47425), .b(n47423), .c(n44557), .o(n47426) );
ao12f01 g43635 ( .a(n47424), .b(n47422), .c(n44566), .o(n47427) );
oa12f01 g43636 ( .a(n32734), .b(n47427), .c(n47426), .o(n47428) );
na02f01 g43637 ( .a(n47428), .b(n47421), .o(n6121) );
ao12f01 g43638 ( .a(n39466), .b(n40032), .c(n39452), .o(n47430) );
in01f01 g43639 ( .a(n47430), .o(n47431) );
no02f01 g43640 ( .a(n39469), .b(n39372), .o(n47432) );
na02f01 g43641 ( .a(n47432), .b(n47431), .o(n47433) );
in01f01 g43642 ( .a(n47432), .o(n47434) );
na02f01 g43643 ( .a(n47434), .b(n47430), .o(n47435) );
na02f01 g43644 ( .a(n47435), .b(n47433), .o(n6130) );
na03f01 g43645 ( .a(n27357), .b(n27657), .c(n27649), .o(n47437) );
oa12f01 g43646 ( .a(n27356), .b(n27658), .c(n27334), .o(n47438) );
na02f01 g43647 ( .a(n47438), .b(n47437), .o(n6135) );
na02f01 g43648 ( .a(n3762), .b(n8066), .o(n47440) );
na03f01 g43649 ( .a(n45248), .b(n45245), .c(n1821), .o(n47441) );
na02f01 g43650 ( .a(n47441), .b(n47440), .o(n6140) );
na02f01 g43651 ( .a(n44136), .b(n5799), .o(n47443) );
na02f01 g43652 ( .a(n2941), .b(n911), .o(n47444) );
na02f01 g43653 ( .a(n47444), .b(n47443), .o(n6145) );
no02f01 g43654 ( .a(n40301), .b(n38143), .o(n47446) );
no02f01 g43655 ( .a(n47446), .b(n40307), .o(n47447) );
no02f01 g43656 ( .a(n46993), .b(n40293), .o(n47448) );
na02f01 g43657 ( .a(n47448), .b(n47447), .o(n47449) );
in01f01 g43658 ( .a(n47448), .o(n47450) );
oa12f01 g43659 ( .a(n47450), .b(n47446), .c(n40307), .o(n47451) );
na02f01 g43660 ( .a(n47451), .b(n47449), .o(n6154) );
na02f01 g43661 ( .a(n32732), .b(cos_out_9), .o(n47453) );
in01f01 g43662 ( .a(n36279), .o(n47454) );
ao12f01 g43663 ( .a(n47239), .b(n47454), .c(n39661), .o(n47455) );
in01f01 g43664 ( .a(n47455), .o(n47456) );
no02f01 g43665 ( .a(n36288), .b(n35944), .o(n47457) );
no02f01 g43666 ( .a(n47457), .b(n36290), .o(n47458) );
in01f01 g43667 ( .a(n47458), .o(n47459) );
no02f01 g43668 ( .a(n47459), .b(n47456), .o(n47460) );
no02f01 g43669 ( .a(n47458), .b(n47455), .o(n47461) );
oa12f01 g43670 ( .a(n32734), .b(n47461), .c(n47460), .o(n47462) );
na02f01 g43671 ( .a(n47462), .b(n47453), .o(n6159) );
na03f01 g43672 ( .a(n27035), .b(n27034), .c(n26946), .o(n47464) );
oa12f01 g43673 ( .a(n27231), .b(n27036), .c(n26945), .o(n47465) );
na02f01 g43674 ( .a(n47465), .b(n47464), .o(n6163) );
na02f01 g43675 ( .a(n32732), .b(sin_out_31), .o(n47467) );
in01f01 g43676 ( .a(n44801), .o(n47468) );
no02f01 g43677 ( .a(n35911), .b(n34267), .o(n47469) );
no02f01 g43678 ( .a(n35931), .b(n34307), .o(n47470) );
no02f01 g43679 ( .a(n47470), .b(n47469), .o(n47471) );
in01f01 g43680 ( .a(n47471), .o(n47472) );
no03f01 g43681 ( .a(n46319), .b(n46309), .c(n44798), .o(n47473) );
in01f01 g43682 ( .a(n47473), .o(n47474) );
ao12f01 g43683 ( .a(n47474), .b(n41371), .c(n41353), .o(n47475) );
ao12f01 g43684 ( .a(n34307), .b(n46316), .c(n46310), .o(n47476) );
no04f01 g43685 ( .a(n47476), .b(n47475), .c(n47472), .d(n47468), .o(n47477) );
oa12f01 g43686 ( .a(n47473), .b(n46337), .c(n46336), .o(n47478) );
no02f01 g43687 ( .a(n47476), .b(n47468), .o(n47479) );
ao12f01 g43688 ( .a(n47471), .b(n47479), .c(n47478), .o(n47480) );
oa12f01 g43689 ( .a(n32734), .b(n47480), .c(n47477), .o(n47481) );
na02f01 g43690 ( .a(n47481), .b(n47467), .o(n6168) );
na02f01 g43691 ( .a(n22489), .b(n22488), .o(n6172) );
in01f01 g43692 ( .a(n40171), .o(n47484) );
ao12f01 g43693 ( .a(n40168), .b(n47484), .c(n40158), .o(n47485) );
in01f01 g43694 ( .a(n47485), .o(n47486) );
no02f01 g43695 ( .a(n40169), .b(n40156), .o(n47487) );
na02f01 g43696 ( .a(n47487), .b(n47486), .o(n47488) );
oa12f01 g43697 ( .a(n47485), .b(n40169), .c(n40156), .o(n47489) );
na02f01 g43698 ( .a(n47489), .b(n47488), .o(n6177) );
in01f01 g43699 ( .a(n45796), .o(n47491) );
na03f01 g43700 ( .a(n10985), .b(n10981), .c(n43057), .o(n47492) );
no02f01 g43701 ( .a(n10756), .b(n3521), .o(n47493) );
no02f01 g43702 ( .a(n47493), .b(n10984), .o(n47494) );
na04f01 g43703 ( .a(n47494), .b(n47492), .c(n45793), .d(n47491), .o(n47495) );
na03f01 g43704 ( .a(n47492), .b(n45793), .c(n47491), .o(n47496) );
in01f01 g43705 ( .a(n47494), .o(n47497) );
na02f01 g43706 ( .a(n47497), .b(n47496), .o(n47498) );
na02f01 g43707 ( .a(n47498), .b(n47495), .o(n6182) );
no02f01 g43708 ( .a(n27636), .b(n47286), .o(n47500) );
no02f01 g43709 ( .a(n47289), .b(n27621), .o(n47501) );
na02f01 g43710 ( .a(n47501), .b(n47500), .o(n47502) );
in01f01 g43711 ( .a(n47501), .o(n47503) );
oa12f01 g43712 ( .a(n47503), .b(n27636), .c(n47286), .o(n47504) );
na02f01 g43713 ( .a(n47504), .b(n47502), .o(n6187) );
na03f01 g43714 ( .a(n40997), .b(n40994), .c(n1821), .o(n47506) );
na02f01 g43715 ( .a(n1210), .b(n8066), .o(n47507) );
na02f01 g43716 ( .a(n47507), .b(n47506), .o(n6192) );
na03f01 g43717 ( .a(n42116), .b(n42114), .c(n6037), .o(n47509) );
no03f01 g43718 ( .a(n42115), .b(n42110), .c(n25181), .o(n47510) );
ao12f01 g43719 ( .a(n42111), .b(n42113), .c(n25180), .o(n47511) );
oa12f01 g43720 ( .a(n5873), .b(n47511), .c(n47510), .o(n47512) );
na02f01 g43721 ( .a(n47512), .b(n47509), .o(n6197) );
no02f01 g43722 ( .a(n42644), .b(n42643), .o(n47514) );
oa12f01 g43723 ( .a(n47514), .b(n8584), .c(n8578), .o(n47515) );
in01f01 g43724 ( .a(n47514), .o(n47516) );
na02f01 g43725 ( .a(n47516), .b(n42642), .o(n47517) );
na02f01 g43726 ( .a(n47517), .b(n47515), .o(n6202) );
no02f01 g43727 ( .a(n44347), .b(n44028), .o(n47519) );
no02f01 g43728 ( .a(n10815), .b(n3521), .o(n47520) );
no02f01 g43729 ( .a(n47520), .b(n10861), .o(n47521) );
na02f01 g43730 ( .a(n47521), .b(n47519), .o(n47522) );
in01f01 g43731 ( .a(n47521), .o(n47523) );
oa12f01 g43732 ( .a(n47523), .b(n44347), .c(n44028), .o(n47524) );
na02f01 g43733 ( .a(n47524), .b(n47522), .o(n6207) );
in01f01 g43734 ( .a(n40440), .o(n47526) );
ao12f01 g43735 ( .a(n40439), .b(n47526), .c(n21374), .o(n47527) );
no02f01 g43736 ( .a(n16479), .b(n16329), .o(n47528) );
no02f01 g43737 ( .a(n16480), .b(n16155), .o(n47529) );
no02f01 g43738 ( .a(n47529), .b(n47528), .o(n47530) );
na02f01 g43739 ( .a(n47530), .b(n47527), .o(n47531) );
in01f01 g43740 ( .a(n47527), .o(n47532) );
in01f01 g43741 ( .a(n47530), .o(n47533) );
na02f01 g43742 ( .a(n47533), .b(n47532), .o(n47534) );
na02f01 g43743 ( .a(n47534), .b(n47531), .o(n6212) );
na02f01 g43744 ( .a(n43993), .b(n43988), .o(n6217) );
no02f01 g43745 ( .a(n44759), .b(n44758), .o(n47537) );
na03f01 g43746 ( .a(n47537), .b(n29720), .c(n29719), .o(n47538) );
in01f01 g43747 ( .a(n47537), .o(n47539) );
na02f01 g43748 ( .a(n47539), .b(n44757), .o(n47540) );
na02f01 g43749 ( .a(n47540), .b(n47538), .o(n6227) );
na03f01 g43750 ( .a(n38036), .b(n37966), .c(n37965), .o(n47542) );
oa12f01 g43751 ( .a(n38035), .b(n37970), .c(n37964), .o(n47543) );
na02f01 g43752 ( .a(n47543), .b(n47542), .o(n6236) );
na03f01 g43753 ( .a(n29691), .b(n29361), .c(n29684), .o(n47545) );
oa12f01 g43754 ( .a(n29383), .b(n29685), .c(n29360), .o(n47546) );
na02f01 g43755 ( .a(n47546), .b(n47545), .o(n6241) );
na02f01 g43756 ( .a(n9642), .b(n9641), .o(n47548) );
in01f01 g43757 ( .a(n42532), .o(n47549) );
no02f01 g43758 ( .a(n9555), .b(n9225), .o(n47550) );
no02f01 g43759 ( .a(n47550), .b(n9557), .o(n47551) );
na03f01 g43760 ( .a(n47551), .b(n47549), .c(n47548), .o(n47552) );
na02f01 g43761 ( .a(n47549), .b(n47548), .o(n47553) );
in01f01 g43762 ( .a(n47551), .o(n47554) );
na02f01 g43763 ( .a(n47554), .b(n47553), .o(n47555) );
na02f01 g43764 ( .a(n47555), .b(n47552), .o(n6246) );
na03f01 g43765 ( .a(n41659), .b(n41655), .c(n3633), .o(n47557) );
na02f01 g43766 ( .a(n1396), .b(n6203), .o(n47558) );
na02f01 g43767 ( .a(n47558), .b(n47557), .o(n6251) );
no02f01 g43768 ( .a(n14158), .b(n14088), .o(n47560) );
na02f01 g43769 ( .a(n47560), .b(n14157), .o(n47561) );
in01f01 g43770 ( .a(n14157), .o(n47562) );
in01f01 g43771 ( .a(n47560), .o(n47563) );
na02f01 g43772 ( .a(n47563), .b(n47562), .o(n47564) );
na02f01 g43773 ( .a(n47564), .b(n47561), .o(n6256) );
oa12f01 g43774 ( .a(n27353), .b(n27654), .c(n27653), .o(n47566) );
na03f01 g43775 ( .a(n27352), .b(n27347), .c(n27346), .o(n47567) );
na02f01 g43776 ( .a(n47567), .b(n47566), .o(n6265) );
bf01f01 g43777 ( .a(cordic_combinational_sub_ln23_0_unr20_z_0_), .o(n203) );
bf01f01 g43778 ( .a(n_27923), .o(n218) );
bf01f01 g43779 ( .a(n_186), .o(n765) );
bf01f01 g43780 ( .a(cordic_combinational_sub_ln23_0_unr12_z_0_), .o(n818) );
no02f01 g43781 ( .a(n9646), .b(n9645), .o(n1540) );
no02f01 g43782 ( .a(n9646), .b(n9645), .o(n1664) );
bf01f01 g43783 ( .a(cordic_combinational_sub_ln23_0_unr16_z_0_), .o(n1763) );
na02f01 g43784 ( .a(n40561), .b(n40559), .o(n2072) );
no02f01 g43785 ( .a(n9646), .b(n9645), .o(n3994) );
bf01f01 g43786 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_0_), .o(n4443) );
bf01f01 g43787 ( .a(rst), .o(n4843) );
bf01f01 g43788 ( .a(beta_31), .o(n5026) );
bf01f01 g43789 ( .a(delay_sub_ln23_0_unr27_stage10_stallmux_z), .o(n5070) );
bf01f01 g43790 ( .a(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .o(n6051) );
in01f01 g43791 ( .a(n3707), .o(n6149) );
no02f01 g43792 ( .a(n9646), .b(n9645), .o(n6231) );
bf01f01 g43793 ( .a(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .o(n6260) );
ms00f80 l0001 ( .d(n198), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_4_), .ck(clk) );
ms00f80 l0002 ( .d(n203), .o(n_186), .ck(clk) );
ms00f80 l0003 ( .d(n208), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_19_), .ck(clk) );
ms00f80 l0004 ( .d(n213), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_10_), .ck(clk) );
ms00f80 l0005 ( .d(n218), .o(n_44962), .ck(clk) );
ms00f80 l0006 ( .d(n223), .o(delay_add_ln22_unr23_stage9_stallmux_q_5_), .ck(clk) );
ms00f80 l0007 ( .d(n228), .o(delay_sub_ln23_unr17_stage6_stallmux_q_1_), .ck(clk) );
ms00f80 l0008 ( .d(n233), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_5_), .ck(clk) );
ms00f80 l0009 ( .d(n238), .o(delay_xor_ln21_unr3_stage2_stallmux_q_9_), .ck(clk) );
ms00f80 l0010 ( .d(n243), .o(delay_sub_ln23_unr21_stage7_stallmux_q_1_), .ck(clk) );
ms00f80 l0011 ( .d(n248), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_22_), .ck(clk) );
ms00f80 l0012 ( .d(n253), .o(delay_xor_ln21_unr6_stage3_stallmux_q_15_), .ck(clk) );
ms00f80 l0013 ( .d(n258), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_19_), .ck(clk) );
ms00f80 l0014 ( .d(n263), .o(delay_add_ln22_unr14_stage6_stallmux_q_3_), .ck(clk) );
ms00f80 l0015 ( .d(n268), .o(delay_add_ln22_unr23_stage9_stallmux_q_4_), .ck(clk) );
ms00f80 l0016 ( .d(n273), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_24_), .ck(clk) );
ms00f80 l0017 ( .d(n278), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_12_), .ck(clk) );
ms00f80 l0018 ( .d(n283), .o(delay_xor_ln22_unr28_stage10_stallmux_q_1_), .ck(clk) );
ms00f80 l0019 ( .d(n288), .o(delay_xor_ln22_unr6_stage3_stallmux_q_24_), .ck(clk) );
ms00f80 l0020 ( .d(n293), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_20_), .ck(clk) );
ms00f80 l0021 ( .d(n298), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_16_), .ck(clk) );
ms00f80 l0022 ( .d(n303), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_30_), .ck(clk) );
ms00f80 l0023 ( .d(n308), .o(delay_xor_ln21_unr6_stage3_stallmux_q_17_), .ck(clk) );
ms00f80 l0024 ( .d(n313), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_10_), .ck(clk) );
ms00f80 l0025 ( .d(n318), .o(delay_xor_ln22_unr6_stage3_stallmux_q_20_), .ck(clk) );
ms00f80 l0026 ( .d(n323), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_21_), .ck(clk) );
ms00f80 l0027 ( .d(n328), .o(n_44847), .ck(clk) );
ms00f80 l0028 ( .d(n333), .o(delay_add_ln22_unr5_stage3_stallmux_q_3_), .ck(clk) );
ms00f80 l0029 ( .d(n338), .o(delay_add_ln22_unr5_stage3_stallmux_q_0_), .ck(clk) );
ms00f80 l0030 ( .d(n343), .o(delay_xor_ln21_unr15_stage6_stallmux_q_15_), .ck(clk) );
ms00f80 l0031 ( .d(n348), .o(delay_add_ln22_unr27_stage10_stallmux_q_28_), .ck(clk) );
ms00f80 l0032 ( .d(n353), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_21_), .ck(clk) );
ms00f80 l0033 ( .d(n358), .o(delay_add_ln22_unr14_stage6_stallmux_q_4_), .ck(clk) );
ms00f80 l0034 ( .d(n363), .o(delay_add_ln22_unr27_stage10_stallmux_q_20_), .ck(clk) );
ms00f80 l0035 ( .d(n368), .o(delay_add_ln22_unr8_stage4_stallmux_q_5_), .ck(clk) );
ms00f80 l0036 ( .d(n373), .o(delay_add_ln22_unr14_stage6_stallmux_q_14_), .ck(clk) );
ms00f80 l0037 ( .d(n378), .o(delay_xor_ln22_unr3_stage2_stallmux_q_20_), .ck(clk) );
ms00f80 l0038 ( .d(n383), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_23_), .ck(clk) );
ms00f80 l0039 ( .d(n388), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_3_), .ck(clk) );
ms00f80 l0040 ( .d(n393), .o(delay_xor_ln21_unr12_stage5_stallmux_q_16_), .ck(clk) );
ms00f80 l0041 ( .d(n398), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_28_), .ck(clk) );
ms00f80 l0042 ( .d(n403), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_24_), .ck(clk) );
ms00f80 l0043 ( .d(n408), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_26_), .ck(clk) );
ms00f80 l0044 ( .d(n413), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_9_), .ck(clk) );
ms00f80 l0045 ( .d(n418), .o(sin_out_5), .ck(clk) );
ms00f80 l0046 ( .d(n422), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_27_), .ck(clk) );
ms00f80 l0047 ( .d(n427), .o(delay_xor_ln23_unr3_stage2_stallmux_q), .ck(clk) );
ms00f80 l0048 ( .d(n432), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_16_), .ck(clk) );
ms00f80 l0049 ( .d(n437), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_24_), .ck(clk) );
ms00f80 l0050 ( .d(n442), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_14_), .ck(clk) );
ms00f80 l0051 ( .d(n447), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_26_), .ck(clk) );
ms00f80 l0052 ( .d(n452), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_0_), .ck(clk) );
ms00f80 l0053 ( .d(n457), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_5_), .ck(clk) );
ms00f80 l0054 ( .d(n462), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_2_), .ck(clk) );
ms00f80 l0055 ( .d(n467), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_16_), .ck(clk) );
ms00f80 l0056 ( .d(n472), .o(cos_out_4), .ck(clk) );
ms00f80 l0057 ( .d(n476), .o(delay_add_ln22_unr23_stage9_stallmux_q_19_), .ck(clk) );
ms00f80 l0058 ( .d(n481), .o(cos_out_17), .ck(clk) );
ms00f80 l0059 ( .d(n485), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_29_), .ck(clk) );
ms00f80 l0060 ( .d(n490), .o(delay_add_ln22_unr5_stage3_stallmux_q_27_), .ck(clk) );
ms00f80 l0061 ( .d(n495), .o(delay_add_ln22_unr11_stage5_stallmux_q_25_), .ck(clk) );
ms00f80 l0062 ( .d(n500), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_16_), .ck(clk) );
ms00f80 l0063 ( .d(n505), .o(sin_out_9), .ck(clk) );
ms00f80 l0064 ( .d(n509), .o(delay_xor_ln22_unr12_stage5_stallmux_q_0_), .ck(clk) );
ms00f80 l0065 ( .d(n514), .o(delay_xor_ln21_unr6_stage3_stallmux_q_0_), .ck(clk) );
ms00f80 l0066 ( .d(n519), .o(delay_xor_ln22_unr21_stage8_stallmux_q_6_), .ck(clk) );
ms00f80 l0067 ( .d(n524), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_29_), .ck(clk) );
ms00f80 l0068 ( .d(n529), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_17_), .ck(clk) );
ms00f80 l0069 ( .d(n534), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_22_), .ck(clk) );
ms00f80 l0070 ( .d(n539), .o(delay_sub_ln22_unr24_stage9_stallmux_q_6_), .ck(clk) );
ms00f80 l0071 ( .d(n544), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_8_), .ck(clk) );
ms00f80 l0072 ( .d(n549), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_2_), .ck(clk) );
ms00f80 l0073 ( .d(n554), .o(delay_add_ln22_unr2_stage2_stallmux_q_27_), .ck(clk) );
ms00f80 l0074 ( .d(n559), .o(delay_add_ln22_unr2_stage2_stallmux_q_6_), .ck(clk) );
ms00f80 l0075 ( .d(n564), .o(delay_xor_ln21_unr15_stage6_stallmux_q_10_), .ck(clk) );
ms00f80 l0076 ( .d(n569), .o(delay_sub_ln23_0_unr30_stage10_stallmux_q), .ck(clk) );
ms00f80 l0077 ( .d(n574), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_11_), .ck(clk) );
ms00f80 l0078 ( .d(n579), .o(delay_xor_ln22_unr15_stage6_stallmux_q_7_), .ck(clk) );
ms00f80 l0079 ( .d(n584), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_23_), .ck(clk) );
ms00f80 l0080 ( .d(n589), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_18_), .ck(clk) );
ms00f80 l0081 ( .d(n594), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_24_), .ck(clk) );
ms00f80 l0082 ( .d(n599), .o(delay_add_ln22_unr2_stage2_stallmux_q_25_), .ck(clk) );
ms00f80 l0083 ( .d(n604), .o(delay_add_ln22_unr5_stage3_stallmux_q_12_), .ck(clk) );
ms00f80 l0084 ( .d(n609), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_18_), .ck(clk) );
ms00f80 l0085 ( .d(n614), .o(delay_add_ln22_unr27_stage10_stallmux_q_30_), .ck(clk) );
ms00f80 l0086 ( .d(n619), .o(delay_add_ln22_unr17_stage7_stallmux_q_14_), .ck(clk) );
ms00f80 l0087 ( .d(n624), .o(delay_add_ln22_unr14_stage6_stallmux_q_21_), .ck(clk) );
ms00f80 l0088 ( .d(n629), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_2_), .ck(clk) );
ms00f80 l0089 ( .d(n634), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_16_), .ck(clk) );
ms00f80 l0090 ( .d(n639), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_27_), .ck(clk) );
ms00f80 l0091 ( .d(n644), .o(delay_xor_ln22_unr6_stage3_stallmux_q_1_), .ck(clk) );
ms00f80 l0092 ( .d(n649), .o(sin_out_11), .ck(clk) );
ms00f80 l0093 ( .d(n653), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_13_), .ck(clk) );
ms00f80 l0094 ( .d(n658), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_5_), .ck(clk) );
ms00f80 l0095 ( .d(n663), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_13_), .ck(clk) );
ms00f80 l0096 ( .d(n668), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_13_), .ck(clk) );
ms00f80 l0097 ( .d(n673), .o(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .ck(clk) );
ms00f80 l0098 ( .d(n678), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_18_), .ck(clk) );
ms00f80 l0099 ( .d(n683), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_15_), .ck(clk) );
ms00f80 l0100 ( .d(n688), .o(delay_add_ln22_unr14_stage6_stallmux_q_24_), .ck(clk) );
ms00f80 l0101 ( .d(n693), .o(delay_add_ln22_unr23_stage9_stallmux_q_18_), .ck(clk) );
ms00f80 l0102 ( .d(n698), .o(delay_xor_ln22_unr9_stage4_stallmux_q_10_), .ck(clk) );
ms00f80 l0103 ( .d(n703), .o(delay_add_ln22_unr23_stage9_stallmux_q_29_), .ck(clk) );
ms00f80 l0104 ( .d(n708), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_2_), .ck(clk) );
ms00f80 l0105 ( .d(n713), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_10_), .ck(clk) );
ms00f80 l0106 ( .d(n718), .o(delay_xor_ln22_unr3_stage2_stallmux_q_14_), .ck(clk) );
ms00f80 l0107 ( .d(n723), .o(sin_out_6), .ck(clk) );
ms00f80 l0108 ( .d(n727), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_22_), .ck(clk) );
ms00f80 l0109 ( .d(n732), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_17_), .ck(clk) );
ms00f80 l0110 ( .d(n737), .o(delay_xor_ln22_unr12_stage5_stallmux_q_7_), .ck(clk) );
ms00f80 l0111 ( .d(n742), .o(delay_add_ln22_unr5_stage3_stallmux_q_15_), .ck(clk) );
ms00f80 l0112 ( .d(n747), .o(delay_xor_ln22_unr3_stage2_stallmux_q_9_), .ck(clk) );
ms00f80 l0113 ( .d(n752), .o(cos_out_12), .ck(clk) );
ms00f80 l0114 ( .d(n756), .o(delay_add_ln22_unr17_stage7_stallmux_q_24_), .ck(clk) );
ms00f80 l0115 ( .d(n761), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_21_), .ck(clk) );
ms00f80 l0116 ( .d(n765), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_0_), .ck(clk) );
ms00f80 l0117 ( .d(n770), .o(delay_xor_ln22_unr18_stage7_stallmux_q_12_), .ck(clk) );
ms00f80 l0118 ( .d(n775), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_23_), .ck(clk) );
ms00f80 l0119 ( .d(n780), .o(delay_add_ln22_unr20_stage8_stallmux_q_10_), .ck(clk) );
ms00f80 l0120 ( .d(n785), .o(delay_add_ln22_unr5_stage3_stallmux_q_20_), .ck(clk) );
ms00f80 l0121 ( .d(n790), .o(sin_out_12), .ck(clk) );
ms00f80 l0122 ( .d(n794), .o(delay_xor_ln22_unr18_stage7_stallmux_q_0_), .ck(clk) );
ms00f80 l0123 ( .d(n799), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_10_), .ck(clk) );
ms00f80 l0124 ( .d(n804), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_26_), .ck(clk) );
ms00f80 l0125 ( .d(n809), .o(delay_xor_ln22_unr3_stage2_stallmux_q_15_), .ck(clk) );
ms00f80 l0126 ( .d(n814), .o(sin_out_17), .ck(clk) );
ms00f80 l0127 ( .d(n818), .o(cordic_combinational_sub_ln23_0_unr16_z_0_), .ck(clk) );
ms00f80 l0128 ( .d(n823), .o(delay_xor_ln21_unr3_stage2_stallmux_q_27_), .ck(clk) );
ms00f80 l0129 ( .d(n828), .o(delay_add_ln22_unr14_stage6_stallmux_q_30_), .ck(clk) );
ms00f80 l0130 ( .d(n833), .o(delay_xor_ln22_unr3_stage2_stallmux_q_10_), .ck(clk) );
ms00f80 l0131 ( .d(n838), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_29_), .ck(clk) );
ms00f80 l0132 ( .d(n843), .o(cos_out_20), .ck(clk) );
ms00f80 l0133 ( .d(n847), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_15_), .ck(clk) );
ms00f80 l0134 ( .d(n852), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_10_), .ck(clk) );
ms00f80 l0135 ( .d(n857), .o(delay_sub_ln23_0_unr1_stage2_stallmux_q_1_), .ck(clk) );
ms00f80 l0136 ( .d(n862), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_4_), .ck(clk) );
ms00f80 l0137 ( .d(n867), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_12_), .ck(clk) );
ms00f80 l0138 ( .d(n872), .o(cos_out_14), .ck(clk) );
ms00f80 l0139 ( .d(n876), .o(delay_xor_ln21_unr15_stage6_stallmux_q_5_), .ck(clk) );
ms00f80 l0140 ( .d(n881), .o(delay_xor_ln22_unr9_stage4_stallmux_q_13_), .ck(clk) );
ms00f80 l0141 ( .d(n886), .o(delay_xor_ln21_unr6_stage3_stallmux_q_4_), .ck(clk) );
ms00f80 l0142 ( .d(n891), .o(delay_add_ln22_unr17_stage7_stallmux_q_25_), .ck(clk) );
ms00f80 l0143 ( .d(n896), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_24_), .ck(clk) );
ms00f80 l0144 ( .d(n901), .o(delay_add_ln22_unr27_stage10_stallmux_q_31_), .ck(clk) );
ms00f80 l0145 ( .d(n906), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_14_), .ck(clk) );
ms00f80 l0146 ( .d(n911), .o(delay_sub_ln23_unr9_stage4_stallmux_q_3_), .ck(clk) );
ms00f80 l0147 ( .d(n916), .o(delay_add_ln22_unr17_stage7_stallmux_q_8_), .ck(clk) );
ms00f80 l0148 ( .d(n921), .o(delay_add_ln22_unr2_stage2_stallmux_q_20_), .ck(clk) );
ms00f80 l0149 ( .d(n926), .o(delay_add_ln22_unr20_stage8_stallmux_q_26_), .ck(clk) );
ms00f80 l0150 ( .d(n931), .o(delay_add_ln22_unr11_stage5_stallmux_q_30_), .ck(clk) );
ms00f80 l0151 ( .d(n936), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_12_), .ck(clk) );
ms00f80 l0152 ( .d(n941), .o(delay_xor_ln21_unr12_stage5_stallmux_q_18_), .ck(clk) );
ms00f80 l0153 ( .d(n946), .o(delay_add_ln22_unr20_stage8_stallmux_q_13_), .ck(clk) );
ms00f80 l0154 ( .d(n951), .o(delay_add_ln22_unr8_stage4_stallmux_q_12_), .ck(clk) );
ms00f80 l0155 ( .d(n956), .o(delay_add_ln22_unr20_stage8_stallmux_q_14_), .ck(clk) );
ms00f80 l0156 ( .d(n961), .o(delay_xor_ln21_unr12_stage5_stallmux_q_12_), .ck(clk) );
ms00f80 l0157 ( .d(n966), .o(delay_add_ln22_unr23_stage9_stallmux_q_0_), .ck(clk) );
ms00f80 l0158 ( .d(n971), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_27_), .ck(clk) );
ms00f80 l0159 ( .d(n976), .o(delay_add_ln22_unr11_stage5_stallmux_q_17_), .ck(clk) );
ms00f80 l0160 ( .d(n981), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_12_), .ck(clk) );
ms00f80 l0161 ( .d(n986), .o(delay_xor_ln21_unr6_stage3_stallmux_q_18_), .ck(clk) );
ms00f80 l0162 ( .d(n991), .o(n_17093), .ck(clk) );
ms00f80 l0163 ( .d(n996), .o(delay_add_ln22_unr20_stage8_stallmux_q_24_), .ck(clk) );
ms00f80 l0164 ( .d(n1001), .o(delay_xor_ln21_unr6_stage3_stallmux_q_8_), .ck(clk) );
ms00f80 l0165 ( .d(n1006), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_20_), .ck(clk) );
ms00f80 l0166 ( .d(n1011), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_25_), .ck(clk) );
ms00f80 l0167 ( .d(n1016), .o(delay_xor_ln21_unr15_stage6_stallmux_q_11_), .ck(clk) );
ms00f80 l0168 ( .d(n1021), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_26_), .ck(clk) );
ms00f80 l0169 ( .d(n1026), .o(delay_xor_ln21_unr9_stage4_stallmux_q_3_), .ck(clk) );
ms00f80 l0170 ( .d(n1031), .o(sin_out_3), .ck(clk) );
ms00f80 l0171 ( .d(n1035), .o(delay_add_ln22_unr20_stage8_stallmux_q_15_), .ck(clk) );
ms00f80 l0172 ( .d(n1040), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_29_), .ck(clk) );
ms00f80 l0173 ( .d(n1045), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_14_), .ck(clk) );
ms00f80 l0174 ( .d(n1050), .o(delay_add_ln22_unr2_stage2_stallmux_q_5_), .ck(clk) );
ms00f80 l0175 ( .d(n1055), .o(delay_add_ln22_unr20_stage8_stallmux_q_18_), .ck(clk) );
ms00f80 l0176 ( .d(n1060), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_2_), .ck(clk) );
ms00f80 l0177 ( .d(n1065), .o(delay_add_ln22_unr23_stage9_stallmux_q_21_), .ck(clk) );
ms00f80 l0178 ( .d(n1070), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_16_), .ck(clk) );
ms00f80 l0179 ( .d(n1075), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_24_), .ck(clk) );
ms00f80 l0180 ( .d(n1080), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_9_), .ck(clk) );
ms00f80 l0181 ( .d(n1085), .o(delay_xor_ln21_unr3_stage2_stallmux_q_0_), .ck(clk) );
ms00f80 l0182 ( .d(n1090), .o(delay_add_ln22_unr5_stage3_stallmux_q_25_), .ck(clk) );
ms00f80 l0183 ( .d(n1095), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_16_), .ck(clk) );
ms00f80 l0184 ( .d(n1100), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_7_), .ck(clk) );
ms00f80 l0185 ( .d(n1105), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_28_), .ck(clk) );
ms00f80 l0186 ( .d(n1110), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_9_), .ck(clk) );
ms00f80 l0187 ( .d(n1115), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_12_), .ck(clk) );
ms00f80 l0188 ( .d(n1120), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_11_), .ck(clk) );
ms00f80 l0189 ( .d(n1125), .o(delay_xor_ln21_unr15_stage6_stallmux_q_12_), .ck(clk) );
ms00f80 l0190 ( .d(n1130), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_18_), .ck(clk) );
ms00f80 l0191 ( .d(n1135), .o(n_27923), .ck(clk) );
ms00f80 l0192 ( .d(n1140), .o(delay_add_ln22_unr27_stage10_stallmux_q_25_), .ck(clk) );
ms00f80 l0193 ( .d(n1145), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_8_), .ck(clk) );
ms00f80 l0194 ( .d(n1150), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_15_), .ck(clk) );
ms00f80 l0195 ( .d(n1155), .o(delay_add_ln22_unr11_stage5_stallmux_q_0_), .ck(clk) );
ms00f80 l0196 ( .d(n1160), .o(delay_xor_ln22_unr3_stage2_stallmux_q_3_), .ck(clk) );
ms00f80 l0197 ( .d(n1165), .o(delay_xor_ln21_unr21_stage8_stallmux_q_9_), .ck(clk) );
ms00f80 l0198 ( .d(n1170), .o(delay_xor_ln21_unr3_stage2_stallmux_q_21_), .ck(clk) );
ms00f80 l0199 ( .d(n1175), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_30_), .ck(clk) );
ms00f80 l0200 ( .d(n1180), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_0_), .ck(clk) );
ms00f80 l0201 ( .d(n1185), .o(delay_xor_ln21_unr9_stage4_stallmux_q_15_), .ck(clk) );
ms00f80 l0202 ( .d(n1190), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_15_), .ck(clk) );
ms00f80 l0203 ( .d(n1195), .o(delay_add_ln22_unr2_stage2_stallmux_q_26_), .ck(clk) );
ms00f80 l0204 ( .d(n1200), .o(delay_xor_ln21_unr9_stage4_stallmux_q_5_), .ck(clk) );
ms00f80 l0205 ( .d(n1205), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_26_), .ck(clk) );
ms00f80 l0206 ( .d(n1210), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_24_), .ck(clk) );
ms00f80 l0207 ( .d(n1215), .o(delay_xor_ln22_unr3_stage2_stallmux_q_1_), .ck(clk) );
ms00f80 l0208 ( .d(n1220), .o(delay_xor_ln22_unr9_stage4_stallmux_q_15_), .ck(clk) );
ms00f80 l0209 ( .d(n1225), .o(delay_xor_ln21_unr18_stage7_stallmux_q_13_), .ck(clk) );
ms00f80 l0210 ( .d(n1230), .o(delay_add_ln22_unr23_stage9_stallmux_q_23_), .ck(clk) );
ms00f80 l0211 ( .d(n1235), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_28_), .ck(clk) );
ms00f80 l0212 ( .d(n1240), .o(delay_xor_ln22_unr12_stage5_stallmux_q_1_), .ck(clk) );
ms00f80 l0213 ( .d(n1245), .o(delay_xor_ln21_unr12_stage5_stallmux_q_11_), .ck(clk) );
ms00f80 l0214 ( .d(n1250), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_31_), .ck(clk) );
ms00f80 l0215 ( .d(n1255), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_8_), .ck(clk) );
ms00f80 l0216 ( .d(n1260), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_1_), .ck(clk) );
ms00f80 l0217 ( .d(n1265), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_12_), .ck(clk) );
ms00f80 l0218 ( .d(n1270), .o(delay_add_ln22_unr27_stage10_stallmux_q_9_), .ck(clk) );
ms00f80 l0219 ( .d(n1275), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_27_), .ck(clk) );
ms00f80 l0220 ( .d(n1280), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_21_), .ck(clk) );
ms00f80 l0221 ( .d(n1285), .o(delay_add_ln22_unr11_stage5_stallmux_q_12_), .ck(clk) );
ms00f80 l0222 ( .d(n1290), .o(delay_add_ln22_unr5_stage3_stallmux_q_17_), .ck(clk) );
ms00f80 l0223 ( .d(n1295), .o(delay_add_ln22_unr17_stage7_stallmux_q_27_), .ck(clk) );
ms00f80 l0224 ( .d(n1300), .o(delay_xor_ln21_unr9_stage4_stallmux_q_21_), .ck(clk) );
ms00f80 l0225 ( .d(n1305), .o(delay_xor_ln22_unr15_stage6_stallmux_q_16_), .ck(clk) );
ms00f80 l0226 ( .d(n1310), .o(delay_xor_ln21_unr12_stage5_stallmux_q_7_), .ck(clk) );
ms00f80 l0227 ( .d(n1315), .o(sin_out_25), .ck(clk) );
ms00f80 l0228 ( .d(n1319), .o(delay_xor_ln22_unr9_stage4_stallmux_q_19_), .ck(clk) );
ms00f80 l0229 ( .d(n1324), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_6_), .ck(clk) );
ms00f80 l0230 ( .d(n1329), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_9_), .ck(clk) );
ms00f80 l0231 ( .d(n1334), .o(mux_while_ln12_psv_q_7_), .ck(clk) );
ms00f80 l0232 ( .d(n1339), .o(delay_add_ln22_unr23_stage9_stallmux_q_16_), .ck(clk) );
ms00f80 l0233 ( .d(n1344), .o(cos_out_2), .ck(clk) );
ms00f80 l0234 ( .d(n1348), .o(delay_xor_ln22_unr3_stage2_stallmux_q_19_), .ck(clk) );
ms00f80 l0235 ( .d(n1353), .o(delay_add_ln22_unr20_stage8_stallmux_q_5_), .ck(clk) );
ms00f80 l0236 ( .d(n1358), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_9_), .ck(clk) );
ms00f80 l0237 ( .d(n1363), .o(delay_xor_ln21_unr3_stage2_stallmux_q_5_), .ck(clk) );
ms00f80 l0238 ( .d(n1368), .o(delay_add_ln22_unr11_stage5_stallmux_q_4_), .ck(clk) );
ms00f80 l0239 ( .d(n1373), .o(cos_out_22), .ck(clk) );
ms00f80 l0240 ( .d(n1377), .o(delay_add_ln22_unr17_stage7_stallmux_q_3_), .ck(clk) );
ms00f80 l0241 ( .d(n1382), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_26_), .ck(clk) );
ms00f80 l0242 ( .d(n1387), .o(delay_xor_ln22_unr6_stage3_stallmux_q_18_), .ck(clk) );
ms00f80 l0243 ( .d(n1392), .o(cos_out_31), .ck(clk) );
ms00f80 l0244 ( .d(n1396), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_26_), .ck(clk) );
ms00f80 l0245 ( .d(n1401), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_2_), .ck(clk) );
ms00f80 l0246 ( .d(n1406), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_23_), .ck(clk) );
ms00f80 l0247 ( .d(n1411), .o(delay_xor_ln21_unr6_stage3_stallmux_q_25_), .ck(clk) );
ms00f80 l0248 ( .d(n1416), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_8_), .ck(clk) );
ms00f80 l0249 ( .d(n1421), .o(delay_xor_ln22_unr21_stage8_stallmux_q_10_), .ck(clk) );
ms00f80 l0250 ( .d(n1426), .o(delay_add_ln22_unr17_stage7_stallmux_q_1_), .ck(clk) );
ms00f80 l0251 ( .d(n1431), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_5_), .ck(clk) );
ms00f80 l0252 ( .d(n1436), .o(delay_add_ln22_unr23_stage9_stallmux_q_11_), .ck(clk) );
ms00f80 l0253 ( .d(n1441), .o(delay_xor_ln21_unr3_stage2_stallmux_q_10_), .ck(clk) );
ms00f80 l0254 ( .d(n1446), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_27_), .ck(clk) );
ms00f80 l0255 ( .d(n1451), .o(delay_xor_ln22_unr6_stage3_stallmux_q_3_), .ck(clk) );
ms00f80 l0256 ( .d(n1456), .o(delay_xor_ln21_unr15_stage6_stallmux_q_8_), .ck(clk) );
ms00f80 l0257 ( .d(n1461), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_8_), .ck(clk) );
ms00f80 l0258 ( .d(n1466), .o(delay_add_ln22_unr23_stage9_stallmux_q_1_), .ck(clk) );
ms00f80 l0259 ( .d(n1471), .o(delay_xor_ln21_unr18_stage7_stallmux_q_10_), .ck(clk) );
ms00f80 l0260 ( .d(n1476), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_19_), .ck(clk) );
ms00f80 l0261 ( .d(n1481), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_21_), .ck(clk) );
ms00f80 l0262 ( .d(n1486), .o(delay_add_ln22_unr14_stage6_stallmux_q_1_), .ck(clk) );
ms00f80 l0263 ( .d(n1491), .o(delay_xor_ln21_unr18_stage7_stallmux_q_12_), .ck(clk) );
ms00f80 l0264 ( .d(n1496), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_29_), .ck(clk) );
ms00f80 l0265 ( .d(n1501), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_10_), .ck(clk) );
ms00f80 l0266 ( .d(n1506), .o(delay_xor_ln21_unr6_stage3_stallmux_q_7_), .ck(clk) );
ms00f80 l0267 ( .d(n1511), .o(delay_add_ln22_unr14_stage6_stallmux_q_29_), .ck(clk) );
ms00f80 l0268 ( .d(n1516), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_20_), .ck(clk) );
ms00f80 l0269 ( .d(n1521), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_3_), .ck(clk) );
ms00f80 l0270 ( .d(n1526), .o(delay_xor_ln22_unr3_stage2_stallmux_q_28_), .ck(clk) );
ms00f80 l0271 ( .d(n1531), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_7_), .ck(clk) );
ms00f80 l0272 ( .d(n1536), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_15_), .ck(clk) );
ms00f80 l0273 ( .d(n1540), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .ck(clk) );
ms00f80 l0274 ( .d(n1545), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_11_), .ck(clk) );
ms00f80 l0275 ( .d(n1550), .o(delay_xor_ln22_unr6_stage3_stallmux_q_25_), .ck(clk) );
ms00f80 l0276 ( .d(n1555), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_26_), .ck(clk) );
ms00f80 l0277 ( .d(n1560), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_12_), .ck(clk) );
ms00f80 l0278 ( .d(n1565), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_0_), .ck(clk) );
ms00f80 l0279 ( .d(n1570), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_18_), .ck(clk) );
ms00f80 l0280 ( .d(n1575), .o(delay_add_ln22_unr5_stage3_stallmux_q_2_), .ck(clk) );
ms00f80 l0281 ( .d(n1580), .o(delay_add_ln22_unr8_stage4_stallmux_q_18_), .ck(clk) );
ms00f80 l0282 ( .d(n1585), .o(delay_add_ln22_unr17_stage7_stallmux_q_10_), .ck(clk) );
ms00f80 l0283 ( .d(n1590), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_21_), .ck(clk) );
ms00f80 l0284 ( .d(n1595), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_29_), .ck(clk) );
ms00f80 l0285 ( .d(n1600), .o(delay_add_ln22_unr14_stage6_stallmux_q_5_), .ck(clk) );
ms00f80 l0286 ( .d(n1605), .o(delay_xor_ln21_unr6_stage3_stallmux_q_2_), .ck(clk) );
ms00f80 l0287 ( .d(n1610), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_23_), .ck(clk) );
ms00f80 l0288 ( .d(n1615), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_4_), .ck(clk) );
ms00f80 l0289 ( .d(n1620), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_27_), .ck(clk) );
ms00f80 l0290 ( .d(n1625), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_25_), .ck(clk) );
ms00f80 l0291 ( .d(n1630), .o(delay_add_ln22_unr8_stage4_stallmux_q_3_), .ck(clk) );
ms00f80 l0292 ( .d(n1635), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_19_), .ck(clk) );
ms00f80 l0293 ( .d(n1640), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_13_), .ck(clk) );
ms00f80 l0294 ( .d(n1645), .o(delay_add_ln22_unr2_stage2_stallmux_q_8_), .ck(clk) );
ms00f80 l0295 ( .d(n1650), .o(mux_while_ln12_psv_q_8_), .ck(clk) );
ms00f80 l0296 ( .d(n1655), .o(delay_xor_ln21_unr9_stage4_stallmux_q_7_), .ck(clk) );
ms00f80 l0297 ( .d(n1660), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_28_), .ck(clk) );
ms00f80 l0298 ( .d(n1664), .o(delay_xor_ln22_unr3_stage2_stallmux_q_27_), .ck(clk) );
ms00f80 l0299 ( .d(n1669), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_21_), .ck(clk) );
ms00f80 l0300 ( .d(n1674), .o(delay_add_ln22_unr11_stage5_stallmux_q_7_), .ck(clk) );
ms00f80 l0301 ( .d(n1679), .o(delay_sub_ln22_unr24_stage9_stallmux_q_7_), .ck(clk) );
ms00f80 l0302 ( .d(n1684), .o(delay_xor_ln21_unr9_stage4_stallmux_q_11_), .ck(clk) );
ms00f80 l0303 ( .d(n1689), .o(delay_add_ln22_unr11_stage5_stallmux_q_13_), .ck(clk) );
ms00f80 l0304 ( .d(n1694), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_17_), .ck(clk) );
ms00f80 l0305 ( .d(n1699), .o(delay_xor_ln22_unr3_stage2_stallmux_q_13_), .ck(clk) );
ms00f80 l0306 ( .d(n1704), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_25_), .ck(clk) );
ms00f80 l0307 ( .d(n1709), .o(delay_add_ln22_unr23_stage9_stallmux_q_20_), .ck(clk) );
ms00f80 l0308 ( .d(n1714), .o(delay_add_ln22_unr11_stage5_stallmux_q_26_), .ck(clk) );
ms00f80 l0309 ( .d(n1719), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_18_), .ck(clk) );
ms00f80 l0310 ( .d(n1724), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_4_), .ck(clk) );
ms00f80 l0311 ( .d(n1729), .o(delay_add_ln22_unr5_stage3_stallmux_q_8_), .ck(clk) );
ms00f80 l0312 ( .d(n1734), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_18_), .ck(clk) );
ms00f80 l0313 ( .d(n1739), .o(delay_add_ln22_unr5_stage3_stallmux_q_7_), .ck(clk) );
ms00f80 l0314 ( .d(n1744), .o(delay_xor_ln22_unr12_stage5_stallmux_q_19_), .ck(clk) );
ms00f80 l0315 ( .d(n1749), .o(delay_add_ln22_unr20_stage8_stallmux_q_1_), .ck(clk) );
ms00f80 l0316 ( .d(n1754), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_13_), .ck(clk) );
ms00f80 l0317 ( .d(n1759), .o(delay_xor_ln22_unr12_stage5_stallmux_q_3_), .ck(clk) );
ms00f80 l0318 ( .d(n1763), .o(cordic_combinational_sub_ln23_0_unr20_z_0_), .ck(clk) );
ms00f80 l0319 ( .d(n1767), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_18_), .ck(clk) );
ms00f80 l0320 ( .d(n1772), .o(delay_add_ln22_unr14_stage6_stallmux_q_9_), .ck(clk) );
ms00f80 l0321 ( .d(n1777), .o(delay_xor_ln22_unr18_stage7_stallmux_q_6_), .ck(clk) );
ms00f80 l0322 ( .d(n1782), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_19_), .ck(clk) );
ms00f80 l0323 ( .d(n1787), .o(delay_add_ln22_unr27_stage10_stallmux_q_14_), .ck(clk) );
ms00f80 l0324 ( .d(n1792), .o(cos_out_26), .ck(clk) );
ms00f80 l0325 ( .d(n1796), .o(delay_add_ln22_unr23_stage9_stallmux_q_28_), .ck(clk) );
ms00f80 l0326 ( .d(n1801), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_29_), .ck(clk) );
ms00f80 l0327 ( .d(n1806), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_25_), .ck(clk) );
ms00f80 l0328 ( .d(n1811), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_26_), .ck(clk) );
ms00f80 l0329 ( .d(n1816), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_16_), .ck(clk) );
ms00f80 l0330 ( .d(n1821), .o(n_44061), .ck(clk) );
ms00f80 l0331 ( .d(n1826), .o(delay_add_ln22_unr8_stage4_stallmux_q_2_), .ck(clk) );
ms00f80 l0332 ( .d(n1831), .o(sin_out_10), .ck(clk) );
ms00f80 l0333 ( .d(n1835), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_28_), .ck(clk) );
ms00f80 l0334 ( .d(n1840), .o(delay_sub_ln21_unr24_stage9_stallmux_q_6_), .ck(clk) );
ms00f80 l0335 ( .d(n1845), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_22_), .ck(clk) );
ms00f80 l0336 ( .d(n1850), .o(delay_add_ln22_unr27_stage10_stallmux_q_21_), .ck(clk) );
ms00f80 l0337 ( .d(n1855), .o(delay_xor_ln21_unr3_stage2_stallmux_q_4_), .ck(clk) );
ms00f80 l0338 ( .d(n1860), .o(delay_xor_ln21_unr9_stage4_stallmux_q_13_), .ck(clk) );
ms00f80 l0339 ( .d(n1865), .o(cos_out_30), .ck(clk) );
ms00f80 l0340 ( .d(n1869), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_0_), .ck(clk) );
ms00f80 l0341 ( .d(n1874), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_13_), .ck(clk) );
ms00f80 l0342 ( .d(n1879), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_3_), .ck(clk) );
ms00f80 l0343 ( .d(n1884), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_24_), .ck(clk) );
ms00f80 l0344 ( .d(n1889), .o(delay_add_ln22_unr14_stage6_stallmux_q_20_), .ck(clk) );
ms00f80 l0345 ( .d(n1894), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_20_), .ck(clk) );
ms00f80 l0346 ( .d(n1899), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_14_), .ck(clk) );
ms00f80 l0347 ( .d(n1904), .o(delay_add_ln22_unr11_stage5_stallmux_q_6_), .ck(clk) );
ms00f80 l0348 ( .d(n1909), .o(delay_xor_ln22_unr12_stage5_stallmux_q_16_), .ck(clk) );
ms00f80 l0349 ( .d(n1914), .o(delay_add_ln22_unr8_stage4_stallmux_q_13_), .ck(clk) );
ms00f80 l0350 ( .d(n1919), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_2_), .ck(clk) );
ms00f80 l0351 ( .d(n1924), .o(delay_xor_ln21_unr21_stage8_stallmux_q_0_), .ck(clk) );
ms00f80 l0352 ( .d(n1929), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_14_), .ck(clk) );
ms00f80 l0353 ( .d(n1934), .o(delay_add_ln22_unr8_stage4_stallmux_q_23_), .ck(clk) );
ms00f80 l0354 ( .d(n1939), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_19_), .ck(clk) );
ms00f80 l0355 ( .d(n1944), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_26_), .ck(clk) );
ms00f80 l0356 ( .d(n1949), .o(delay_xor_ln21_unr15_stage6_stallmux_q_14_), .ck(clk) );
ms00f80 l0357 ( .d(n1954), .o(delay_add_ln22_unr27_stage10_stallmux_q_13_), .ck(clk) );
ms00f80 l0358 ( .d(n1959), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_17_), .ck(clk) );
ms00f80 l0359 ( .d(n1964), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_7_), .ck(clk) );
ms00f80 l0360 ( .d(n1969), .o(delay_add_ln22_unr17_stage7_stallmux_q_13_), .ck(clk) );
ms00f80 l0361 ( .d(n1974), .o(delay_xor_ln22_unr15_stage6_stallmux_q_13_), .ck(clk) );
ms00f80 l0362 ( .d(n1979), .o(sin_out_1), .ck(clk) );
ms00f80 l0363 ( .d(n1983), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_20_), .ck(clk) );
ms00f80 l0364 ( .d(n1988), .o(delay_xor_ln22_unr9_stage4_stallmux_q_18_), .ck(clk) );
ms00f80 l0365 ( .d(n1993), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_10_), .ck(clk) );
ms00f80 l0366 ( .d(n1998), .o(delay_xor_ln22_unr18_stage7_stallmux_q_5_), .ck(clk) );
ms00f80 l0367 ( .d(n2003), .o(delay_add_ln22_unr11_stage5_stallmux_q_24_), .ck(clk) );
ms00f80 l0368 ( .d(n2008), .o(delay_add_ln22_unr27_stage10_stallmux_q_5_), .ck(clk) );
ms00f80 l0369 ( .d(n2013), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_22_), .ck(clk) );
ms00f80 l0370 ( .d(n2018), .o(delay_add_ln22_unr20_stage8_stallmux_q_30_), .ck(clk) );
ms00f80 l0371 ( .d(n2023), .o(delay_add_ln22_unr27_stage10_stallmux_q_11_), .ck(clk) );
ms00f80 l0372 ( .d(n2028), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_3_), .ck(clk) );
ms00f80 l0373 ( .d(n2033), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_16_), .ck(clk) );
ms00f80 l0374 ( .d(n2038), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_7_), .ck(clk) );
ms00f80 l0375 ( .d(n2043), .o(delay_xor_ln21_unr3_stage2_stallmux_q_25_), .ck(clk) );
ms00f80 l0376 ( .d(n2048), .o(delay_add_ln22_unr8_stage4_stallmux_q_14_), .ck(clk) );
ms00f80 l0377 ( .d(n2053), .o(delay_sub_ln21_unr24_stage9_stallmux_q_5_), .ck(clk) );
ms00f80 l0378 ( .d(n2058), .o(delay_add_ln22_unr11_stage5_stallmux_q_14_), .ck(clk) );
ms00f80 l0379 ( .d(n2063), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_16_), .ck(clk) );
ms00f80 l0380 ( .d(n2068), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_9_), .ck(clk) );
ms00f80 l0381 ( .d(n2072), .o(delay_xor_ln22_unr3_stage2_stallmux_q_6_), .ck(clk) );
ms00f80 l0382 ( .d(n2077), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_30_), .ck(clk) );
ms00f80 l0383 ( .d(n2082), .o(delay_add_ln22_unr14_stage6_stallmux_q_15_), .ck(clk) );
ms00f80 l0384 ( .d(n2087), .o(delay_xor_ln21_unr21_stage8_stallmux_q_2_), .ck(clk) );
ms00f80 l0385 ( .d(n2092), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_25_), .ck(clk) );
ms00f80 l0386 ( .d(n2097), .o(delay_xor_ln22_unr18_stage7_stallmux_q_4_), .ck(clk) );
ms00f80 l0387 ( .d(n2102), .o(delay_add_ln22_unr2_stage2_stallmux_q_12_), .ck(clk) );
ms00f80 l0388 ( .d(n2107), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_9_), .ck(clk) );
ms00f80 l0389 ( .d(n2112), .o(delay_xor_ln21_unr9_stage4_stallmux_q_2_), .ck(clk) );
ms00f80 l0390 ( .d(n2117), .o(cos_out_27), .ck(clk) );
ms00f80 l0391 ( .d(n2121), .o(delay_xor_ln21_unr12_stage5_stallmux_q_4_), .ck(clk) );
ms00f80 l0392 ( .d(n2126), .o(delay_xor_ln22_unr12_stage5_stallmux_q_18_), .ck(clk) );
ms00f80 l0393 ( .d(n2131), .o(n_22641), .ck(clk) );
ms00f80 l0394 ( .d(n2136), .o(delay_add_ln22_unr27_stage10_stallmux_q_19_), .ck(clk) );
ms00f80 l0395 ( .d(n2141), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_27_), .ck(clk) );
ms00f80 l0396 ( .d(n2146), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_3_), .ck(clk) );
ms00f80 l0397 ( .d(n2151), .o(cos_out_25), .ck(clk) );
ms00f80 l0398 ( .d(n2155), .o(delay_xor_ln22_unr21_stage8_stallmux_q_5_), .ck(clk) );
ms00f80 l0399 ( .d(n2160), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_18_), .ck(clk) );
ms00f80 l0400 ( .d(n2165), .o(cos_out_7), .ck(clk) );
ms00f80 l0401 ( .d(n2169), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_16_), .ck(clk) );
ms00f80 l0402 ( .d(n2174), .o(delay_xor_ln21_unr18_stage7_stallmux_q_8_), .ck(clk) );
ms00f80 l0403 ( .d(n2179), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_25_), .ck(clk) );
ms00f80 l0404 ( .d(n2184), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_4_), .ck(clk) );
ms00f80 l0405 ( .d(n2189), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_2_), .ck(clk) );
ms00f80 l0406 ( .d(n2194), .o(sin_out_15), .ck(clk) );
ms00f80 l0407 ( .d(n2198), .o(delay_xor_ln22_unr9_stage4_stallmux_q_22_), .ck(clk) );
ms00f80 l0408 ( .d(n2203), .o(delay_xor_ln21_unr9_stage4_stallmux_q_20_), .ck(clk) );
ms00f80 l0409 ( .d(n2208), .o(delay_add_ln22_unr17_stage7_stallmux_q_4_), .ck(clk) );
ms00f80 l0410 ( .d(n2213), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_26_), .ck(clk) );
ms00f80 l0411 ( .d(n2218), .o(delay_xor_ln22_unr12_stage5_stallmux_q_10_), .ck(clk) );
ms00f80 l0412 ( .d(n2223), .o(cos_out_6), .ck(clk) );
ms00f80 l0413 ( .d(n2227), .o(delay_xor_ln21_unr6_stage3_stallmux_q_6_), .ck(clk) );
ms00f80 l0414 ( .d(n2232), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_8_), .ck(clk) );
ms00f80 l0415 ( .d(n2237), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_31_), .ck(clk) );
ms00f80 l0416 ( .d(n2242), .o(delay_add_ln22_unr20_stage8_stallmux_q_4_), .ck(clk) );
ms00f80 l0417 ( .d(n2247), .o(delay_add_ln22_unr23_stage9_stallmux_q_8_), .ck(clk) );
ms00f80 l0418 ( .d(n2252), .o(delay_add_ln22_unr23_stage9_stallmux_q_17_), .ck(clk) );
ms00f80 l0419 ( .d(n2257), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_20_), .ck(clk) );
ms00f80 l0420 ( .d(n2262), .o(delay_add_ln22_unr27_stage10_stallmux_q_18_), .ck(clk) );
ms00f80 l0421 ( .d(n2267), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_14_), .ck(clk) );
ms00f80 l0422 ( .d(n2272), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_2_), .ck(clk) );
ms00f80 l0423 ( .d(n2277), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_7_), .ck(clk) );
ms00f80 l0424 ( .d(n2282), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_10_), .ck(clk) );
ms00f80 l0425 ( .d(n2287), .o(delay_add_ln22_unr2_stage2_stallmux_q_17_), .ck(clk) );
ms00f80 l0426 ( .d(n2292), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_12_), .ck(clk) );
ms00f80 l0427 ( .d(n2297), .o(delay_xor_ln21_unr15_stage6_stallmux_q_6_), .ck(clk) );
ms00f80 l0428 ( .d(n2302), .o(delay_add_ln22_unr2_stage2_stallmux_q_16_), .ck(clk) );
ms00f80 l0429 ( .d(n2307), .o(delay_xor_ln21_unr3_stage2_stallmux_q_13_), .ck(clk) );
ms00f80 l0430 ( .d(n2312), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_31_), .ck(clk) );
ms00f80 l0431 ( .d(n2317), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_19_), .ck(clk) );
ms00f80 l0432 ( .d(n2322), .o(delay_xor_ln21_unr6_stage3_stallmux_q_22_), .ck(clk) );
ms00f80 l0433 ( .d(n2327), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_29_), .ck(clk) );
ms00f80 l0434 ( .d(n2332), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_28_), .ck(clk) );
ms00f80 l0435 ( .d(n2337), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_9_), .ck(clk) );
ms00f80 l0436 ( .d(n2342), .o(n_44695), .ck(clk) );
ms00f80 l0437 ( .d(n2347), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_22_), .ck(clk) );
ms00f80 l0438 ( .d(n2352), .o(delay_xor_ln21_unr21_stage8_stallmux_q_7_), .ck(clk) );
ms00f80 l0439 ( .d(n2357), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_5_), .ck(clk) );
ms00f80 l0440 ( .d(n2362), .o(delay_xor_ln22_unr9_stage4_stallmux_q_3_), .ck(clk) );
ms00f80 l0441 ( .d(n2367), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_8_), .ck(clk) );
ms00f80 l0442 ( .d(n2372), .o(delay_sub_ln23_0_unr26_stage9_stallmux_q_1_), .ck(clk) );
ms00f80 l0443 ( .d(n2377), .o(delay_sub_ln23_0_unr29_stage10_stallmux_q), .ck(clk) );
ms00f80 l0444 ( .d(n2382), .o(delay_xor_ln21_unr9_stage4_stallmux_q_19_), .ck(clk) );
ms00f80 l0445 ( .d(n2387), .o(delay_xor_ln21_unr3_stage2_stallmux_q_17_), .ck(clk) );
ms00f80 l0446 ( .d(n2392), .o(delay_add_ln22_unr2_stage2_stallmux_q_2_), .ck(clk) );
ms00f80 l0447 ( .d(n2397), .o(delay_xor_ln22_unr6_stage3_stallmux_q_0_), .ck(clk) );
ms00f80 l0448 ( .d(n2402), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_9_), .ck(clk) );
ms00f80 l0449 ( .d(n2407), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_28_), .ck(clk) );
ms00f80 l0450 ( .d(n2412), .o(delay_xor_ln22_unr15_stage6_stallmux_q_3_), .ck(clk) );
ms00f80 l0451 ( .d(n2417), .o(mux_while_ln12_psv_q_5_), .ck(clk) );
ms00f80 l0452 ( .d(n2422), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_5_), .ck(clk) );
ms00f80 l0453 ( .d(n2427), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_23_), .ck(clk) );
ms00f80 l0454 ( .d(n2432), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_2_), .ck(clk) );
ms00f80 l0455 ( .d(n2437), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_9_), .ck(clk) );
ms00f80 l0456 ( .d(n2442), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_7_), .ck(clk) );
ms00f80 l0457 ( .d(n2447), .o(sin_out_22), .ck(clk) );
ms00f80 l0458 ( .d(n2451), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_8_), .ck(clk) );
ms00f80 l0459 ( .d(n2456), .o(delay_xor_ln22_unr12_stage5_stallmux_q_14_), .ck(clk) );
ms00f80 l0460 ( .d(n2461), .o(delay_xor_ln22_unr15_stage6_stallmux_q_10_), .ck(clk) );
ms00f80 l0461 ( .d(n2466), .o(delay_xor_ln21_unr15_stage6_stallmux_q_7_), .ck(clk) );
ms00f80 l0462 ( .d(n2471), .o(delay_xor_ln22_unr12_stage5_stallmux_q_12_), .ck(clk) );
ms00f80 l0463 ( .d(n2476), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_7_), .ck(clk) );
ms00f80 l0464 ( .d(n2481), .o(delay_add_ln22_unr11_stage5_stallmux_q_21_), .ck(clk) );
ms00f80 l0465 ( .d(n2486), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_28_), .ck(clk) );
ms00f80 l0466 ( .d(n2491), .o(delay_xor_ln21_unr3_stage2_stallmux_q_1_), .ck(clk) );
ms00f80 l0467 ( .d(n2496), .o(delay_xor_ln22_unr6_stage3_stallmux_q_16_), .ck(clk) );
ms00f80 l0468 ( .d(n2501), .o(delay_xor_ln21_unr18_stage7_stallmux_q_9_), .ck(clk) );
ms00f80 l0469 ( .d(n2506), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_22_), .ck(clk) );
ms00f80 l0470 ( .d(n2511), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_7_), .ck(clk) );
ms00f80 l0471 ( .d(n2516), .o(delay_add_ln22_unr2_stage2_stallmux_q_18_), .ck(clk) );
ms00f80 l0472 ( .d(n2521), .o(sin_out_23), .ck(clk) );
ms00f80 l0473 ( .d(n2525), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_10_), .ck(clk) );
ms00f80 l0474 ( .d(n2530), .o(delay_xor_ln22_unr3_stage2_stallmux_q_0_), .ck(clk) );
ms00f80 l0475 ( .d(n2535), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_1_), .ck(clk) );
ms00f80 l0476 ( .d(n2540), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_6_), .ck(clk) );
ms00f80 l0477 ( .d(n2545), .o(delay_xor_ln22_unr12_stage5_stallmux_q_9_), .ck(clk) );
ms00f80 l0478 ( .d(n2550), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_12_), .ck(clk) );
ms00f80 l0479 ( .d(n2555), .o(delay_add_ln22_unr23_stage9_stallmux_q_30_), .ck(clk) );
ms00f80 l0480 ( .d(n2560), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_5_), .ck(clk) );
ms00f80 l0481 ( .d(n2565), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_28_), .ck(clk) );
ms00f80 l0482 ( .d(n2570), .o(delay_add_ln22_unr11_stage5_stallmux_q_1_), .ck(clk) );
ms00f80 l0483 ( .d(n2575), .o(sin_out_4), .ck(clk) );
ms00f80 l0484 ( .d(n2579), .o(delay_sub_ln22_unr24_stage9_stallmux_q_1_), .ck(clk) );
ms00f80 l0485 ( .d(n2584), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_5_), .ck(clk) );
ms00f80 l0486 ( .d(n2589), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .ck(clk) );
ms00f80 l0487 ( .d(n2594), .o(delay_xor_ln22_unr18_stage7_stallmux_q_7_), .ck(clk) );
ms00f80 l0488 ( .d(n2599), .o(delay_xor_ln21_unr9_stage4_stallmux_q_6_), .ck(clk) );
ms00f80 l0489 ( .d(n2604), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_11_), .ck(clk) );
ms00f80 l0490 ( .d(n2609), .o(delay_xor_ln22_unr18_stage7_stallmux_q_13_), .ck(clk) );
ms00f80 l0491 ( .d(n2614), .o(cos_out_18), .ck(clk) );
ms00f80 l0492 ( .d(n2618), .o(delay_xor_ln22_unr6_stage3_stallmux_q_19_), .ck(clk) );
ms00f80 l0493 ( .d(n2623), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_3_), .ck(clk) );
ms00f80 l0494 ( .d(n2628), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_12_), .ck(clk) );
ms00f80 l0495 ( .d(n2633), .o(sin_out_2), .ck(clk) );
ms00f80 l0496 ( .d(n2637), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_8_), .ck(clk) );
ms00f80 l0497 ( .d(n2642), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_2_), .ck(clk) );
ms00f80 l0498 ( .d(n2647), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_7_), .ck(clk) );
ms00f80 l0499 ( .d(n2652), .o(mux_while_ln12_psv_q_4_), .ck(clk) );
ms00f80 l0500 ( .d(n2657), .o(delay_add_ln22_unr17_stage7_stallmux_q_7_), .ck(clk) );
ms00f80 l0501 ( .d(n2662), .o(delay_add_ln22_unr20_stage8_stallmux_q_25_), .ck(clk) );
ms00f80 l0502 ( .d(n2667), .o(delay_xor_ln22_unr3_stage2_stallmux_q_24_), .ck(clk) );
ms00f80 l0503 ( .d(n2672), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_22_), .ck(clk) );
ms00f80 l0504 ( .d(n2677), .o(delay_xor_ln21_unr12_stage5_stallmux_q_3_), .ck(clk) );
ms00f80 l0505 ( .d(n2682), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_13_), .ck(clk) );
ms00f80 l0506 ( .d(n2687), .o(delay_add_ln22_unr23_stage9_stallmux_q_31_), .ck(clk) );
ms00f80 l0507 ( .d(n2692), .o(delay_xor_ln22_unr21_stage8_stallmux_q_1_), .ck(clk) );
ms00f80 l0508 ( .d(n2697), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_27_), .ck(clk) );
ms00f80 l0509 ( .d(n2702), .o(delay_add_ln22_unr5_stage3_stallmux_q_1_), .ck(clk) );
ms00f80 l0510 ( .d(n2707), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_7_), .ck(clk) );
ms00f80 l0511 ( .d(n2712), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_15_), .ck(clk) );
ms00f80 l0512 ( .d(n2717), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_30_), .ck(clk) );
ms00f80 l0513 ( .d(n2722), .o(delay_add_ln22_unr23_stage9_stallmux_q_6_), .ck(clk) );
ms00f80 l0514 ( .d(n2727), .o(cos_out_15), .ck(clk) );
ms00f80 l0515 ( .d(n2731), .o(delay_xor_ln22_unr12_stage5_stallmux_q_17_), .ck(clk) );
ms00f80 l0516 ( .d(n2736), .o(delay_add_ln22_unr27_stage10_stallmux_q_12_), .ck(clk) );
ms00f80 l0517 ( .d(n2741), .o(delay_xor_ln21_unr15_stage6_stallmux_q_4_), .ck(clk) );
ms00f80 l0518 ( .d(n2746), .o(delay_xor_ln22_unr15_stage6_stallmux_q_6_), .ck(clk) );
ms00f80 l0519 ( .d(n2751), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_14_), .ck(clk) );
ms00f80 l0520 ( .d(n2756), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_20_), .ck(clk) );
ms00f80 l0521 ( .d(n2761), .o(delay_xor_ln21_unr3_stage2_stallmux_q_12_), .ck(clk) );
ms00f80 l0522 ( .d(n2766), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_24_), .ck(clk) );
ms00f80 l0523 ( .d(n2771), .o(delay_xor_ln21_unr28_stage10_stallmux_q_2_), .ck(clk) );
ms00f80 l0524 ( .d(n2776), .o(delay_xor_ln22_unr3_stage2_stallmux_q_23_), .ck(clk) );
ms00f80 l0525 ( .d(n2781), .o(delay_add_ln22_unr14_stage6_stallmux_q_25_), .ck(clk) );
ms00f80 l0526 ( .d(n2786), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_25_), .ck(clk) );
ms00f80 l0527 ( .d(n2791), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_22_), .ck(clk) );
ms00f80 l0528 ( .d(n2796), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_13_), .ck(clk) );
ms00f80 l0529 ( .d(n2801), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_22_), .ck(clk) );
ms00f80 l0530 ( .d(n2806), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_16_), .ck(clk) );
ms00f80 l0531 ( .d(n2811), .o(delay_xor_ln22_unr15_stage6_stallmux_q_5_), .ck(clk) );
ms00f80 l0532 ( .d(n2816), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_5_), .ck(clk) );
ms00f80 l0533 ( .d(n2821), .o(delay_xor_ln22_unr6_stage3_stallmux_q_8_), .ck(clk) );
ms00f80 l0534 ( .d(n2826), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_11_), .ck(clk) );
ms00f80 l0535 ( .d(n2831), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_20_), .ck(clk) );
ms00f80 l0536 ( .d(n2836), .o(delay_xor_ln21_unr21_stage8_stallmux_q_6_), .ck(clk) );
ms00f80 l0537 ( .d(n2841), .o(delay_add_ln22_unr27_stage10_stallmux_q_7_), .ck(clk) );
ms00f80 l0538 ( .d(n2846), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_29_), .ck(clk) );
ms00f80 l0539 ( .d(n2851), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_21_), .ck(clk) );
ms00f80 l0540 ( .d(n2856), .o(delay_xor_ln21_unr3_stage2_stallmux_q_24_), .ck(clk) );
ms00f80 l0541 ( .d(n2861), .o(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .ck(clk) );
ms00f80 l0542 ( .d(n2866), .o(delay_add_ln22_unr14_stage6_stallmux_q_27_), .ck(clk) );
ms00f80 l0543 ( .d(n2871), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_6_), .ck(clk) );
ms00f80 l0544 ( .d(n2876), .o(delay_xor_ln21_unr12_stage5_stallmux_q_17_), .ck(clk) );
ms00f80 l0545 ( .d(n2881), .o(delay_xor_ln21_unr6_stage3_stallmux_q_14_), .ck(clk) );
ms00f80 l0546 ( .d(n2886), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_2_), .ck(clk) );
ms00f80 l0547 ( .d(n2891), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_25_), .ck(clk) );
ms00f80 l0548 ( .d(n2896), .o(delay_xor_ln22_unr3_stage2_stallmux_q_18_), .ck(clk) );
ms00f80 l0549 ( .d(n2901), .o(delay_add_ln22_unr27_stage10_stallmux_q_1_), .ck(clk) );
ms00f80 l0550 ( .d(n2906), .o(delay_add_ln22_unr8_stage4_stallmux_q_19_), .ck(clk) );
ms00f80 l0551 ( .d(n2911), .o(delay_add_ln22_unr8_stage4_stallmux_q_4_), .ck(clk) );
ms00f80 l0552 ( .d(n2916), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_12_), .ck(clk) );
ms00f80 l0553 ( .d(n2921), .o(delay_add_ln22_unr14_stage6_stallmux_q_8_), .ck(clk) );
ms00f80 l0554 ( .d(n2926), .o(delay_xor_ln21_unr21_stage8_stallmux_q_10_), .ck(clk) );
ms00f80 l0555 ( .d(n2931), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_30_), .ck(clk) );
ms00f80 l0556 ( .d(n2936), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_1_), .ck(clk) );
ms00f80 l0557 ( .d(n2941), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_15_), .ck(clk) );
ms00f80 l0558 ( .d(n2946), .o(delay_xor_ln21_unr28_stage10_stallmux_q_1_), .ck(clk) );
ms00f80 l0559 ( .d(n2951), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_14_), .ck(clk) );
ms00f80 l0560 ( .d(n2956), .o(delay_xor_ln22_unr28_stage10_stallmux_q_3_), .ck(clk) );
ms00f80 l0561 ( .d(n2961), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_17_), .ck(clk) );
ms00f80 l0562 ( .d(n2966), .o(delay_xor_ln21_unr3_stage2_stallmux_q_18_), .ck(clk) );
ms00f80 l0563 ( .d(n2971), .o(delay_add_ln22_unr17_stage7_stallmux_q_5_), .ck(clk) );
ms00f80 l0564 ( .d(n2976), .o(delay_add_ln22_unr17_stage7_stallmux_q_16_), .ck(clk) );
ms00f80 l0565 ( .d(n2981), .o(delay_xor_ln22_unr9_stage4_stallmux_q_2_), .ck(clk) );
ms00f80 l0566 ( .d(n2986), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_31_), .ck(clk) );
ms00f80 l0567 ( .d(n2991), .o(delay_xor_ln21_unr3_stage2_stallmux_q_16_), .ck(clk) );
ms00f80 l0568 ( .d(n2996), .o(delay_add_ln22_unr8_stage4_stallmux_q_26_), .ck(clk) );
ms00f80 l0569 ( .d(n3001), .o(cos_out_11), .ck(clk) );
ms00f80 l0570 ( .d(n3005), .o(delay_xor_ln22_unr9_stage4_stallmux_q_11_), .ck(clk) );
ms00f80 l0571 ( .d(n3010), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_21_), .ck(clk) );
ms00f80 l0572 ( .d(n3015), .o(delay_xor_ln21_unr15_stage6_stallmux_q_9_), .ck(clk) );
ms00f80 l0573 ( .d(n3020), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_7_), .ck(clk) );
ms00f80 l0574 ( .d(n3025), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_2_), .ck(clk) );
ms00f80 l0575 ( .d(n3030), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_16_), .ck(clk) );
ms00f80 l0576 ( .d(n3035), .o(delay_xor_ln21_unr3_stage2_stallmux_q_19_), .ck(clk) );
ms00f80 l0577 ( .d(n3040), .o(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .ck(clk) );
ms00f80 l0578 ( .d(n3045), .o(n_45622), .ck(clk) );
ms00f80 l0579 ( .d(n3050), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_10_), .ck(clk) );
ms00f80 l0580 ( .d(n3055), .o(delay_sub_ln23_0_unr25_stage9_stallmux_q), .ck(clk) );
ms00f80 l0581 ( .d(n3060), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_6_), .ck(clk) );
ms00f80 l0582 ( .d(n3065), .o(delay_add_ln22_unr2_stage2_stallmux_q_3_), .ck(clk) );
ms00f80 l0583 ( .d(n3070), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_21_), .ck(clk) );
ms00f80 l0584 ( .d(n3075), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_1_), .ck(clk) );
ms00f80 l0585 ( .d(n3080), .o(delay_add_ln22_unr8_stage4_stallmux_q_0_), .ck(clk) );
ms00f80 l0586 ( .d(n3085), .o(delay_xor_ln21_unr18_stage7_stallmux_q_2_), .ck(clk) );
ms00f80 l0587 ( .d(n3090), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_4_), .ck(clk) );
ms00f80 l0588 ( .d(n3095), .o(delay_xor_ln21_unr21_stage8_stallmux_q_5_), .ck(clk) );
ms00f80 l0589 ( .d(n3100), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_8_), .ck(clk) );
ms00f80 l0590 ( .d(n3105), .o(delay_xor_ln21_unr9_stage4_stallmux_q_16_), .ck(clk) );
ms00f80 l0591 ( .d(n3110), .o(delay_xor_ln21_unr3_stage2_stallmux_q_26_), .ck(clk) );
ms00f80 l0592 ( .d(n3115), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_13_), .ck(clk) );
ms00f80 l0593 ( .d(n3120), .o(delay_add_ln22_unr5_stage3_stallmux_q_28_), .ck(clk) );
ms00f80 l0594 ( .d(n3125), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_20_), .ck(clk) );
ms00f80 l0595 ( .d(n3130), .o(delay_sub_ln22_unr24_stage9_stallmux_q_0_), .ck(clk) );
ms00f80 l0596 ( .d(n3135), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_5_), .ck(clk) );
ms00f80 l0597 ( .d(n3140), .o(delay_xor_ln21_unr28_stage10_stallmux_q_3_), .ck(clk) );
ms00f80 l0598 ( .d(n3145), .o(delay_xor_ln21_unr21_stage8_stallmux_q_1_), .ck(clk) );
ms00f80 l0599 ( .d(n3150), .o(delay_add_ln22_unr11_stage5_stallmux_q_18_), .ck(clk) );
ms00f80 l0600 ( .d(n3155), .o(delay_xor_ln22_unr6_stage3_stallmux_q_2_), .ck(clk) );
ms00f80 l0601 ( .d(n3160), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_14_), .ck(clk) );
ms00f80 l0602 ( .d(n3165), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_1_), .ck(clk) );
ms00f80 l0603 ( .d(n3170), .o(delay_add_ln22_unr23_stage9_stallmux_q_12_), .ck(clk) );
ms00f80 l0604 ( .d(n3175), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_28_), .ck(clk) );
ms00f80 l0605 ( .d(n3180), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_24_), .ck(clk) );
ms00f80 l0606 ( .d(n3185), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_4_), .ck(clk) );
ms00f80 l0607 ( .d(n3190), .o(sin_out_0), .ck(clk) );
ms00f80 l0608 ( .d(n3194), .o(delay_xor_ln22_unr6_stage3_stallmux_q_5_), .ck(clk) );
ms00f80 l0609 ( .d(n3199), .o(delay_add_ln22_unr8_stage4_stallmux_q_22_), .ck(clk) );
ms00f80 l0610 ( .d(n3204), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_4_), .ck(clk) );
ms00f80 l0611 ( .d(n3209), .o(delay_add_ln22_unr8_stage4_stallmux_q_29_), .ck(clk) );
ms00f80 l0612 ( .d(n3214), .o(delay_xor_ln22_unr15_stage6_stallmux_q_12_), .ck(clk) );
ms00f80 l0613 ( .d(n3219), .o(delay_xor_ln21_unr6_stage3_stallmux_q_24_), .ck(clk) );
ms00f80 l0614 ( .d(n3224), .o(cos_out_23), .ck(clk) );
ms00f80 l0615 ( .d(n3228), .o(delay_add_ln22_unr2_stage2_stallmux_q_28_), .ck(clk) );
ms00f80 l0616 ( .d(n3233), .o(delay_add_ln22_unr20_stage8_stallmux_q_21_), .ck(clk) );
ms00f80 l0617 ( .d(n3238), .o(delay_xor_ln22_unr12_stage5_stallmux_q_6_), .ck(clk) );
ms00f80 l0618 ( .d(n3243), .o(delay_add_ln22_unr23_stage9_stallmux_q_26_), .ck(clk) );
ms00f80 l0619 ( .d(n3248), .o(sin_out_27), .ck(clk) );
ms00f80 l0620 ( .d(n3252), .o(delay_xor_ln22_unr21_stage8_stallmux_q_9_), .ck(clk) );
ms00f80 l0621 ( .d(n3257), .o(delay_sub_ln21_unr24_stage9_stallmux_q_4_), .ck(clk) );
ms00f80 l0622 ( .d(n3262), .o(delay_add_ln22_unr27_stage10_stallmux_q_22_), .ck(clk) );
ms00f80 l0623 ( .d(n3267), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_2_), .ck(clk) );
ms00f80 l0624 ( .d(n3272), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_4_), .ck(clk) );
ms00f80 l0625 ( .d(n3277), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_8_), .ck(clk) );
ms00f80 l0626 ( .d(n3282), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_23_), .ck(clk) );
ms00f80 l0627 ( .d(n3287), .o(delay_add_ln22_unr2_stage2_stallmux_q_24_), .ck(clk) );
ms00f80 l0628 ( .d(n3292), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_9_), .ck(clk) );
ms00f80 l0629 ( .d(n3297), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_12_), .ck(clk) );
ms00f80 l0630 ( .d(n3302), .o(delay_xor_ln21_unr6_stage3_stallmux_q_13_), .ck(clk) );
ms00f80 l0631 ( .d(n3307), .o(delay_xor_ln21_unr6_stage3_stallmux_q_11_), .ck(clk) );
ms00f80 l0632 ( .d(n3312), .o(delay_sub_ln21_unr24_stage9_stallmux_q_7_), .ck(clk) );
ms00f80 l0633 ( .d(n3317), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_23_), .ck(clk) );
ms00f80 l0634 ( .d(n3322), .o(delay_xor_ln21_unr9_stage4_stallmux_q_18_), .ck(clk) );
ms00f80 l0635 ( .d(n3327), .o(delay_xor_ln22_unr15_stage6_stallmux_q_14_), .ck(clk) );
ms00f80 l0636 ( .d(n3332), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_28_), .ck(clk) );
ms00f80 l0637 ( .d(n3337), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_21_), .ck(clk) );
ms00f80 l0638 ( .d(n3342), .o(delay_add_ln22_unr14_stage6_stallmux_q_31_), .ck(clk) );
ms00f80 l0639 ( .d(n3347), .o(delay_xor_ln21_unr9_stage4_stallmux_q_0_), .ck(clk) );
ms00f80 l0640 ( .d(n3352), .o(delay_xor_ln22_unr21_stage8_stallmux_q_0_), .ck(clk) );
ms00f80 l0641 ( .d(n3357), .o(delay_add_ln22_unr23_stage9_stallmux_q_27_), .ck(clk) );
ms00f80 l0642 ( .d(n3362), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_0_), .ck(clk) );
ms00f80 l0643 ( .d(n3367), .o(delay_add_ln22_unr17_stage7_stallmux_q_22_), .ck(clk) );
ms00f80 l0644 ( .d(n3372), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_1_), .ck(clk) );
ms00f80 l0645 ( .d(n3377), .o(delay_add_ln22_unr8_stage4_stallmux_q_8_), .ck(clk) );
ms00f80 l0646 ( .d(n3382), .o(delay_add_ln22_unr27_stage10_stallmux_q_10_), .ck(clk) );
ms00f80 l0647 ( .d(n3387), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_17_), .ck(clk) );
ms00f80 l0648 ( .d(n3392), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_3_), .ck(clk) );
ms00f80 l0649 ( .d(n3397), .o(delay_xor_ln21_unr15_stage6_stallmux_q_0_), .ck(clk) );
ms00f80 l0650 ( .d(n3402), .o(delay_sub_ln22_unr24_stage9_stallmux_q_5_), .ck(clk) );
ms00f80 l0651 ( .d(n3407), .o(sin_out_29), .ck(clk) );
ms00f80 l0652 ( .d(n3411), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_24_), .ck(clk) );
ms00f80 l0653 ( .d(n3416), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_6_), .ck(clk) );
ms00f80 l0654 ( .d(n3421), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_4_), .ck(clk) );
ms00f80 l0655 ( .d(n3426), .o(delay_add_ln22_unr23_stage9_stallmux_q_24_), .ck(clk) );
ms00f80 l0656 ( .d(n3431), .o(delay_xor_ln21_unr3_stage2_stallmux_q_22_), .ck(clk) );
ms00f80 l0657 ( .d(n3436), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_3_), .ck(clk) );
ms00f80 l0658 ( .d(n3441), .o(delay_xor_ln22_unr21_stage8_stallmux_q_3_), .ck(clk) );
ms00f80 l0659 ( .d(n3446), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_25_), .ck(clk) );
ms00f80 l0660 ( .d(n3451), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_11_), .ck(clk) );
ms00f80 l0661 ( .d(n3456), .o(delay_add_ln22_unr2_stage2_stallmux_q_22_), .ck(clk) );
ms00f80 l0662 ( .d(n3461), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_0_), .ck(clk) );
ms00f80 l0663 ( .d(n3466), .o(delay_add_ln22_unr2_stage2_stallmux_q_21_), .ck(clk) );
ms00f80 l0664 ( .d(n3471), .o(delay_add_ln22_unr23_stage9_stallmux_q_7_), .ck(clk) );
ms00f80 l0665 ( .d(n3476), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_3_), .ck(clk) );
ms00f80 l0666 ( .d(n3481), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_22_), .ck(clk) );
ms00f80 l0667 ( .d(n3486), .o(delay_add_ln22_unr20_stage8_stallmux_q_23_), .ck(clk) );
ms00f80 l0668 ( .d(n3491), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_6_), .ck(clk) );
ms00f80 l0669 ( .d(n3496), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_7_), .ck(clk) );
ms00f80 l0670 ( .d(n3501), .o(delay_xor_ln21_unr6_stage3_stallmux_q_16_), .ck(clk) );
ms00f80 l0671 ( .d(n3506), .o(delay_xor_ln21_unr9_stage4_stallmux_q_1_), .ck(clk) );
ms00f80 l0672 ( .d(n3511), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_6_), .ck(clk) );
ms00f80 l0673 ( .d(n3516), .o(delay_xor_ln22_unr6_stage3_stallmux_q_17_), .ck(clk) );
ms00f80 l0674 ( .d(n3521), .o(delay_sub_ln23_0_unr27_stage10_stallmux_z), .ck(clk) );
ms00f80 l0675 ( .d(n3526), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_20_), .ck(clk) );
ms00f80 l0676 ( .d(n3531), .o(sin_out_14), .ck(clk) );
ms00f80 l0677 ( .d(n3535), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_25_), .ck(clk) );
ms00f80 l0678 ( .d(n3540), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_1_), .ck(clk) );
ms00f80 l0679 ( .d(n3545), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_16_), .ck(clk) );
ms00f80 l0680 ( .d(n3550), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_14_), .ck(clk) );
ms00f80 l0681 ( .d(n3555), .o(delay_xor_ln22_unr6_stage3_stallmux_q_15_), .ck(clk) );
ms00f80 l0682 ( .d(n3560), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_22_), .ck(clk) );
ms00f80 l0683 ( .d(n3565), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_10_), .ck(clk) );
ms00f80 l0684 ( .d(n3570), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_28_), .ck(clk) );
ms00f80 l0685 ( .d(n3575), .o(n_45202), .ck(clk) );
ms00f80 l0686 ( .d(n3580), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_15_), .ck(clk) );
ms00f80 l0687 ( .d(n3585), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_22_), .ck(clk) );
ms00f80 l0688 ( .d(n3590), .o(delay_xor_ln22_unr12_stage5_stallmux_q_4_), .ck(clk) );
ms00f80 l0689 ( .d(n3595), .o(delay_add_ln22_unr14_stage6_stallmux_q_2_), .ck(clk) );
ms00f80 l0690 ( .d(n3600), .o(cos_out_21), .ck(clk) );
ms00f80 l0691 ( .d(n3604), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_14_), .ck(clk) );
ms00f80 l0692 ( .d(n3609), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_30_), .ck(clk) );
ms00f80 l0693 ( .d(n3614), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_1_), .ck(clk) );
ms00f80 l0694 ( .d(n3619), .o(sin_out_19), .ck(clk) );
ms00f80 l0695 ( .d(n3623), .o(delay_add_ln22_unr2_stage2_stallmux_q_1_), .ck(clk) );
ms00f80 l0696 ( .d(n3628), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_27_), .ck(clk) );
ms00f80 l0697 ( .d(n3633), .o(n_44722), .ck(clk) );
ms00f80 l0698 ( .d(n3638), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_23_), .ck(clk) );
ms00f80 l0699 ( .d(n3643), .o(delay_add_ln22_unr27_stage10_stallmux_q_6_), .ck(clk) );
ms00f80 l0700 ( .d(n3648), .o(delay_add_ln22_unr11_stage5_stallmux_q_10_), .ck(clk) );
ms00f80 l0701 ( .d(n3653), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_12_), .ck(clk) );
ms00f80 l0702 ( .d(n3658), .o(delay_add_ln22_unr5_stage3_stallmux_q_31_), .ck(clk) );
ms00f80 l0703 ( .d(n3663), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_27_), .ck(clk) );
ms00f80 l0704 ( .d(n3668), .o(delay_add_ln22_unr27_stage10_stallmux_q_29_), .ck(clk) );
ms00f80 l0705 ( .d(n3673), .o(delay_add_ln22_unr8_stage4_stallmux_q_25_), .ck(clk) );
ms00f80 l0706 ( .d(n3678), .o(delay_xor_ln22_unr6_stage3_stallmux_q_12_), .ck(clk) );
ms00f80 l0707 ( .d(n3683), .o(delay_xor_ln21_unr12_stage5_stallmux_q_10_), .ck(clk) );
ms00f80 l0708 ( .d(n3688), .o(delay_add_ln22_unr27_stage10_stallmux_q_16_), .ck(clk) );
ms00f80 l0709 ( .d(n3693), .o(delay_xor_ln21_unr12_stage5_stallmux_q_2_), .ck(clk) );
ms00f80 l0710 ( .d(n3698), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_13_), .ck(clk) );
ms00f80 l0711 ( .d(n3703), .o(cos_out_13), .ck(clk) );
ms00f80 l0712 ( .d(n3707), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_28_), .ck(clk) );
ms00f80 l0713 ( .d(n3712), .o(delay_xor_ln21_unr9_stage4_stallmux_q_17_), .ck(clk) );
ms00f80 l0714 ( .d(n3717), .o(delay_add_ln22_unr11_stage5_stallmux_q_3_), .ck(clk) );
ms00f80 l0715 ( .d(n3722), .o(delay_add_ln22_unr20_stage8_stallmux_q_17_), .ck(clk) );
ms00f80 l0716 ( .d(n3727), .o(delay_xor_ln22_unr9_stage4_stallmux_q_16_), .ck(clk) );
ms00f80 l0717 ( .d(n3732), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_14_), .ck(clk) );
ms00f80 l0718 ( .d(n3737), .o(delay_add_ln22_unr17_stage7_stallmux_q_9_), .ck(clk) );
ms00f80 l0719 ( .d(n3742), .o(delay_add_ln22_unr23_stage9_stallmux_q_13_), .ck(clk) );
ms00f80 l0720 ( .d(n3747), .o(delay_add_ln22_unr5_stage3_stallmux_q_21_), .ck(clk) );
ms00f80 l0721 ( .d(n3752), .o(delay_add_ln22_unr17_stage7_stallmux_q_6_), .ck(clk) );
ms00f80 l0722 ( .d(n3757), .o(n_44422), .ck(clk) );
ms00f80 l0723 ( .d(n3762), .o(delay_add_ln22_unr14_stage6_stallmux_q_17_), .ck(clk) );
ms00f80 l0724 ( .d(n3767), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_8_), .ck(clk) );
ms00f80 l0725 ( .d(n3772), .o(delay_xor_ln22_unr28_stage10_stallmux_q_2_), .ck(clk) );
ms00f80 l0726 ( .d(n3777), .o(delay_xor_ln21_unr21_stage8_stallmux_q_4_), .ck(clk) );
ms00f80 l0727 ( .d(n3782), .o(delay_add_ln22_unr11_stage5_stallmux_q_28_), .ck(clk) );
ms00f80 l0728 ( .d(n3787), .o(delay_add_ln22_unr8_stage4_stallmux_q_1_), .ck(clk) );
ms00f80 l0729 ( .d(n3792), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_6_), .ck(clk) );
ms00f80 l0730 ( .d(n3797), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_1_), .ck(clk) );
ms00f80 l0731 ( .d(n3802), .o(cos_out_5), .ck(clk) );
ms00f80 l0732 ( .d(n3806), .o(delay_xor_ln21_unr12_stage5_stallmux_q_8_), .ck(clk) );
ms00f80 l0733 ( .d(n3811), .o(delay_sub_ln21_unr24_stage9_stallmux_q_1_), .ck(clk) );
ms00f80 l0734 ( .d(n3816), .o(delay_xor_ln22_unr12_stage5_stallmux_q_5_), .ck(clk) );
ms00f80 l0735 ( .d(n3821), .o(delay_add_ln22_unr23_stage9_stallmux_q_22_), .ck(clk) );
ms00f80 l0736 ( .d(n3826), .o(delay_add_ln22_unr5_stage3_stallmux_q_26_), .ck(clk) );
ms00f80 l0737 ( .d(n3831), .o(delay_add_ln22_unr17_stage7_stallmux_q_17_), .ck(clk) );
ms00f80 l0738 ( .d(n3836), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_17_), .ck(clk) );
ms00f80 l0739 ( .d(n3841), .o(delay_add_ln22_unr20_stage8_stallmux_q_22_), .ck(clk) );
ms00f80 l0740 ( .d(n3846), .o(cos_out_0), .ck(clk) );
ms00f80 l0741 ( .d(n3850), .o(delay_add_ln22_unr20_stage8_stallmux_q_8_), .ck(clk) );
ms00f80 l0742 ( .d(n3855), .o(delay_add_ln22_unr2_stage2_stallmux_q_29_), .ck(clk) );
ms00f80 l0743 ( .d(n3860), .o(delay_xor_ln22_unr9_stage4_stallmux_q_7_), .ck(clk) );
ms00f80 l0744 ( .d(n3865), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_13_), .ck(clk) );
ms00f80 l0745 ( .d(n3870), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_20_), .ck(clk) );
ms00f80 l0746 ( .d(n3875), .o(delay_xor_ln22_unr18_stage7_stallmux_q_9_), .ck(clk) );
ms00f80 l0747 ( .d(n3880), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_3_), .ck(clk) );
ms00f80 l0748 ( .d(n3885), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_13_), .ck(clk) );
ms00f80 l0749 ( .d(n3890), .o(delay_xor_ln22_unr9_stage4_stallmux_q_20_), .ck(clk) );
ms00f80 l0750 ( .d(n3895), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_13_), .ck(clk) );
ms00f80 l0751 ( .d(n3900), .o(delay_add_ln22_unr8_stage4_stallmux_q_31_), .ck(clk) );
ms00f80 l0752 ( .d(n3905), .o(delay_xor_ln21_unr6_stage3_stallmux_q_23_), .ck(clk) );
ms00f80 l0753 ( .d(n3910), .o(delay_add_ln22_unr2_stage2_stallmux_q_9_), .ck(clk) );
ms00f80 l0754 ( .d(n3915), .o(delay_xor_ln22_unr9_stage4_stallmux_q_17_), .ck(clk) );
ms00f80 l0755 ( .d(n3920), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_4_), .ck(clk) );
ms00f80 l0756 ( .d(n3925), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_9_), .ck(clk) );
ms00f80 l0757 ( .d(n3930), .o(delay_xor_ln21_unr6_stage3_stallmux_q_9_), .ck(clk) );
ms00f80 l0758 ( .d(n3935), .o(delay_add_ln22_unr2_stage2_stallmux_q_30_), .ck(clk) );
ms00f80 l0759 ( .d(n3940), .o(delay_xor_ln21_unr6_stage3_stallmux_q_10_), .ck(clk) );
ms00f80 l0760 ( .d(n3945), .o(delay_xor_ln21_unr21_stage8_stallmux_q_3_), .ck(clk) );
ms00f80 l0761 ( .d(n3950), .o(delay_xor_ln22_unr3_stage2_stallmux_q_5_), .ck(clk) );
ms00f80 l0762 ( .d(n3955), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_11_), .ck(clk) );
ms00f80 l0763 ( .d(n3960), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_13_), .ck(clk) );
ms00f80 l0764 ( .d(n3965), .o(delay_add_ln22_unr20_stage8_stallmux_q_20_), .ck(clk) );
ms00f80 l0765 ( .d(n3970), .o(delay_add_ln22_unr11_stage5_stallmux_q_2_), .ck(clk) );
ms00f80 l0766 ( .d(n3975), .o(delay_add_ln22_unr17_stage7_stallmux_q_30_), .ck(clk) );
ms00f80 l0767 ( .d(n3980), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_6_), .ck(clk) );
ms00f80 l0768 ( .d(n3985), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_6_), .ck(clk) );
ms00f80 l0769 ( .d(n3990), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_28_), .ck(clk) );
ms00f80 l0770 ( .d(n3994), .o(delay_xor_ln22_unr3_stage2_stallmux_q_8_), .ck(clk) );
ms00f80 l0771 ( .d(n3999), .o(delay_add_ln22_unr20_stage8_stallmux_q_0_), .ck(clk) );
ms00f80 l0772 ( .d(n4004), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_18_), .ck(clk) );
ms00f80 l0773 ( .d(n4009), .o(delay_sub_ln22_unr24_stage9_stallmux_q_3_), .ck(clk) );
ms00f80 l0774 ( .d(n4014), .o(delay_add_ln22_unr11_stage5_stallmux_q_31_), .ck(clk) );
ms00f80 l0775 ( .d(n4019), .o(delay_xor_ln22_unr18_stage7_stallmux_q_1_), .ck(clk) );
ms00f80 l0776 ( .d(n4024), .o(cos_out_10), .ck(clk) );
ms00f80 l0777 ( .d(n4028), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_17_), .ck(clk) );
ms00f80 l0778 ( .d(n4033), .o(delay_xor_ln21_unr12_stage5_stallmux_q_13_), .ck(clk) );
ms00f80 l0779 ( .d(n4038), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_14_), .ck(clk) );
ms00f80 l0780 ( .d(n4043), .o(n_25834), .ck(clk) );
ms00f80 l0781 ( .d(n4048), .o(mux_while_ln12_psv_q_1_), .ck(clk) );
ms00f80 l0782 ( .d(n4053), .o(delay_add_ln22_unr2_stage2_stallmux_q_11_), .ck(clk) );
ms00f80 l0783 ( .d(n4058), .o(delay_xor_ln22_unr6_stage3_stallmux_q_14_), .ck(clk) );
ms00f80 l0784 ( .d(n4063), .o(delay_add_ln22_unr14_stage6_stallmux_q_12_), .ck(clk) );
ms00f80 l0785 ( .d(n4068), .o(delay_add_ln22_unr17_stage7_stallmux_q_15_), .ck(clk) );
ms00f80 l0786 ( .d(n4073), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_11_), .ck(clk) );
ms00f80 l0787 ( .d(n4078), .o(delay_xor_ln22_unr6_stage3_stallmux_q_13_), .ck(clk) );
ms00f80 l0788 ( .d(n4083), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_4_), .ck(clk) );
ms00f80 l0789 ( .d(n4088), .o(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .ck(clk) );
ms00f80 l0790 ( .d(n4093), .o(delay_xor_ln22_unr15_stage6_stallmux_q_0_), .ck(clk) );
ms00f80 l0791 ( .d(n4098), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_23_), .ck(clk) );
ms00f80 l0792 ( .d(n4103), .o(sin_out_13), .ck(clk) );
ms00f80 l0793 ( .d(n4107), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_7_), .ck(clk) );
ms00f80 l0794 ( .d(n4112), .o(cos_out_3), .ck(clk) );
ms00f80 l0795 ( .d(n4116), .o(delay_xor_ln23_unr6_stage3_stallmux_q), .ck(clk) );
ms00f80 l0796 ( .d(n4121), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_19_), .ck(clk) );
ms00f80 l0797 ( .d(n4126), .o(delay_add_ln22_unr8_stage4_stallmux_q_28_), .ck(clk) );
ms00f80 l0798 ( .d(n4131), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_19_), .ck(clk) );
ms00f80 l0799 ( .d(n4136), .o(delay_xor_ln21_unr9_stage4_stallmux_q_4_), .ck(clk) );
ms00f80 l0800 ( .d(n4141), .o(delay_add_ln22_unr17_stage7_stallmux_q_19_), .ck(clk) );
ms00f80 l0801 ( .d(n4146), .o(delay_xor_ln21_unr3_stage2_stallmux_q_2_), .ck(clk) );
ms00f80 l0802 ( .d(n4151), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_8_), .ck(clk) );
ms00f80 l0803 ( .d(n4156), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_12_), .ck(clk) );
ms00f80 l0804 ( .d(n4161), .o(delay_xor_ln21_unr6_stage3_stallmux_q_19_), .ck(clk) );
ms00f80 l0805 ( .d(n4166), .o(delay_xor_ln21_unr3_stage2_stallmux_q_6_), .ck(clk) );
ms00f80 l0806 ( .d(n4171), .o(delay_add_ln22_unr5_stage3_stallmux_q_18_), .ck(clk) );
ms00f80 l0807 ( .d(n4176), .o(delay_sub_ln23_0_unr23_stage8_stallmux_q), .ck(clk) );
ms00f80 l0808 ( .d(n4181), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_6_), .ck(clk) );
ms00f80 l0809 ( .d(n4186), .o(delay_add_ln22_unr11_stage5_stallmux_q_29_), .ck(clk) );
ms00f80 l0810 ( .d(n4191), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_27_), .ck(clk) );
ms00f80 l0811 ( .d(n4196), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_17_), .ck(clk) );
ms00f80 l0812 ( .d(n4201), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_13_), .ck(clk) );
ms00f80 l0813 ( .d(n4206), .o(delay_xor_ln22_unr21_stage8_stallmux_q_7_), .ck(clk) );
ms00f80 l0814 ( .d(n4211), .o(mux_while_ln12_psv_q_6_), .ck(clk) );
ms00f80 l0815 ( .d(n4216), .o(delay_xor_ln22_unr3_stage2_stallmux_q_4_), .ck(clk) );
ms00f80 l0816 ( .d(n4221), .o(delay_xor_ln21_unr12_stage5_stallmux_q_6_), .ck(clk) );
ms00f80 l0817 ( .d(n4226), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_7_), .ck(clk) );
ms00f80 l0818 ( .d(n4231), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_29_), .ck(clk) );
ms00f80 l0819 ( .d(n4236), .o(delay_add_ln22_unr11_stage5_stallmux_q_11_), .ck(clk) );
ms00f80 l0820 ( .d(n4241), .o(delay_add_ln22_unr8_stage4_stallmux_q_11_), .ck(clk) );
ms00f80 l0821 ( .d(n4246), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_6_), .ck(clk) );
ms00f80 l0822 ( .d(n4251), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_10_), .ck(clk) );
ms00f80 l0823 ( .d(n4256), .o(delay_add_ln22_unr5_stage3_stallmux_q_6_), .ck(clk) );
ms00f80 l0824 ( .d(n4261), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_31_), .ck(clk) );
ms00f80 l0825 ( .d(n4266), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_23_), .ck(clk) );
ms00f80 l0826 ( .d(n4271), .o(sin_out_20), .ck(clk) );
ms00f80 l0827 ( .d(n4275), .o(delay_add_ln22_unr17_stage7_stallmux_q_18_), .ck(clk) );
ms00f80 l0828 ( .d(n4280), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_3_), .ck(clk) );
ms00f80 l0829 ( .d(n4285), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_18_), .ck(clk) );
ms00f80 l0830 ( .d(n4290), .o(delay_xor_ln22_unr3_stage2_stallmux_q_12_), .ck(clk) );
ms00f80 l0831 ( .d(n4295), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_3_), .ck(clk) );
ms00f80 l0832 ( .d(n4300), .o(delay_xor_ln22_unr6_stage3_stallmux_q_23_), .ck(clk) );
ms00f80 l0833 ( .d(n4305), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_29_), .ck(clk) );
ms00f80 l0834 ( .d(n4310), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_11_), .ck(clk) );
ms00f80 l0835 ( .d(n4315), .o(delay_add_ln22_unr14_stage6_stallmux_q_23_), .ck(clk) );
ms00f80 l0836 ( .d(n4320), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_6_), .ck(clk) );
ms00f80 l0837 ( .d(n4325), .o(delay_add_ln22_unr8_stage4_stallmux_q_27_), .ck(clk) );
ms00f80 l0838 ( .d(n4330), .o(cos_out_28), .ck(clk) );
ms00f80 l0839 ( .d(n4334), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_25_), .ck(clk) );
ms00f80 l0840 ( .d(n4339), .o(delay_xor_ln22_unr9_stage4_stallmux_q_12_), .ck(clk) );
ms00f80 l0841 ( .d(n4344), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_30_), .ck(clk) );
ms00f80 l0842 ( .d(n4349), .o(delay_add_ln22_unr8_stage4_stallmux_q_10_), .ck(clk) );
ms00f80 l0843 ( .d(n4354), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_10_), .ck(clk) );
ms00f80 l0844 ( .d(n4359), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_1_), .ck(clk) );
ms00f80 l0845 ( .d(n4364), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_30_), .ck(clk) );
ms00f80 l0846 ( .d(n4369), .o(delay_add_ln22_unr17_stage7_stallmux_q_11_), .ck(clk) );
ms00f80 l0847 ( .d(n4374), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_31_), .ck(clk) );
ms00f80 l0848 ( .d(n4379), .o(delay_add_ln22_unr5_stage3_stallmux_q_30_), .ck(clk) );
ms00f80 l0849 ( .d(n4384), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_17_), .ck(clk) );
ms00f80 l0850 ( .d(n4389), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_21_), .ck(clk) );
ms00f80 l0851 ( .d(n4394), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_1_), .ck(clk) );
ms00f80 l0852 ( .d(n4399), .o(delay_add_ln22_unr20_stage8_stallmux_q_28_), .ck(clk) );
ms00f80 l0853 ( .d(n4404), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_15_), .ck(clk) );
ms00f80 l0854 ( .d(n4409), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_5_), .ck(clk) );
ms00f80 l0855 ( .d(n4414), .o(delay_xor_ln22_unr6_stage3_stallmux_q_11_), .ck(clk) );
ms00f80 l0856 ( .d(n4419), .o(delay_add_ln22_unr20_stage8_stallmux_q_2_), .ck(clk) );
ms00f80 l0857 ( .d(n4424), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_26_), .ck(clk) );
ms00f80 l0858 ( .d(n4429), .o(delay_add_ln22_unr27_stage10_stallmux_q_15_), .ck(clk) );
ms00f80 l0859 ( .d(n4434), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_11_), .ck(clk) );
ms00f80 l0860 ( .d(n4439), .o(delay_add_ln22_unr11_stage5_stallmux_q_5_), .ck(clk) );
ms00f80 l0861 ( .d(n4443), .o(delay_sub_ln23_0_unr26_stage9_stallmux_q_0_), .ck(clk) );
ms00f80 l0862 ( .d(n4448), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_0_), .ck(clk) );
ms00f80 l0863 ( .d(n4453), .o(delay_xor_ln22_unr9_stage4_stallmux_q_21_), .ck(clk) );
ms00f80 l0864 ( .d(n4458), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_23_), .ck(clk) );
ms00f80 l0865 ( .d(n4463), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_12_), .ck(clk) );
ms00f80 l0866 ( .d(n4468), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_27_), .ck(clk) );
ms00f80 l0867 ( .d(n4473), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_10_), .ck(clk) );
ms00f80 l0868 ( .d(n4478), .o(n_46254), .ck(clk) );
ms00f80 l0869 ( .d(n4483), .o(delay_add_ln22_unr23_stage9_stallmux_q_9_), .ck(clk) );
ms00f80 l0870 ( .d(n4488), .o(delay_add_ln22_unr8_stage4_stallmux_q_16_), .ck(clk) );
ms00f80 l0871 ( .d(n4493), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_17_), .ck(clk) );
ms00f80 l0872 ( .d(n4498), .o(cordic_combinational_sub_ln23_0_unr12_z_0_), .ck(clk) );
ms00f80 l0873 ( .d(n4503), .o(delay_xor_ln22_unr12_stage5_stallmux_q_11_), .ck(clk) );
ms00f80 l0874 ( .d(n4508), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_26_), .ck(clk) );
ms00f80 l0875 ( .d(n4513), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_6_), .ck(clk) );
ms00f80 l0876 ( .d(n4518), .o(delay_xor_ln22_unr3_stage2_stallmux_q_2_), .ck(clk) );
ms00f80 l0877 ( .d(n4523), .o(delay_add_ln22_unr14_stage6_stallmux_q_7_), .ck(clk) );
ms00f80 l0878 ( .d(n4528), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_9_), .ck(clk) );
ms00f80 l0879 ( .d(n4533), .o(delay_xor_ln21_unr6_stage3_stallmux_q_5_), .ck(clk) );
ms00f80 l0880 ( .d(n4538), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_17_), .ck(clk) );
ms00f80 l0881 ( .d(n4543), .o(delay_xor_ln22_unr18_stage7_stallmux_q_2_), .ck(clk) );
ms00f80 l0882 ( .d(n4548), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_13_), .ck(clk) );
ms00f80 l0883 ( .d(n4553), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_30_), .ck(clk) );
ms00f80 l0884 ( .d(n4558), .o(delay_add_ln22_unr11_stage5_stallmux_q_20_), .ck(clk) );
ms00f80 l0885 ( .d(n4563), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_8_), .ck(clk) );
ms00f80 l0886 ( .d(n4568), .o(delay_add_ln22_unr5_stage3_stallmux_q_10_), .ck(clk) );
ms00f80 l0887 ( .d(n4573), .o(delay_add_ln22_unr8_stage4_stallmux_q_9_), .ck(clk) );
ms00f80 l0888 ( .d(n4578), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_5_), .ck(clk) );
ms00f80 l0889 ( .d(n4583), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_23_), .ck(clk) );
ms00f80 l0890 ( .d(n4588), .o(delay_xor_ln22_unr3_stage2_stallmux_q_16_), .ck(clk) );
ms00f80 l0891 ( .d(n4593), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_2_), .ck(clk) );
ms00f80 l0892 ( .d(n4598), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_27_), .ck(clk) );
ms00f80 l0893 ( .d(n4603), .o(delay_add_ln22_unr2_stage2_stallmux_q_23_), .ck(clk) );
ms00f80 l0894 ( .d(n4608), .o(delay_add_ln22_unr5_stage3_stallmux_q_9_), .ck(clk) );
ms00f80 l0895 ( .d(n4613), .o(delay_add_ln22_unr5_stage3_stallmux_q_22_), .ck(clk) );
ms00f80 l0896 ( .d(n4618), .o(delay_xor_ln21_unr12_stage5_stallmux_q_19_), .ck(clk) );
ms00f80 l0897 ( .d(n4623), .o(delay_add_ln22_unr27_stage10_stallmux_q_23_), .ck(clk) );
ms00f80 l0898 ( .d(n4628), .o(delay_add_ln22_unr17_stage7_stallmux_q_31_), .ck(clk) );
ms00f80 l0899 ( .d(n4633), .o(delay_add_ln22_unr27_stage10_stallmux_q_17_), .ck(clk) );
ms00f80 l0900 ( .d(n4638), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_5_), .ck(clk) );
ms00f80 l0901 ( .d(n4643), .o(delay_add_ln22_unr14_stage6_stallmux_q_28_), .ck(clk) );
ms00f80 l0902 ( .d(n4648), .o(sin_out_8), .ck(clk) );
ms00f80 l0903 ( .d(n4652), .o(delay_add_ln22_unr14_stage6_stallmux_q_0_), .ck(clk) );
ms00f80 l0904 ( .d(n4657), .o(n_44721), .ck(clk) );
ms00f80 l0905 ( .d(n4662), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_15_), .ck(clk) );
ms00f80 l0906 ( .d(n4667), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_25_), .ck(clk) );
ms00f80 l0907 ( .d(n4672), .o(delay_xor_ln22_unr3_stage2_stallmux_q_25_), .ck(clk) );
ms00f80 l0908 ( .d(n4677), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_4_), .ck(clk) );
ms00f80 l0909 ( .d(n4682), .o(delay_xor_ln22_unr6_stage3_stallmux_q_6_), .ck(clk) );
ms00f80 l0910 ( .d(n4687), .o(delay_xor_ln21_unr6_stage3_stallmux_q_1_), .ck(clk) );
ms00f80 l0911 ( .d(n4692), .o(delay_xor_ln22_unr21_stage8_stallmux_q_4_), .ck(clk) );
ms00f80 l0912 ( .d(n4697), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_9_), .ck(clk) );
ms00f80 l0913 ( .d(n4702), .o(delay_add_ln22_unr20_stage8_stallmux_q_16_), .ck(clk) );
ms00f80 l0914 ( .d(n4707), .o(delay_add_ln22_unr23_stage9_stallmux_q_10_), .ck(clk) );
ms00f80 l0915 ( .d(n4712), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_8_), .ck(clk) );
ms00f80 l0916 ( .d(n4717), .o(delay_add_ln22_unr17_stage7_stallmux_q_29_), .ck(clk) );
ms00f80 l0917 ( .d(n4722), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_20_), .ck(clk) );
ms00f80 l0918 ( .d(n4727), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_11_), .ck(clk) );
ms00f80 l0919 ( .d(n4732), .o(cos_out_19), .ck(clk) );
ms00f80 l0920 ( .d(n4736), .o(delay_add_ln22_unr8_stage4_stallmux_q_15_), .ck(clk) );
ms00f80 l0921 ( .d(n4741), .o(delay_xor_ln22_unr9_stage4_stallmux_q_9_), .ck(clk) );
ms00f80 l0922 ( .d(n4746), .o(delay_add_ln22_unr23_stage9_stallmux_q_3_), .ck(clk) );
ms00f80 l0923 ( .d(n4751), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_1_), .ck(clk) );
ms00f80 l0924 ( .d(n4756), .o(delay_add_ln22_unr27_stage10_stallmux_q_24_), .ck(clk) );
ms00f80 l0925 ( .d(n4761), .o(delay_add_ln22_unr2_stage2_stallmux_q_15_), .ck(clk) );
ms00f80 l0926 ( .d(n4766), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_14_), .ck(clk) );
ms00f80 l0927 ( .d(n4771), .o(delay_xor_ln22_unr18_stage7_stallmux_q_10_), .ck(clk) );
ms00f80 l0928 ( .d(n4776), .o(mux_while_ln12_psv_q_3_), .ck(clk) );
ms00f80 l0929 ( .d(n4781), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_31_), .ck(clk) );
ms00f80 l0930 ( .d(n4786), .o(delay_add_ln22_unr11_stage5_stallmux_q_23_), .ck(clk) );
ms00f80 l0931 ( .d(n4791), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_3_), .ck(clk) );
ms00f80 l0932 ( .d(n4796), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_30_), .ck(clk) );
ms00f80 l0933 ( .d(n4801), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_19_), .ck(clk) );
ms00f80 l0934 ( .d(n4806), .o(sin_out_30), .ck(clk) );
ms00f80 l0935 ( .d(n4810), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_1_), .ck(clk) );
ms00f80 l0936 ( .d(n4815), .o(delay_add_ln22_unr20_stage8_stallmux_q_3_), .ck(clk) );
ms00f80 l0937 ( .d(n4820), .o(delay_xor_ln22_unr9_stage4_stallmux_q_5_), .ck(clk) );
ms00f80 l0938 ( .d(n4825), .o(sin_out_24), .ck(clk) );
ms00f80 l0939 ( .d(n4829), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_1_), .ck(clk) );
ms00f80 l0940 ( .d(n4834), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_11_), .ck(clk) );
ms00f80 l0941 ( .d(n4839), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_20_), .ck(clk) );
ms00f80 l0942 ( .d(n4843), .o(state_cordic_1_), .ck(clk) );
ms00f80 l0943 ( .d(n4848), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_24_), .ck(clk) );
ms00f80 l0944 ( .d(n4853), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_0_), .ck(clk) );
ms00f80 l0945 ( .d(n4858), .o(delay_xor_ln21_unr3_stage2_stallmux_q_8_), .ck(clk) );
ms00f80 l0946 ( .d(n4863), .o(delay_xor_ln21_unr28_stage10_stallmux_q_0_), .ck(clk) );
ms00f80 l0947 ( .d(n4868), .o(delay_xor_ln21_unr12_stage5_stallmux_q_5_), .ck(clk) );
ms00f80 l0948 ( .d(n4873), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_25_), .ck(clk) );
ms00f80 l0949 ( .d(n4878), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_31_), .ck(clk) );
ms00f80 l0950 ( .d(n4883), .o(delay_add_ln22_unr23_stage9_stallmux_q_25_), .ck(clk) );
ms00f80 l0951 ( .d(n4888), .o(delay_xor_ln21_unr15_stage6_stallmux_q_16_), .ck(clk) );
ms00f80 l0952 ( .d(n4893), .o(sin_out_7), .ck(clk) );
ms00f80 l0953 ( .d(n4897), .o(delay_add_ln22_unr20_stage8_stallmux_q_31_), .ck(clk) );
ms00f80 l0954 ( .d(n4902), .o(delay_xor_ln21_unr6_stage3_stallmux_q_12_), .ck(clk) );
ms00f80 l0955 ( .d(n4907), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_18_), .ck(clk) );
ms00f80 l0956 ( .d(n4912), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_15_), .ck(clk) );
ms00f80 l0957 ( .d(n4917), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_22_), .ck(clk) );
ms00f80 l0958 ( .d(n4922), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_23_), .ck(clk) );
ms00f80 l0959 ( .d(n4927), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_18_), .ck(clk) );
ms00f80 l0960 ( .d(n4932), .o(delay_sub_ln23_0_unr1_stage2_stallmux_q_0_), .ck(clk) );
ms00f80 l0961 ( .d(n4937), .o(delay_xor_ln22_unr6_stage3_stallmux_q_7_), .ck(clk) );
ms00f80 l0962 ( .d(n4942), .o(delay_xor_ln22_unr6_stage3_stallmux_q_10_), .ck(clk) );
ms00f80 l0963 ( .d(n4947), .o(delay_xor_ln22_unr21_stage8_stallmux_q_8_), .ck(clk) );
ms00f80 l0964 ( .d(n4952), .o(delay_sub_ln23_unr25_stage8_stallmux_q_1_), .ck(clk) );
ms00f80 l0965 ( .d(n4957), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_1_), .ck(clk) );
ms00f80 l0966 ( .d(n4962), .o(n_45204), .ck(clk) );
ms00f80 l0967 ( .d(n4967), .o(delay_xor_ln22_unr3_stage2_stallmux_q_26_), .ck(clk) );
ms00f80 l0968 ( .d(n4972), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_21_), .ck(clk) );
ms00f80 l0969 ( .d(n4977), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_10_), .ck(clk) );
ms00f80 l0970 ( .d(n4982), .o(delay_sub_ln22_unr24_stage9_stallmux_q_4_), .ck(clk) );
ms00f80 l0971 ( .d(n4987), .o(delay_add_ln22_unr11_stage5_stallmux_q_8_), .ck(clk) );
ms00f80 l0972 ( .d(n4992), .o(delay_add_ln22_unr2_stage2_stallmux_q_14_), .ck(clk) );
ms00f80 l0973 ( .d(n4997), .o(cos_out_29), .ck(clk) );
ms00f80 l0974 ( .d(n5001), .o(n_27014), .ck(clk) );
ms00f80 l0975 ( .d(n5006), .o(delay_xor_ln21_unr9_stage4_stallmux_q_12_), .ck(clk) );
ms00f80 l0976 ( .d(n5011), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_24_), .ck(clk) );
ms00f80 l0977 ( .d(n5016), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_29_), .ck(clk) );
ms00f80 l0978 ( .d(n5021), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_18_), .ck(clk) );
ms00f80 l0979 ( .d(n5026), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_0_), .ck(clk) );
ms00f80 l0980 ( .d(n5031), .o(delay_add_ln22_unr14_stage6_stallmux_q_22_), .ck(clk) );
ms00f80 l0981 ( .d(n5036), .o(delay_add_ln22_unr5_stage3_stallmux_q_14_), .ck(clk) );
ms00f80 l0982 ( .d(n5041), .o(delay_add_ln22_unr8_stage4_stallmux_q_17_), .ck(clk) );
ms00f80 l0983 ( .d(n5046), .o(mux_while_ln12_psv_q_2_), .ck(clk) );
ms00f80 l0984 ( .d(n5051), .o(delay_add_ln22_unr2_stage2_stallmux_q_7_), .ck(clk) );
ms00f80 l0985 ( .d(n5056), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_12_), .ck(clk) );
ms00f80 l0986 ( .d(n5061), .o(delay_xor_ln22_unr9_stage4_stallmux_q_4_), .ck(clk) );
ms00f80 l0987 ( .d(n5066), .o(delay_add_ln22_unr14_stage6_stallmux_q_11_), .ck(clk) );
ms00f80 l0988 ( .d(n5070), .o(n_44610), .ck(clk) );
ms00f80 l0989 ( .d(n5075), .o(delay_add_ln22_unr5_stage3_stallmux_q_4_), .ck(clk) );
ms00f80 l0990 ( .d(n5080), .o(delay_add_ln22_unr5_stage3_stallmux_q_16_), .ck(clk) );
ms00f80 l0991 ( .d(n5085), .o(delay_xor_ln22_unr15_stage6_stallmux_q_4_), .ck(clk) );
ms00f80 l0992 ( .d(n5090), .o(delay_xor_ln21_unr3_stage2_stallmux_q_23_), .ck(clk) );
ms00f80 l0993 ( .d(n5095), .o(delay_xor_ln21_unr3_stage2_stallmux_q_7_), .ck(clk) );
ms00f80 l0994 ( .d(n5100), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_18_), .ck(clk) );
ms00f80 l0995 ( .d(n5105), .o(delay_xor_ln22_unr12_stage5_stallmux_q_13_), .ck(clk) );
ms00f80 l0996 ( .d(n5110), .o(delay_xor_ln21_unr9_stage4_stallmux_q_9_), .ck(clk) );
ms00f80 l0997 ( .d(n5115), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_15_), .ck(clk) );
ms00f80 l0998 ( .d(n5120), .o(delay_add_ln22_unr20_stage8_stallmux_q_11_), .ck(clk) );
ms00f80 l0999 ( .d(n5125), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_9_), .ck(clk) );
ms00f80 l1000 ( .d(n5130), .o(delay_xor_ln21_unr6_stage3_stallmux_q_20_), .ck(clk) );
ms00f80 l1001 ( .d(n5135), .o(delay_add_ln22_unr23_stage9_stallmux_q_15_), .ck(clk) );
ms00f80 l1002 ( .d(n5140), .o(delay_add_ln22_unr17_stage7_stallmux_q_21_), .ck(clk) );
ms00f80 l1003 ( .d(n5145), .o(delay_add_ln22_unr20_stage8_stallmux_q_9_), .ck(clk) );
ms00f80 l1004 ( .d(n5150), .o(delay_xor_ln21_unr3_stage2_stallmux_q_20_), .ck(clk) );
ms00f80 l1005 ( .d(n5155), .o(delay_xor_ln22_unr15_stage6_stallmux_q_11_), .ck(clk) );
ms00f80 l1006 ( .d(n5160), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_24_), .ck(clk) );
ms00f80 l1007 ( .d(n5165), .o(delay_xor_ln21_unr6_stage3_stallmux_q_3_), .ck(clk) );
ms00f80 l1008 ( .d(n5170), .o(delay_xor_ln22_unr28_stage10_stallmux_q_0_), .ck(clk) );
ms00f80 l1009 ( .d(n5175), .o(delay_add_ln22_unr14_stage6_stallmux_q_16_), .ck(clk) );
ms00f80 l1010 ( .d(n5180), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_26_), .ck(clk) );
ms00f80 l1011 ( .d(n5185), .o(delay_xor_ln22_unr15_stage6_stallmux_q_15_), .ck(clk) );
ms00f80 l1012 ( .d(n5190), .o(delay_xor_ln21_unr9_stage4_stallmux_q_8_), .ck(clk) );
ms00f80 l1013 ( .d(n5195), .o(delay_add_ln22_unr8_stage4_stallmux_q_24_), .ck(clk) );
ms00f80 l1014 ( .d(n5200), .o(delay_xor_ln21_unr21_stage8_stallmux_q_8_), .ck(clk) );
ms00f80 l1015 ( .d(n5205), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_19_), .ck(clk) );
ms00f80 l1016 ( .d(n5210), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_19_), .ck(clk) );
ms00f80 l1017 ( .d(n5215), .o(delay_add_ln22_unr2_stage2_stallmux_q_13_), .ck(clk) );
ms00f80 l1018 ( .d(n5220), .o(delay_add_ln22_unr5_stage3_stallmux_q_11_), .ck(clk) );
ms00f80 l1019 ( .d(n5225), .o(delay_sub_ln22_unr24_stage9_stallmux_q_2_), .ck(clk) );
ms00f80 l1020 ( .d(n5230), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_3_), .ck(clk) );
ms00f80 l1021 ( .d(n5235), .o(delay_xor_ln21_unr3_stage2_stallmux_q_15_), .ck(clk) );
ms00f80 l1022 ( .d(n5240), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_1_), .ck(clk) );
ms00f80 l1023 ( .d(n5245), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_8_), .ck(clk) );
ms00f80 l1024 ( .d(n5250), .o(delay_add_ln22_unr2_stage2_stallmux_q_10_), .ck(clk) );
ms00f80 l1025 ( .d(n5255), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_0_), .ck(clk) );
ms00f80 l1026 ( .d(n5260), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_17_), .ck(clk) );
ms00f80 l1027 ( .d(n5265), .o(delay_add_ln22_unr27_stage10_stallmux_q_4_), .ck(clk) );
ms00f80 l1028 ( .d(n5270), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_0_), .ck(clk) );
ms00f80 l1029 ( .d(n5275), .o(delay_add_ln22_unr23_stage9_stallmux_q_14_), .ck(clk) );
ms00f80 l1030 ( .d(n5280), .o(delay_xor_ln22_unr3_stage2_stallmux_q_21_), .ck(clk) );
ms00f80 l1031 ( .d(n5285), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_13_), .ck(clk) );
ms00f80 l1032 ( .d(n5290), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_21_), .ck(clk) );
ms00f80 l1033 ( .d(n5295), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_11_), .ck(clk) );
ms00f80 l1034 ( .d(n5300), .o(delay_xor_ln22_unr6_stage3_stallmux_q_22_), .ck(clk) );
ms00f80 l1035 ( .d(n5305), .o(delay_add_ln22_unr20_stage8_stallmux_q_19_), .ck(clk) );
ms00f80 l1036 ( .d(n5310), .o(delay_xor_ln21_unr3_stage2_stallmux_q_3_), .ck(clk) );
ms00f80 l1037 ( .d(n5315), .o(delay_xor_ln21_unr3_stage2_stallmux_q_28_), .ck(clk) );
ms00f80 l1038 ( .d(n5320), .o(delay_xor_ln21_unr6_stage3_stallmux_q_21_), .ck(clk) );
ms00f80 l1039 ( .d(n5325), .o(delay_add_ln22_unr20_stage8_stallmux_q_6_), .ck(clk) );
ms00f80 l1040 ( .d(n5330), .o(delay_add_ln22_unr17_stage7_stallmux_q_28_), .ck(clk) );
ms00f80 l1041 ( .d(n5335), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_25_), .ck(clk) );
ms00f80 l1042 ( .d(n5340), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_26_), .ck(clk) );
ms00f80 l1043 ( .d(n5345), .o(delay_add_ln22_unr2_stage2_stallmux_q_4_), .ck(clk) );
ms00f80 l1044 ( .d(n5350), .o(delay_xor_ln22_unr3_stage2_stallmux_q_17_), .ck(clk) );
ms00f80 l1045 ( .d(n5355), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_14_), .ck(clk) );
ms00f80 l1046 ( .d(n5360), .o(delay_xor_ln22_unr21_stage8_stallmux_q_2_), .ck(clk) );
ms00f80 l1047 ( .d(n5365), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_27_), .ck(clk) );
ms00f80 l1048 ( .d(n5370), .o(delay_xor_ln21_unr12_stage5_stallmux_q_15_), .ck(clk) );
ms00f80 l1049 ( .d(n5375), .o(delay_xor_ln22_unr3_stage2_stallmux_q_7_), .ck(clk) );
ms00f80 l1050 ( .d(n5380), .o(delay_sub_ln23_0_unr21_stage8_stallmux_q), .ck(clk) );
ms00f80 l1051 ( .d(n5385), .o(delay_add_ln22_unr14_stage6_stallmux_q_26_), .ck(clk) );
ms00f80 l1052 ( .d(n5390), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_20_), .ck(clk) );
ms00f80 l1053 ( .d(n5395), .o(delay_add_ln22_unr8_stage4_stallmux_q_30_), .ck(clk) );
ms00f80 l1054 ( .d(n5400), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_17_), .ck(clk) );
ms00f80 l1055 ( .d(n5405), .o(delay_add_ln22_unr11_stage5_stallmux_q_27_), .ck(clk) );
ms00f80 l1056 ( .d(n5410), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_25_), .ck(clk) );
ms00f80 l1057 ( .d(n5415), .o(delay_add_ln22_unr27_stage10_stallmux_q_8_), .ck(clk) );
ms00f80 l1058 ( .d(n5420), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_11_), .ck(clk) );
ms00f80 l1059 ( .d(n5425), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_28_), .ck(clk) );
ms00f80 l1060 ( .d(n5430), .o(delay_add_ln22_unr5_stage3_stallmux_q_13_), .ck(clk) );
ms00f80 l1061 ( .d(n5435), .o(delay_add_ln22_unr27_stage10_stallmux_q_3_), .ck(clk) );
ms00f80 l1062 ( .d(n5440), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_23_), .ck(clk) );
ms00f80 l1063 ( .d(n5445), .o(delay_xor_ln22_unr18_stage7_stallmux_q_3_), .ck(clk) );
ms00f80 l1064 ( .d(n5450), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_14_), .ck(clk) );
ms00f80 l1065 ( .d(n5455), .o(cos_out_24), .ck(clk) );
ms00f80 l1066 ( .d(n5459), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_27_), .ck(clk) );
ms00f80 l1067 ( .d(n5464), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_28_), .ck(clk) );
ms00f80 l1068 ( .d(n5469), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_29_), .ck(clk) );
ms00f80 l1069 ( .d(n5474), .o(delay_add_ln22_unr8_stage4_stallmux_q_20_), .ck(clk) );
ms00f80 l1070 ( .d(n5479), .o(sin_out_21), .ck(clk) );
ms00f80 l1071 ( .d(n5483), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_1_), .ck(clk) );
ms00f80 l1072 ( .d(n5488), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_15_), .ck(clk) );
ms00f80 l1073 ( .d(n5493), .o(delay_add_ln22_unr11_stage5_stallmux_q_19_), .ck(clk) );
ms00f80 l1074 ( .d(n5498), .o(delay_xor_ln22_unr12_stage5_stallmux_q_2_), .ck(clk) );
ms00f80 l1075 ( .d(n5503), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_23_), .ck(clk) );
ms00f80 l1076 ( .d(n5508), .o(delay_xor_ln21_unr9_stage4_stallmux_q_22_), .ck(clk) );
ms00f80 l1077 ( .d(n5513), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_10_), .ck(clk) );
ms00f80 l1078 ( .d(n5518), .o(delay_add_ln22_unr20_stage8_stallmux_q_12_), .ck(clk) );
ms00f80 l1079 ( .d(n5523), .o(delay_xor_ln22_unr15_stage6_stallmux_q_8_), .ck(clk) );
ms00f80 l1080 ( .d(n5528), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_28_), .ck(clk) );
ms00f80 l1081 ( .d(n5533), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_27_), .ck(clk) );
ms00f80 l1082 ( .d(n5538), .o(delay_add_ln22_unr17_stage7_stallmux_q_0_), .ck(clk) );
ms00f80 l1083 ( .d(n5543), .o(delay_add_ln22_unr17_stage7_stallmux_q_12_), .ck(clk) );
ms00f80 l1084 ( .d(n5548), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_19_), .ck(clk) );
ms00f80 l1085 ( .d(n5553), .o(delay_xor_ln21_unr12_stage5_stallmux_q_14_), .ck(clk) );
ms00f80 l1086 ( .d(n5558), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_4_), .ck(clk) );
ms00f80 l1087 ( .d(n5563), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_22_), .ck(clk) );
ms00f80 l1088 ( .d(n5568), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_7_), .ck(clk) );
ms00f80 l1089 ( .d(n5573), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_3_), .ck(clk) );
ms00f80 l1090 ( .d(n5578), .o(delay_add_ln22_unr17_stage7_stallmux_q_26_), .ck(clk) );
ms00f80 l1091 ( .d(n5583), .o(delay_add_ln22_unr5_stage3_stallmux_q_29_), .ck(clk) );
ms00f80 l1092 ( .d(n5588), .o(delay_sub_ln21_unr24_stage9_stallmux_q_3_), .ck(clk) );
ms00f80 l1093 ( .d(n5593), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_4_), .ck(clk) );
ms00f80 l1094 ( .d(n5598), .o(delay_xor_ln22_unr9_stage4_stallmux_q_14_), .ck(clk) );
ms00f80 l1095 ( .d(n5603), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_15_), .ck(clk) );
ms00f80 l1096 ( .d(n5608), .o(delay_xor_ln22_unr15_stage6_stallmux_q_2_), .ck(clk) );
ms00f80 l1097 ( .d(n5613), .o(delay_add_ln22_unr23_stage9_stallmux_q_2_), .ck(clk) );
ms00f80 l1098 ( .d(n5618), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_0_), .ck(clk) );
ms00f80 l1099 ( .d(n5623), .o(delay_sub_ln21_unr24_stage9_stallmux_q_2_), .ck(clk) );
ms00f80 l1100 ( .d(n5628), .o(delay_add_ln22_unr2_stage2_stallmux_q_19_), .ck(clk) );
ms00f80 l1101 ( .d(n5633), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_19_), .ck(clk) );
ms00f80 l1102 ( .d(n5638), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_4_), .ck(clk) );
ms00f80 l1103 ( .d(n5643), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_22_), .ck(clk) );
ms00f80 l1104 ( .d(n5648), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_19_), .ck(clk) );
ms00f80 l1105 ( .d(n5653), .o(cos_out_1), .ck(clk) );
ms00f80 l1106 ( .d(n5657), .o(delay_xor_ln21_unr15_stage6_stallmux_q_13_), .ck(clk) );
ms00f80 l1107 ( .d(n5662), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_20_), .ck(clk) );
ms00f80 l1108 ( .d(n5667), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_24_), .ck(clk) );
ms00f80 l1109 ( .d(n5672), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_2_), .ck(clk) );
ms00f80 l1110 ( .d(n5677), .o(delay_xor_ln21_unr3_stage2_stallmux_q_14_), .ck(clk) );
ms00f80 l1111 ( .d(n5682), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_15_), .ck(clk) );
ms00f80 l1112 ( .d(n5687), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_23_), .ck(clk) );
ms00f80 l1113 ( .d(n5692), .o(delay_add_ln22_unr11_stage5_stallmux_q_16_), .ck(clk) );
ms00f80 l1114 ( .d(n5697), .o(sin_out_16), .ck(clk) );
ms00f80 l1115 ( .d(n5701), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_29_), .ck(clk) );
ms00f80 l1116 ( .d(n5706), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_5_), .ck(clk) );
ms00f80 l1117 ( .d(n5711), .o(delay_xor_ln22_unr3_stage2_stallmux_q_22_), .ck(clk) );
ms00f80 l1118 ( .d(n5716), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_6_), .ck(clk) );
ms00f80 l1119 ( .d(n5721), .o(delay_xor_ln21_unr9_stage4_stallmux_q_10_), .ck(clk) );
ms00f80 l1120 ( .d(n5726), .o(sin_out_28), .ck(clk) );
ms00f80 l1121 ( .d(n5730), .o(delay_add_ln22_unr5_stage3_stallmux_q_24_), .ck(clk) );
ms00f80 l1122 ( .d(n5735), .o(delay_add_ln22_unr11_stage5_stallmux_q_15_), .ck(clk) );
ms00f80 l1123 ( .d(n5740), .o(delay_xor_ln22_unr6_stage3_stallmux_q_4_), .ck(clk) );
ms00f80 l1124 ( .d(n5745), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_30_), .ck(clk) );
ms00f80 l1125 ( .d(n5750), .o(delay_xor_ln21_unr3_stage2_stallmux_q_11_), .ck(clk) );
ms00f80 l1126 ( .d(n5755), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_7_), .ck(clk) );
ms00f80 l1127 ( .d(n5760), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_19_), .ck(clk) );
ms00f80 l1128 ( .d(n5765), .o(sin_out_18), .ck(clk) );
ms00f80 l1129 ( .d(n5769), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_6_), .ck(clk) );
ms00f80 l1130 ( .d(n5774), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_21_), .ck(clk) );
ms00f80 l1131 ( .d(n5779), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_3_), .ck(clk) );
ms00f80 l1132 ( .d(n5784), .o(delay_xor_ln22_unr6_stage3_stallmux_q_21_), .ck(clk) );
ms00f80 l1133 ( .d(n5789), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_29_), .ck(clk) );
ms00f80 l1134 ( .d(n5794), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_12_), .ck(clk) );
ms00f80 l1135 ( .d(n5799), .o(n_45224), .ck(clk) );
ms00f80 l1136 ( .d(n5804), .o(delay_xor_ln21_unr18_stage7_stallmux_q_5_), .ck(clk) );
ms00f80 l1137 ( .d(n5809), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_8_), .ck(clk) );
ms00f80 l1138 ( .d(n5814), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_9_), .ck(clk) );
ms00f80 l1139 ( .d(n5819), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_11_), .ck(clk) );
ms00f80 l1140 ( .d(n5824), .o(delay_xor_ln21_unr18_stage7_stallmux_q_7_), .ck(clk) );
ms00f80 l1141 ( .d(n5829), .o(delay_xor_ln22_unr18_stage7_stallmux_q_11_), .ck(clk) );
ms00f80 l1142 ( .d(n5834), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_18_), .ck(clk) );
ms00f80 l1143 ( .d(n5839), .o(n_45209), .ck(clk) );
ms00f80 l1144 ( .d(n5844), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_24_), .ck(clk) );
ms00f80 l1145 ( .d(n5849), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_17_), .ck(clk) );
ms00f80 l1146 ( .d(n5854), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_6_), .ck(clk) );
ms00f80 l1147 ( .d(n5859), .o(delay_add_ln22_unr14_stage6_stallmux_q_13_), .ck(clk) );
ms00f80 l1148 ( .d(n5864), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_30_), .ck(clk) );
ms00f80 l1149 ( .d(n5869), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_11_), .ck(clk) );
ms00f80 l1150 ( .d(n5874), .o(cos_out_8), .ck(clk) );
ms00f80 l1151 ( .d(n5878), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_5_), .ck(clk) );
ms00f80 l1152 ( .d(n5883), .o(delay_add_ln22_unr20_stage8_stallmux_q_29_), .ck(clk) );
ms00f80 l1153 ( .d(n5888), .o(delay_add_ln22_unr2_stage2_stallmux_q_31_), .ck(clk) );
ms00f80 l1154 ( .d(n5893), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_27_), .ck(clk) );
ms00f80 l1155 ( .d(n5898), .o(delay_add_ln22_unr17_stage7_stallmux_q_2_), .ck(clk) );
ms00f80 l1156 ( .d(n5903), .o(delay_add_ln22_unr11_stage5_stallmux_q_22_), .ck(clk) );
ms00f80 l1157 ( .d(n5908), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_26_), .ck(clk) );
ms00f80 l1158 ( .d(n5913), .o(delay_add_ln22_unr8_stage4_stallmux_q_21_), .ck(clk) );
ms00f80 l1159 ( .d(n5918), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_7_), .ck(clk) );
ms00f80 l1160 ( .d(n5923), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_21_), .ck(clk) );
ms00f80 l1161 ( .d(n5928), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_21_), .ck(clk) );
ms00f80 l1162 ( .d(n5933), .o(delay_add_ln22_unr27_stage10_stallmux_q_27_), .ck(clk) );
ms00f80 l1163 ( .d(n5938), .o(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .ck(clk) );
ms00f80 l1164 ( .d(n5943), .o(delay_xor_ln22_unr6_stage3_stallmux_q_9_), .ck(clk) );
ms00f80 l1165 ( .d(n5948), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_20_), .ck(clk) );
ms00f80 l1166 ( .d(n5953), .o(delay_add_ln22_unr14_stage6_stallmux_q_6_), .ck(clk) );
ms00f80 l1167 ( .d(n5958), .o(delay_xor_ln21_unr15_stage6_stallmux_q_1_), .ck(clk) );
ms00f80 l1168 ( .d(n5963), .o(delay_xor_ln22_unr9_stage4_stallmux_q_8_), .ck(clk) );
ms00f80 l1169 ( .d(n5968), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_4_), .ck(clk) );
ms00f80 l1170 ( .d(n5973), .o(delay_sub_ln23_0_unr15_stage6_stallmux_q), .ck(clk) );
ms00f80 l1171 ( .d(n5978), .o(delay_sub_ln23_0_unr22_stage8_stallmux_q), .ck(clk) );
ms00f80 l1172 ( .d(n5983), .o(delay_xor_ln21_unr18_stage7_stallmux_q_3_), .ck(clk) );
ms00f80 l1173 ( .d(n5988), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_24_), .ck(clk) );
ms00f80 l1174 ( .d(n5993), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_0_), .ck(clk) );
ms00f80 l1175 ( .d(n5998), .o(delay_xor_ln21_unr18_stage7_stallmux_q_11_), .ck(clk) );
ms00f80 l1176 ( .d(n6003), .o(cos_out_16), .ck(clk) );
ms00f80 l1177 ( .d(n6007), .o(delay_xor_ln21_unr18_stage7_stallmux_q_6_), .ck(clk) );
ms00f80 l1178 ( .d(n6012), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_20_), .ck(clk) );
ms00f80 l1179 ( .d(n6017), .o(delay_add_ln22_unr17_stage7_stallmux_q_20_), .ck(clk) );
ms00f80 l1180 ( .d(n6022), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_22_), .ck(clk) );
ms00f80 l1181 ( .d(n6027), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_5_), .ck(clk) );
ms00f80 l1182 ( .d(n6032), .o(delay_xor_ln22_unr12_stage5_stallmux_q_8_), .ck(clk) );
ms00f80 l1183 ( .d(n6037), .o(n_44365), .ck(clk) );
ms00f80 l1184 ( .d(n6042), .o(delay_add_ln22_unr8_stage4_stallmux_q_6_), .ck(clk) );
ms00f80 l1185 ( .d(n6047), .o(delay_add_ln22_unr5_stage3_stallmux_q_23_), .ck(clk) );
ms00f80 l1186 ( .d(n6051), .o(delay_sub_ln23_0_unr28_stage10_stallmux_q), .ck(clk) );
ms00f80 l1187 ( .d(n6056), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_17_), .ck(clk) );
ms00f80 l1188 ( .d(n6061), .o(delay_add_ln22_unr5_stage3_stallmux_q_19_), .ck(clk) );
ms00f80 l1189 ( .d(n6066), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_3_), .ck(clk) );
ms00f80 l1190 ( .d(n6071), .o(delay_xor_ln21_unr15_stage6_stallmux_q_3_), .ck(clk) );
ms00f80 l1191 ( .d(n6076), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_18_), .ck(clk) );
ms00f80 l1192 ( .d(n6081), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_16_), .ck(clk) );
ms00f80 l1193 ( .d(n6086), .o(delay_xor_ln21_unr12_stage5_stallmux_q_9_), .ck(clk) );
ms00f80 l1194 ( .d(n6091), .o(delay_xor_ln21_unr9_stage4_stallmux_q_14_), .ck(clk) );
ms00f80 l1195 ( .d(n6096), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_15_), .ck(clk) );
ms00f80 l1196 ( .d(n6101), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_15_), .ck(clk) );
ms00f80 l1197 ( .d(n6106), .o(delay_add_ln22_unr17_stage7_stallmux_q_23_), .ck(clk) );
ms00f80 l1198 ( .d(n6111), .o(delay_add_ln22_unr11_stage5_stallmux_q_9_), .ck(clk) );
ms00f80 l1199 ( .d(n6116), .o(delay_add_ln22_unr14_stage6_stallmux_q_19_), .ck(clk) );
ms00f80 l1200 ( .d(n6121), .o(sin_out_26), .ck(clk) );
ms00f80 l1201 ( .d(n6125), .o(delay_add_ln22_unr14_stage6_stallmux_q_18_), .ck(clk) );
ms00f80 l1202 ( .d(n6130), .o(delay_add_ln22_unr20_stage8_stallmux_q_7_), .ck(clk) );
ms00f80 l1203 ( .d(n6135), .o(delay_add_ln22_unr27_stage10_stallmux_q_2_), .ck(clk) );
ms00f80 l1204 ( .d(n6140), .o(delay_xor_ln21_unr15_stage6_stallmux_q_2_), .ck(clk) );
ms00f80 l1205 ( .d(n6145), .o(delay_xor_ln22_unr9_stage4_stallmux_q_6_), .ck(clk) );
ms00f80 l1206 ( .d(n6149), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_9_), .ck(clk) );
ms00f80 l1207 ( .d(n6154), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_26_), .ck(clk) );
ms00f80 l1208 ( .d(n6159), .o(cos_out_9), .ck(clk) );
ms00f80 l1209 ( .d(n6163), .o(delay_add_ln22_unr14_stage6_stallmux_q_10_), .ck(clk) );
ms00f80 l1210 ( .d(n6168), .o(sin_out_31), .ck(clk) );
ms00f80 l1211 ( .d(n6172), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_30_), .ck(clk) );
ms00f80 l1212 ( .d(n6177), .o(delay_add_ln22_unr8_stage4_stallmux_q_7_), .ck(clk) );
ms00f80 l1213 ( .d(n6182), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_19_), .ck(clk) );
ms00f80 l1214 ( .d(n6187), .o(delay_add_ln22_unr27_stage10_stallmux_q_26_), .ck(clk) );
ms00f80 l1215 ( .d(n6192), .o(delay_xor_ln22_unr15_stage6_stallmux_q_9_), .ck(clk) );
ms00f80 l1216 ( .d(n6197), .o(delay_xor_ln22_unr12_stage5_stallmux_q_15_), .ck(clk) );
ms00f80 l1217 ( .d(n6202), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_16_), .ck(clk) );
ms00f80 l1218 ( .d(n6207), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_5_), .ck(clk) );
ms00f80 l1219 ( .d(n6212), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_17_), .ck(clk) );
ms00f80 l1220 ( .d(n6217), .o(delay_add_ln22_unr20_stage8_stallmux_q_27_), .ck(clk) );
ms00f80 l1221 ( .d(n6222), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_25_), .ck(clk) );
ms00f80 l1222 ( .d(n6227), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_16_), .ck(clk) );
ms00f80 l1223 ( .d(n6231), .o(delay_xor_ln22_unr3_stage2_stallmux_q_11_), .ck(clk) );
ms00f80 l1224 ( .d(n6236), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_10_), .ck(clk) );
ms00f80 l1225 ( .d(n6241), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_2_), .ck(clk) );
ms00f80 l1226 ( .d(n6246), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_25_), .ck(clk) );
ms00f80 l1227 ( .d(n6251), .o(delay_xor_ln22_unr18_stage7_stallmux_q_8_), .ck(clk) );
ms00f80 l1228 ( .d(n6256), .o(delay_add_ln22_unr5_stage3_stallmux_q_5_), .ck(clk) );
ms00f80 l1229 ( .d(n6260), .o(delay_sub_ln23_0_unr24_stage9_stallmux_q), .ck(clk) );
ms00f80 l1230 ( .d(n6265), .o(delay_add_ln22_unr27_stage10_stallmux_q_0_), .ck(clk) );

endmodule
