../libs/open_design_flow.lef