// Latch-mapped netlist written by map_latches.py, 2019-06-04 13:24:08
// Written ISPD/ICCAD/TAU contest Verilog format. 
//    Input file:  ac97_ctrl/ac97_ctrl_remapped.v
//    Latch cell:  ms00f80
//    Clock port:  clk
//    Output file: ac97_ctrl/ac97_ctrl_remapped.v

module ac97_ctrl (
clk,
x1006,
x1034,
x1062,
x1101,
x1126,
x1155,
x1193,
x1203,
x1209,
x1215,
x1231,
x1261,
x1286,
x130629,
x130630,
x130631,
x130632,
x130633,
x130634,
x130635,
x130636,
x130637,
x130638,
x130639,
x130640,
x130641,
x130642,
x130643,
x130644,
x130645,
x130646,
x130647,
x130648,
x130649,
x130650,
x130651,
x130652,
x130653,
x130654,
x130655,
x130656,
x130657,
x1322,
x1345,
x1351,
x1358,
x1366,
x1374,
x1382,
x1390,
x1398,
x1406,
x1417,
x1424,
x1432,
x1443,
x1451,
x1459,
x1467,
x1479,
x1486,
x1494,
x1501,
x1511,
x1519,
x1527,
x1534,
x1542,
x1550,
x1557,
x1564,
x1572,
x1580,
x1587,
x1595,
x1822,
x806,
x821,
x837,
x868,
x889,
x906,
x940,
x977,
x0,
x101,
x106,
x114,
x124,
x131,
x138,
x14,
x145,
x149,
x172,
x179,
x187,
x195,
x217,
x234,
x249,
x264,
x287,
x30,
x315,
x342,
x361,
x379,
x38,
x390,
x397,
x420,
x447,
x476,
x494,
x522,
x538,
x561,
x589,
x620,
x63,
x638,
x657,
x681,
x699,
x718,
x744,
x765,
x77,
x786,
x84,
x96
);

// Start PIs
input clk;
input x1006;
input x1034;
input x1062;
input x1101;
input x1126;
input x1155;
input x1193;
input x1203;
input x1209;
input x1215;
input x1231;
input x1261;
input x1286;
input x130629;
input x130630;
input x130631;
input x130632;
input x130633;
input x130634;
input x130635;
input x130636;
input x130637;
input x130638;
input x130639;
input x130640;
input x130641;
input x130642;
input x130643;
input x130644;
input x130645;
input x130646;
input x130647;
input x130648;
input x130649;
input x130650;
input x130651;
input x130652;
input x130653;
input x130654;
input x130655;
input x130656;
input x130657;
input x1322;
input x1345;
input x1351;
input x1358;
input x1366;
input x1374;
input x1382;
input x1390;
input x1398;
input x1406;
input x1417;
input x1424;
input x1432;
input x1443;
input x1451;
input x1459;
input x1467;
input x1479;
input x1486;
input x1494;
input x1501;
input x1511;
input x1519;
input x1527;
input x1534;
input x1542;
input x1550;
input x1557;
input x1564;
input x1572;
input x1580;
input x1587;
input x1595;
input x1822;
input x806;
input x821;
input x837;
input x868;
input x889;
input x906;
input x940;
input x977;

// Start POs
output x0;
output x101;
output x106;
output x114;
output x124;
output x131;
output x138;
output x14;
output x145;
output x149;
output x172;
output x179;
output x187;
output x195;
output x217;
output x234;
output x249;
output x264;
output x287;
output x30;
output x315;
output x342;
output x361;
output x379;
output x38;
output x390;
output x397;
output x420;
output x447;
output x476;
output x494;
output x522;
output x538;
output x561;
output x589;
output x620;
output x63;
output x638;
output x657;
output x681;
output x699;
output x718;
output x744;
output x765;
output x77;
output x786;
output x84;
output x96;

// Start wires
wire clk;
wire x1006;
wire x1034;
wire x1062;
wire x1101;
wire x1126;
wire x1155;
wire x1193;
wire x1203;
wire x1209;
wire x1215;
wire x1231;
wire x1261;
wire x1286;
wire x130629;
wire x130630;
wire x130631;
wire x130632;
wire x130633;
wire x130634;
wire x130635;
wire x130636;
wire x130637;
wire x130638;
wire x130639;
wire x130640;
wire x130641;
wire x130642;
wire x130643;
wire x130644;
wire x130645;
wire x130646;
wire x130647;
wire x130648;
wire x130649;
wire x130650;
wire x130651;
wire x130652;
wire x130653;
wire x130654;
wire x130655;
wire x130656;
wire x130657;
wire x1322;
wire x1345;
wire x1351;
wire x1358;
wire x1366;
wire x1374;
wire x1382;
wire x1390;
wire x1398;
wire x1406;
wire x1417;
wire x1424;
wire x1432;
wire x1443;
wire x1451;
wire x1459;
wire x1467;
wire x1479;
wire x1486;
wire x1494;
wire x1501;
wire x1511;
wire x1519;
wire x1527;
wire x1534;
wire x1542;
wire x1550;
wire x1557;
wire x1564;
wire x1572;
wire x1580;
wire x1587;
wire x1595;
wire x1822;
wire x806;
wire x821;
wire x837;
wire x868;
wire x889;
wire x906;
wire x940;
wire x977;
wire x0;
wire x101;
wire x106;
wire x114;
wire x124;
wire x131;
wire x138;
wire x14;
wire x145;
wire x149;
wire x172;
wire x179;
wire x187;
wire x195;
wire x217;
wire x234;
wire x249;
wire x264;
wire x287;
wire x30;
wire x315;
wire x342;
wire x361;
wire x379;
wire x38;
wire x390;
wire x397;
wire x420;
wire x447;
wire x476;
wire x494;
wire x522;
wire x538;
wire x561;
wire x589;
wire x620;
wire x63;
wire x638;
wire x657;
wire x681;
wire x699;
wire x718;
wire x744;
wire x765;
wire x77;
wire x786;
wire x84;
wire x96;
wire _net_113;
wire _net_114;
wire _net_115;
wire _net_116;
wire _net_117;
wire _net_118;
wire _net_119;
wire _net_120;
wire _net_121;
wire _net_122;
wire _net_123;
wire _net_124;
wire _net_125;
wire _net_126;
wire _net_127;
wire _net_128;
wire _net_129;
wire _net_154;
wire _net_172;
wire _net_173;
wire _net_174;
wire _net_175;
wire _net_176;
wire _net_177;
wire _net_178;
wire _net_180;
wire _net_184;
wire _net_188;
wire _net_189;
wire _net_190;
wire _net_191;
wire _net_192;
wire _net_193;
wire _net_201;
wire _net_209;
wire _net_210;
wire _net_211;
wire _net_212;
wire _net_213;
wire _net_214;
wire _net_215;
wire _net_217;
wire _net_221;
wire _net_225;
wire _net_226;
wire _net_227;
wire _net_228;
wire _net_229;
wire _net_262;
wire _net_263;
wire _net_264;
wire _net_265;
wire _net_266;
wire _net_267;
wire _net_268;
wire _net_269;
wire _net_270;
wire _net_271;
wire _net_272;
wire _net_273;
wire _net_276;
wire _net_277;
wire _net_278;
wire _net_279;
wire _net_280;
wire _net_281;
wire _net_282;
wire _net_283;
wire _net_284;
wire _net_287;
wire _net_288;
wire _net_289;
wire _net_290;
wire _net_291;
wire _net_292;
wire _net_293;
wire _net_294;
wire _net_295;
wire _net_298;
wire _net_299;
wire _net_392;
wire _net_5848;
wire _net_5850;
wire _net_5851;
wire _net_5852;
wire _net_5853;
wire _net_5854;
wire _net_5855;
wire _net_5856;
wire _net_5857;
wire _net_5859;
wire _net_5920;
wire _net_5922;
wire _net_5924;
wire _net_5960;
wire _net_5961;
wire _net_5962;
wire _net_5963;
wire _net_5964;
wire _net_5965;
wire _net_5966;
wire _net_5967;
wire _net_5968;
wire _net_5969;
wire _net_5970;
wire _net_5971;
wire _net_5972;
wire _net_5973;
wire _net_5974;
wire _net_5975;
wire _net_5976;
wire _net_5977;
wire _net_5978;
wire _net_5979;
wire _net_5980;
wire _net_5981;
wire _net_5982;
wire _net_5983;
wire _net_5984;
wire _net_5985;
wire _net_5986;
wire _net_5987;
wire _net_5988;
wire _net_5989;
wire _net_5990;
wire _net_5991;
wire _net_5993;
wire _net_5994;
wire _net_5995;
wire _net_5996;
wire _net_5997;
wire _net_5998;
wire _net_5999;
wire _net_6000;
wire _net_6001;
wire _net_6002;
wire _net_6004;
wire _net_6005;
wire _net_6006;
wire _net_6007;
wire _net_6008;
wire _net_6009;
wire _net_6010;
wire _net_6011;
wire _net_6012;
wire _net_6015;
wire _net_6016;
wire _net_6017;
wire _net_6018;
wire _net_6019;
wire _net_6020;
wire _net_6021;
wire _net_6022;
wire _net_6023;
wire _net_6026;
wire _net_6027;
wire _net_6028;
wire _net_6029;
wire _net_6030;
wire _net_6031;
wire _net_6032;
wire _net_6033;
wire _net_6034;
wire _net_6037;
wire _net_6038;
wire _net_6039;
wire _net_6040;
wire _net_6041;
wire _net_6042;
wire _net_6043;
wire _net_6044;
wire _net_6045;
wire _net_6048;
wire _net_6049;
wire _net_6050;
wire _net_6051;
wire _net_6052;
wire _net_6062;
wire _net_6063;
wire _net_6064;
wire _net_6065;
wire _net_6066;
wire _net_6067;
wire _net_6068;
wire _net_6069;
wire _net_6070;
wire _net_6071;
wire _net_6072;
wire _net_6073;
wire _net_6074;
wire _net_6075;
wire _net_6076;
wire _net_6077;
wire _net_6078;
wire _net_6079;
wire _net_6080;
wire _net_6081;
wire _net_6082;
wire _net_6083;
wire _net_6084;
wire _net_6085;
wire _net_6086;
wire _net_6087;
wire _net_6088;
wire _net_6089;
wire _net_6090;
wire _net_6091;
wire _net_6092;
wire _net_6093;
wire _net_6094;
wire _net_6095;
wire _net_6096;
wire _net_6097;
wire _net_6098;
wire _net_6099;
wire _net_6100;
wire _net_6101;
wire _net_6102;
wire _net_6103;
wire _net_6104;
wire _net_6105;
wire _net_6106;
wire _net_6107;
wire _net_6108;
wire _net_6109;
wire _net_6110;
wire _net_6111;
wire _net_6112;
wire _net_6113;
wire _net_6114;
wire _net_6115;
wire _net_6116;
wire _net_6117;
wire _net_6118;
wire _net_6119;
wire _net_6120;
wire _net_6121;
wire _net_6122;
wire _net_6123;
wire _net_6124;
wire _net_6125;
wire _net_6126;
wire _net_6127;
wire _net_6128;
wire _net_6129;
wire _net_6130;
wire _net_6131;
wire _net_6132;
wire _net_6133;
wire _net_6134;
wire _net_6135;
wire _net_6136;
wire _net_6137;
wire _net_6138;
wire _net_6139;
wire _net_6140;
wire _net_6141;
wire _net_6142;
wire _net_6143;
wire _net_6144;
wire _net_6145;
wire _net_6146;
wire _net_6147;
wire _net_6148;
wire _net_6149;
wire _net_6150;
wire _net_6151;
wire _net_6152;
wire _net_6153;
wire _net_6154;
wire _net_6155;
wire _net_6156;
wire _net_6157;
wire _net_6158;
wire _net_6159;
wire _net_6160;
wire _net_6161;
wire _net_6162;
wire _net_6163;
wire _net_6164;
wire _net_6165;
wire _net_6166;
wire _net_6167;
wire _net_6168;
wire _net_6169;
wire _net_6170;
wire _net_6171;
wire _net_6172;
wire _net_6173;
wire _net_6174;
wire _net_6175;
wire _net_6176;
wire _net_6177;
wire _net_6178;
wire _net_6179;
wire _net_6180;
wire _net_6181;
wire _net_6182;
wire _net_6183;
wire _net_6184;
wire _net_6185;
wire _net_6186;
wire _net_6187;
wire _net_6188;
wire _net_6189;
wire _net_6194;
wire _net_6199;
wire _net_6200;
wire _net_6201;
wire _net_6202;
wire _net_6203;
wire _net_6204;
wire _net_6205;
wire _net_6206;
wire _net_6207;
wire _net_6208;
wire _net_6209;
wire _net_6210;
wire _net_6219;
wire _net_6220;
wire _net_6221;
wire _net_6222;
wire _net_6239;
wire _net_6259;
wire _net_6280;
wire _net_6281;
wire _net_6282;
wire _net_6283;
wire _net_6284;
wire _net_6285;
wire _net_6286;
wire _net_6287;
wire _net_6288;
wire _net_6289;
wire _net_6290;
wire _net_6291;
wire _net_6292;
wire _net_6293;
wire _net_6294;
wire _net_6295;
wire _net_6296;
wire _net_6297;
wire _net_6298;
wire _net_6319;
wire _net_6401;
wire _net_6402;
wire _net_6404;
wire _net_6405;
wire _net_6406;
wire _net_6407;
wire _net_6408;
wire _net_6409;
wire _net_6410;
wire _net_6411;
wire _net_6413;
wire _net_6414;
wire _net_6415;
wire _net_6418;
wire _net_6419;
wire _net_6420;
wire _net_6421;
wire _net_6422;
wire _net_6423;
wire _net_6552;
wire _net_6553;
wire _net_6554;
wire _net_6555;
wire _net_6557;
wire _net_6558;
wire _net_6687;
wire _net_6688;
wire _net_6689;
wire _net_6690;
wire _net_6692;
wire _net_6693;
wire _net_6822;
wire _net_6823;
wire _net_6824;
wire _net_6825;
wire _net_6827;
wire _net_6828;
wire _net_6957;
wire _net_6958;
wire _net_6959;
wire _net_6960;
wire _net_6962;
wire _net_6963;
wire _net_7092;
wire _net_7093;
wire _net_7094;
wire _net_7095;
wire _net_7097;
wire _net_7098;
wire _net_7227;
wire _net_7228;
wire _net_7229;
wire _net_7230;
wire _net_7232;
wire _net_7233;
wire _net_7250;
wire _net_7251;
wire _net_7252;
wire _net_7253;
wire _net_7254;
wire _net_7255;
wire _net_7256;
wire _net_7257;
wire _net_7258;
wire _net_7259;
wire _net_7260;
wire _net_7261;
wire _net_7262;
wire _net_7263;
wire _net_7264;
wire _net_7265;
wire _net_7266;
wire _net_7267;
wire _net_7268;
wire _net_7269;
wire _net_7270;
wire _net_7271;
wire _net_7272;
wire _net_7273;
wire _net_7274;
wire _net_7275;
wire _net_7276;
wire _net_7277;
wire _net_7278;
wire _net_7279;
wire _net_7280;
wire _net_7281;
wire _net_7282;
wire _net_7283;
wire _net_7284;
wire _net_7285;
wire _net_7286;
wire _net_7287;
wire _net_7288;
wire _net_7289;
wire _net_7290;
wire _net_7291;
wire _net_7292;
wire _net_7293;
wire _net_7294;
wire _net_7295;
wire _net_7296;
wire _net_7297;
wire _net_7298;
wire _net_7299;
wire _net_7300;
wire _net_7301;
wire _net_7314;
wire _net_7315;
wire _net_7316;
wire _net_7317;
wire _net_7318;
wire _net_7319;
wire _net_7320;
wire _net_7321;
wire _net_7322;
wire _net_7323;
wire _net_7324;
wire _net_7325;
wire _net_7326;
wire _net_7327;
wire _net_7328;
wire _net_7329;
wire _net_7330;
wire _net_7331;
wire _net_7332;
wire _net_7333;
wire _net_7346;
wire _net_7347;
wire _net_7348;
wire _net_7349;
wire _net_7350;
wire _net_7351;
wire _net_7352;
wire _net_7353;
wire _net_7354;
wire _net_7355;
wire _net_7356;
wire _net_7357;
wire _net_7358;
wire _net_7359;
wire _net_7360;
wire _net_7361;
wire _net_7362;
wire _net_7363;
wire _net_7364;
wire _net_7365;
wire _net_7379;
wire _net_7380;
wire _net_7381;
wire _net_7382;
wire _net_7383;
wire _net_7384;
wire _net_7401;
wire _net_7402;
wire _net_7403;
wire _net_7404;
wire _net_7405;
wire _net_7406;
wire _net_7407;
wire _net_7408;
wire _net_7409;
wire _net_7410;
wire _net_7411;
wire _net_7412;
wire _net_7413;
wire _net_7414;
wire _net_7415;
wire _net_7416;
wire _net_7417;
wire _net_7418;
wire _net_7419;
wire _net_7420;
wire _net_7421;
wire _net_7422;
wire _net_7423;
wire _net_7424;
wire _net_7425;
wire _net_7426;
wire _net_7427;
wire _net_7428;
wire _net_7429;
wire _net_7430;
wire _net_7431;
wire _net_7432;
wire _net_7433;
wire _net_7434;
wire _net_7435;
wire _net_7436;
wire _net_7437;
wire _net_7438;
wire _net_7439;
wire _net_7440;
wire _net_7441;
wire _net_7442;
wire _net_7443;
wire _net_7444;
wire _net_7445;
wire _net_7446;
wire _net_7447;
wire _net_7448;
wire _net_7449;
wire _net_7450;
wire _net_7451;
wire _net_7452;
wire _net_7465;
wire _net_7466;
wire _net_7467;
wire _net_7468;
wire _net_7469;
wire _net_7470;
wire _net_7471;
wire _net_7472;
wire _net_7473;
wire _net_7474;
wire _net_7475;
wire _net_7476;
wire _net_7477;
wire _net_7478;
wire _net_7479;
wire _net_7480;
wire _net_7481;
wire _net_7482;
wire _net_7483;
wire _net_7484;
wire _net_7497;
wire _net_7498;
wire _net_7499;
wire _net_7500;
wire _net_7501;
wire _net_7502;
wire _net_7503;
wire _net_7504;
wire _net_7505;
wire _net_7506;
wire _net_7507;
wire _net_7508;
wire _net_7509;
wire _net_7510;
wire _net_7511;
wire _net_7512;
wire _net_7513;
wire _net_7514;
wire _net_7515;
wire _net_7516;
wire _net_7530;
wire _net_7531;
wire _net_7532;
wire _net_7533;
wire _net_7534;
wire _net_7535;
wire _net_7552;
wire _net_7553;
wire _net_7554;
wire _net_7555;
wire _net_7556;
wire _net_7557;
wire _net_7558;
wire _net_7559;
wire _net_7560;
wire _net_7561;
wire _net_7562;
wire _net_7563;
wire _net_7564;
wire _net_7565;
wire _net_7566;
wire _net_7567;
wire _net_7568;
wire _net_7569;
wire _net_7570;
wire _net_7571;
wire _net_7572;
wire _net_7573;
wire _net_7574;
wire _net_7575;
wire _net_7576;
wire _net_7577;
wire _net_7578;
wire _net_7579;
wire _net_7580;
wire _net_7581;
wire _net_7582;
wire _net_7583;
wire _net_7584;
wire _net_7585;
wire _net_7586;
wire _net_7587;
wire _net_7588;
wire _net_7589;
wire _net_7590;
wire _net_7591;
wire _net_7592;
wire _net_7593;
wire _net_7594;
wire _net_7595;
wire _net_7596;
wire _net_7597;
wire _net_7598;
wire _net_7599;
wire _net_7600;
wire _net_7601;
wire _net_7602;
wire _net_7603;
wire _net_7616;
wire _net_7617;
wire _net_7618;
wire _net_7619;
wire _net_7620;
wire _net_7621;
wire _net_7622;
wire _net_7623;
wire _net_7624;
wire _net_7625;
wire _net_7626;
wire _net_7627;
wire _net_7628;
wire _net_7629;
wire _net_7630;
wire _net_7631;
wire _net_7632;
wire _net_7633;
wire _net_7634;
wire _net_7635;
wire _net_7648;
wire _net_7649;
wire _net_7650;
wire _net_7651;
wire _net_7652;
wire _net_7653;
wire _net_7654;
wire _net_7655;
wire _net_7656;
wire _net_7657;
wire _net_7658;
wire _net_7659;
wire _net_7660;
wire _net_7661;
wire _net_7662;
wire _net_7663;
wire _net_7664;
wire _net_7665;
wire _net_7666;
wire _net_7667;
wire _net_7681;
wire _net_7682;
wire _net_7683;
wire _net_7684;
wire _net_7685;
wire _net_7686;
wire _net_7687;
wire _net_7688;
wire _net_7689;
wire _net_7690;
wire _net_7692;
wire _net_7693;
wire _net_7694;
wire _net_7695;
wire _net_7696;
wire _net_7697;
wire _net_7698;
wire _net_7699;
wire _net_7700;
wire _net_7701;
wire _net_7702;
wire _net_7703;
wire _net_7704;
wire _net_7705;
wire _net_7706;
wire _net_7707;
wire _net_7716;
wire _net_7717;
wire _net_7718;
wire _net_7719;
wire _net_7720;
wire _net_7721;
wire _net_7722;
wire _net_7723;
wire _net_7724;
wire _net_7725;
wire _net_7726;
wire _net_7727;
wire _net_7728;
wire _net_7729;
wire _net_7730;
wire _net_7731;
wire _net_7732;
wire _net_7733;
wire _net_7734;
wire _net_7735;
wire _net_7736;
wire _net_7745;
wire _net_7746;
wire _net_7747;
wire _net_7748;
wire _net_7749;
wire _net_7751;
wire _net_7753;
wire _net_7755;
wire _net_7757;
wire _net_7759;
wire _net_7761;
wire _net_7763;
wire _net_7765;
wire _net_7768;
wire _net_7781;
wire _net_7782;
wire _net_7783;
wire _net_7784;
wire _net_7785;
wire _net_7786;
wire _net_7787;
wire _net_7788;
wire _net_7789;
wire _net_7791;
wire _net_7793;
wire _net_7794;
wire _net_7795;
wire _net_7796;
wire _net_7797;
wire _net_7798;
wire _net_7800;
wire _net_7801;
wire _net_7803;
wire _net_7804;
wire _net_7805;
wire _net_7806;
wire _net_7808;
wire _net_7809;
wire _net_7810;
wire _net_7811;
wire _net_7812;
wire _net_7813;
wire _net_7814;
wire _net_7815;
wire _net_7816;
wire _net_7817;
wire _net_7818;
wire _net_7819;
wire _net_7820;
wire _net_7821;
wire _net_7822;
wire _net_7823;
wire _net_7824;
wire n1000;
wire n10000;
wire n10001;
wire n10001_1;
wire n10002;
wire n10003;
wire n10004;
wire n10005;
wire n10006;
wire n10006_1;
wire n10007;
wire n10009;
wire n10010;
wire n10010_1;
wire n10012;
wire n10013;
wire n10014;
wire n10014_1;
wire n10015;
wire n10016;
wire n10017;
wire n10018;
wire n10019;
wire n10019_1;
wire n10020;
wire n10021;
wire n10022;
wire n10023;
wire n10024;
wire n10026;
wire n10028;
wire n10028_1;
wire n10029;
wire n10031;
wire n10032;
wire n10032_1;
wire n10034;
wire n10035;
wire n10037;
wire n10037_1;
wire n10038;
wire n10040;
wire n10041;
wire n10042;
wire n10043;
wire n10044;
wire n10045;
wire n10046;
wire n10047;
wire n10047_1;
wire n10048;
wire n10049;
wire n1005;
wire n10050;
wire n10051;
wire n10052;
wire n10052_1;
wire n10053;
wire n10055;
wire n10056;
wire n10056_1;
wire n10057;
wire n10058;
wire n10059;
wire n10060;
wire n10061;
wire n10061_1;
wire n10062;
wire n10063;
wire n10064;
wire n10065;
wire n10066;
wire n10066_1;
wire n10068;
wire n10069;
wire n10070;
wire n10070_1;
wire n10071;
wire n10072;
wire n10074;
wire n10074_1;
wire n10075;
wire n10077;
wire n10078;
wire n10079;
wire n10080;
wire n10081;
wire n10083;
wire n10084;
wire n10084_1;
wire n10086;
wire n10087;
wire n10088;
wire n10089;
wire n10089_1;
wire n10090;
wire n10092;
wire n10093;
wire n10094;
wire n10095;
wire n10097;
wire n10098;
wire n10099;
wire n1010;
wire n10100;
wire n10101;
wire n10103;
wire n10103_1;
wire n10104;
wire n10106;
wire n10107;
wire n10107_1;
wire n10108;
wire n10109;
wire n10110;
wire n10112;
wire n10112_1;
wire n10113;
wire n10115;
wire n10116;
wire n10116_1;
wire n10117;
wire n10119;
wire n10120;
wire n10120_1;
wire n10122;
wire n10123;
wire n10124;
wire n10125;
wire n10126;
wire n10127;
wire n10128;
wire n10128_1;
wire n10129;
wire n10130;
wire n10131;
wire n10132;
wire n10132_1;
wire n10133;
wire n10134;
wire n10135;
wire n10136;
wire n10137;
wire n10137_1;
wire n10138;
wire n10139;
wire n10140;
wire n10141;
wire n10141_1;
wire n10142;
wire n10143;
wire n10145;
wire n10145_1;
wire n10146;
wire n10148;
wire n10149;
wire n1015;
wire n10150;
wire n10151;
wire n10152;
wire n10154;
wire n10154_1;
wire n10155;
wire n10157;
wire n10158;
wire n10158_1;
wire n10160;
wire n10161;
wire n10163;
wire n10164;
wire n10166;
wire n10167;
wire n10169;
wire n10170;
wire n10172;
wire n10174;
wire n10175;
wire n10177;
wire n10178;
wire n10179;
wire n10180;
wire n10181;
wire n10182;
wire n10183;
wire n10184;
wire n10186;
wire n10187;
wire n10188;
wire n10189;
wire n10191;
wire n10192;
wire n10193;
wire n10194;
wire n10195;
wire n10196;
wire n10197;
wire n10198;
wire n10199;
wire n1020;
wire n10200;
wire n10201;
wire n10202;
wire n10203;
wire n10204;
wire n10206;
wire n10207;
wire n10208;
wire n10210;
wire n10211;
wire n10214;
wire n10215;
wire n10217;
wire n10219;
wire n10220;
wire n10222;
wire n10223;
wire n10225;
wire n10226;
wire n10227;
wire n10228;
wire n10229;
wire n10230;
wire n10231;
wire n10232;
wire n10233;
wire n10234;
wire n10235;
wire n10236;
wire n10237;
wire n10239;
wire n1024;
wire n10240;
wire n10242;
wire n10243;
wire n10244;
wire n10245;
wire n10246;
wire n10247;
wire n10248;
wire n10249;
wire n10250;
wire n10251;
wire n10252;
wire n10253;
wire n10254;
wire n10255;
wire n10256;
wire n10257;
wire n10258;
wire n10259;
wire n10260;
wire n10262;
wire n10264;
wire n10266;
wire n10267;
wire n10270;
wire n10271;
wire n10272;
wire n10274;
wire n10275;
wire n10277;
wire n10279;
wire n10280;
wire n10283;
wire n10284;
wire n10286;
wire n10287;
wire n10289;
wire n1029;
wire n10290;
wire n10291;
wire n10292;
wire n10293;
wire n10294;
wire n10295;
wire n10297;
wire n10298;
wire n10299;
wire n10301;
wire n10302;
wire n10303;
wire n10304;
wire n10305;
wire n10306;
wire n10307;
wire n10308;
wire n10309;
wire n10310;
wire n10311;
wire n10312;
wire n10314;
wire n10315;
wire n10317;
wire n10319;
wire n10320;
wire n10322;
wire n10323;
wire n10325;
wire n10326;
wire n10328;
wire n10329;
wire n10331;
wire n10332;
wire n10333;
wire n10334;
wire n10336;
wire n10337;
wire n10338;
wire n10339;
wire n1034;
wire n10340;
wire n10341;
wire n10342;
wire n10343;
wire n10344;
wire n10346;
wire n10348;
wire n10349;
wire n10351;
wire n10352;
wire n10354;
wire n10355;
wire n10357;
wire n10359;
wire n10360;
wire n10362;
wire n10363;
wire n10364;
wire n10365;
wire n10366;
wire n10367;
wire n10369;
wire n10371;
wire n10372;
wire n10374;
wire n10375;
wire n10377;
wire n10378;
wire n10380;
wire n10381;
wire n10382;
wire n10383;
wire n10384;
wire n10385;
wire n10386;
wire n10387;
wire n10388;
wire n10389;
wire n1039;
wire n10390;
wire n10391;
wire n10393;
wire n10394;
wire n10396;
wire n10397;
wire n10398;
wire n10399;
wire n10400;
wire n10401;
wire n10402;
wire n10403;
wire n10404;
wire n10405;
wire n10406;
wire n10407;
wire n10409;
wire n10410;
wire n10412;
wire n10413;
wire n10414;
wire n10415;
wire n10416;
wire n10418;
wire n10419;
wire n10421;
wire n10422;
wire n10423;
wire n10424;
wire n10426;
wire n10427;
wire n10429;
wire n10430;
wire n10431;
wire n10432;
wire n10433;
wire n10434;
wire n10435;
wire n10436;
wire n10437;
wire n10438;
wire n10439;
wire n1044;
wire n10440;
wire n10441;
wire n10442;
wire n10443;
wire n10444;
wire n10445;
wire n10446;
wire n10447;
wire n10448;
wire n10450;
wire n10452;
wire n10453;
wire n10455;
wire n10456;
wire n10458;
wire n10460;
wire n10462;
wire n10463;
wire n10464;
wire n10465;
wire n10466;
wire n10468;
wire n10469;
wire n10471;
wire n10472;
wire n10473;
wire n10474;
wire n10475;
wire n10476;
wire n10477;
wire n10479;
wire n10480;
wire n10482;
wire n10483;
wire n10485;
wire n10486;
wire n10487;
wire n10488;
wire n10489;
wire n1049;
wire n10490;
wire n10491;
wire n10492;
wire n10493;
wire n10494;
wire n10495;
wire n10496;
wire n10497;
wire n10498;
wire n10499;
wire n10500;
wire n10501;
wire n10502;
wire n10503;
wire n10505;
wire n10506;
wire n10508;
wire n10509;
wire n10511;
wire n10512;
wire n10514;
wire n10515;
wire n10517;
wire n10518;
wire n10520;
wire n10521;
wire n10523;
wire n10524;
wire n10525;
wire n10526;
wire n10527;
wire n10528;
wire n10529;
wire n1053;
wire n10530;
wire n10532;
wire n10533;
wire n10534;
wire n10535;
wire n10536;
wire n10537;
wire n10539;
wire n10540;
wire n10541;
wire n10543;
wire n10544;
wire n10546;
wire n10547;
wire n10548;
wire n10549;
wire n10550;
wire n10551;
wire n10552;
wire n10553;
wire n10554;
wire n10555;
wire n10556;
wire n10557;
wire n10558;
wire n10559;
wire n10560;
wire n10561;
wire n10562;
wire n10563;
wire n10564;
wire n10565;
wire n10567;
wire n10568;
wire n10570;
wire n10571;
wire n10573;
wire n10574;
wire n10575;
wire n10576;
wire n10577;
wire n10578;
wire n1058;
wire n10580;
wire n10581;
wire n10583;
wire n10584;
wire n10585;
wire n10586;
wire n10587;
wire n10588;
wire n10589;
wire n10590;
wire n10591;
wire n10592;
wire n10593;
wire n10594;
wire n10595;
wire n10596;
wire n10597;
wire n10598;
wire n10599;
wire n10600;
wire n10601;
wire n10603;
wire n10604;
wire n10606;
wire n10607;
wire n10609;
wire n10610;
wire n10611;
wire n10613;
wire n10614;
wire n10616;
wire n10617;
wire n10619;
wire n1062;
wire n10620;
wire n10621;
wire n10622;
wire n10623;
wire n10624;
wire n10625;
wire n10626;
wire n10627;
wire n10628;
wire n10629;
wire n10630;
wire n10631;
wire n10632;
wire n10633;
wire n10634;
wire n10636;
wire n10637;
wire n10639;
wire n10640;
wire n10642;
wire n10643;
wire n10645;
wire n10646;
wire n10648;
wire n10649;
wire n10651;
wire n10652;
wire n10654;
wire n10655;
wire n10656;
wire n10657;
wire n10658;
wire n10659;
wire n10660;
wire n10661;
wire n10662;
wire n10663;
wire n10664;
wire n10665;
wire n10666;
wire n10667;
wire n10668;
wire n10669;
wire n1067;
wire n10670;
wire n10671;
wire n10672;
wire n10674;
wire n10675;
wire n10677;
wire n10678;
wire n10679;
wire n10680;
wire n10681;
wire n10682;
wire n10683;
wire n10684;
wire n10686;
wire n10687;
wire n10689;
wire n10690;
wire n10691;
wire n10692;
wire n10694;
wire n10695;
wire n10696;
wire n10697;
wire n10698;
wire n10699;
wire n10701;
wire n10702;
wire n10704;
wire n10705;
wire n10706;
wire n10707;
wire n10708;
wire n10709;
wire n10710;
wire n10711;
wire n10712;
wire n10713;
wire n10714;
wire n10715;
wire n10716;
wire n10717;
wire n10719;
wire n1072;
wire n10721;
wire n10722;
wire n10723;
wire n10724;
wire n10725;
wire n10726;
wire n10727;
wire n10728;
wire n10730;
wire n10731;
wire n10733;
wire n10734;
wire n10736;
wire n10737;
wire n10738;
wire n10739;
wire n10740;
wire n10741;
wire n10742;
wire n10743;
wire n10744;
wire n10745;
wire n10746;
wire n10747;
wire n10748;
wire n10749;
wire n10750;
wire n10751;
wire n10752;
wire n10753;
wire n10754;
wire n10755;
wire n10756;
wire n10757;
wire n10758;
wire n10759;
wire n10760;
wire n10761;
wire n10762;
wire n10763;
wire n10765;
wire n10766;
wire n10768;
wire n10769;
wire n1077;
wire n10770;
wire n10771;
wire n10772;
wire n10773;
wire n10774;
wire n10775;
wire n10776;
wire n10777;
wire n10778;
wire n10779;
wire n10781;
wire n10782;
wire n10783;
wire n10784;
wire n10785;
wire n10786;
wire n10787;
wire n10788;
wire n10789;
wire n10790;
wire n10791;
wire n10792;
wire n10794;
wire n10795;
wire n10797;
wire n10798;
wire n10800;
wire n10801;
wire n10803;
wire n10804;
wire n10806;
wire n10807;
wire n1081;
wire n10810;
wire n10811;
wire n10813;
wire n10814;
wire n10816;
wire n10817;
wire n10819;
wire n10820;
wire n10822;
wire n10823;
wire n10824;
wire n10825;
wire n10826;
wire n10827;
wire n10828;
wire n10829;
wire n10830;
wire n10831;
wire n10832;
wire n10833;
wire n10835;
wire n10836;
wire n10838;
wire n10839;
wire n10841;
wire n10842;
wire n10844;
wire n10845;
wire n10847;
wire n10848;
wire n1085;
wire n10850;
wire n10851;
wire n10853;
wire n10854;
wire n10856;
wire n10857;
wire n10858;
wire n10859;
wire n10860;
wire n10861;
wire n10862;
wire n10863;
wire n10864;
wire n10865;
wire n10866;
wire n10867;
wire n10869;
wire n10870;
wire n10872;
wire n10873;
wire n10875;
wire n10877;
wire n10878;
wire n10880;
wire n10881;
wire n10882;
wire n10883;
wire n10884;
wire n10885;
wire n10886;
wire n10887;
wire n10888;
wire n10889;
wire n1089;
wire n10890;
wire n10891;
wire n10893;
wire n10894;
wire n10896;
wire n10897;
wire n10899;
wire n10900;
wire n10902;
wire n10903;
wire n10905;
wire n10906;
wire n10907;
wire n10908;
wire n10909;
wire n10910;
wire n10911;
wire n10912;
wire n10913;
wire n10914;
wire n10915;
wire n10916;
wire n10917;
wire n10920;
wire n10922;
wire n10923;
wire n10925;
wire n10926;
wire n10928;
wire n10929;
wire n1093;
wire n10931;
wire n10933;
wire n10934;
wire n10935;
wire n10936;
wire n10938;
wire n10940;
wire n10941;
wire n10943;
wire n10944;
wire n10945;
wire n10947;
wire n10948;
wire n10949;
wire n10950;
wire n10951;
wire n10952;
wire n10953;
wire n10954;
wire n10955;
wire n10956;
wire n10957;
wire n10958;
wire n10960;
wire n10961;
wire n10963;
wire n10965;
wire n10967;
wire n10969;
wire n1097;
wire n10970;
wire n10972;
wire n10973;
wire n10974;
wire n10977;
wire n10978;
wire n10979;
wire n10980;
wire n10982;
wire n10985;
wire n10987;
wire n10989;
wire n10990;
wire n10992;
wire n10993;
wire n10995;
wire n10996;
wire n10997;
wire n10998;
wire n10999;
wire n11000;
wire n11001;
wire n11002;
wire n11003;
wire n11004;
wire n11005;
wire n11006;
wire n11008;
wire n11009;
wire n11011;
wire n11012;
wire n11014;
wire n11015;
wire n11017;
wire n11018;
wire n1102;
wire n11020;
wire n11021;
wire n11023;
wire n11024;
wire n11026;
wire n11027;
wire n11028;
wire n11029;
wire n11030;
wire n11031;
wire n11034;
wire n11035;
wire n11036;
wire n11037;
wire n11039;
wire n11040;
wire n11042;
wire n11043;
wire n11045;
wire n11047;
wire n11048;
wire n11050;
wire n11051;
wire n11052;
wire n11054;
wire n11055;
wire n11056;
wire n11057;
wire n1106;
wire n11060;
wire n11061;
wire n11063;
wire n11064;
wire n11065;
wire n11066;
wire n11067;
wire n11068;
wire n11069;
wire n11070;
wire n11072;
wire n11073;
wire n11075;
wire n11076;
wire n11078;
wire n11079;
wire n11080;
wire n11081;
wire n11083;
wire n11084;
wire n11086;
wire n11087;
wire n11089;
wire n11090;
wire n11092;
wire n11093;
wire n11095;
wire n11096;
wire n11097;
wire n11099;
wire n11100;
wire n11101;
wire n11103;
wire n11104;
wire n11106;
wire n11108;
wire n11109;
wire n1111;
wire n11111;
wire n11113;
wire n11115;
wire n11116;
wire n11118;
wire n11119;
wire n11120;
wire n11121;
wire n11122;
wire n11123;
wire n11124;
wire n11125;
wire n11126;
wire n11127;
wire n11128;
wire n11129;
wire n11130;
wire n11131;
wire n11133;
wire n11134;
wire n11135;
wire n11136;
wire n11137;
wire n11138;
wire n11139;
wire n11140;
wire n11141;
wire n11142;
wire n11143;
wire n11144;
wire n11146;
wire n11147;
wire n11149;
wire n11150;
wire n11152;
wire n11154;
wire n11155;
wire n11156;
wire n11157;
wire n11158;
wire n11159;
wire n1116;
wire n11161;
wire n11162;
wire n11164;
wire n11165;
wire n11167;
wire n11168;
wire n11169;
wire n11170;
wire n11171;
wire n11172;
wire n11173;
wire n11174;
wire n11177;
wire n11178;
wire n11179;
wire n11181;
wire n11182;
wire n11184;
wire n11185;
wire n11187;
wire n11188;
wire n11189;
wire n11190;
wire n11191;
wire n11192;
wire n11193;
wire n11194;
wire n11196;
wire n11197;
wire n11198;
wire n11199;
wire n11200;
wire n11201;
wire n11202;
wire n11203;
wire n11204;
wire n11205;
wire n11206;
wire n11207;
wire n11209;
wire n1121;
wire n11210;
wire n11211;
wire n11212;
wire n11214;
wire n11215;
wire n11217;
wire n11218;
wire n11219;
wire n11220;
wire n11221;
wire n11222;
wire n11223;
wire n11224;
wire n11225;
wire n11226;
wire n11227;
wire n11229;
wire n11231;
wire n11232;
wire n11234;
wire n11235;
wire n11236;
wire n11237;
wire n11239;
wire n11240;
wire n11243;
wire n11244;
wire n11246;
wire n11247;
wire n11249;
wire n1125;
wire n11250;
wire n11251;
wire n11253;
wire n11254;
wire n11256;
wire n11257;
wire n11258;
wire n11259;
wire n11261;
wire n11262;
wire n11264;
wire n11265;
wire n11267;
wire n11268;
wire n11269;
wire n11271;
wire n11272;
wire n11274;
wire n11275;
wire n11277;
wire n11278;
wire n11279;
wire n11280;
wire n11281;
wire n11282;
wire n11283;
wire n11284;
wire n11285;
wire n11286;
wire n11287;
wire n11288;
wire n11289;
wire n11290;
wire n11291;
wire n11293;
wire n11294;
wire n11296;
wire n11298;
wire n11299;
wire n1130;
wire n11300;
wire n11301;
wire n11302;
wire n11303;
wire n11304;
wire n11305;
wire n11306;
wire n11307;
wire n11308;
wire n11309;
wire n11311;
wire n11312;
wire n11314;
wire n11315;
wire n11317;
wire n11318;
wire n11320;
wire n11321;
wire n11323;
wire n11324;
wire n11325;
wire n11326;
wire n11327;
wire n11328;
wire n11329;
wire n11330;
wire n11331;
wire n11332;
wire n11333;
wire n11334;
wire n11336;
wire n11337;
wire n11339;
wire n11340;
wire n11342;
wire n11343;
wire n11346;
wire n11347;
wire n11349;
wire n1135;
wire n11350;
wire n11352;
wire n11353;
wire n11355;
wire n11356;
wire n11358;
wire n11359;
wire n11360;
wire n11361;
wire n11362;
wire n11363;
wire n11365;
wire n11366;
wire n11367;
wire n11368;
wire n11369;
wire n11370;
wire n11371;
wire n11372;
wire n11373;
wire n11374;
wire n11375;
wire n11376;
wire n11378;
wire n11379;
wire n11380;
wire n11381;
wire n11382;
wire n11383;
wire n11384;
wire n11385;
wire n11386;
wire n11388;
wire n11389;
wire n11392;
wire n11393;
wire n11395;
wire n11396;
wire n11398;
wire n11399;
wire n1140;
wire n11401;
wire n11402;
wire n11404;
wire n11405;
wire n11407;
wire n11408;
wire n11410;
wire n11412;
wire n11413;
wire n11414;
wire n11415;
wire n11416;
wire n11417;
wire n11418;
wire n11419;
wire n11420;
wire n11421;
wire n11422;
wire n11423;
wire n11424;
wire n11425;
wire n11426;
wire n11428;
wire n11429;
wire n11431;
wire n11433;
wire n11434;
wire n11435;
wire n11436;
wire n11438;
wire n1144;
wire n11440;
wire n11441;
wire n11443;
wire n11444;
wire n11445;
wire n11447;
wire n11448;
wire n11450;
wire n11451;
wire n11453;
wire n11454;
wire n11456;
wire n11457;
wire n11458;
wire n11459;
wire n11461;
wire n11462;
wire n11463;
wire n11464;
wire n11465;
wire n11466;
wire n11467;
wire n11468;
wire n11471;
wire n11472;
wire n11474;
wire n11475;
wire n11476;
wire n11477;
wire n11478;
wire n11479;
wire n1148;
wire n11480;
wire n11481;
wire n11482;
wire n11483;
wire n11484;
wire n11485;
wire n11486;
wire n11487;
wire n11488;
wire n11489;
wire n11490;
wire n11491;
wire n11492;
wire n11494;
wire n11495;
wire n11497;
wire n11498;
wire n11499;
wire n11501;
wire n11502;
wire n11504;
wire n11505;
wire n11507;
wire n11508;
wire n11510;
wire n11511;
wire n11513;
wire n11514;
wire n11516;
wire n11517;
wire n11519;
wire n11521;
wire n11523;
wire n11524;
wire n11526;
wire n11527;
wire n11529;
wire n1153;
wire n11530;
wire n11532;
wire n11534;
wire n11536;
wire n11537;
wire n11538;
wire n11539;
wire n11540;
wire n11541;
wire n11542;
wire n11543;
wire n11544;
wire n11545;
wire n11546;
wire n11547;
wire n11548;
wire n11550;
wire n11551;
wire n11553;
wire n11554;
wire n11556;
wire n11558;
wire n11559;
wire n11561;
wire n11562;
wire n11564;
wire n11566;
wire n11567;
wire n11568;
wire n11569;
wire n11570;
wire n11571;
wire n11572;
wire n11573;
wire n11575;
wire n11576;
wire n11578;
wire n11579;
wire n1158;
wire n11580;
wire n11582;
wire n11583;
wire n11584;
wire n11585;
wire n11586;
wire n11588;
wire n11589;
wire n11591;
wire n11592;
wire n11594;
wire n11595;
wire n11597;
wire n11599;
wire n11600;
wire n11602;
wire n11603;
wire n11604;
wire n11605;
wire n11606;
wire n11608;
wire n11609;
wire n11612;
wire n11613;
wire n11615;
wire n11616;
wire n11618;
wire n11619;
wire n11621;
wire n11623;
wire n11624;
wire n11626;
wire n11627;
wire n11629;
wire n1163;
wire n11631;
wire n11633;
wire n11634;
wire n11636;
wire n11637;
wire n11639;
wire n11640;
wire n11642;
wire n11643;
wire n11645;
wire n11646;
wire n11648;
wire n11649;
wire n11651;
wire n11652;
wire n11654;
wire n11656;
wire n11658;
wire n11659;
wire n11660;
wire n11662;
wire n11663;
wire n11664;
wire n11665;
wire n11667;
wire n11668;
wire n11670;
wire n11671;
wire n11673;
wire n11674;
wire n11676;
wire n11677;
wire n11679;
wire n1168;
wire n11681;
wire n11682;
wire n11684;
wire n11686;
wire n11687;
wire n11689;
wire n11690;
wire n11692;
wire n11693;
wire n11695;
wire n11696;
wire n11698;
wire n11700;
wire n11701;
wire n11703;
wire n11704;
wire n11706;
wire n11707;
wire n11708;
wire n11710;
wire n11711;
wire n11713;
wire n11715;
wire n11716;
wire n11717;
wire n11718;
wire n11719;
wire n11720;
wire n11721;
wire n11722;
wire n11723;
wire n11724;
wire n11725;
wire n11726;
wire n11728;
wire n11729;
wire n1173;
wire n11731;
wire n11733;
wire n11734;
wire n11736;
wire n11738;
wire n11739;
wire n11741;
wire n11742;
wire n11743;
wire n11744;
wire n11745;
wire n11746;
wire n11747;
wire n11748;
wire n11749;
wire n11750;
wire n11751;
wire n11752;
wire n11754;
wire n11755;
wire n11757;
wire n11759;
wire n11760;
wire n11763;
wire n11764;
wire n11766;
wire n11767;
wire n11769;
wire n11770;
wire n11772;
wire n11773;
wire n11775;
wire n11776;
wire n11778;
wire n11779;
wire n1178;
wire n11781;
wire n11782;
wire n11783;
wire n11784;
wire n11785;
wire n11786;
wire n11787;
wire n11788;
wire n11790;
wire n11792;
wire n11793;
wire n11794;
wire n11796;
wire n11797;
wire n11799;
wire n11800;
wire n11802;
wire n11803;
wire n11805;
wire n11806;
wire n11808;
wire n11809;
wire n11811;
wire n11812;
wire n11814;
wire n11815;
wire n11816;
wire n11817;
wire n11818;
wire n11819;
wire n11820;
wire n11821;
wire n11822;
wire n11823;
wire n11824;
wire n11825;
wire n11826;
wire n11827;
wire n11828;
wire n11829;
wire n1183;
wire n11830;
wire n11831;
wire n11832;
wire n11833;
wire n11834;
wire n11836;
wire n11837;
wire n11840;
wire n11842;
wire n11843;
wire n11845;
wire n11846;
wire n11847;
wire n11848;
wire n11849;
wire n11850;
wire n11852;
wire n11853;
wire n11855;
wire n11856;
wire n11857;
wire n11858;
wire n11859;
wire n11860;
wire n11862;
wire n11863;
wire n11864;
wire n11865;
wire n11866;
wire n11867;
wire n11868;
wire n11869;
wire n1187;
wire n11870;
wire n11871;
wire n11872;
wire n11873;
wire n11875;
wire n11876;
wire n11878;
wire n11880;
wire n11881;
wire n11883;
wire n11884;
wire n11886;
wire n11887;
wire n11889;
wire n11890;
wire n11892;
wire n11893;
wire n11896;
wire n11897;
wire n11899;
wire n11900;
wire n11901;
wire n11902;
wire n11903;
wire n11904;
wire n11905;
wire n11906;
wire n11908;
wire n1191;
wire n11910;
wire n11911;
wire n11912;
wire n11913;
wire n11914;
wire n11915;
wire n11916;
wire n11917;
wire n11918;
wire n11919;
wire n11920;
wire n11921;
wire n11922;
wire n11923;
wire n11924;
wire n11926;
wire n11927;
wire n11928;
wire n11929;
wire n11930;
wire n11931;
wire n11932;
wire n11933;
wire n11934;
wire n11935;
wire n11936;
wire n11937;
wire n11939;
wire n11940;
wire n11941;
wire n11942;
wire n11943;
wire n11944;
wire n11945;
wire n11947;
wire n11948;
wire n1195;
wire n11950;
wire n11951;
wire n11953;
wire n11954;
wire n11956;
wire n11957;
wire n11959;
wire n11960;
wire n11962;
wire n11964;
wire n11965;
wire n11966;
wire n11967;
wire n11968;
wire n11969;
wire n11970;
wire n11971;
wire n11972;
wire n11974;
wire n11975;
wire n11976;
wire n11978;
wire n11979;
wire n11980;
wire n11981;
wire n11982;
wire n11984;
wire n11985;
wire n11986;
wire n11987;
wire n11989;
wire n11990;
wire n11992;
wire n11993;
wire n11995;
wire n11996;
wire n11997;
wire n11999;
wire n1200;
wire n12000;
wire n12001;
wire n12003;
wire n12004;
wire n12005;
wire n12006;
wire n12008;
wire n12009;
wire n12011;
wire n12012;
wire n12013;
wire n12014;
wire n12015;
wire n12016;
wire n12017;
wire n12018;
wire n12021;
wire n12022;
wire n12024;
wire n12025;
wire n12027;
wire n12028;
wire n12029;
wire n12030;
wire n12031;
wire n12032;
wire n12033;
wire n12034;
wire n12035;
wire n12036;
wire n12037;
wire n12038;
wire n12040;
wire n12042;
wire n12043;
wire n12045;
wire n12047;
wire n12048;
wire n1205;
wire n12050;
wire n12052;
wire n12054;
wire n12055;
wire n12057;
wire n12059;
wire n12060;
wire n12061;
wire n12062;
wire n12063;
wire n12064;
wire n12065;
wire n12066;
wire n12068;
wire n12069;
wire n12071;
wire n12072;
wire n12073;
wire n12074;
wire n12075;
wire n12077;
wire n12078;
wire n12079;
wire n12080;
wire n12082;
wire n12083;
wire n12084;
wire n12085;
wire n12086;
wire n12087;
wire n12088;
wire n12089;
wire n12090;
wire n12091;
wire n12092;
wire n12093;
wire n12094;
wire n12096;
wire n12097;
wire n12099;
wire n1210;
wire n12100;
wire n12102;
wire n12103;
wire n12105;
wire n12106;
wire n12108;
wire n12109;
wire n12110;
wire n12111;
wire n12112;
wire n12113;
wire n12114;
wire n12115;
wire n12116;
wire n12117;
wire n12118;
wire n12119;
wire n12121;
wire n1214;
wire n1219;
wire n1224;
wire n1228;
wire n1232;
wire n1236;
wire n1240;
wire n1244;
wire n1248;
wire n1253;
wire n1258;
wire n1262;
wire n1267;
wire n1272;
wire n1277;
wire n1282;
wire n1287;
wire n1291;
wire n1295;
wire n1300;
wire n1305;
wire n1309;
wire n1314;
wire n1318;
wire n1322;
wire n1326;
wire n1331;
wire n1335;
wire n1340;
wire n1345;
wire n1350;
wire n1355;
wire n1359;
wire n1363;
wire n1368;
wire n1373;
wire n1378;
wire n1383;
wire n1386;
wire n1391;
wire n1396;
wire n1400;
wire n1405;
wire n1410;
wire n1414;
wire n1419;
wire n1423;
wire n1428;
wire n1433;
wire n1438;
wire n1442;
wire n1446;
wire n1451;
wire n1455;
wire n1460;
wire n1465;
wire n1469;
wire n1474;
wire n1478;
wire n1482;
wire n1487;
wire n1491;
wire n1496;
wire n1501;
wire n1506;
wire n1510;
wire n1515;
wire n1519;
wire n1524;
wire n1528;
wire n1533;
wire n1538;
wire n1542;
wire n1546;
wire n1551;
wire n1555;
wire n1560;
wire n1564;
wire n1568;
wire n1572;
wire n1577;
wire n1582;
wire n1587;
wire n1591;
wire n1596;
wire n1600;
wire n1605;
wire n1610;
wire n1615;
wire n1619;
wire n1624;
wire n1629;
wire n1634;
wire n1639;
wire n1644;
wire n1649;
wire n1653;
wire n1658;
wire n1663;
wire n1668;
wire n1673;
wire n1677;
wire n1681;
wire n1686;
wire n1691;
wire n1696;
wire n1701;
wire n1704;
wire n1709;
wire n1714;
wire n1718;
wire n1722;
wire n1727;
wire n1732;
wire n1737;
wire n1742;
wire n1747;
wire n1752;
wire n1756;
wire n1761;
wire n1765;
wire n1770;
wire n1775;
wire n1779;
wire n1782;
wire n1787;
wire n1792;
wire n1797;
wire n1802;
wire n1807;
wire n1812;
wire n1817;
wire n1822;
wire n1827;
wire n1832;
wire n1836;
wire n1841;
wire n1846;
wire n1851;
wire n1855;
wire n1860;
wire n1865;
wire n1869;
wire n1874;
wire n1878;
wire n1883;
wire n1888;
wire n1893;
wire n1898;
wire n1903;
wire n1908;
wire n1913;
wire n1918;
wire n1922;
wire n1927;
wire n1932;
wire n1936;
wire n1941;
wire n1945;
wire n1950;
wire n1954;
wire n1959;
wire n1964;
wire n1969;
wire n1973;
wire n1978;
wire n1983;
wire n1988;
wire n1993;
wire n1998;
wire n2002;
wire n2007;
wire n2011;
wire n2016;
wire n2021;
wire n2026;
wire n2031;
wire n2036;
wire n2041;
wire n2046;
wire n2051;
wire n2055;
wire n2060;
wire n2065;
wire n2070;
wire n2074;
wire n2079;
wire n2084;
wire n2088;
wire n2093;
wire n2098;
wire n2102;
wire n2106;
wire n2111;
wire n2115;
wire n2119;
wire n2122;
wire n2127;
wire n2132;
wire n2136;
wire n2140;
wire n2144;
wire n2149;
wire n2152;
wire n2157;
wire n2162;
wire n2167;
wire n2172;
wire n2177;
wire n2181;
wire n2186;
wire n2189;
wire n2194;
wire n2199;
wire n2203;
wire n2208;
wire n2213;
wire n2218;
wire n2222;
wire n2227;
wire n2232;
wire n2237;
wire n2242;
wire n2247;
wire n2251;
wire n2256;
wire n2260;
wire n2265;
wire n2270;
wire n2275;
wire n2280;
wire n2284;
wire n2288;
wire n2293;
wire n2298;
wire n2303;
wire n2307;
wire n2312;
wire n2316;
wire n2321;
wire n2324;
wire n2329;
wire n2334;
wire n2338;
wire n2342;
wire n2347;
wire n2350;
wire n2355;
wire n2360;
wire n2365;
wire n2370;
wire n2373;
wire n2377;
wire n2381;
wire n2386;
wire n2391;
wire n2395;
wire n2399;
wire n2404;
wire n2409;
wire n2414;
wire n2417;
wire n2422;
wire n2426;
wire n2430;
wire n2435;
wire n2440;
wire n2444;
wire n2448;
wire n2452;
wire n2457;
wire n2462;
wire n2465;
wire n2470;
wire n2474;
wire n2479;
wire n2484;
wire n2488;
wire n2493;
wire n2496;
wire n2500;
wire n2505;
wire n2510;
wire n2515;
wire n2519;
wire n2524;
wire n2529;
wire n2534;
wire n2539;
wire n2543;
wire n2547;
wire n2552;
wire n2556;
wire n2561;
wire n2566;
wire n2570;
wire n2575;
wire n2580;
wire n2585;
wire n2590;
wire n2594;
wire n2597;
wire n2601;
wire n2605;
wire n2610;
wire n2615;
wire n2618;
wire n2622;
wire n2627;
wire n2632;
wire n2637;
wire n2642;
wire n2647;
wire n2651;
wire n2656;
wire n266;
wire n2660;
wire n2665;
wire n2670;
wire n2675;
wire n2679;
wire n2682;
wire n2687;
wire n2692;
wire n2696;
wire n2701;
wire n2705;
wire n2709;
wire n271;
wire n2713;
wire n2718;
wire n2723;
wire n2727;
wire n2732;
wire n2737;
wire n2741;
wire n2745;
wire n2748;
wire n2753;
wire n2758;
wire n276;
wire n2762;
wire n2767;
wire n2771;
wire n2776;
wire n2781;
wire n2784;
wire n2788;
wire n2792;
wire n2797;
wire n2801;
wire n2805;
wire n281;
wire n2810;
wire n2814;
wire n2819;
wire n2823;
wire n2827;
wire n2831;
wire n2836;
wire n2840;
wire n2845;
wire n2850;
wire n2855;
wire n286;
wire n2860;
wire n2864;
wire n2869;
wire n2873;
wire n2877;
wire n2882;
wire n2885;
wire n2890;
wire n2895;
wire n2900;
wire n2904;
wire n2908;
wire n291;
wire n2913;
wire n2918;
wire n2922;
wire n2926;
wire n2930;
wire n2935;
wire n2939;
wire n2944;
wire n2948;
wire n295;
wire n2953;
wire n2958;
wire n2963;
wire n2967;
wire n2972;
wire n2976;
wire n2981;
wire n2986;
wire n2991;
wire n2996;
wire n300;
wire n3000;
wire n3005;
wire n3010;
wire n3015;
wire n3020;
wire n3025;
wire n3030;
wire n3033;
wire n3037;
wire n3042;
wire n3047;
wire n305;
wire n3052;
wire n3056;
wire n3061;
wire n3065;
wire n3069;
wire n3074;
wire n3078;
wire n3082;
wire n3087;
wire n3092;
wire n3097;
wire n310;
wire n3102;
wire n3105;
wire n3110;
wire n3114;
wire n3117;
wire n3121;
wire n3126;
wire n3130;
wire n3134;
wire n3139;
wire n314;
wire n3143;
wire n3148;
wire n3152;
wire n3157;
wire n3162;
wire n3165;
wire n3170;
wire n3174;
wire n3178;
wire n3182;
wire n3186;
wire n319;
wire n3190;
wire n3194;
wire n3199;
wire n3203;
wire n3207;
wire n3212;
wire n3217;
wire n3222;
wire n3226;
wire n3231;
wire n3235;
wire n324;
wire n3240;
wire n3244;
wire n3249;
wire n3254;
wire n3258;
wire n3263;
wire n3268;
wire n3272;
wire n3276;
wire n3280;
wire n3285;
wire n329;
wire n3290;
wire n3294;
wire n3299;
wire n3303;
wire n3308;
wire n3313;
wire n3318;
wire n3322;
wire n3325;
wire n3330;
wire n3333;
wire n3338;
wire n334;
wire n3343;
wire n3348;
wire n3352;
wire n3356;
wire n3361;
wire n3365;
wire n3370;
wire n3374;
wire n3379;
wire n3383;
wire n3386;
wire n339;
wire n3390;
wire n3395;
wire n3400;
wire n3404;
wire n3408;
wire n3413;
wire n3418;
wire n3422;
wire n3427;
wire n3431;
wire n3436;
wire n344;
wire n3440;
wire n3445;
wire n3450;
wire n3455;
wire n3459;
wire n3464;
wire n3469;
wire n3474;
wire n3479;
wire n3484;
wire n3489;
wire n349;
wire n3494;
wire n3497;
wire n3502;
wire n3507;
wire n3511;
wire n3516;
wire n352;
wire n3520;
wire n3524;
wire n3528;
wire n3532;
wire n3537;
wire n3542;
wire n3546;
wire n3551;
wire n3555;
wire n3559;
wire n3564;
wire n3567;
wire n357;
wire n3572;
wire n3577;
wire n3582;
wire n3587;
wire n3590;
wire n3595;
wire n3600;
wire n3604;
wire n3609;
wire n361;
wire n3614;
wire n3618;
wire n3623;
wire n3628;
wire n3633;
wire n3638;
wire n3642;
wire n3647;
wire n3651;
wire n3655;
wire n3658;
wire n366;
wire n3661;
wire n3666;
wire n3670;
wire n3675;
wire n3679;
wire n3684;
wire n3689;
wire n3693;
wire n3698;
wire n370;
wire n3703;
wire n3707;
wire n3711;
wire n3716;
wire n3720;
wire n3725;
wire n3729;
wire n3733;
wire n3737;
wire n3742;
wire n3747;
wire n375;
wire n3752;
wire n3756;
wire n3761;
wire n3765;
wire n3770;
wire n3773;
wire n3777;
wire n3782;
wire n3787;
wire n3791;
wire n3796;
wire n380;
wire n3801;
wire n3805;
wire n3809;
wire n3813;
wire n3817;
wire n3822;
wire n3827;
wire n3831;
wire n3836;
wire n3841;
wire n3846;
wire n385;
wire n3851;
wire n3855;
wire n3859;
wire n3864;
wire n3867;
wire n3872;
wire n3877;
wire n3881;
wire n3886;
wire n3891;
wire n3896;
wire n3899;
wire n390;
wire n3904;
wire n3908;
wire n3913;
wire n3917;
wire n3922;
wire n3927;
wire n3932;
wire n3936;
wire n3941;
wire n3945;
wire n3949;
wire n395;
wire n3953;
wire n3957;
wire n3962;
wire n3967;
wire n3972;
wire n3976;
wire n3981;
wire n3985;
wire n3989;
wire n3993;
wire n3998;
wire n400;
wire n4002;
wire n4007;
wire n4011;
wire n4016;
wire n4020;
wire n4024;
wire n4029;
wire n4033;
wire n4037;
wire n4042;
wire n4046;
wire n405;
wire n4051;
wire n4055;
wire n4059;
wire n4063;
wire n4068;
wire n4071;
wire n4075;
wire n4079;
wire n4084;
wire n4089;
wire n4094;
wire n4098;
wire n410;
wire n4102;
wire n4107;
wire n4112;
wire n4116;
wire n4121;
wire n4126;
wire n4131;
wire n4135;
wire n4140;
wire n4145;
wire n4148;
wire n415;
wire n4153;
wire n4158;
wire n4161;
wire n4166;
wire n4171;
wire n4176;
wire n4181;
wire n4186;
wire n4191;
wire n4194;
wire n4199;
wire n420;
wire n4203;
wire n4207;
wire n4212;
wire n4217;
wire n4221;
wire n4226;
wire n4231;
wire n4235;
wire n424;
wire n4240;
wire n4245;
wire n4249;
wire n4253;
wire n4258;
wire n4263;
wire n4267;
wire n4271;
wire n4276;
wire n4280;
wire n4284;
wire n4289;
wire n429;
wire n4294;
wire n4299;
wire n4304;
wire n4309;
wire n4313;
wire n4318;
wire n4322;
wire n4326;
wire n4330;
wire n4333;
wire n4338;
wire n434;
wire n4343;
wire n4348;
wire n4352;
wire n4357;
wire n4362;
wire n4365;
wire n4370;
wire n4374;
wire n4379;
wire n438;
wire n4384;
wire n4388;
wire n4392;
wire n4397;
wire n4401;
wire n4405;
wire n4410;
wire n4414;
wire n4419;
wire n4424;
wire n4428;
wire n443;
wire n4433;
wire n4438;
wire n4443;
wire n4448;
wire n4451;
wire n4456;
wire n4459;
wire n4464;
wire n4469;
wire n447;
wire n4473;
wire n4478;
wire n4482;
wire n4487;
wire n4491;
wire n4496;
wire n4501;
wire n4505;
wire n451;
wire n4510;
wire n4515;
wire n4520;
wire n4524;
wire n4529;
wire n4534;
wire n4539;
wire n4544;
wire n4548;
wire n455;
wire n4553;
wire n4558;
wire n4562;
wire n4567;
wire n4572;
wire n4577;
wire n4581;
wire n4586;
wire n4591;
wire n4596;
wire n460;
wire n4600;
wire n4604;
wire n4609;
wire n4613;
wire n4617;
wire n4622;
wire n4627;
wire n4631;
wire n4636;
wire n4641;
wire n4646;
wire n465;
wire n4651;
wire n4656;
wire n4660;
wire n4665;
wire n4669;
wire n4673;
wire n4678;
wire n4681;
wire n4686;
wire n4690;
wire n4694;
wire n4699;
wire n470;
wire n4703;
wire n4708;
wire n4713;
wire n4717;
wire n4722;
wire n4727;
wire n4732;
wire n4737;
wire n474;
wire n4742;
wire n4745;
wire n4750;
wire n4755;
wire n4760;
wire n4765;
wire n4769;
wire n4774;
wire n4778;
wire n4782;
wire n4787;
wire n479;
wire n4791;
wire n4795;
wire n4800;
wire n4805;
wire n4809;
wire n4814;
wire n4818;
wire n4822;
wire n4827;
wire n4831;
wire n4834;
wire n4838;
wire n484;
wire n4843;
wire n4848;
wire n4853;
wire n4857;
wire n4862;
wire n4867;
wire n4872;
wire n4877;
wire n488;
wire n4881;
wire n4886;
wire n4890;
wire n4895;
wire n4899;
wire n4904;
wire n4908;
wire n4913;
wire n4917;
wire n4922;
wire n4927;
wire n493;
wire n4931;
wire n4936;
wire n4940;
wire n4944;
wire n4947;
wire n4952;
wire n4957;
wire n4961;
wire n4965;
wire n4969;
wire n4974;
wire n4979;
wire n498;
wire n4983;
wire n4987;
wire n4992;
wire n4996;
wire n5001;
wire n5005;
wire n5008;
wire n5013;
wire n5018;
wire n5023;
wire n5027;
wire n503;
wire n5031;
wire n5035;
wire n5040;
wire n5045;
wire n5048;
wire n5053;
wire n5056;
wire n5061;
wire n5066;
wire n5070;
wire n5075;
wire n508;
wire n5080;
wire n5085;
wire n5090;
wire n5094;
wire n5098;
wire n5103;
wire n5107;
wire n5112;
wire n5117;
wire n5121;
wire n5126;
wire n513;
wire n5130;
wire n5134;
wire n5139;
wire n5143;
wire n5148;
wire n5151;
wire n5156;
wire n5159;
wire n5164;
wire n5169;
wire n5173;
wire n5178;
wire n518;
wire n5181;
wire n5186;
wire n5189;
wire n5193;
wire n5198;
wire n5202;
wire n5207;
wire n5212;
wire n5217;
wire n5221;
wire n5225;
wire n523;
wire n5230;
wire n5234;
wire n5239;
wire n5242;
wire n5246;
wire n5251;
wire n5256;
wire n5261;
wire n5265;
wire n5269;
wire n5274;
wire n5279;
wire n528;
wire n5284;
wire n5288;
wire n5293;
wire n5298;
wire n5302;
wire n5307;
wire n5312;
wire n5316;
wire n5321;
wire n5326;
wire n533;
wire n5330;
wire n5335;
wire n5339;
wire n5344;
wire n5349;
wire n5353;
wire n5358;
wire n5362;
wire n5366;
wire n5370;
wire n5375;
wire n538;
wire n5380;
wire n5383;
wire n5388;
wire n5393;
wire n5397;
wire n5402;
wire n5406;
wire n5411;
wire n5415;
wire n5420;
wire n5424;
wire n5429;
wire n543;
wire n5433;
wire n5437;
wire n5441;
wire n5446;
wire n5451;
wire n5455;
wire n5460;
wire n5464;
wire n5469;
wire n5472;
wire n5477;
wire n548;
wire n5481;
wire n5486;
wire n5490;
wire n5495;
wire n5500;
wire n5504;
wire n5508;
wire n5513;
wire n5517;
wire n5521;
wire n5525;
wire n5529;
wire n553;
wire n5534;
wire n5539;
wire n5543;
wire n5547;
wire n5552;
wire n5556;
wire n556;
wire n5560;
wire n5565;
wire n5570;
wire n5575;
wire n5579;
wire n5584;
wire n5588;
wire n5591;
wire n5596;
wire n5601;
wire n5606;
wire n561;
wire n5610;
wire n5613;
wire n5618;
wire n5623;
wire n5628;
wire n5633;
wire n5638;
wire n5643;
wire n5648;
wire n5651;
wire n5655;
wire n566;
wire n5660;
wire n5664;
wire n5669;
wire n5674;
wire n5679;
wire n5682;
wire n5686;
wire n5691;
wire n5696;
wire n5700;
wire n5704;
wire n5709;
wire n571;
wire n5713;
wire n5717;
wire n5722;
wire n5727;
wire n5731;
wire n5735;
wire n5739;
wire n5744;
wire n5748;
wire n5753;
wire n5758;
wire n576;
wire n5763;
wire n5767;
wire n5771;
wire n5775;
wire n5779;
wire n5783;
wire n5787;
wire n5792;
wire n5796;
wire n580;
wire n5801;
wire n5805;
wire n5809;
wire n5814;
wire n5819;
wire n5824;
wire n5828;
wire n5833;
wire n5836;
wire n5840;
wire n5845;
wire n585;
wire n5850;
wire n5855;
wire n5860;
wire n5864;
wire n5867;
wire n5872;
wire n5876;
wire n5881;
wire n5885;
wire n5890;
wire n5894;
wire n5899;
wire n590;
wire n5903;
wire n5908;
wire n5912;
wire n5917;
wire n5920;
wire n5925;
wire n5930;
wire n5934;
wire n5938;
wire n5943;
wire n5947;
wire n595;
wire n5951;
wire n5955;
wire n5960;
wire n5964;
wire n5968;
wire n5973;
wire n5978;
wire n5982;
wire n5987;
wire n5992;
wire n5997;
wire n600;
wire n6002;
wire n6006;
wire n6009;
wire n6014;
wire n6019;
wire n6024;
wire n6029;
wire n6034;
wire n6038;
wire n6043;
wire n6047;
wire n605;
wire n6052;
wire n6056;
wire n6061;
wire n6066;
wire n6069;
wire n6074;
wire n6078;
wire n6083;
wire n6088;
wire n6093;
wire n6098;
wire n610;
wire n6102;
wire n6106;
wire n6110;
wire n6114;
wire n6119;
wire n6124;
wire n6128;
wire n6132;
wire n6136;
wire n6140;
wire n6145;
wire n6148;
wire n615;
wire n6153;
wire n6158;
wire n6161;
wire n6166;
wire n6171;
wire n6176;
wire n6181;
wire n6186;
wire n6191;
wire n6195;
wire n620;
wire n6200;
wire n6204;
wire n6209;
wire n6214;
wire n6218;
wire n6222;
wire n6227;
wire n6231;
wire n6235;
wire n6239;
wire n6244;
wire n6249;
wire n625;
wire n6254;
wire n6258;
wire n6261;
wire n6266;
wire n6271;
wire n6276;
wire n6281;
wire n6285;
wire n629;
wire n6290;
wire n6294;
wire n6299;
wire n6302;
wire n6306;
wire n6311;
wire n6316;
wire n6319;
wire n6324;
wire n6329;
wire n6332;
wire n6337;
wire n634;
wire n6342;
wire n6346;
wire n6350;
wire n6354;
wire n6357;
wire n6362;
wire n6367;
wire n6371;
wire n6376;
wire n6381;
wire n6386;
wire n639;
wire n6390;
wire n6395;
wire n6399;
wire n6403;
wire n6407;
wire n6411;
wire n6415;
wire n6419;
wire n6423;
wire n6427;
wire n6432;
wire n6437;
wire n644;
wire n6441;
wire n6446;
wire n6450;
wire n6455;
wire n6460;
wire n6464;
wire n6469;
wire n6472;
wire n6477;
wire n6480;
wire n6485;
wire n6489;
wire n649;
wire n6493;
wire n6498;
wire n6502;
wire n6507;
wire n6511;
wire n6515;
wire n6519;
wire n6522;
wire n6527;
wire n6531;
wire n6535;
wire n654;
wire n6540;
wire n6545;
wire n6550;
wire n6554;
wire n6558;
wire n6563;
wire n6566;
wire n6570;
wire n6574;
wire n6578;
wire n6583;
wire n6586;
wire n659;
wire n6591;
wire n6596;
wire n6601;
wire n6606;
wire n6611;
wire n6615;
wire n6619;
wire n6624;
wire n6629;
wire n6634;
wire n6638;
wire n664;
wire n6643;
wire n6648;
wire n6652;
wire n6656;
wire n6661;
wire n6665;
wire n6669;
wire n6674;
wire n6678;
wire n6682;
wire n6687;
wire n669;
wire n6691;
wire n6695;
wire n6700;
wire n6704;
wire n6709;
wire n6713;
wire n6717;
wire n6722;
wire n6727;
wire n673;
wire n6730;
wire n6731;
wire n6732;
wire n6733;
wire n6734;
wire n6735;
wire n6736;
wire n6736_1;
wire n6737;
wire n6738;
wire n6739;
wire n6740;
wire n6741;
wire n6742;
wire n6743;
wire n6745;
wire n6746;
wire n6746_1;
wire n6747;
wire n6748;
wire n6749;
wire n6749_1;
wire n6750;
wire n6751;
wire n6752;
wire n6752_1;
wire n6753;
wire n6754;
wire n6755;
wire n6756;
wire n6756_1;
wire n6757;
wire n6758;
wire n6759;
wire n6760;
wire n6761;
wire n6761_1;
wire n6762;
wire n6763;
wire n6764;
wire n6765;
wire n6765_1;
wire n6766;
wire n6767;
wire n6768;
wire n6769;
wire n6770;
wire n6770_1;
wire n6771;
wire n6772;
wire n6773;
wire n6774;
wire n6774_1;
wire n6775;
wire n6776;
wire n6777;
wire n6778;
wire n6779;
wire n6779_1;
wire n678;
wire n6780;
wire n6781;
wire n6782;
wire n6783;
wire n6783_1;
wire n6784;
wire n6785;
wire n6786;
wire n6787;
wire n6788;
wire n6788_1;
wire n6789;
wire n6790;
wire n6791;
wire n6792;
wire n6793;
wire n6793_1;
wire n6794;
wire n6795;
wire n6796;
wire n6796_1;
wire n6797;
wire n6799;
wire n6800;
wire n6801;
wire n6801_1;
wire n6802;
wire n6803;
wire n6804;
wire n6806;
wire n6806_1;
wire n6807;
wire n6808;
wire n6809;
wire n6809_1;
wire n6810;
wire n6811;
wire n6812;
wire n6813;
wire n6813_1;
wire n6814;
wire n6815;
wire n6816;
wire n6817;
wire n6818;
wire n6818_1;
wire n6819;
wire n6820;
wire n6821;
wire n6822;
wire n6822_1;
wire n6823;
wire n6824;
wire n6825;
wire n6826;
wire n6826_1;
wire n6827;
wire n6828;
wire n6829;
wire n683;
wire n6830;
wire n6831;
wire n6831_1;
wire n6832;
wire n6833;
wire n6834;
wire n6835;
wire n6836;
wire n6836_1;
wire n6837;
wire n6838;
wire n6839;
wire n6840;
wire n6840_1;
wire n6841;
wire n6842;
wire n6843;
wire n6844;
wire n6845;
wire n6845_1;
wire n6846;
wire n6847;
wire n6848;
wire n6849;
wire n6850;
wire n6850_1;
wire n6851;
wire n6852;
wire n6853;
wire n6854;
wire n6855;
wire n6855_1;
wire n6856;
wire n6857;
wire n6859;
wire n6860;
wire n6860_1;
wire n6861;
wire n6862;
wire n6863;
wire n6863_1;
wire n6864;
wire n6865;
wire n6866;
wire n6867;
wire n6867_1;
wire n6868;
wire n6869;
wire n6870;
wire n6871;
wire n6872;
wire n6872_1;
wire n6873;
wire n6875;
wire n6876;
wire n6876_1;
wire n6877;
wire n6878;
wire n6879;
wire n688;
wire n6880;
wire n6881;
wire n6881_1;
wire n6882;
wire n6884;
wire n6885;
wire n6886;
wire n6886_1;
wire n6888;
wire n6889;
wire n6890;
wire n6890_1;
wire n6891;
wire n6892;
wire n6894;
wire n6895;
wire n6895_1;
wire n6896;
wire n6897;
wire n6898;
wire n6899;
wire n6899_1;
wire n6900;
wire n6901;
wire n6902;
wire n6902_1;
wire n6903;
wire n6904;
wire n6905;
wire n6906;
wire n6907;
wire n6908;
wire n6910;
wire n6910_1;
wire n6912;
wire n6913;
wire n6914;
wire n6915;
wire n6915_1;
wire n6916;
wire n6917;
wire n6918;
wire n6919;
wire n6919_1;
wire n6920;
wire n6921;
wire n6922;
wire n6923;
wire n6924;
wire n6924_1;
wire n6925;
wire n6926;
wire n6927;
wire n6928;
wire n6929;
wire n6929_1;
wire n693;
wire n6930;
wire n6931;
wire n6932;
wire n6933;
wire n6934;
wire n6934_1;
wire n6935;
wire n6936;
wire n6937;
wire n6938;
wire n6938_1;
wire n6939;
wire n6940;
wire n6941;
wire n6942;
wire n6943;
wire n6943_1;
wire n6944;
wire n6945;
wire n6946;
wire n6947;
wire n6947_1;
wire n6948;
wire n6949;
wire n6950;
wire n6951;
wire n6952;
wire n6952_1;
wire n6953;
wire n6954;
wire n6955;
wire n6956;
wire n6957;
wire n6958;
wire n6959;
wire n6960;
wire n6960_1;
wire n6961;
wire n6962;
wire n6963;
wire n6964;
wire n6964_1;
wire n6965;
wire n6966;
wire n6967;
wire n6968;
wire n6969;
wire n6969_1;
wire n6970;
wire n6971;
wire n6972;
wire n6974;
wire n6974_1;
wire n6976;
wire n6977;
wire n6977_1;
wire n6978;
wire n6979;
wire n698;
wire n6980;
wire n6981;
wire n6982;
wire n6982_1;
wire n6983;
wire n6984;
wire n6985;
wire n6986;
wire n6986_1;
wire n6987;
wire n6988;
wire n6989;
wire n6990;
wire n6990_1;
wire n6991;
wire n6992;
wire n6993;
wire n6994;
wire n6995;
wire n6995_1;
wire n6996;
wire n6997;
wire n6998;
wire n6999;
wire n7000;
wire n7000_1;
wire n7001;
wire n7002;
wire n7003;
wire n7004;
wire n7005;
wire n7005_1;
wire n7006;
wire n7007;
wire n7008;
wire n7009;
wire n7009_1;
wire n7010;
wire n7011;
wire n7012;
wire n7013;
wire n7013_1;
wire n7014;
wire n7015;
wire n7016;
wire n7017;
wire n7018;
wire n7018_1;
wire n7019;
wire n7020;
wire n7021;
wire n7022;
wire n7023;
wire n7023_1;
wire n7025;
wire n7026;
wire n7027;
wire n7027_1;
wire n7028;
wire n7029;
wire n703;
wire n7030;
wire n7031;
wire n7032;
wire n7032_1;
wire n7033;
wire n7034;
wire n7036;
wire n7036_1;
wire n7037;
wire n7038;
wire n7039;
wire n7040;
wire n7041;
wire n7041_1;
wire n7042;
wire n7043;
wire n7044;
wire n7045;
wire n7045_1;
wire n7046;
wire n7047;
wire n7048;
wire n7049;
wire n7049_1;
wire n7050;
wire n7051;
wire n7052;
wire n7053;
wire n7053_1;
wire n7054;
wire n7055;
wire n7056;
wire n7057;
wire n7058;
wire n7058_1;
wire n7059;
wire n7060;
wire n7061;
wire n7062;
wire n7062_1;
wire n7063;
wire n7064;
wire n7065;
wire n7067;
wire n7067_1;
wire n7069;
wire n7071;
wire n7072;
wire n7072_1;
wire n7073;
wire n7074;
wire n7075;
wire n7076;
wire n7077;
wire n7077_1;
wire n7078;
wire n7079;
wire n708;
wire n7080;
wire n7081;
wire n7082;
wire n7082_1;
wire n7083;
wire n7084;
wire n7085;
wire n7085_1;
wire n7086;
wire n7087;
wire n7088;
wire n7089;
wire n7089_1;
wire n7090;
wire n7091;
wire n7092;
wire n7093;
wire n7093_1;
wire n7094;
wire n7095;
wire n7096;
wire n7097;
wire n7098;
wire n7098_1;
wire n7099;
wire n7100;
wire n7101;
wire n7102;
wire n7102_1;
wire n7103;
wire n7105;
wire n7106;
wire n7107;
wire n7107_1;
wire n7108;
wire n7109;
wire n7110;
wire n7111;
wire n7111_1;
wire n7112;
wire n7113;
wire n7114;
wire n7116;
wire n7116_1;
wire n7117;
wire n7118;
wire n7119;
wire n7120;
wire n7120_1;
wire n7121;
wire n7122;
wire n7123;
wire n7124;
wire n7125;
wire n7125_1;
wire n7126;
wire n7127;
wire n7128;
wire n7128_1;
wire n7129;
wire n713;
wire n7130;
wire n7131;
wire n7132;
wire n7133;
wire n7133_1;
wire n7134;
wire n7135;
wire n7136;
wire n7137;
wire n7138;
wire n7138_1;
wire n7140;
wire n7141;
wire n7142;
wire n7142_1;
wire n7143;
wire n7144;
wire n7145;
wire n7147;
wire n7147_1;
wire n7148;
wire n7149;
wire n7150;
wire n7151;
wire n7151_1;
wire n7153;
wire n7154;
wire n7155;
wire n7155_1;
wire n7156;
wire n7158;
wire n7159;
wire n7160;
wire n7160_1;
wire n7161;
wire n7162;
wire n7163;
wire n7164;
wire n7164_1;
wire n7165;
wire n7166;
wire n7167;
wire n7167_1;
wire n7168;
wire n7169;
wire n7171;
wire n7172;
wire n7173;
wire n7175;
wire n7177;
wire n7177_1;
wire n7178;
wire n7179;
wire n718;
wire n7180;
wire n7181;
wire n7182;
wire n7182_1;
wire n7183;
wire n7184;
wire n7185;
wire n7186;
wire n7188;
wire n7190;
wire n7190_1;
wire n7191;
wire n7193;
wire n7194;
wire n7194_1;
wire n7195;
wire n7196;
wire n7197;
wire n7198;
wire n7199;
wire n7199_1;
wire n7200;
wire n7201;
wire n7203;
wire n7203_1;
wire n7205;
wire n7206;
wire n7207;
wire n7207_1;
wire n7208;
wire n7210;
wire n7211;
wire n7212;
wire n7212_1;
wire n7213;
wire n7214;
wire n7215;
wire n7216;
wire n7216_1;
wire n7217;
wire n7218;
wire n7219;
wire n722;
wire n7220;
wire n7221;
wire n7221_1;
wire n7223;
wire n7224;
wire n7225;
wire n7226;
wire n7226_1;
wire n7227;
wire n7228;
wire n7229;
wire n7230;
wire n7230_1;
wire n7232;
wire n7234;
wire n7235;
wire n7235_1;
wire n7237;
wire n7239;
wire n7240;
wire n7240_1;
wire n7241;
wire n7242;
wire n7243;
wire n7245;
wire n7245_1;
wire n7246;
wire n7248;
wire n7249;
wire n7250;
wire n7252;
wire n7252_1;
wire n7253;
wire n7254;
wire n7255;
wire n7256;
wire n7256_1;
wire n7257;
wire n7259;
wire n7260;
wire n7260_1;
wire n7261;
wire n7262;
wire n7263;
wire n7264;
wire n7265;
wire n7265_1;
wire n7266;
wire n7267;
wire n7268;
wire n7269;
wire n727;
wire n7270;
wire n7270_1;
wire n7271;
wire n7272;
wire n7273;
wire n7274;
wire n7275;
wire n7276;
wire n7278;
wire n7279;
wire n7280;
wire n7281;
wire n7282;
wire n7283;
wire n7284;
wire n7284_1;
wire n7285;
wire n7286;
wire n7287;
wire n7288;
wire n7288_1;
wire n7289;
wire n7290;
wire n7291;
wire n7292;
wire n7292_1;
wire n7293;
wire n7294;
wire n7295;
wire n7296;
wire n7297;
wire n7297_1;
wire n7298;
wire n7299;
wire n7300;
wire n7301;
wire n7302;
wire n7302_1;
wire n7303;
wire n7304;
wire n7305;
wire n7306;
wire n7307;
wire n7307_1;
wire n7308;
wire n7309;
wire n7310;
wire n7311;
wire n7312;
wire n7312_1;
wire n7313;
wire n7315;
wire n7316;
wire n7316_1;
wire n7318;
wire n7319;
wire n732;
wire n7321;
wire n7321_1;
wire n7322;
wire n7323;
wire n7324;
wire n7325;
wire n7326;
wire n7326_1;
wire n7327;
wire n7328;
wire n7330;
wire n7330_1;
wire n7331;
wire n7332;
wire n7334;
wire n7335;
wire n7335_1;
wire n7336;
wire n7337;
wire n7338;
wire n7339;
wire n7340;
wire n7340_1;
wire n7341;
wire n7342;
wire n7343;
wire n7344;
wire n7345;
wire n7346;
wire n7347;
wire n7348;
wire n7349;
wire n7349_1;
wire n7351;
wire n7353;
wire n7354;
wire n7354_1;
wire n7355;
wire n7356;
wire n7357;
wire n7358;
wire n7359;
wire n7359_1;
wire n736;
wire n7360;
wire n7361;
wire n7362;
wire n7363;
wire n7363_1;
wire n7365;
wire n7366;
wire n7368;
wire n7368_1;
wire n7369;
wire n7371;
wire n7372;
wire n7372_1;
wire n7374;
wire n7375;
wire n7376;
wire n7377;
wire n7378;
wire n7381;
wire n7381_1;
wire n7382;
wire n7384;
wire n7385;
wire n7386;
wire n7386_1;
wire n7387;
wire n7388;
wire n7390;
wire n7391;
wire n7391_1;
wire n7392;
wire n7393;
wire n7394;
wire n7395;
wire n7396;
wire n7397;
wire n7398;
wire n7399;
wire n7400;
wire n7400_1;
wire n7401;
wire n7402;
wire n7403;
wire n7404;
wire n7404_1;
wire n7406;
wire n7407;
wire n7408;
wire n7408_1;
wire n7409;
wire n741;
wire n7410;
wire n7411;
wire n7412;
wire n7413;
wire n7413_1;
wire n7414;
wire n7415;
wire n7416;
wire n7417;
wire n7417_1;
wire n7418;
wire n7419;
wire n7420;
wire n7421;
wire n7422;
wire n7422_1;
wire n7423;
wire n7425;
wire n7426;
wire n7427;
wire n7427_1;
wire n7428;
wire n7429;
wire n7431;
wire n7432;
wire n7432_1;
wire n7434;
wire n7435;
wire n7436;
wire n7437;
wire n7437_1;
wire n7438;
wire n7440;
wire n7441;
wire n7442;
wire n7443;
wire n7444;
wire n7445;
wire n7446;
wire n7446_1;
wire n7447;
wire n7448;
wire n7449;
wire n7450;
wire n7450_1;
wire n7452;
wire n7453;
wire n7454;
wire n7454_1;
wire n7456;
wire n7457;
wire n7459;
wire n7459_1;
wire n746;
wire n7460;
wire n7461;
wire n7462;
wire n7463;
wire n7463_1;
wire n7464;
wire n7465;
wire n7466;
wire n7467;
wire n7468;
wire n7468_1;
wire n7469;
wire n7470;
wire n7471;
wire n7472;
wire n7473;
wire n7473_1;
wire n7474;
wire n7475;
wire n7476;
wire n7477;
wire n7478;
wire n7478_1;
wire n7479;
wire n7480;
wire n7481;
wire n7482;
wire n7482_1;
wire n7483;
wire n7484;
wire n7485;
wire n7486;
wire n7487;
wire n7487_1;
wire n7488;
wire n7489;
wire n7490;
wire n7491;
wire n7492;
wire n7492_1;
wire n7493;
wire n7494;
wire n7495;
wire n7496;
wire n7496_1;
wire n7497;
wire n7498;
wire n7499;
wire n7501;
wire n7501_1;
wire n7502;
wire n7503;
wire n7504;
wire n7505;
wire n7505_1;
wire n7507;
wire n7509;
wire n7509_1;
wire n751;
wire n7511;
wire n7513;
wire n7513_1;
wire n7514;
wire n7516;
wire n7518;
wire n7518_1;
wire n7519;
wire n7520;
wire n7522;
wire n7522_1;
wire n7524;
wire n7525;
wire n7526;
wire n7527;
wire n7527_1;
wire n7528;
wire n7529;
wire n7530;
wire n7530_1;
wire n7531;
wire n7533;
wire n7534;
wire n7535;
wire n7535_1;
wire n7536;
wire n7537;
wire n7538;
wire n7539;
wire n7539_1;
wire n7540;
wire n7541;
wire n7542;
wire n7543;
wire n7543_1;
wire n7544;
wire n7545;
wire n7547;
wire n7548;
wire n7549;
wire n7550;
wire n7551;
wire n7552;
wire n7553;
wire n7553_1;
wire n7554;
wire n7556;
wire n7557;
wire n7558;
wire n7559;
wire n756;
wire n7560;
wire n7562;
wire n7563;
wire n7564;
wire n7565;
wire n7566;
wire n7567;
wire n7567_1;
wire n7568;
wire n7570;
wire n7571;
wire n7572;
wire n7572_1;
wire n7573;
wire n7574;
wire n7575;
wire n7576;
wire n7577;
wire n7577_1;
wire n7578;
wire n7579;
wire n7580;
wire n7581;
wire n7581_1;
wire n7582;
wire n7583;
wire n7584;
wire n7585;
wire n7586;
wire n7586_1;
wire n7587;
wire n7588;
wire n7589;
wire n7590;
wire n7591;
wire n7591_1;
wire n7592;
wire n7593;
wire n7594;
wire n7595;
wire n7596;
wire n7596_1;
wire n7597;
wire n7599;
wire n7599_1;
wire n7601;
wire n7603;
wire n7604;
wire n7604_1;
wire n7605;
wire n7606;
wire n7607;
wire n7608;
wire n7608_1;
wire n7609;
wire n761;
wire n7610;
wire n7611;
wire n7612;
wire n7613;
wire n7613_1;
wire n7614;
wire n7615;
wire n7616;
wire n7617;
wire n7618;
wire n7618_1;
wire n7619;
wire n7620;
wire n7621;
wire n7622;
wire n7623;
wire n7624;
wire n7625;
wire n7626;
wire n7626_1;
wire n7627;
wire n7629;
wire n7630;
wire n7631;
wire n7632;
wire n7633;
wire n7635;
wire n7635_1;
wire n7636;
wire n7637;
wire n7638;
wire n7639;
wire n7640;
wire n7641;
wire n7642;
wire n7643;
wire n7644;
wire n7644_1;
wire n7645;
wire n7647;
wire n7648;
wire n7649;
wire n765;
wire n7650;
wire n7652;
wire n7653;
wire n7654;
wire n7654_1;
wire n7656;
wire n7657;
wire n7658;
wire n7658_1;
wire n7659;
wire n7660;
wire n7661;
wire n7662;
wire n7663;
wire n7664;
wire n7665;
wire n7666;
wire n7666_1;
wire n7667;
wire n7668;
wire n7669;
wire n7670;
wire n7671;
wire n7671_1;
wire n7673;
wire n7674;
wire n7676;
wire n7676_1;
wire n7677;
wire n7679;
wire n7680;
wire n7681;
wire n7682;
wire n7684;
wire n7685;
wire n7686;
wire n7687;
wire n7688;
wire n7689;
wire n7690;
wire n7691;
wire n7691_1;
wire n7692;
wire n7693;
wire n7694;
wire n7695;
wire n7695_1;
wire n7696;
wire n7697;
wire n7698;
wire n7699;
wire n770;
wire n7700;
wire n7701;
wire n7702;
wire n7704;
wire n7704_1;
wire n7705;
wire n7706;
wire n7707;
wire n7708;
wire n7709;
wire n7710;
wire n7712;
wire n7713;
wire n7714;
wire n7714_1;
wire n7715;
wire n7716;
wire n7717;
wire n7718;
wire n7719;
wire n7719_1;
wire n7720;
wire n7721;
wire n7722;
wire n7723;
wire n7723_1;
wire n7724;
wire n7725;
wire n7726;
wire n7727;
wire n7728;
wire n7728_1;
wire n7729;
wire n7730;
wire n7731;
wire n7732;
wire n7732_1;
wire n7733;
wire n7734;
wire n7735;
wire n7736;
wire n7737;
wire n7737_1;
wire n7738;
wire n7739;
wire n774;
wire n7740;
wire n7741;
wire n7741_1;
wire n7742;
wire n7743;
wire n7744;
wire n7745;
wire n7746;
wire n7746_1;
wire n7747;
wire n7749;
wire n7750;
wire n7751;
wire n7751_1;
wire n7752;
wire n7753;
wire n7754;
wire n7755;
wire n7756;
wire n7756_1;
wire n7757;
wire n7758;
wire n7759;
wire n7760;
wire n7760_1;
wire n7761;
wire n7762;
wire n7763;
wire n7764;
wire n7764_1;
wire n7765;
wire n7766;
wire n7767;
wire n7768;
wire n7768_1;
wire n7769;
wire n7770;
wire n7771;
wire n7773;
wire n7773_1;
wire n7774;
wire n7776;
wire n7776_1;
wire n7777;
wire n7778;
wire n7779;
wire n7779_1;
wire n7780;
wire n7782;
wire n7784;
wire n7784_1;
wire n7785;
wire n7787;
wire n7788;
wire n7788_1;
wire n779;
wire n7790;
wire n7791;
wire n7793;
wire n7793_1;
wire n7794;
wire n7796;
wire n7797;
wire n7798;
wire n7799;
wire n7800;
wire n7801;
wire n7802;
wire n7802_1;
wire n7803;
wire n7804;
wire n7805;
wire n7806;
wire n7806_1;
wire n7807;
wire n7808;
wire n7809;
wire n7810;
wire n7810_1;
wire n7811;
wire n7812;
wire n7813;
wire n7814;
wire n7815;
wire n7815_1;
wire n7816;
wire n7817;
wire n7818;
wire n7818_1;
wire n7819;
wire n7820;
wire n7821;
wire n7822;
wire n7822_1;
wire n7823;
wire n7824;
wire n7825;
wire n7826;
wire n7826_1;
wire n7827;
wire n7828;
wire n7829;
wire n783;
wire n7830;
wire n7831;
wire n7831_1;
wire n7833;
wire n7834;
wire n7835;
wire n7836;
wire n7837;
wire n7838;
wire n7839;
wire n7840;
wire n7840_1;
wire n7841;
wire n7842;
wire n7844;
wire n7845;
wire n7845_1;
wire n7846;
wire n7847;
wire n7848;
wire n7848_1;
wire n7849;
wire n7850;
wire n7851;
wire n7852;
wire n7853;
wire n7853_1;
wire n7854;
wire n7855;
wire n7857;
wire n7858;
wire n7858_1;
wire n7859;
wire n7860;
wire n7861;
wire n7863;
wire n7863_1;
wire n7864;
wire n7866;
wire n7867;
wire n7867_1;
wire n7868;
wire n7869;
wire n7870;
wire n7871;
wire n7871_1;
wire n7872;
wire n7873;
wire n7874;
wire n7875;
wire n7877;
wire n7878;
wire n7878_1;
wire n788;
wire n7880;
wire n7881;
wire n7882;
wire n7883;
wire n7883_1;
wire n7884;
wire n7886;
wire n7887;
wire n7888;
wire n7889;
wire n7890;
wire n7891;
wire n7892;
wire n7893;
wire n7893_1;
wire n7895;
wire n7897;
wire n7897_1;
wire n7898;
wire n7900;
wire n7901;
wire n7902;
wire n7903;
wire n7904;
wire n7906;
wire n7906_1;
wire n7907;
wire n7908;
wire n7909;
wire n7910;
wire n7911;
wire n7911_1;
wire n7912;
wire n7913;
wire n7914;
wire n7915;
wire n7916;
wire n7916_1;
wire n7917;
wire n7918;
wire n7919;
wire n7920;
wire n7920_1;
wire n7921;
wire n7923;
wire n7924;
wire n7924_1;
wire n7925;
wire n7926;
wire n7927;
wire n7929;
wire n7929_1;
wire n793;
wire n7930;
wire n7931;
wire n7932;
wire n7933;
wire n7933_1;
wire n7934;
wire n7935;
wire n7936;
wire n7937;
wire n7937_1;
wire n7938;
wire n7939;
wire n7940;
wire n7941;
wire n7942;
wire n7942_1;
wire n7943;
wire n7944;
wire n7945;
wire n7945_1;
wire n7946;
wire n7947;
wire n7949;
wire n7950;
wire n7950_1;
wire n7951;
wire n7952;
wire n7953;
wire n7955;
wire n7955_1;
wire n7956;
wire n7958;
wire n7958_1;
wire n7959;
wire n7960;
wire n7961;
wire n7962;
wire n7962_1;
wire n7963;
wire n7964;
wire n7965;
wire n7966;
wire n7967;
wire n7967_1;
wire n7968;
wire n7969;
wire n7970;
wire n7970_1;
wire n7971;
wire n7972;
wire n7973;
wire n7974;
wire n7975;
wire n7975_1;
wire n7976;
wire n7978;
wire n798;
wire n7980;
wire n7980_1;
wire n7981;
wire n7983;
wire n7985;
wire n7986;
wire n7988;
wire n7989;
wire n7989_1;
wire n7991;
wire n7992;
wire n7993;
wire n7994;
wire n7994_1;
wire n7995;
wire n7997;
wire n7997_1;
wire n7998;
wire n7999;
wire n8000;
wire n8001;
wire n8002;
wire n8003;
wire n8004;
wire n8005;
wire n8005_1;
wire n8006;
wire n8007;
wire n8008;
wire n8009;
wire n8010;
wire n8010_1;
wire n8012;
wire n8014;
wire n8015;
wire n8016;
wire n8017;
wire n8019;
wire n8019_1;
wire n802;
wire n8020;
wire n8021;
wire n8022;
wire n8023;
wire n8024;
wire n8025;
wire n8026;
wire n8028;
wire n8028_1;
wire n8029;
wire n8030;
wire n8031;
wire n8032;
wire n8033;
wire n8033_1;
wire n8034;
wire n8035;
wire n8036;
wire n8037;
wire n8038;
wire n8038_1;
wire n8040;
wire n8041;
wire n8042;
wire n8042_1;
wire n8043;
wire n8044;
wire n8046;
wire n8047;
wire n8047_1;
wire n8048;
wire n8049;
wire n8050;
wire n8051;
wire n8051_1;
wire n8052;
wire n8053;
wire n8054;
wire n8055;
wire n8056;
wire n8056_1;
wire n8057;
wire n8058;
wire n8059;
wire n8059_1;
wire n806;
wire n8060;
wire n8061;
wire n8062;
wire n8063;
wire n8064;
wire n8064_1;
wire n8065;
wire n8066;
wire n8067;
wire n8067_1;
wire n8068;
wire n8069;
wire n8070;
wire n8071;
wire n8072;
wire n8072_1;
wire n8073;
wire n8074;
wire n8075;
wire n8075_1;
wire n8076;
wire n8077;
wire n8078;
wire n8079;
wire n8080;
wire n8080_1;
wire n8081;
wire n8082;
wire n8084;
wire n8085;
wire n8085_1;
wire n8086;
wire n8087;
wire n8088;
wire n8088_1;
wire n8089;
wire n8090;
wire n8092;
wire n8092_1;
wire n8093;
wire n8094;
wire n8096;
wire n8097;
wire n8097_1;
wire n8099;
wire n8100;
wire n8101;
wire n8102;
wire n8102_1;
wire n8103;
wire n8104;
wire n8105;
wire n8106;
wire n8107;
wire n8107_1;
wire n8108;
wire n8109;
wire n811;
wire n8110;
wire n8111;
wire n8112;
wire n8112_1;
wire n8113;
wire n8114;
wire n8115;
wire n8116;
wire n8116_1;
wire n8117;
wire n8119;
wire n8120;
wire n8121;
wire n8121_1;
wire n8122;
wire n8123;
wire n8124;
wire n8125;
wire n8125_1;
wire n8126;
wire n8127;
wire n8128;
wire n8129;
wire n8130;
wire n8130_1;
wire n8131;
wire n8132;
wire n8133;
wire n8135;
wire n8135_1;
wire n8136;
wire n8138;
wire n8139;
wire n8140;
wire n8140_1;
wire n8141;
wire n8142;
wire n8144;
wire n8144_1;
wire n8145;
wire n8146;
wire n8147;
wire n8147_1;
wire n8149;
wire n815;
wire n8150;
wire n8152;
wire n8152_1;
wire n8153;
wire n8155;
wire n8156;
wire n8156_1;
wire n8157;
wire n8158;
wire n8159;
wire n8160;
wire n8161;
wire n8161_1;
wire n8162;
wire n8163;
wire n8164;
wire n8165;
wire n8166;
wire n8166_1;
wire n8167;
wire n8168;
wire n8170;
wire n8170_1;
wire n8172;
wire n8173;
wire n8174;
wire n8175;
wire n8177;
wire n8178;
wire n8179;
wire n8179_1;
wire n8181;
wire n8182;
wire n8183;
wire n8183_1;
wire n8184;
wire n8185;
wire n8186;
wire n8187;
wire n8188;
wire n8188_1;
wire n8190;
wire n8191;
wire n8192;
wire n8192_1;
wire n8193;
wire n8194;
wire n8196;
wire n8197;
wire n8197_1;
wire n8198;
wire n8199;
wire n820;
wire n8200;
wire n8202;
wire n8202_1;
wire n8203;
wire n8205;
wire n8206;
wire n8206_1;
wire n8207;
wire n8208;
wire n8209;
wire n8211;
wire n8211_1;
wire n8212;
wire n8213;
wire n8214;
wire n8215;
wire n8216;
wire n8216_1;
wire n8217;
wire n8219;
wire n8220;
wire n8220_1;
wire n8221;
wire n8222;
wire n8223;
wire n8224;
wire n8224_1;
wire n8226;
wire n8227;
wire n8228;
wire n8229;
wire n8231;
wire n8232;
wire n8232_1;
wire n8233;
wire n8234;
wire n8235;
wire n8236;
wire n8237;
wire n8237_1;
wire n8238;
wire n8240;
wire n8241;
wire n8241_1;
wire n8243;
wire n8244;
wire n8245;
wire n8245_1;
wire n8246;
wire n8247;
wire n8249;
wire n8249_1;
wire n825;
wire n8250;
wire n8251;
wire n8252;
wire n8253;
wire n8253_1;
wire n8254;
wire n8255;
wire n8256;
wire n8258;
wire n8258_1;
wire n8259;
wire n8260;
wire n8261;
wire n8262;
wire n8262_1;
wire n8263;
wire n8264;
wire n8265;
wire n8266;
wire n8268;
wire n8269;
wire n8270;
wire n8271;
wire n8271_1;
wire n8272;
wire n8273;
wire n8274;
wire n8275;
wire n8276;
wire n8276_1;
wire n8277;
wire n8278;
wire n8279;
wire n8280;
wire n8280_1;
wire n8281;
wire n8282;
wire n8283;
wire n8284;
wire n8284_1;
wire n8285;
wire n8286;
wire n8287;
wire n8288;
wire n8289;
wire n8289_1;
wire n8290;
wire n8291;
wire n8292;
wire n8293;
wire n8294;
wire n8294_1;
wire n8295;
wire n8296;
wire n8297;
wire n8298;
wire n8299;
wire n8299_1;
wire n830;
wire n8300;
wire n8302;
wire n8303;
wire n8303_1;
wire n8304;
wire n8305;
wire n8306;
wire n8307;
wire n8307_1;
wire n8308;
wire n8309;
wire n8310;
wire n8311;
wire n8311_1;
wire n8312;
wire n8313;
wire n8315;
wire n8316;
wire n8316_1;
wire n8317;
wire n8319;
wire n8320;
wire n8320_1;
wire n8321;
wire n8322;
wire n8323;
wire n8324;
wire n8324_1;
wire n8325;
wire n8326;
wire n8328;
wire n8329;
wire n8330;
wire n8332;
wire n8333;
wire n8334;
wire n8334_1;
wire n8335;
wire n8336;
wire n8337;
wire n8337_1;
wire n8338;
wire n8339;
wire n834;
wire n8340;
wire n8340_1;
wire n8341;
wire n8342;
wire n8343;
wire n8344;
wire n8345;
wire n8345_1;
wire n8346;
wire n8348;
wire n8349;
wire n8350;
wire n8350_1;
wire n8351;
wire n8352;
wire n8353;
wire n8354;
wire n8354_1;
wire n8355;
wire n8356;
wire n8358;
wire n8359;
wire n8359_1;
wire n8360;
wire n8361;
wire n8362;
wire n8362_1;
wire n8365;
wire n8366;
wire n8367;
wire n8368;
wire n8369;
wire n8370;
wire n8371;
wire n8372;
wire n8372_1;
wire n8373;
wire n8374;
wire n8375;
wire n8377;
wire n8377_1;
wire n8378;
wire n8379;
wire n8380;
wire n8382;
wire n8382_1;
wire n8383;
wire n8385;
wire n8386;
wire n8387;
wire n8387_1;
wire n8388;
wire n839;
wire n8390;
wire n8391;
wire n8392;
wire n8392_1;
wire n8393;
wire n8394;
wire n8395;
wire n8396;
wire n8396_1;
wire n8397;
wire n8398;
wire n8399;
wire n8400;
wire n8401;
wire n8401_1;
wire n8402;
wire n8403;
wire n8404;
wire n8405;
wire n8405_1;
wire n8406;
wire n8407;
wire n8408;
wire n8409;
wire n8410;
wire n8410_1;
wire n8411;
wire n8412;
wire n8413;
wire n8414;
wire n8415;
wire n8415_1;
wire n8417;
wire n8418;
wire n8419;
wire n8421;
wire n8422;
wire n8423;
wire n8424;
wire n8425;
wire n8426;
wire n8426_1;
wire n8427;
wire n8429;
wire n8430;
wire n8430_1;
wire n8431;
wire n8432;
wire n8433;
wire n8434;
wire n8435;
wire n8435_1;
wire n8436;
wire n8437;
wire n8438;
wire n8438_1;
wire n8439;
wire n844;
wire n8440;
wire n8441;
wire n8442;
wire n8443;
wire n8443_1;
wire n8444;
wire n8445;
wire n8446;
wire n8447;
wire n8447_1;
wire n8448;
wire n8449;
wire n8450;
wire n8451;
wire n8451_1;
wire n8452;
wire n8453;
wire n8454;
wire n8455;
wire n8455_1;
wire n8456;
wire n8457;
wire n8458;
wire n8459;
wire n8459_1;
wire n8460;
wire n8461;
wire n8463;
wire n8464;
wire n8465;
wire n8466;
wire n8467;
wire n8467_1;
wire n8468;
wire n8469;
wire n8470;
wire n8471;
wire n8472;
wire n8472_1;
wire n8473;
wire n8474;
wire n8475;
wire n8476;
wire n8477;
wire n8477_1;
wire n8478;
wire n8479;
wire n8480;
wire n8481;
wire n8481_1;
wire n8482;
wire n8483;
wire n8484;
wire n8485;
wire n8486;
wire n8486_1;
wire n8487;
wire n8488;
wire n8489;
wire n849;
wire n8490;
wire n8491;
wire n8491_1;
wire n8492;
wire n8493;
wire n8494;
wire n8495;
wire n8497;
wire n8498;
wire n8499;
wire n8499_1;
wire n8500;
wire n8501;
wire n8502;
wire n8503;
wire n8504;
wire n8504_1;
wire n8505;
wire n8506;
wire n8507;
wire n8508;
wire n8508_1;
wire n8509;
wire n8511;
wire n8512;
wire n8513;
wire n8514;
wire n8516;
wire n8517;
wire n8517_1;
wire n8519;
wire n8520;
wire n8521;
wire n8522;
wire n8522_1;
wire n8523;
wire n8524;
wire n8525;
wire n8526;
wire n8526_1;
wire n8528;
wire n8529;
wire n8531;
wire n8531_1;
wire n8532;
wire n8534;
wire n8535;
wire n8535_1;
wire n8536;
wire n8537;
wire n8538;
wire n8539;
wire n854;
wire n8540;
wire n8540_1;
wire n8541;
wire n8542;
wire n8543;
wire n8544;
wire n8544_1;
wire n8545;
wire n8546;
wire n8547;
wire n8549;
wire n8549_1;
wire n8551;
wire n8552;
wire n8552_1;
wire n8553;
wire n8554;
wire n8555;
wire n8556;
wire n8557;
wire n8557_1;
wire n8558;
wire n8559;
wire n8560;
wire n8561;
wire n8561_1;
wire n8562;
wire n8563;
wire n8564;
wire n8565;
wire n8565_1;
wire n8566;
wire n8567;
wire n8568;
wire n8569;
wire n857;
wire n8570;
wire n8571;
wire n8572;
wire n8574;
wire n8575;
wire n8575_1;
wire n8577;
wire n8578;
wire n8578_1;
wire n8580;
wire n8581;
wire n8583;
wire n8583_1;
wire n8584;
wire n8585;
wire n8586;
wire n8587;
wire n8588;
wire n8588_1;
wire n8590;
wire n8591;
wire n8593;
wire n8593_1;
wire n8594;
wire n8596;
wire n8597;
wire n8598;
wire n8598_1;
wire n8599;
wire n8600;
wire n8601;
wire n8602;
wire n8602_1;
wire n8603;
wire n8604;
wire n8605;
wire n8606;
wire n8607;
wire n8607_1;
wire n8608;
wire n8609;
wire n8610;
wire n8611;
wire n8612;
wire n8612_1;
wire n8613;
wire n8614;
wire n8615;
wire n8616;
wire n8616_1;
wire n8617;
wire n8618;
wire n8619;
wire n862;
wire n8620;
wire n8621;
wire n8621_1;
wire n8622;
wire n8623;
wire n8624;
wire n8625;
wire n8625_1;
wire n8626;
wire n8627;
wire n8628;
wire n8628_1;
wire n8630;
wire n8631;
wire n8632;
wire n8632_1;
wire n8633;
wire n8634;
wire n8636;
wire n8637;
wire n8637_1;
wire n8638;
wire n8639;
wire n8640;
wire n8641;
wire n8642;
wire n8643;
wire n8645;
wire n8645_1;
wire n8646;
wire n8648;
wire n8650;
wire n8650_1;
wire n8653;
wire n8654;
wire n8654_1;
wire n8656;
wire n8657;
wire n8658;
wire n8659;
wire n8660;
wire n8661;
wire n8662;
wire n8662_1;
wire n8663;
wire n8664;
wire n8665;
wire n8666;
wire n8666_1;
wire n8667;
wire n8668;
wire n8669;
wire n867;
wire n8670;
wire n8671;
wire n8671_1;
wire n8672;
wire n8673;
wire n8674;
wire n8675;
wire n8676;
wire n8676_1;
wire n8677;
wire n8678;
wire n8679;
wire n8680;
wire n8681;
wire n8681_1;
wire n8682;
wire n8683;
wire n8684;
wire n8685;
wire n8685_1;
wire n8686;
wire n8687;
wire n8688;
wire n8689;
wire n8689_1;
wire n8690;
wire n8691;
wire n8693;
wire n8694;
wire n8694_1;
wire n8695;
wire n8696;
wire n8697;
wire n8698;
wire n8698_1;
wire n8699;
wire n870;
wire n8700;
wire n8701;
wire n8702;
wire n8703;
wire n8703_1;
wire n8704;
wire n8705;
wire n8706;
wire n8707;
wire n8708;
wire n8708_1;
wire n8710;
wire n8711;
wire n8711_1;
wire n8712;
wire n8713;
wire n8714;
wire n8715;
wire n8715_1;
wire n8716;
wire n8717;
wire n8719;
wire n8720;
wire n8720_1;
wire n8722;
wire n8723;
wire n8725;
wire n8725_1;
wire n8726;
wire n8728;
wire n8729;
wire n8730;
wire n8730_1;
wire n8731;
wire n8732;
wire n8734;
wire n8734_1;
wire n8735;
wire n8737;
wire n8738;
wire n8739;
wire n8739_1;
wire n8740;
wire n8741;
wire n8742;
wire n8743;
wire n8743_1;
wire n8744;
wire n8745;
wire n8746;
wire n8747;
wire n8748;
wire n8748_1;
wire n8749;
wire n875;
wire n8750;
wire n8751;
wire n8752;
wire n8753;
wire n8753_1;
wire n8754;
wire n8755;
wire n8757;
wire n8757_1;
wire n8759;
wire n8760;
wire n8761;
wire n8762;
wire n8762_1;
wire n8763;
wire n8764;
wire n8765;
wire n8766;
wire n8767;
wire n8767_1;
wire n8768;
wire n8770;
wire n8771;
wire n8771_1;
wire n8773;
wire n8774;
wire n8775;
wire n8776;
wire n8777;
wire n8778;
wire n8779;
wire n8780;
wire n8780_1;
wire n8781;
wire n8782;
wire n8783;
wire n8784;
wire n8784_1;
wire n8785;
wire n8786;
wire n8787;
wire n8788;
wire n8788_1;
wire n8789;
wire n8790;
wire n8791;
wire n8792;
wire n8793;
wire n8793_1;
wire n8794;
wire n8795;
wire n8796;
wire n8797;
wire n8797_1;
wire n8798;
wire n8799;
wire n880;
wire n8800;
wire n8800_1;
wire n8801;
wire n8803;
wire n8804;
wire n8805;
wire n8806;
wire n8807;
wire n8808;
wire n8809;
wire n8809_1;
wire n8810;
wire n8812;
wire n8813;
wire n8814;
wire n8815;
wire n8816;
wire n8817;
wire n8818;
wire n8818_1;
wire n8820;
wire n8821;
wire n8823;
wire n8823_1;
wire n8824;
wire n8826;
wire n8826_1;
wire n8828;
wire n8829;
wire n8830;
wire n8831;
wire n8831_1;
wire n8832;
wire n8833;
wire n8834;
wire n8835;
wire n8835_1;
wire n8837;
wire n8839;
wire n8840;
wire n8840_1;
wire n8841;
wire n8842;
wire n8843;
wire n8845;
wire n8845_1;
wire n8847;
wire n8848;
wire n8849;
wire n885;
wire n8850;
wire n8850_1;
wire n8851;
wire n8852;
wire n8853;
wire n8855;
wire n8855_1;
wire n8856;
wire n8857;
wire n8858;
wire n8859;
wire n8860;
wire n8860_1;
wire n8861;
wire n8862;
wire n8863;
wire n8864;
wire n8866;
wire n8867;
wire n8868;
wire n8869;
wire n8869_1;
wire n8870;
wire n8872;
wire n8873;
wire n8873_1;
wire n8875;
wire n8876;
wire n8877;
wire n8877_1;
wire n8878;
wire n8880;
wire n8881;
wire n8882;
wire n8882_1;
wire n8883;
wire n8884;
wire n8885;
wire n8886;
wire n8886_1;
wire n8887;
wire n8888;
wire n8889;
wire n8890;
wire n8891;
wire n8891_1;
wire n8892;
wire n8893;
wire n8894;
wire n8895;
wire n8895_1;
wire n8896;
wire n8899;
wire n8899_1;
wire n890;
wire n8901;
wire n8902;
wire n8903;
wire n8904;
wire n8905;
wire n8907;
wire n8908;
wire n8908_1;
wire n8910;
wire n8911;
wire n8912;
wire n8913;
wire n8914;
wire n8915;
wire n8916;
wire n8917;
wire n8917_1;
wire n8918;
wire n8919;
wire n8921;
wire n8922;
wire n8922_1;
wire n8923;
wire n8924;
wire n8925;
wire n8926;
wire n8927;
wire n8928;
wire n8930;
wire n8931;
wire n8931_1;
wire n8933;
wire n8934;
wire n8934_1;
wire n8935;
wire n8936;
wire n8937;
wire n8939;
wire n8939_1;
wire n894;
wire n8941;
wire n8942;
wire n8943;
wire n8944;
wire n8945;
wire n8947;
wire n8948;
wire n8948_1;
wire n8950;
wire n8951;
wire n8953;
wire n8954;
wire n8955;
wire n8957;
wire n8958;
wire n8958_1;
wire n8959;
wire n8960;
wire n8961;
wire n8963;
wire n8963_1;
wire n8964;
wire n8966;
wire n8967;
wire n8968;
wire n8969;
wire n8971;
wire n8971_1;
wire n8972;
wire n8974;
wire n8975;
wire n8976;
wire n8976_1;
wire n8977;
wire n8978;
wire n8979;
wire n8980;
wire n8981;
wire n8981_1;
wire n8982;
wire n8983;
wire n8984;
wire n8985;
wire n8986;
wire n8986_1;
wire n8987;
wire n8988;
wire n8989;
wire n899;
wire n8990;
wire n8991;
wire n8992;
wire n8993;
wire n8994;
wire n8995;
wire n8995_1;
wire n8997;
wire n8999;
wire n9000;
wire n9000_1;
wire n9001;
wire n9002;
wire n9003;
wire n9004;
wire n9005;
wire n9005_1;
wire n9006;
wire n9007;
wire n9008;
wire n9009;
wire n9010;
wire n9010_1;
wire n9011;
wire n9012;
wire n9013;
wire n9014;
wire n9014_1;
wire n9015;
wire n9016;
wire n9017;
wire n9017_1;
wire n9019;
wire n9020;
wire n9022;
wire n9022_1;
wire n9023;
wire n9025;
wire n9025_1;
wire n9026;
wire n9027;
wire n9028;
wire n9029;
wire n903;
wire n9030;
wire n9030_1;
wire n9031;
wire n9032;
wire n9033;
wire n9034;
wire n9034_1;
wire n9035;
wire n9036;
wire n9037;
wire n9038;
wire n9040;
wire n9041;
wire n9042;
wire n9042_1;
wire n9043;
wire n9044;
wire n9045;
wire n9046;
wire n9047;
wire n9047_1;
wire n9048;
wire n9049;
wire n9050;
wire n9051;
wire n9052;
wire n9052_1;
wire n9053;
wire n9054;
wire n9055;
wire n9056;
wire n9057;
wire n9057_1;
wire n9058;
wire n9059;
wire n9060;
wire n9060_1;
wire n9061;
wire n9063;
wire n9064;
wire n9065;
wire n9066;
wire n9067;
wire n9068;
wire n9069;
wire n9069_1;
wire n907;
wire n9070;
wire n9071;
wire n9072;
wire n9073;
wire n9074;
wire n9074_1;
wire n9075;
wire n9077;
wire n9078;
wire n9079;
wire n9079_1;
wire n9080;
wire n9081;
wire n9082;
wire n9082_1;
wire n9083;
wire n9084;
wire n9086;
wire n9086_1;
wire n9087;
wire n9089;
wire n9090;
wire n9091;
wire n9091_1;
wire n9092;
wire n9093;
wire n9094;
wire n9095;
wire n9096;
wire n9096_1;
wire n9098;
wire n9100;
wire n9101;
wire n9102;
wire n9103;
wire n9104;
wire n9105;
wire n9106;
wire n9106_1;
wire n9107;
wire n9108;
wire n9109;
wire n911;
wire n9110;
wire n9110_1;
wire n9111;
wire n9112;
wire n9113;
wire n9114;
wire n9115;
wire n9115_1;
wire n9116;
wire n9117;
wire n9118;
wire n9119;
wire n9120;
wire n9121;
wire n9122;
wire n9123;
wire n9124;
wire n9124_1;
wire n9125;
wire n9126;
wire n9127;
wire n9128;
wire n9129;
wire n9129_1;
wire n9130;
wire n9131;
wire n9132;
wire n9133;
wire n9134;
wire n9134_1;
wire n9135;
wire n9136;
wire n9137;
wire n9138;
wire n9138_1;
wire n9139;
wire n9140;
wire n9141;
wire n9142;
wire n9143;
wire n9143_1;
wire n9144;
wire n9145;
wire n9146;
wire n9146_1;
wire n9147;
wire n9148;
wire n9149;
wire n9151;
wire n9151_1;
wire n9152;
wire n9153;
wire n9154;
wire n9155;
wire n9156;
wire n9157;
wire n9158;
wire n916;
wire n9160;
wire n9160_1;
wire n9161;
wire n9163;
wire n9164;
wire n9164_1;
wire n9166;
wire n9167;
wire n9168;
wire n9169;
wire n9169_1;
wire n9170;
wire n9171;
wire n9172;
wire n9173;
wire n9173_1;
wire n9175;
wire n9176;
wire n9177;
wire n9178;
wire n9178_1;
wire n9179;
wire n9180;
wire n9181;
wire n9182;
wire n9182_1;
wire n9183;
wire n9184;
wire n9185;
wire n9186;
wire n9187;
wire n9187_1;
wire n9188;
wire n9189;
wire n9190;
wire n9191;
wire n9192;
wire n9192_1;
wire n9193;
wire n9195;
wire n9196;
wire n9196_1;
wire n9197;
wire n9199;
wire n920;
wire n9200;
wire n9201;
wire n9201_1;
wire n9202;
wire n9203;
wire n9204;
wire n9205;
wire n9206;
wire n9206_1;
wire n9207;
wire n9208;
wire n9209;
wire n9210;
wire n9211;
wire n9211_1;
wire n9212;
wire n9214;
wire n9215;
wire n9216;
wire n9217;
wire n9219;
wire n9220;
wire n9220_1;
wire n9221;
wire n9222;
wire n9223;
wire n9224;
wire n9225;
wire n9225_1;
wire n9226;
wire n9227;
wire n9228;
wire n9228_1;
wire n9229;
wire n9230;
wire n9231;
wire n9232;
wire n9233;
wire n9233_1;
wire n9234;
wire n9235;
wire n9236;
wire n9237;
wire n9238;
wire n9238_1;
wire n9239;
wire n9240;
wire n9241;
wire n9242;
wire n9242_1;
wire n9243;
wire n9244;
wire n9245;
wire n9246;
wire n9247;
wire n9248;
wire n9249;
wire n925;
wire n9250;
wire n9250_1;
wire n9251;
wire n9253;
wire n9254;
wire n9255;
wire n9256;
wire n9258;
wire n9258_1;
wire n9259;
wire n9260;
wire n9261;
wire n9262;
wire n9263;
wire n9264;
wire n9265;
wire n9267;
wire n9267_1;
wire n9268;
wire n9269;
wire n9270;
wire n9271;
wire n9272;
wire n9272_1;
wire n9273;
wire n9274;
wire n9275;
wire n9276;
wire n9277;
wire n9277_1;
wire n9279;
wire n9282;
wire n9282_1;
wire n9283;
wire n9284;
wire n9285;
wire n9286;
wire n9287;
wire n9287_1;
wire n9288;
wire n9289;
wire n9290;
wire n9290_1;
wire n9291;
wire n9292;
wire n9293;
wire n9294;
wire n9294_1;
wire n9295;
wire n9296;
wire n9297;
wire n9298;
wire n9298_1;
wire n9299;
wire n930;
wire n9300;
wire n9301;
wire n9302;
wire n9303;
wire n9305;
wire n9306;
wire n9307;
wire n9307_1;
wire n9308;
wire n9309;
wire n9310;
wire n9311;
wire n9312;
wire n9312_1;
wire n9313;
wire n9315;
wire n9316;
wire n9316_1;
wire n9317;
wire n9318;
wire n9319;
wire n9321;
wire n9321_1;
wire n9322;
wire n9323;
wire n9324;
wire n9326;
wire n9326_1;
wire n9327;
wire n9329;
wire n9330;
wire n9330_1;
wire n9332;
wire n9333;
wire n9334;
wire n9335;
wire n9335_1;
wire n9336;
wire n9337;
wire n9338;
wire n9339;
wire n9339_1;
wire n9340;
wire n9341;
wire n9342;
wire n9343;
wire n9343_1;
wire n9344;
wire n9345;
wire n9346;
wire n9347;
wire n9348;
wire n9348_1;
wire n935;
wire n9350;
wire n9351;
wire n9352;
wire n9353;
wire n9354;
wire n9355;
wire n9356;
wire n9357;
wire n9358;
wire n9359;
wire n9360;
wire n9361;
wire n9361_1;
wire n9362;
wire n9363;
wire n9364;
wire n9365;
wire n9365_1;
wire n9367;
wire n9368;
wire n9370;
wire n9370_1;
wire n9371;
wire n9372;
wire n9373;
wire n9373_1;
wire n9374;
wire n9376;
wire n9377;
wire n9377_1;
wire n9379;
wire n9380;
wire n9381;
wire n9382;
wire n9383;
wire n9384;
wire n9385;
wire n9385_1;
wire n9386;
wire n9387;
wire n9389;
wire n9390;
wire n9391;
wire n9392;
wire n9393;
wire n9394;
wire n9395;
wire n9396;
wire n9397;
wire n9398;
wire n9398_1;
wire n9399;
wire n940;
wire n9401;
wire n9402;
wire n9402_1;
wire n9403;
wire n9404;
wire n9405;
wire n9405_1;
wire n9406;
wire n9407;
wire n9409;
wire n9410;
wire n9410_1;
wire n9411;
wire n9412;
wire n9413;
wire n9414;
wire n9415;
wire n9416;
wire n9417;
wire n9419;
wire n9420;
wire n9420_1;
wire n9421;
wire n9422;
wire n9423;
wire n9424;
wire n9425;
wire n9425_1;
wire n9426;
wire n9427;
wire n9428;
wire n9428_1;
wire n9429;
wire n9430;
wire n9431;
wire n9432;
wire n9433;
wire n9435;
wire n9436;
wire n9436_1;
wire n9437;
wire n9438;
wire n9439;
wire n944;
wire n9440;
wire n9441;
wire n9441_1;
wire n9442;
wire n9443;
wire n9444;
wire n9445;
wire n9446;
wire n9447;
wire n9449;
wire n9449_1;
wire n9450;
wire n9452;
wire n9453;
wire n9454;
wire n9455;
wire n9456;
wire n9458;
wire n9459;
wire n9459_1;
wire n9461;
wire n9462;
wire n9462_1;
wire n9463;
wire n9464;
wire n9465;
wire n9466;
wire n9467;
wire n9467_1;
wire n9468;
wire n9469;
wire n9470;
wire n9470_1;
wire n9471;
wire n9472;
wire n9473;
wire n9474;
wire n9475;
wire n9475_1;
wire n9476;
wire n9477;
wire n9478;
wire n9478_1;
wire n9479;
wire n948;
wire n9481;
wire n9482;
wire n9483;
wire n9484;
wire n9485;
wire n9486;
wire n9487;
wire n9487_1;
wire n9488;
wire n9490;
wire n9491;
wire n9492;
wire n9492_1;
wire n9493;
wire n9494;
wire n9496;
wire n9497;
wire n9497_1;
wire n9499;
wire n9501;
wire n9502;
wire n9502_1;
wire n9503;
wire n9504;
wire n9505;
wire n9506;
wire n9507;
wire n9507_1;
wire n9508;
wire n9509;
wire n9510;
wire n9511;
wire n9512;
wire n9512_1;
wire n9513;
wire n9515;
wire n9516;
wire n9517;
wire n9517_1;
wire n9518;
wire n9519;
wire n9520;
wire n9520_1;
wire n9521;
wire n9522;
wire n9523;
wire n9525;
wire n9525_1;
wire n9526;
wire n9528;
wire n9528_1;
wire n9529;
wire n953;
wire n9531;
wire n9532;
wire n9533;
wire n9534;
wire n9535;
wire n9536;
wire n9537;
wire n9537_1;
wire n9538;
wire n9540;
wire n9541;
wire n9541_1;
wire n9543;
wire n9544;
wire n9545;
wire n9546;
wire n9546_1;
wire n9547;
wire n9549;
wire n9549_1;
wire n9550;
wire n9552;
wire n9553;
wire n9554;
wire n9555;
wire n9556;
wire n9558;
wire n9559;
wire n9559_1;
wire n956;
wire n9561;
wire n9562;
wire n9563;
wire n9564;
wire n9564_1;
wire n9565;
wire n9566;
wire n9568;
wire n9569;
wire n9569_1;
wire n9570;
wire n9571;
wire n9572;
wire n9574;
wire n9574_1;
wire n9575;
wire n9577;
wire n9578;
wire n9579;
wire n9581;
wire n9582;
wire n9583;
wire n9584;
wire n9585;
wire n9586;
wire n9587;
wire n9588;
wire n9588_1;
wire n9590;
wire n9591;
wire n9592;
wire n9592_1;
wire n9594;
wire n9595;
wire n9597;
wire n9597_1;
wire n9598;
wire n9600;
wire n9601;
wire n9602;
wire n9602_1;
wire n9603;
wire n9604;
wire n9605;
wire n9606;
wire n9606_1;
wire n9607;
wire n9608;
wire n9609;
wire n961;
wire n9610;
wire n9611;
wire n9611_1;
wire n9612;
wire n9613;
wire n9614;
wire n9615;
wire n9616;
wire n9616_1;
wire n9617;
wire n9618;
wire n9619;
wire n9620;
wire n9620_1;
wire n9622;
wire n9623;
wire n9624;
wire n9625;
wire n9626;
wire n9627;
wire n9628;
wire n9628_1;
wire n9629;
wire n9630;
wire n9631;
wire n9632;
wire n9633;
wire n9633_1;
wire n9634;
wire n9635;
wire n9636;
wire n9637;
wire n9638;
wire n9639;
wire n9640;
wire n9641;
wire n9642;
wire n9643;
wire n9644;
wire n9645;
wire n9646;
wire n9647;
wire n9647_1;
wire n9648;
wire n9649;
wire n9651;
wire n9651_1;
wire n9652;
wire n9654;
wire n9655;
wire n9655_1;
wire n9656;
wire n9657;
wire n9658;
wire n9659;
wire n966;
wire n9660;
wire n9660_1;
wire n9663;
wire n9664;
wire n9664_1;
wire n9665;
wire n9666;
wire n9667;
wire n9668;
wire n9668_1;
wire n9670;
wire n9671;
wire n9672;
wire n9673;
wire n9674;
wire n9675;
wire n9677;
wire n9678;
wire n9678_1;
wire n9680;
wire n9681;
wire n9683;
wire n9683_1;
wire n9684;
wire n9685;
wire n9686;
wire n9687;
wire n9688;
wire n9689;
wire n9691;
wire n9692;
wire n9692_1;
wire n9694;
wire n9695;
wire n9695_1;
wire n9697;
wire n9698;
wire n9699;
wire n9700;
wire n9700_1;
wire n9701;
wire n9703;
wire n9704;
wire n9705;
wire n9706;
wire n9707;
wire n9708;
wire n9709;
wire n9709_1;
wire n971;
wire n9710;
wire n9712;
wire n9713;
wire n9714;
wire n9715;
wire n9716;
wire n9717;
wire n9718;
wire n9719;
wire n9719_1;
wire n9720;
wire n9721;
wire n9723;
wire n9724;
wire n9724_1;
wire n9727;
wire n9728;
wire n9729;
wire n9730;
wire n9731;
wire n9732;
wire n9733;
wire n9733_1;
wire n9734;
wire n9735;
wire n9736;
wire n9737;
wire n9737_1;
wire n9738;
wire n9739;
wire n9740;
wire n9741;
wire n9742;
wire n9743;
wire n9744;
wire n9746;
wire n9746_1;
wire n9748;
wire n9750;
wire n9750_1;
wire n9751;
wire n9752;
wire n9753;
wire n9754;
wire n9754_1;
wire n9755;
wire n9756;
wire n9757;
wire n9758;
wire n9758_1;
wire n9759;
wire n976;
wire n9760;
wire n9761;
wire n9762;
wire n9763;
wire n9763_1;
wire n9764;
wire n9765;
wire n9766;
wire n9767;
wire n9768;
wire n9768_1;
wire n9769;
wire n9770;
wire n9771;
wire n9772;
wire n9773;
wire n9773_1;
wire n9774;
wire n9775;
wire n9777;
wire n9778;
wire n9778_1;
wire n9780;
wire n9781;
wire n9783;
wire n9783_1;
wire n9784;
wire n9785;
wire n9786;
wire n9787;
wire n9787_1;
wire n9789;
wire n9791;
wire n9792;
wire n9792_1;
wire n9793;
wire n9795;
wire n9796;
wire n9796_1;
wire n9798;
wire n9799;
wire n9801;
wire n9801_1;
wire n9802;
wire n9804;
wire n9805;
wire n9805_1;
wire n9807;
wire n9808;
wire n9809;
wire n9809_1;
wire n981;
wire n9810;
wire n9811;
wire n9813;
wire n9814;
wire n9814_1;
wire n9816;
wire n9817;
wire n9819;
wire n9819_1;
wire n9821;
wire n9822;
wire n9823;
wire n9824;
wire n9824_1;
wire n9825;
wire n9826;
wire n9827;
wire n9828;
wire n9828_1;
wire n9831;
wire n9832;
wire n9833;
wire n9833_1;
wire n9834;
wire n9835;
wire n9836;
wire n9837;
wire n9837_1;
wire n9838;
wire n9839;
wire n9840;
wire n9840_1;
wire n9841;
wire n9842;
wire n9843;
wire n9844;
wire n9844_1;
wire n9846;
wire n9847;
wire n9849;
wire n9849_1;
wire n985;
wire n9850;
wire n9852;
wire n9853;
wire n9853_1;
wire n9854;
wire n9855;
wire n9856;
wire n9857;
wire n9858;
wire n9858_1;
wire n9859;
wire n9860;
wire n9861;
wire n9863;
wire n9863_1;
wire n9864;
wire n9866;
wire n9867;
wire n9867_1;
wire n9869;
wire n9870;
wire n9871;
wire n9871_1;
wire n9872;
wire n9873;
wire n9875;
wire n9875_1;
wire n9876;
wire n9878;
wire n9879;
wire n9880;
wire n9880_1;
wire n9881;
wire n9882;
wire n9884;
wire n9885;
wire n9885_1;
wire n9886;
wire n9887;
wire n9889;
wire n9889_1;
wire n9890;
wire n9892;
wire n9893;
wire n9894;
wire n9895;
wire n9896;
wire n9898;
wire n9899;
wire n990;
wire n9900;
wire n9901;
wire n9902;
wire n9904;
wire n9906;
wire n9907;
wire n9907_1;
wire n9908;
wire n9909;
wire n9910;
wire n9911;
wire n9911_1;
wire n9913;
wire n9914;
wire n9914_1;
wire n9915;
wire n9916;
wire n9918;
wire n9918_1;
wire n9919;
wire n9921;
wire n9922;
wire n9923;
wire n9924;
wire n9925;
wire n9926;
wire n9927;
wire n9928;
wire n9929;
wire n9930;
wire n9930_1;
wire n9931;
wire n9932;
wire n9933;
wire n9934;
wire n9935;
wire n9935_1;
wire n9936;
wire n9937;
wire n9938;
wire n9939;
wire n9939_1;
wire n9940;
wire n9941;
wire n9942;
wire n9943;
wire n9944;
wire n9944_1;
wire n9945;
wire n9947;
wire n9948;
wire n9949;
wire n995;
wire n9950;
wire n9951;
wire n9952;
wire n9953;
wire n9953_1;
wire n9954;
wire n9955;
wire n9956;
wire n9957;
wire n9957_1;
wire n9958;
wire n9959;
wire n9960;
wire n9961;
wire n9961_1;
wire n9962;
wire n9963;
wire n9964;
wire n9965;
wire n9966;
wire n9966_1;
wire n9967;
wire n9968;
wire n9970;
wire n9971;
wire n9971_1;
wire n9973;
wire n9974;
wire n9975;
wire n9976;
wire n9976_1;
wire n9977;
wire n9978;
wire n9980;
wire n9981;
wire n9982;
wire n9983;
wire n9985;
wire n9985_1;
wire n9986;
wire n9988;
wire n9988_1;
wire n9989;
wire n9991;
wire n9992;
wire n9992_1;
wire n9994;
wire n9995;
wire n9997;
wire n9997_1;
wire n9998;
wire net_130;
wire net_131;
wire net_132;
wire net_133;
wire net_134;
wire net_135;
wire net_136;
wire net_137;
wire net_138;
wire net_139;
wire net_140;
wire net_141;
wire net_142;
wire net_143;
wire net_144;
wire net_145;
wire net_146;
wire net_147;
wire net_148;
wire net_149;
wire net_150;
wire net_151;
wire net_152;
wire net_153;
wire net_155;
wire net_156;
wire net_157;
wire net_158;
wire net_159;
wire net_160;
wire net_161;
wire net_162;
wire net_163;
wire net_164;
wire net_165;
wire net_166;
wire net_167;
wire net_168;
wire net_169;
wire net_170;
wire net_171;
wire net_179;
wire net_181;
wire net_182;
wire net_183;
wire net_185;
wire net_186;
wire net_187;
wire net_194;
wire net_195;
wire net_196;
wire net_197;
wire net_198;
wire net_199;
wire net_200;
wire net_202;
wire net_203;
wire net_204;
wire net_205;
wire net_206;
wire net_207;
wire net_208;
wire net_216;
wire net_218;
wire net_219;
wire net_220;
wire net_222;
wire net_223;
wire net_224;
wire net_230;
wire net_231;
wire net_232;
wire net_233;
wire net_234;
wire net_235;
wire net_236;
wire net_237;
wire net_238;
wire net_239;
wire net_240;
wire net_241;
wire net_242;
wire net_243;
wire net_244;
wire net_245;
wire net_246;
wire net_247;
wire net_248;
wire net_249;
wire net_250;
wire net_251;
wire net_252;
wire net_253;
wire net_254;
wire net_255;
wire net_256;
wire net_257;
wire net_258;
wire net_259;
wire net_260;
wire net_261;
wire net_274;
wire net_275;
wire net_285;
wire net_286;
wire net_296;
wire net_297;
wire net_300;
wire net_301;
wire net_302;
wire net_303;
wire net_304;
wire net_305;
wire net_306;
wire net_307;
wire net_308;
wire net_309;
wire net_310;
wire net_311;
wire net_312;
wire net_313;
wire net_314;
wire net_315;
wire net_316;
wire net_317;
wire net_318;
wire net_319;
wire net_320;
wire net_321;
wire net_322;
wire net_323;
wire net_324;
wire net_325;
wire net_326;
wire net_327;
wire net_328;
wire net_329;
wire net_330;
wire net_331;
wire net_332;
wire net_333;
wire net_334;
wire net_335;
wire net_336;
wire net_337;
wire net_338;
wire net_339;
wire net_340;
wire net_341;
wire net_342;
wire net_343;
wire net_344;
wire net_345;
wire net_346;
wire net_347;
wire net_348;
wire net_349;
wire net_350;
wire net_351;
wire net_352;
wire net_353;
wire net_354;
wire net_355;
wire net_356;
wire net_357;
wire net_358;
wire net_359;
wire net_360;
wire net_361;
wire net_362;
wire net_363;
wire net_364;
wire net_365;
wire net_366;
wire net_367;
wire net_368;
wire net_369;
wire net_370;
wire net_371;
wire net_372;
wire net_373;
wire net_374;
wire net_375;
wire net_376;
wire net_377;
wire net_378;
wire net_379;
wire net_380;
wire net_381;
wire net_382;
wire net_383;
wire net_384;
wire net_385;
wire net_386;
wire net_387;
wire net_388;
wire net_389;
wire net_390;
wire net_391;
wire net_5849;
wire net_5858;
wire net_5860;
wire net_5861;
wire net_5992;
wire net_6003;
wire net_6013;
wire net_6014;
wire net_6024;
wire net_6025;
wire net_6035;
wire net_6036;
wire net_6046;
wire net_6047;
wire net_6053;
wire net_6054;
wire net_6055;
wire net_6056;
wire net_6057;
wire net_6058;
wire net_6059;
wire net_6060;
wire net_6061;
wire net_6190;
wire net_6191;
wire net_6192;
wire net_6193;
wire net_6195;
wire net_6196;
wire net_6197;
wire net_6198;
wire net_6211;
wire net_6212;
wire net_6213;
wire net_6214;
wire net_6215;
wire net_6216;
wire net_6217;
wire net_6218;
wire net_6223;
wire net_6224;
wire net_6225;
wire net_6226;
wire net_6227;
wire net_6228;
wire net_6229;
wire net_6230;
wire net_6231;
wire net_6232;
wire net_6233;
wire net_6234;
wire net_6235;
wire net_6236;
wire net_6237;
wire net_6238;
wire net_6240;
wire net_6241;
wire net_6242;
wire net_6243;
wire net_6244;
wire net_6245;
wire net_6246;
wire net_6247;
wire net_6248;
wire net_6249;
wire net_6250;
wire net_6251;
wire net_6252;
wire net_6253;
wire net_6254;
wire net_6255;
wire net_6256;
wire net_6257;
wire net_6258;
wire net_6260;
wire net_6261;
wire net_6262;
wire net_6263;
wire net_6264;
wire net_6265;
wire net_6266;
wire net_6267;
wire net_6268;
wire net_6269;
wire net_6270;
wire net_6271;
wire net_6272;
wire net_6273;
wire net_6274;
wire net_6275;
wire net_6276;
wire net_6277;
wire net_6278;
wire net_6279;
wire net_6299;
wire net_6300;
wire net_6301;
wire net_6302;
wire net_6303;
wire net_6304;
wire net_6305;
wire net_6306;
wire net_6307;
wire net_6308;
wire net_6309;
wire net_6310;
wire net_6311;
wire net_6312;
wire net_6313;
wire net_6314;
wire net_6315;
wire net_6316;
wire net_6317;
wire net_6318;
wire net_6320;
wire net_6321;
wire net_6322;
wire net_6323;
wire net_6324;
wire net_6325;
wire net_6326;
wire net_6327;
wire net_6328;
wire net_6329;
wire net_6330;
wire net_6331;
wire net_6332;
wire net_6333;
wire net_6334;
wire net_6335;
wire net_6336;
wire net_6337;
wire net_6338;
wire net_6339;
wire net_6340;
wire net_6341;
wire net_6342;
wire net_6343;
wire net_6344;
wire net_6345;
wire net_6346;
wire net_6347;
wire net_6348;
wire net_6349;
wire net_6350;
wire net_6351;
wire net_6352;
wire net_6353;
wire net_6354;
wire net_6355;
wire net_6356;
wire net_6357;
wire net_6358;
wire net_6359;
wire net_6360;
wire net_6361;
wire net_6362;
wire net_6363;
wire net_6364;
wire net_6365;
wire net_6366;
wire net_6367;
wire net_6368;
wire net_6369;
wire net_6370;
wire net_6371;
wire net_6372;
wire net_6373;
wire net_6374;
wire net_6375;
wire net_6376;
wire net_6377;
wire net_6378;
wire net_6379;
wire net_6380;
wire net_6381;
wire net_6382;
wire net_6383;
wire net_6384;
wire net_6385;
wire net_6386;
wire net_6387;
wire net_6388;
wire net_6389;
wire net_6390;
wire net_6391;
wire net_6392;
wire net_6393;
wire net_6394;
wire net_6395;
wire net_6396;
wire net_6397;
wire net_6398;
wire net_6399;
wire net_6400;
wire net_6403;
wire net_6412;
wire net_6416;
wire net_6417;
wire net_6424;
wire net_6425;
wire net_6426;
wire net_6427;
wire net_6428;
wire net_6429;
wire net_6430;
wire net_6431;
wire net_6432;
wire net_6433;
wire net_6434;
wire net_6435;
wire net_6436;
wire net_6437;
wire net_6438;
wire net_6439;
wire net_6440;
wire net_6441;
wire net_6442;
wire net_6443;
wire net_6444;
wire net_6445;
wire net_6446;
wire net_6447;
wire net_6448;
wire net_6449;
wire net_6450;
wire net_6451;
wire net_6452;
wire net_6453;
wire net_6454;
wire net_6455;
wire net_6456;
wire net_6457;
wire net_6458;
wire net_6459;
wire net_6460;
wire net_6461;
wire net_6462;
wire net_6463;
wire net_6464;
wire net_6465;
wire net_6466;
wire net_6467;
wire net_6468;
wire net_6469;
wire net_6470;
wire net_6471;
wire net_6472;
wire net_6473;
wire net_6474;
wire net_6475;
wire net_6476;
wire net_6477;
wire net_6478;
wire net_6479;
wire net_6480;
wire net_6481;
wire net_6482;
wire net_6483;
wire net_6484;
wire net_6485;
wire net_6486;
wire net_6487;
wire net_6488;
wire net_6489;
wire net_6490;
wire net_6491;
wire net_6492;
wire net_6493;
wire net_6494;
wire net_6495;
wire net_6496;
wire net_6497;
wire net_6498;
wire net_6499;
wire net_6500;
wire net_6501;
wire net_6502;
wire net_6503;
wire net_6504;
wire net_6505;
wire net_6506;
wire net_6507;
wire net_6508;
wire net_6509;
wire net_6510;
wire net_6511;
wire net_6512;
wire net_6513;
wire net_6514;
wire net_6515;
wire net_6516;
wire net_6517;
wire net_6518;
wire net_6519;
wire net_6520;
wire net_6521;
wire net_6522;
wire net_6523;
wire net_6524;
wire net_6525;
wire net_6526;
wire net_6527;
wire net_6528;
wire net_6529;
wire net_6530;
wire net_6531;
wire net_6532;
wire net_6533;
wire net_6534;
wire net_6535;
wire net_6536;
wire net_6537;
wire net_6538;
wire net_6539;
wire net_6540;
wire net_6541;
wire net_6542;
wire net_6543;
wire net_6544;
wire net_6545;
wire net_6546;
wire net_6547;
wire net_6548;
wire net_6549;
wire net_6550;
wire net_6551;
wire net_6556;
wire net_6559;
wire net_6560;
wire net_6561;
wire net_6562;
wire net_6563;
wire net_6564;
wire net_6565;
wire net_6566;
wire net_6567;
wire net_6568;
wire net_6569;
wire net_6570;
wire net_6571;
wire net_6572;
wire net_6573;
wire net_6574;
wire net_6575;
wire net_6576;
wire net_6577;
wire net_6578;
wire net_6579;
wire net_6580;
wire net_6581;
wire net_6582;
wire net_6583;
wire net_6584;
wire net_6585;
wire net_6586;
wire net_6587;
wire net_6588;
wire net_6589;
wire net_6590;
wire net_6591;
wire net_6592;
wire net_6593;
wire net_6594;
wire net_6595;
wire net_6596;
wire net_6597;
wire net_6598;
wire net_6599;
wire net_6600;
wire net_6601;
wire net_6602;
wire net_6603;
wire net_6604;
wire net_6605;
wire net_6606;
wire net_6607;
wire net_6608;
wire net_6609;
wire net_6610;
wire net_6611;
wire net_6612;
wire net_6613;
wire net_6614;
wire net_6615;
wire net_6616;
wire net_6617;
wire net_6618;
wire net_6619;
wire net_6620;
wire net_6621;
wire net_6622;
wire net_6623;
wire net_6624;
wire net_6625;
wire net_6626;
wire net_6627;
wire net_6628;
wire net_6629;
wire net_6630;
wire net_6631;
wire net_6632;
wire net_6633;
wire net_6634;
wire net_6635;
wire net_6636;
wire net_6637;
wire net_6638;
wire net_6639;
wire net_6640;
wire net_6641;
wire net_6642;
wire net_6643;
wire net_6644;
wire net_6645;
wire net_6646;
wire net_6647;
wire net_6648;
wire net_6649;
wire net_6650;
wire net_6651;
wire net_6652;
wire net_6653;
wire net_6654;
wire net_6655;
wire net_6656;
wire net_6657;
wire net_6658;
wire net_6659;
wire net_6660;
wire net_6661;
wire net_6662;
wire net_6663;
wire net_6664;
wire net_6665;
wire net_6666;
wire net_6667;
wire net_6668;
wire net_6669;
wire net_6670;
wire net_6671;
wire net_6672;
wire net_6673;
wire net_6674;
wire net_6675;
wire net_6676;
wire net_6677;
wire net_6678;
wire net_6679;
wire net_6680;
wire net_6681;
wire net_6682;
wire net_6683;
wire net_6684;
wire net_6685;
wire net_6686;
wire net_6691;
wire net_6694;
wire net_6695;
wire net_6696;
wire net_6697;
wire net_6698;
wire net_6699;
wire net_6700;
wire net_6701;
wire net_6702;
wire net_6703;
wire net_6704;
wire net_6705;
wire net_6706;
wire net_6707;
wire net_6708;
wire net_6709;
wire net_6710;
wire net_6711;
wire net_6712;
wire net_6713;
wire net_6714;
wire net_6715;
wire net_6716;
wire net_6717;
wire net_6718;
wire net_6719;
wire net_6720;
wire net_6721;
wire net_6722;
wire net_6723;
wire net_6724;
wire net_6725;
wire net_6726;
wire net_6727;
wire net_6728;
wire net_6729;
wire net_6730;
wire net_6731;
wire net_6732;
wire net_6733;
wire net_6734;
wire net_6735;
wire net_6736;
wire net_6737;
wire net_6738;
wire net_6739;
wire net_6740;
wire net_6741;
wire net_6742;
wire net_6743;
wire net_6744;
wire net_6745;
wire net_6746;
wire net_6747;
wire net_6748;
wire net_6749;
wire net_6750;
wire net_6751;
wire net_6752;
wire net_6753;
wire net_6754;
wire net_6755;
wire net_6756;
wire net_6757;
wire net_6758;
wire net_6759;
wire net_6760;
wire net_6761;
wire net_6762;
wire net_6763;
wire net_6764;
wire net_6765;
wire net_6766;
wire net_6767;
wire net_6768;
wire net_6769;
wire net_6770;
wire net_6771;
wire net_6772;
wire net_6773;
wire net_6774;
wire net_6775;
wire net_6776;
wire net_6777;
wire net_6778;
wire net_6779;
wire net_6780;
wire net_6781;
wire net_6782;
wire net_6783;
wire net_6784;
wire net_6785;
wire net_6786;
wire net_6787;
wire net_6788;
wire net_6789;
wire net_6790;
wire net_6791;
wire net_6792;
wire net_6793;
wire net_6794;
wire net_6795;
wire net_6796;
wire net_6797;
wire net_6798;
wire net_6799;
wire net_6800;
wire net_6801;
wire net_6802;
wire net_6803;
wire net_6804;
wire net_6805;
wire net_6806;
wire net_6807;
wire net_6808;
wire net_6809;
wire net_6810;
wire net_6811;
wire net_6812;
wire net_6813;
wire net_6814;
wire net_6815;
wire net_6816;
wire net_6817;
wire net_6818;
wire net_6819;
wire net_6820;
wire net_6821;
wire net_6826;
wire net_6829;
wire net_6830;
wire net_6831;
wire net_6832;
wire net_6833;
wire net_6834;
wire net_6835;
wire net_6836;
wire net_6837;
wire net_6838;
wire net_6839;
wire net_6840;
wire net_6841;
wire net_6842;
wire net_6843;
wire net_6844;
wire net_6845;
wire net_6846;
wire net_6847;
wire net_6848;
wire net_6849;
wire net_6850;
wire net_6851;
wire net_6852;
wire net_6853;
wire net_6854;
wire net_6855;
wire net_6856;
wire net_6857;
wire net_6858;
wire net_6859;
wire net_6860;
wire net_6861;
wire net_6862;
wire net_6863;
wire net_6864;
wire net_6865;
wire net_6866;
wire net_6867;
wire net_6868;
wire net_6869;
wire net_6870;
wire net_6871;
wire net_6872;
wire net_6873;
wire net_6874;
wire net_6875;
wire net_6876;
wire net_6877;
wire net_6878;
wire net_6879;
wire net_6880;
wire net_6881;
wire net_6882;
wire net_6883;
wire net_6884;
wire net_6885;
wire net_6886;
wire net_6887;
wire net_6888;
wire net_6889;
wire net_6890;
wire net_6891;
wire net_6892;
wire net_6893;
wire net_6894;
wire net_6895;
wire net_6896;
wire net_6897;
wire net_6898;
wire net_6899;
wire net_6900;
wire net_6901;
wire net_6902;
wire net_6903;
wire net_6904;
wire net_6905;
wire net_6906;
wire net_6907;
wire net_6908;
wire net_6909;
wire net_6910;
wire net_6911;
wire net_6912;
wire net_6913;
wire net_6914;
wire net_6915;
wire net_6916;
wire net_6917;
wire net_6918;
wire net_6919;
wire net_6920;
wire net_6921;
wire net_6922;
wire net_6923;
wire net_6924;
wire net_6925;
wire net_6926;
wire net_6927;
wire net_6928;
wire net_6929;
wire net_6930;
wire net_6931;
wire net_6932;
wire net_6933;
wire net_6934;
wire net_6935;
wire net_6936;
wire net_6937;
wire net_6938;
wire net_6939;
wire net_6940;
wire net_6941;
wire net_6942;
wire net_6943;
wire net_6944;
wire net_6945;
wire net_6946;
wire net_6947;
wire net_6948;
wire net_6949;
wire net_6950;
wire net_6951;
wire net_6952;
wire net_6953;
wire net_6954;
wire net_6955;
wire net_6956;
wire net_6961;
wire net_6964;
wire net_6965;
wire net_6966;
wire net_6967;
wire net_6968;
wire net_6969;
wire net_6970;
wire net_6971;
wire net_6972;
wire net_6973;
wire net_6974;
wire net_6975;
wire net_6976;
wire net_6977;
wire net_6978;
wire net_6979;
wire net_6980;
wire net_6981;
wire net_6982;
wire net_6983;
wire net_6984;
wire net_6985;
wire net_6986;
wire net_6987;
wire net_6988;
wire net_6989;
wire net_6990;
wire net_6991;
wire net_6992;
wire net_6993;
wire net_6994;
wire net_6995;
wire net_6996;
wire net_6997;
wire net_6998;
wire net_6999;
wire net_7000;
wire net_7001;
wire net_7002;
wire net_7003;
wire net_7004;
wire net_7005;
wire net_7006;
wire net_7007;
wire net_7008;
wire net_7009;
wire net_7010;
wire net_7011;
wire net_7012;
wire net_7013;
wire net_7014;
wire net_7015;
wire net_7016;
wire net_7017;
wire net_7018;
wire net_7019;
wire net_7020;
wire net_7021;
wire net_7022;
wire net_7023;
wire net_7024;
wire net_7025;
wire net_7026;
wire net_7027;
wire net_7028;
wire net_7029;
wire net_7030;
wire net_7031;
wire net_7032;
wire net_7033;
wire net_7034;
wire net_7035;
wire net_7036;
wire net_7037;
wire net_7038;
wire net_7039;
wire net_7040;
wire net_7041;
wire net_7042;
wire net_7043;
wire net_7044;
wire net_7045;
wire net_7046;
wire net_7047;
wire net_7048;
wire net_7049;
wire net_7050;
wire net_7051;
wire net_7052;
wire net_7053;
wire net_7054;
wire net_7055;
wire net_7056;
wire net_7057;
wire net_7058;
wire net_7059;
wire net_7060;
wire net_7061;
wire net_7062;
wire net_7063;
wire net_7064;
wire net_7065;
wire net_7066;
wire net_7067;
wire net_7068;
wire net_7069;
wire net_7070;
wire net_7071;
wire net_7072;
wire net_7073;
wire net_7074;
wire net_7075;
wire net_7076;
wire net_7077;
wire net_7078;
wire net_7079;
wire net_7080;
wire net_7081;
wire net_7082;
wire net_7083;
wire net_7084;
wire net_7085;
wire net_7086;
wire net_7087;
wire net_7088;
wire net_7089;
wire net_7090;
wire net_7091;
wire net_7096;
wire net_7099;
wire net_7100;
wire net_7101;
wire net_7102;
wire net_7103;
wire net_7104;
wire net_7105;
wire net_7106;
wire net_7107;
wire net_7108;
wire net_7109;
wire net_7110;
wire net_7111;
wire net_7112;
wire net_7113;
wire net_7114;
wire net_7115;
wire net_7116;
wire net_7117;
wire net_7118;
wire net_7119;
wire net_7120;
wire net_7121;
wire net_7122;
wire net_7123;
wire net_7124;
wire net_7125;
wire net_7126;
wire net_7127;
wire net_7128;
wire net_7129;
wire net_7130;
wire net_7131;
wire net_7132;
wire net_7133;
wire net_7134;
wire net_7135;
wire net_7136;
wire net_7137;
wire net_7138;
wire net_7139;
wire net_7140;
wire net_7141;
wire net_7142;
wire net_7143;
wire net_7144;
wire net_7145;
wire net_7146;
wire net_7147;
wire net_7148;
wire net_7149;
wire net_7150;
wire net_7151;
wire net_7152;
wire net_7153;
wire net_7154;
wire net_7155;
wire net_7156;
wire net_7157;
wire net_7158;
wire net_7159;
wire net_7160;
wire net_7161;
wire net_7162;
wire net_7163;
wire net_7164;
wire net_7165;
wire net_7166;
wire net_7167;
wire net_7168;
wire net_7169;
wire net_7170;
wire net_7171;
wire net_7172;
wire net_7173;
wire net_7174;
wire net_7175;
wire net_7176;
wire net_7177;
wire net_7178;
wire net_7179;
wire net_7180;
wire net_7181;
wire net_7182;
wire net_7183;
wire net_7184;
wire net_7185;
wire net_7186;
wire net_7187;
wire net_7188;
wire net_7189;
wire net_7190;
wire net_7191;
wire net_7192;
wire net_7193;
wire net_7194;
wire net_7195;
wire net_7196;
wire net_7197;
wire net_7198;
wire net_7199;
wire net_7200;
wire net_7201;
wire net_7202;
wire net_7203;
wire net_7204;
wire net_7205;
wire net_7206;
wire net_7207;
wire net_7208;
wire net_7209;
wire net_7210;
wire net_7211;
wire net_7212;
wire net_7213;
wire net_7214;
wire net_7215;
wire net_7216;
wire net_7217;
wire net_7218;
wire net_7219;
wire net_7220;
wire net_7221;
wire net_7222;
wire net_7223;
wire net_7224;
wire net_7225;
wire net_7226;
wire net_7231;
wire net_7234;
wire net_7235;
wire net_7236;
wire net_7237;
wire net_7238;
wire net_7239;
wire net_7240;
wire net_7241;
wire net_7242;
wire net_7243;
wire net_7244;
wire net_7245;
wire net_7246;
wire net_7247;
wire net_7248;
wire net_7249;
wire net_7302;
wire net_7303;
wire net_7304;
wire net_7305;
wire net_7306;
wire net_7307;
wire net_7308;
wire net_7309;
wire net_7310;
wire net_7311;
wire net_7312;
wire net_7313;
wire net_7334;
wire net_7335;
wire net_7336;
wire net_7337;
wire net_7338;
wire net_7339;
wire net_7340;
wire net_7341;
wire net_7342;
wire net_7343;
wire net_7344;
wire net_7345;
wire net_7366;
wire net_7367;
wire net_7368;
wire net_7369;
wire net_7370;
wire net_7371;
wire net_7372;
wire net_7373;
wire net_7374;
wire net_7375;
wire net_7376;
wire net_7377;
wire net_7378;
wire net_7385;
wire net_7386;
wire net_7387;
wire net_7388;
wire net_7389;
wire net_7390;
wire net_7391;
wire net_7392;
wire net_7393;
wire net_7394;
wire net_7395;
wire net_7396;
wire net_7397;
wire net_7398;
wire net_7399;
wire net_7400;
wire net_7453;
wire net_7454;
wire net_7455;
wire net_7456;
wire net_7457;
wire net_7458;
wire net_7459;
wire net_7460;
wire net_7461;
wire net_7462;
wire net_7463;
wire net_7464;
wire net_7485;
wire net_7486;
wire net_7487;
wire net_7488;
wire net_7489;
wire net_7490;
wire net_7491;
wire net_7492;
wire net_7493;
wire net_7494;
wire net_7495;
wire net_7496;
wire net_7517;
wire net_7518;
wire net_7519;
wire net_7520;
wire net_7521;
wire net_7522;
wire net_7523;
wire net_7524;
wire net_7525;
wire net_7526;
wire net_7527;
wire net_7528;
wire net_7529;
wire net_7536;
wire net_7537;
wire net_7538;
wire net_7539;
wire net_7540;
wire net_7541;
wire net_7542;
wire net_7543;
wire net_7544;
wire net_7545;
wire net_7546;
wire net_7547;
wire net_7548;
wire net_7549;
wire net_7550;
wire net_7551;
wire net_7604;
wire net_7605;
wire net_7606;
wire net_7607;
wire net_7608;
wire net_7609;
wire net_7610;
wire net_7611;
wire net_7612;
wire net_7613;
wire net_7614;
wire net_7615;
wire net_7636;
wire net_7637;
wire net_7638;
wire net_7639;
wire net_7640;
wire net_7641;
wire net_7642;
wire net_7643;
wire net_7644;
wire net_7645;
wire net_7646;
wire net_7647;
wire net_7668;
wire net_7669;
wire net_7670;
wire net_7671;
wire net_7672;
wire net_7673;
wire net_7674;
wire net_7675;
wire net_7676;
wire net_7677;
wire net_7678;
wire net_7679;
wire net_7680;
wire net_7691;
wire net_7708;
wire net_7709;
wire net_7710;
wire net_7711;
wire net_7712;
wire net_7713;
wire net_7714;
wire net_7715;
wire net_7737;
wire net_7738;
wire net_7739;
wire net_7740;
wire net_7741;
wire net_7742;
wire net_7743;
wire net_7744;
wire net_7750;
wire net_7752;
wire net_7754;
wire net_7756;
wire net_7758;
wire net_7760;
wire net_7762;
wire net_7764;
wire net_7766;
wire net_7767;
wire net_7769;
wire net_7770;
wire net_7771;
wire net_7772;
wire net_7773;
wire net_7774;
wire net_7775;
wire net_7776;
wire net_7777;
wire net_7778;
wire net_7779;
wire net_7780;
wire net_7790;
wire net_7792;
wire net_7799;
wire net_7802;
wire net_7807;

// Start cells
in01f01 g0000 ( .a(net_6416), .o(n6730) );
in01f01 g0001 ( .a(net_6417), .o(n6731) );
na02f01 g0002 ( .a(n6731), .b(n6730), .o(x30) );
in01f01 g0003 ( .a(net_7680), .o(n6733) );
no02f01 g0004 ( .a(n6733), .b(_net_7681), .o(n6734) );
in01f01 g0005 ( .a(_net_7681), .o(n6735) );
no02f01 g0006 ( .a(net_7680), .b(n6735), .o(n6736_1) );
ao22f01 g0007 ( .a(n6736_1), .b(_net_7635), .c(n6734), .d(_net_7603), .o(n6737) );
no02f01 g0008 ( .a(net_7680), .b(_net_7681), .o(n6738) );
no02f01 g0009 ( .a(n6733), .b(n6735), .o(n6739) );
ao22f01 g0010 ( .a(n6739), .b(_net_7667), .c(n6738), .d(_net_7571), .o(n6740) );
na02f01 g0011 ( .a(n6740), .b(n6737), .o(n266) );
ao22f01 g0012 ( .a(n6736_1), .b(net_7640), .c(n6734), .d(net_7608), .o(n6742) );
ao22f01 g0013 ( .a(n6739), .b(net_7672), .c(n6738), .d(_net_7576), .o(n6743) );
na02f01 g0014 ( .a(n6743), .b(n6742), .o(n271) );
in01f01 g0015 ( .a(net_6438), .o(n6745) );
in01f01 g0016 ( .a(net_6502), .o(n6746_1) );
in01f01 g0017 ( .a(_net_6553), .o(n6747) );
na02f01 g0018 ( .a(_net_6554), .b(n6747), .o(n6748) );
in01f01 g0019 ( .a(_net_6554), .o(n6749_1) );
na02f01 g0020 ( .a(n6749_1), .b(n6747), .o(n6750) );
oa22f01 g0021 ( .a(n6750), .b(n6745), .c(n6748), .d(n6746_1), .o(n6751) );
in01f01 g0022 ( .a(net_6470), .o(n6752_1) );
in01f01 g0023 ( .a(net_6534), .o(n6753) );
na02f01 g0024 ( .a(_net_6554), .b(_net_6553), .o(n6754) );
na02f01 g0025 ( .a(n6749_1), .b(_net_6553), .o(n6755) );
oa22f01 g0026 ( .a(n6755), .b(n6752_1), .c(n6754), .d(n6753), .o(n6756_1) );
no02f01 g0027 ( .a(n6756_1), .b(n6751), .o(n6757) );
in01f01 g0028 ( .a(_net_6552), .o(n6758) );
in01f01 g0029 ( .a(_net_5984), .o(n6759) );
in01f01 g0030 ( .a(_net_7749), .o(n6760) );
na03f01 g0031 ( .a(_net_7791), .b(net_6061), .c(n6760), .o(n6761_1) );
no02f01 g0032 ( .a(n6761_1), .b(n6759), .o(n6762) );
no02f01 g0033 ( .a(_net_5986), .b(_net_5987), .o(n6763) );
na03f01 g0034 ( .a(n6763), .b(n6762), .c(n6758), .o(n6764) );
no02f01 g0035 ( .a(n6764), .b(n6757), .o(n6765_1) );
na02f01 g0036 ( .a(n6762), .b(_net_5986), .o(n6766) );
in01f01 g0037 ( .a(net_6440), .o(n6767) );
in01f01 g0038 ( .a(net_6504), .o(n6768) );
oa22f01 g0039 ( .a(n6750), .b(n6767), .c(n6748), .d(n6768), .o(n6769) );
in01f01 g0040 ( .a(net_6536), .o(n6770_1) );
in01f01 g0041 ( .a(net_6472), .o(n6771) );
oa22f01 g0042 ( .a(n6755), .b(n6771), .c(n6754), .d(n6770_1), .o(n6772) );
no02f01 g0043 ( .a(n6772), .b(n6769), .o(n6773) );
no02f01 g0044 ( .a(n6773), .b(n6766), .o(n6774_1) );
na02f01 g0045 ( .a(n6762), .b(_net_5987), .o(n6775) );
in01f01 g0046 ( .a(n6748), .o(n6776) );
in01f01 g0047 ( .a(n6750), .o(n6777) );
ao22f01 g0048 ( .a(n6777), .b(net_6442), .c(n6776), .d(net_6506), .o(n6778) );
in01f01 g0049 ( .a(n6754), .o(n6779_1) );
in01f01 g0050 ( .a(n6755), .o(n6780) );
ao22f01 g0051 ( .a(n6780), .b(net_6474), .c(n6779_1), .d(net_6538), .o(n6781) );
ao12f01 g0052 ( .a(n6775), .b(n6781), .c(n6778), .o(n6782) );
in01f01 g0053 ( .a(_net_6082), .o(n6783_1) );
na02f01 g0054 ( .a(n6761_1), .b(_net_5984), .o(n6784) );
no02f01 g0055 ( .a(n6784), .b(n6783_1), .o(n6785) );
no04f01 g0056 ( .a(n6785), .b(n6782), .c(n6774_1), .d(n6765_1), .o(n6786) );
in01f01 g0057 ( .a(net_6486), .o(n6787) );
in01f01 g0058 ( .a(net_6454), .o(n6788_1) );
na04f01 g0059 ( .a(n6763), .b(n6762), .c(n6780), .d(_net_6552), .o(n6789) );
na04f01 g0060 ( .a(n6763), .b(n6762), .c(n6777), .d(_net_6552), .o(n6790) );
oa22f01 g0061 ( .a(n6790), .b(n6788_1), .c(n6789), .d(n6787), .o(n6791) );
in01f01 g0062 ( .a(net_6550), .o(n6792) );
in01f01 g0063 ( .a(net_6518), .o(n6793_1) );
na04f01 g0064 ( .a(n6763), .b(n6762), .c(n6776), .d(_net_6552), .o(n6794) );
na04f01 g0065 ( .a(n6763), .b(n6762), .c(n6779_1), .d(_net_6552), .o(n6795) );
oa22f01 g0066 ( .a(n6795), .b(n6792), .c(n6794), .d(n6793_1), .o(n6796_1) );
no02f01 g0067 ( .a(n6796_1), .b(n6791), .o(n6797) );
na02f01 g0068 ( .a(n6797), .b(n6786), .o(n281) );
in01f01 g0069 ( .a(_net_7797), .o(n6799) );
in01f01 g0070 ( .a(x1322), .o(n6800) );
in01f01 g0071 ( .a(x1286), .o(n6801_1) );
no02f01 g0072 ( .a(n6801_1), .b(x1261), .o(n6802) );
na03f01 g0073 ( .a(n6802), .b(_net_6184), .c(n6800), .o(n6803) );
na02f01 g0074 ( .a(n6803), .b(_net_6032), .o(n6804) );
oa12f01 g0075 ( .a(n6804), .b(n6803), .c(n6799), .o(n295) );
in01f01 g0076 ( .a(_net_6958), .o(n6806_1) );
na02f01 g0077 ( .a(n6806_1), .b(_net_6959), .o(n6807) );
in01f01 g0078 ( .a(n6807), .o(n6808) );
in01f01 g0079 ( .a(_net_6959), .o(n6809_1) );
na02f01 g0080 ( .a(n6806_1), .b(n6809_1), .o(n6810) );
in01f01 g0081 ( .a(n6810), .o(n6811) );
ao22f01 g0082 ( .a(n6811), .b(net_6834), .c(n6808), .d(net_6898), .o(n6812) );
na02f01 g0083 ( .a(_net_6958), .b(_net_6959), .o(n6813_1) );
in01f01 g0084 ( .a(n6813_1), .o(n6814) );
na02f01 g0085 ( .a(_net_6958), .b(n6809_1), .o(n6815) );
in01f01 g0086 ( .a(n6815), .o(n6816) );
ao22f01 g0087 ( .a(n6816), .b(net_6866), .c(n6814), .d(net_6930), .o(n6817) );
in01f01 g0088 ( .a(_net_6957), .o(n6818_1) );
in01f01 g0089 ( .a(_net_6017), .o(n6819) );
in01f01 g0090 ( .a(_net_7755), .o(n6820) );
na03f01 g0091 ( .a(net_6058), .b(n6820), .c(_net_7791), .o(n6821) );
no02f01 g0092 ( .a(n6821), .b(n6819), .o(n6822_1) );
no02f01 g0093 ( .a(_net_6020), .b(_net_6019), .o(n6823) );
na03f01 g0094 ( .a(n6823), .b(n6822_1), .c(n6818_1), .o(n6824) );
ao12f01 g0095 ( .a(n6824), .b(n6817), .c(n6812), .o(n6825) );
na02f01 g0096 ( .a(n6822_1), .b(_net_6019), .o(n6826_1) );
in01f01 g0097 ( .a(net_6900), .o(n6827) );
in01f01 g0098 ( .a(net_6836), .o(n6828) );
oa22f01 g0099 ( .a(n6810), .b(n6828), .c(n6807), .d(n6827), .o(n6829) );
in01f01 g0100 ( .a(net_6868), .o(n6830) );
in01f01 g0101 ( .a(net_6932), .o(n6831_1) );
oa22f01 g0102 ( .a(n6815), .b(n6830), .c(n6813_1), .d(n6831_1), .o(n6832) );
no02f01 g0103 ( .a(n6832), .b(n6829), .o(n6833) );
no02f01 g0104 ( .a(n6833), .b(n6826_1), .o(n6834) );
in01f01 g0105 ( .a(_net_6133), .o(n6835) );
na02f01 g0106 ( .a(n6822_1), .b(_net_6020), .o(n6836_1) );
in01f01 g0107 ( .a(net_6902), .o(n6837) );
in01f01 g0108 ( .a(net_6838), .o(n6838) );
oa22f01 g0109 ( .a(n6810), .b(n6838), .c(n6807), .d(n6837), .o(n6839) );
in01f01 g0110 ( .a(net_6870), .o(n6840_1) );
in01f01 g0111 ( .a(net_6934), .o(n6841) );
oa22f01 g0112 ( .a(n6815), .b(n6840_1), .c(n6813_1), .d(n6841), .o(n6842) );
no02f01 g0113 ( .a(n6842), .b(n6839), .o(n6843) );
na02f01 g0114 ( .a(n6821), .b(_net_6017), .o(n6844) );
oa22f01 g0115 ( .a(n6844), .b(n6835), .c(n6843), .d(n6836_1), .o(n6845_1) );
no03f01 g0116 ( .a(n6845_1), .b(n6834), .c(n6825), .o(n6846) );
in01f01 g0117 ( .a(net_6850), .o(n6847) );
in01f01 g0118 ( .a(net_6882), .o(n6848) );
na04f01 g0119 ( .a(n6823), .b(n6822_1), .c(n6816), .d(_net_6957), .o(n6849) );
na04f01 g0120 ( .a(n6823), .b(n6822_1), .c(n6811), .d(_net_6957), .o(n6850_1) );
oa22f01 g0121 ( .a(n6850_1), .b(n6847), .c(n6849), .d(n6848), .o(n6851) );
in01f01 g0122 ( .a(net_6914), .o(n6852) );
in01f01 g0123 ( .a(net_6946), .o(n6853) );
na04f01 g0124 ( .a(n6823), .b(n6822_1), .c(n6808), .d(_net_6957), .o(n6854) );
na04f01 g0125 ( .a(n6823), .b(n6822_1), .c(n6814), .d(_net_6957), .o(n6855_1) );
oa22f01 g0126 ( .a(n6855_1), .b(n6853), .c(n6854), .d(n6852), .o(n6856) );
no02f01 g0127 ( .a(n6856), .b(n6851), .o(n6857) );
na02f01 g0128 ( .a(n6857), .b(n6846), .o(n300) );
in01f01 g0129 ( .a(_net_7481), .o(n6859) );
in01f01 g0130 ( .a(_net_7534), .o(n6860_1) );
no02f01 g0131 ( .a(_net_7533), .b(n6860_1), .o(n6861) );
in01f01 g0132 ( .a(n6861), .o(n6862) );
in01f01 g0133 ( .a(_net_5920), .o(n6863_1) );
in01f01 g0134 ( .a(net_5860), .o(n6864) );
no03f01 g0135 ( .a(n6864), .b(n6863_1), .c(_net_7763), .o(n6865) );
no02f01 g0136 ( .a(_net_281), .b(_net_280), .o(n6866) );
in01f01 g0137 ( .a(n6866), .o(n6867_1) );
oa12f01 g0138 ( .a(n6865), .b(n6867_1), .c(_net_7532), .o(n6868) );
no02f01 g0139 ( .a(n6868), .b(n6862), .o(n6869) );
na02f01 g0140 ( .a(n6866), .b(net_350), .o(n6870) );
ao22f01 g0141 ( .a(_net_281), .b(net_362), .c(net_364), .d(_net_280), .o(n6871) );
na02f01 g0142 ( .a(n6871), .b(n6870), .o(n6872_1) );
na02f01 g0143 ( .a(n6872_1), .b(n6869), .o(n6873) );
oa12f01 g0144 ( .a(n6873), .b(n6869), .c(n6859), .o(n314) );
in01f01 g0145 ( .a(_net_7379), .o(n6875) );
no02f01 g0146 ( .a(net_7378), .b(n6875), .o(n6876_1) );
no02f01 g0147 ( .a(net_7378), .b(_net_7379), .o(n6877) );
ao22f01 g0148 ( .a(n6877), .b(_net_7269), .c(n6876_1), .d(_net_7333), .o(n6878) );
in01f01 g0149 ( .a(net_7378), .o(n6879) );
no02f01 g0150 ( .a(n6879), .b(n6875), .o(n6880) );
no02f01 g0151 ( .a(n6879), .b(_net_7379), .o(n6881_1) );
ao22f01 g0152 ( .a(n6881_1), .b(_net_7301), .c(n6880), .d(_net_7365), .o(n6882) );
na02f01 g0153 ( .a(n6882), .b(n6878), .o(n319) );
in01f01 g0154 ( .a(_net_6062), .o(n6884) );
in01f01 g0155 ( .a(net_155), .o(n6885) );
oa12f01 g0156 ( .a(_net_7791), .b(net_155), .c(net_7767), .o(n6886_1) );
oa22f01 g0157 ( .a(n6886_1), .b(n6885), .c(_net_7791), .d(n6884), .o(n329) );
in01f01 g0158 ( .a(_net_7474), .o(n6888) );
na02f01 g0159 ( .a(n6866), .b(net_7394), .o(n6889) );
ao22f01 g0160 ( .a(_net_281), .b(net_355), .c(_net_280), .d(net_357), .o(n6890_1) );
na02f01 g0161 ( .a(n6890_1), .b(n6889), .o(n6891) );
na02f01 g0162 ( .a(n6891), .b(n6869), .o(n6892) );
oa12f01 g0163 ( .a(n6892), .b(n6869), .c(n6888), .o(n370) );
in01f01 g0164 ( .a(_net_7252), .o(n6894) );
in01f01 g0165 ( .a(net_5861), .o(n6895_1) );
in01f01 g0166 ( .a(_net_5922), .o(n6896) );
no03f01 g0167 ( .a(_net_7761), .b(n6896), .c(n6895_1), .o(n6897) );
no02f01 g0168 ( .a(_net_269), .b(_net_270), .o(n6898) );
in01f01 g0169 ( .a(n6898), .o(n6899_1) );
oa12f01 g0170 ( .a(n6897), .b(n6899_1), .c(_net_7381), .o(n6900) );
no03f01 g0171 ( .a(n6900), .b(_net_7383), .c(_net_7382), .o(n6901) );
na02f01 g0172 ( .a(n6898), .b(net_7236), .o(n6902_1) );
ao22f01 g0173 ( .a(net_328), .b(_net_270), .c(net_330), .d(_net_269), .o(n6903) );
na02f01 g0174 ( .a(n6903), .b(n6902_1), .o(n6904) );
na02f01 g0175 ( .a(n6904), .b(n6901), .o(n6905) );
oa12f01 g0176 ( .a(n6905), .b(n6901), .c(n6894), .o(n375) );
in01f01 g0177 ( .a(_net_298), .o(n6907) );
na02f01 g0178 ( .a(_net_262), .b(_net_264), .o(n6908) );
na02f01 g0179 ( .a(n6908), .b(n6907), .o(n380) );
in01f01 g0180 ( .a(x38), .o(n6910_1) );
na02f01 g0181 ( .a(n6910_1), .b(_net_6404), .o(n385) );
in01f01 g0182 ( .a(_net_5995), .o(n6912) );
in01f01 g0183 ( .a(_net_7751), .o(n6913) );
na03f01 g0184 ( .a(_net_7791), .b(n6913), .c(net_6060), .o(n6914) );
no02f01 g0185 ( .a(n6914), .b(n6912), .o(n6915_1) );
na02f01 g0186 ( .a(n6915_1), .b(_net_5998), .o(n6916) );
in01f01 g0187 ( .a(n6916), .o(n6917) );
in01f01 g0188 ( .a(_net_6688), .o(n6918) );
na02f01 g0189 ( .a(_net_6689), .b(n6918), .o(n6919_1) );
in01f01 g0190 ( .a(n6919_1), .o(n6920) );
in01f01 g0191 ( .a(_net_6689), .o(n6921) );
na02f01 g0192 ( .a(n6921), .b(n6918), .o(n6922) );
in01f01 g0193 ( .a(n6922), .o(n6923) );
ao22f01 g0194 ( .a(n6923), .b(net_6563), .c(n6920), .d(net_6627), .o(n6924_1) );
na02f01 g0195 ( .a(_net_6689), .b(_net_6688), .o(n6925) );
in01f01 g0196 ( .a(n6925), .o(n6926) );
na02f01 g0197 ( .a(n6921), .b(_net_6688), .o(n6927) );
in01f01 g0198 ( .a(n6927), .o(n6928) );
ao22f01 g0199 ( .a(n6928), .b(net_6595), .c(n6926), .d(net_6659), .o(n6929_1) );
na02f01 g0200 ( .a(n6929_1), .b(n6924_1), .o(n6930) );
na02f01 g0201 ( .a(n6930), .b(n6917), .o(n6931) );
na02f01 g0202 ( .a(n6914), .b(_net_5995), .o(n6932) );
in01f01 g0203 ( .a(n6932), .o(n6933) );
na02f01 g0204 ( .a(n6915_1), .b(_net_5997), .o(n6934_1) );
in01f01 g0205 ( .a(n6934_1), .o(n6935) );
ao22f01 g0206 ( .a(n6923), .b(net_6561), .c(n6920), .d(net_6625), .o(n6936) );
ao22f01 g0207 ( .a(n6928), .b(net_6593), .c(n6926), .d(net_6657), .o(n6937) );
na02f01 g0208 ( .a(n6937), .b(n6936), .o(n6938_1) );
ao22f01 g0209 ( .a(n6938_1), .b(n6935), .c(n6933), .d(_net_6088), .o(n6939) );
ao22f01 g0210 ( .a(n6923), .b(net_6559), .c(n6920), .d(net_6623), .o(n6940) );
ao22f01 g0211 ( .a(n6928), .b(net_6591), .c(n6926), .d(net_6655), .o(n6941) );
na02f01 g0212 ( .a(n6941), .b(n6940), .o(n6942) );
in01f01 g0213 ( .a(_net_6687), .o(n6943_1) );
no02f01 g0214 ( .a(_net_5998), .b(_net_5997), .o(n6944) );
na03f01 g0215 ( .a(n6944), .b(n6915_1), .c(n6943_1), .o(n6945) );
in01f01 g0216 ( .a(n6945), .o(n6946) );
na02f01 g0217 ( .a(n6944), .b(n6915_1), .o(n6947_1) );
in01f01 g0218 ( .a(net_6639), .o(n6948) );
in01f01 g0219 ( .a(net_6575), .o(n6949) );
oa22f01 g0220 ( .a(n6922), .b(n6949), .c(n6919_1), .d(n6948), .o(n6950) );
in01f01 g0221 ( .a(net_6671), .o(n6951) );
in01f01 g0222 ( .a(net_6607), .o(n6952_1) );
oa22f01 g0223 ( .a(n6927), .b(n6952_1), .c(n6925), .d(n6951), .o(n6953) );
no02f01 g0224 ( .a(n6953), .b(n6950), .o(n6954) );
no03f01 g0225 ( .a(n6954), .b(n6947_1), .c(n6943_1), .o(n6955) );
ao12f01 g0226 ( .a(n6955), .b(n6946), .c(n6942), .o(n6956) );
na03f01 g0227 ( .a(n6956), .b(n6939), .c(n6931), .o(n390) );
in01f01 g0228 ( .a(_net_7595), .o(n6958) );
in01f01 g0229 ( .a(_net_7684), .o(n6959) );
no02f01 g0230 ( .a(_net_7685), .b(n6959), .o(n6960_1) );
in01f01 g0231 ( .a(n6960_1), .o(n6961) );
in01f01 g0232 ( .a(net_5858), .o(n6962) );
in01f01 g0233 ( .a(_net_5924), .o(n6963) );
no03f01 g0234 ( .a(n6963), .b(n6962), .c(_net_7765), .o(n6964_1) );
no02f01 g0235 ( .a(_net_292), .b(_net_291), .o(n6965) );
in01f01 g0236 ( .a(n6965), .o(n6966) );
oa12f01 g0237 ( .a(n6964_1), .b(n6966), .c(_net_7683), .o(n6967) );
no02f01 g0238 ( .a(n6967), .b(n6961), .o(n6968) );
na02f01 g0239 ( .a(n6965), .b(net_7547), .o(n6969_1) );
ao22f01 g0240 ( .a(_net_292), .b(net_377), .c(_net_291), .d(net_379), .o(n6970) );
na02f01 g0241 ( .a(n6970), .b(n6969_1), .o(n6971) );
na02f01 g0242 ( .a(n6971), .b(n6968), .o(n6972) );
oa12f01 g0243 ( .a(n6972), .b(n6968), .c(n6958), .o(n400) );
in01f01 g0244 ( .a(net_362), .o(n6974_1) );
no02f01 g0245 ( .a(n6867_1), .b(n6974_1), .o(n420) );
in01f01 g0246 ( .a(_net_6028), .o(n6976) );
in01f01 g0247 ( .a(_net_7757), .o(n6977_1) );
na03f01 g0248 ( .a(n6977_1), .b(_net_7791), .c(net_6057), .o(n6978) );
no02f01 g0249 ( .a(n6978), .b(n6976), .o(n6979) );
na02f01 g0250 ( .a(n6979), .b(_net_6031), .o(n6980) );
in01f01 g0251 ( .a(n6980), .o(n6981) );
in01f01 g0252 ( .a(net_7034), .o(n6982_1) );
in01f01 g0253 ( .a(net_6970), .o(n6983) );
in01f01 g0254 ( .a(_net_7093), .o(n6984) );
na02f01 g0255 ( .a(n6984), .b(_net_7094), .o(n6985) );
in01f01 g0256 ( .a(_net_7094), .o(n6986_1) );
na02f01 g0257 ( .a(n6984), .b(n6986_1), .o(n6987) );
oa22f01 g0258 ( .a(n6987), .b(n6983), .c(n6985), .d(n6982_1), .o(n6988) );
in01f01 g0259 ( .a(net_7066), .o(n6989) );
in01f01 g0260 ( .a(net_7002), .o(n6990_1) );
na02f01 g0261 ( .a(_net_7093), .b(_net_7094), .o(n6991) );
na02f01 g0262 ( .a(_net_7093), .b(n6986_1), .o(n6992) );
oa22f01 g0263 ( .a(n6992), .b(n6990_1), .c(n6991), .d(n6989), .o(n6993) );
oa12f01 g0264 ( .a(n6981), .b(n6993), .c(n6988), .o(n6994) );
na02f01 g0265 ( .a(n6978), .b(_net_6028), .o(n6995_1) );
in01f01 g0266 ( .a(n6995_1), .o(n6996) );
na02f01 g0267 ( .a(n6979), .b(_net_6030), .o(n6997) );
in01f01 g0268 ( .a(n6997), .o(n6998) );
in01f01 g0269 ( .a(n6985), .o(n6999) );
in01f01 g0270 ( .a(n6987), .o(n7000_1) );
ao22f01 g0271 ( .a(n7000_1), .b(net_6968), .c(n6999), .d(net_7032), .o(n7001) );
in01f01 g0272 ( .a(n6991), .o(n7002) );
in01f01 g0273 ( .a(n6992), .o(n7003) );
ao22f01 g0274 ( .a(n7003), .b(net_7000), .c(n7002), .d(net_7064), .o(n7004) );
na02f01 g0275 ( .a(n7004), .b(n7001), .o(n7005_1) );
ao22f01 g0276 ( .a(n7005_1), .b(n6998), .c(n6996), .d(_net_6150), .o(n7006) );
ao22f01 g0277 ( .a(n7000_1), .b(net_6966), .c(n6999), .d(net_7030), .o(n7007) );
ao22f01 g0278 ( .a(n7003), .b(net_6998), .c(n7002), .d(net_7062), .o(n7008) );
na02f01 g0279 ( .a(n7008), .b(n7007), .o(n7009_1) );
in01f01 g0280 ( .a(_net_7092), .o(n7010) );
no02f01 g0281 ( .a(_net_6031), .b(_net_6030), .o(n7011) );
na03f01 g0282 ( .a(n7011), .b(n6979), .c(n7010), .o(n7012) );
in01f01 g0283 ( .a(n7012), .o(n7013_1) );
na02f01 g0284 ( .a(n7013_1), .b(n7009_1), .o(n7014) );
in01f01 g0285 ( .a(net_6982), .o(n7015) );
in01f01 g0286 ( .a(net_7046), .o(n7016) );
oa22f01 g0287 ( .a(n6987), .b(n7015), .c(n6985), .d(n7016), .o(n7017) );
in01f01 g0288 ( .a(net_7014), .o(n7018_1) );
in01f01 g0289 ( .a(net_7078), .o(n7019) );
oa22f01 g0290 ( .a(n6992), .b(n7018_1), .c(n6991), .d(n7019), .o(n7020) );
na02f01 g0291 ( .a(n7011), .b(n6979), .o(n7021) );
no02f01 g0292 ( .a(n7021), .b(n7010), .o(n7022) );
oa12f01 g0293 ( .a(n7022), .b(n7020), .c(n7017), .o(n7023_1) );
na04f01 g0294 ( .a(n7023_1), .b(n7014), .c(n7006), .d(n6994), .o(n447) );
in01f01 g0295 ( .a(_net_7355), .o(n7025) );
in01f01 g0296 ( .a(_net_7382), .o(n7026) );
in01f01 g0297 ( .a(_net_7383), .o(n7027_1) );
no02f01 g0298 ( .a(n7027_1), .b(n7026), .o(n7028) );
in01f01 g0299 ( .a(n7028), .o(n7029) );
no02f01 g0300 ( .a(n7029), .b(n6900), .o(n7030) );
na02f01 g0301 ( .a(n6898), .b(net_7243), .o(n7031) );
ao22f01 g0302 ( .a(net_335), .b(_net_270), .c(_net_269), .d(net_337), .o(n7032_1) );
na02f01 g0303 ( .a(n7032_1), .b(n7031), .o(n7033) );
na02f01 g0304 ( .a(n7033), .b(n7030), .o(n7034) );
oa12f01 g0305 ( .a(n7034), .b(n7030), .c(n7025), .o(n460) );
in01f01 g0306 ( .a(net_6635), .o(n7036_1) );
in01f01 g0307 ( .a(net_6571), .o(n7037) );
oa22f01 g0308 ( .a(n6922), .b(n7037), .c(n6919_1), .d(n7036_1), .o(n7038) );
in01f01 g0309 ( .a(net_6603), .o(n7039) );
in01f01 g0310 ( .a(net_6667), .o(n7040) );
oa22f01 g0311 ( .a(n6927), .b(n7039), .c(n6925), .d(n7040), .o(n7041_1) );
no02f01 g0312 ( .a(n7041_1), .b(n7038), .o(n7042) );
no02f01 g0313 ( .a(n7042), .b(n6945), .o(n7043) );
in01f01 g0314 ( .a(net_6637), .o(n7044) );
in01f01 g0315 ( .a(net_6573), .o(n7045_1) );
oa22f01 g0316 ( .a(n6922), .b(n7045_1), .c(n6919_1), .d(n7044), .o(n7046) );
in01f01 g0317 ( .a(net_6605), .o(n7047) );
in01f01 g0318 ( .a(net_6669), .o(n7048) );
oa22f01 g0319 ( .a(n6927), .b(n7047), .c(n6925), .d(n7048), .o(n7049_1) );
no02f01 g0320 ( .a(n7049_1), .b(n7046), .o(n7050) );
no02f01 g0321 ( .a(n7050), .b(n6934_1), .o(n7051) );
in01f01 g0322 ( .a(_net_6100), .o(n7052) );
oa22f01 g0323 ( .a(n6954), .b(n6916), .c(n6932), .d(n7052), .o(n7053_1) );
no03f01 g0324 ( .a(n7053_1), .b(n7051), .c(n7043), .o(n7054) );
in01f01 g0325 ( .a(net_6619), .o(n7055) );
in01f01 g0326 ( .a(net_6587), .o(n7056) );
na04f01 g0327 ( .a(n6944), .b(n6928), .c(n6915_1), .d(_net_6687), .o(n7057) );
na04f01 g0328 ( .a(n6944), .b(n6923), .c(n6915_1), .d(_net_6687), .o(n7058_1) );
oa22f01 g0329 ( .a(n7058_1), .b(n7056), .c(n7057), .d(n7055), .o(n7059) );
in01f01 g0330 ( .a(net_6651), .o(n7060) );
in01f01 g0331 ( .a(net_6683), .o(n7061) );
na04f01 g0332 ( .a(n6944), .b(n6920), .c(n6915_1), .d(_net_6687), .o(n7062_1) );
na04f01 g0333 ( .a(n6944), .b(n6926), .c(n6915_1), .d(_net_6687), .o(n7063) );
oa22f01 g0334 ( .a(n7063), .b(n7061), .c(n7062_1), .d(n7060), .o(n7064) );
no02f01 g0335 ( .a(n7064), .b(n7059), .o(n7065) );
na02f01 g0336 ( .a(n7065), .b(n7054), .o(n465) );
in01f01 g0337 ( .a(_net_5967), .o(n7067_1) );
no02f01 g0338 ( .a(n6912), .b(n7067_1), .o(n513) );
in01f01 g0339 ( .a(net_337), .o(n7069) );
no02f01 g0340 ( .a(n6899_1), .b(n7069), .o(n518) );
in01f01 g0341 ( .a(net_6435), .o(n7071) );
in01f01 g0342 ( .a(net_6499), .o(n7072_1) );
oa22f01 g0343 ( .a(n6750), .b(n7071), .c(n6748), .d(n7072_1), .o(n7073) );
in01f01 g0344 ( .a(net_6467), .o(n7074) );
in01f01 g0345 ( .a(net_6531), .o(n7075) );
oa22f01 g0346 ( .a(n6755), .b(n7074), .c(n6754), .d(n7075), .o(n7076) );
no02f01 g0347 ( .a(n7076), .b(n7073), .o(n7077_1) );
no02f01 g0348 ( .a(n7077_1), .b(n6764), .o(n7078) );
in01f01 g0349 ( .a(net_6501), .o(n7079) );
in01f01 g0350 ( .a(net_6437), .o(n7080) );
oa22f01 g0351 ( .a(n6750), .b(n7080), .c(n6748), .d(n7079), .o(n7081) );
in01f01 g0352 ( .a(net_6469), .o(n7082_1) );
in01f01 g0353 ( .a(net_6533), .o(n7083) );
oa22f01 g0354 ( .a(n6755), .b(n7082_1), .c(n6754), .d(n7083), .o(n7084) );
no02f01 g0355 ( .a(n7084), .b(n7081), .o(n7085_1) );
no02f01 g0356 ( .a(n7085_1), .b(n6766), .o(n7086) );
in01f01 g0357 ( .a(_net_6079), .o(n7087) );
in01f01 g0358 ( .a(net_6439), .o(n7088) );
in01f01 g0359 ( .a(net_6503), .o(n7089_1) );
oa22f01 g0360 ( .a(n6750), .b(n7088), .c(n6748), .d(n7089_1), .o(n7090) );
in01f01 g0361 ( .a(net_6471), .o(n7091) );
in01f01 g0362 ( .a(net_6535), .o(n7092) );
oa22f01 g0363 ( .a(n6755), .b(n7091), .c(n6754), .d(n7092), .o(n7093_1) );
no02f01 g0364 ( .a(n7093_1), .b(n7090), .o(n7094) );
oa22f01 g0365 ( .a(n7094), .b(n6775), .c(n6784), .d(n7087), .o(n7095) );
no03f01 g0366 ( .a(n7095), .b(n7086), .c(n7078), .o(n7096) );
in01f01 g0367 ( .a(net_6451), .o(n7097) );
in01f01 g0368 ( .a(net_6483), .o(n7098_1) );
oa22f01 g0369 ( .a(n6790), .b(n7097), .c(n6789), .d(n7098_1), .o(n7099) );
in01f01 g0370 ( .a(net_6515), .o(n7100) );
in01f01 g0371 ( .a(net_6547), .o(n7101) );
oa22f01 g0372 ( .a(n6795), .b(n7101), .c(n6794), .d(n7100), .o(n7102_1) );
no02f01 g0373 ( .a(n7102_1), .b(n7099), .o(n7103) );
na02f01 g0374 ( .a(n7103), .b(n7096), .o(n523) );
in01f01 g0375 ( .a(x1155), .o(n7105) );
in01f01 g0376 ( .a(x1101), .o(n7106) );
in01f01 g0377 ( .a(x1126), .o(n7107_1) );
no02f01 g0378 ( .a(n7107_1), .b(n7106), .o(n7108) );
in01f01 g0379 ( .a(_net_7689), .o(n7109) );
no03f01 g0380 ( .a(_net_7690), .b(n7109), .c(n7105), .o(n7110) );
na02f01 g0381 ( .a(n7110), .b(n7108), .o(n7111_1) );
in01f01 g0382 ( .a(n7111_1), .o(n7112) );
no03f01 g0383 ( .a(x1193), .b(x1209), .c(x1203), .o(n7113) );
na02f01 g0384 ( .a(n7113), .b(n7108), .o(n7114) );
no03f01 g0385 ( .a(n7114), .b(n7112), .c(n7105), .o(n528) );
in01f01 g0386 ( .a(_net_7753), .o(n7116_1) );
na03f01 g0387 ( .a(_net_7791), .b(net_6059), .c(n7116_1), .o(n7117) );
na02f01 g0388 ( .a(n7117), .b(_net_6006), .o(n7118) );
in01f01 g0389 ( .a(n7118), .o(n7119) );
na02f01 g0390 ( .a(n7119), .b(_net_6104), .o(n7120_1) );
in01f01 g0391 ( .a(_net_6006), .o(n7121) );
no02f01 g0392 ( .a(n7117), .b(n7121), .o(n7122) );
na02f01 g0393 ( .a(n7122), .b(_net_6009), .o(n7123) );
in01f01 g0394 ( .a(n7123), .o(n7124) );
in01f01 g0395 ( .a(_net_6823), .o(n7125_1) );
na02f01 g0396 ( .a(_net_6824), .b(n7125_1), .o(n7126) );
in01f01 g0397 ( .a(n7126), .o(n7127) );
in01f01 g0398 ( .a(_net_6824), .o(n7128_1) );
na02f01 g0399 ( .a(n7128_1), .b(n7125_1), .o(n7129) );
in01f01 g0400 ( .a(n7129), .o(n7130) );
ao22f01 g0401 ( .a(n7130), .b(net_6694), .c(n7127), .d(net_6758), .o(n7131) );
na02f01 g0402 ( .a(_net_6824), .b(_net_6823), .o(n7132) );
in01f01 g0403 ( .a(n7132), .o(n7133_1) );
na02f01 g0404 ( .a(n7128_1), .b(_net_6823), .o(n7134) );
in01f01 g0405 ( .a(n7134), .o(n7135) );
ao22f01 g0406 ( .a(n7135), .b(net_6726), .c(n7133_1), .d(net_6790), .o(n7136) );
na02f01 g0407 ( .a(n7136), .b(n7131), .o(n7137) );
na02f01 g0408 ( .a(n7137), .b(n7124), .o(n7138_1) );
na02f01 g0409 ( .a(n7138_1), .b(n7120_1), .o(n533) );
in01f01 g0410 ( .a(_net_7603), .o(n7140) );
in01f01 g0411 ( .a(net_373), .o(n7141) );
in01f01 g0412 ( .a(net_385), .o(n7142_1) );
in01f01 g0413 ( .a(_net_292), .o(n7143) );
oa22f01 g0414 ( .a(n6966), .b(n7141), .c(n7143), .d(n7142_1), .o(n7144) );
na02f01 g0415 ( .a(n7144), .b(n6968), .o(n7145) );
oa12f01 g0416 ( .a(n7145), .b(n6968), .c(n7140), .o(n538) );
in01f01 g0417 ( .a(_net_7316), .o(n7147_1) );
no02f01 g0418 ( .a(n7027_1), .b(_net_7382), .o(n7148) );
in01f01 g0419 ( .a(n7148), .o(n7149) );
no02f01 g0420 ( .a(n7149), .b(n6900), .o(n7150) );
na02f01 g0421 ( .a(n7150), .b(n6904), .o(n7151_1) );
oa12f01 g0422 ( .a(n7151_1), .b(n7150), .c(n7147_1), .o(n543) );
in01f01 g0423 ( .a(net_6691), .o(n7153) );
no02f01 g0424 ( .a(n6918), .b(n7153), .o(n7154) );
no02f01 g0425 ( .a(_net_6688), .b(net_6691), .o(n7155_1) );
no02f01 g0426 ( .a(n7155_1), .b(n7154), .o(n7156) );
in01f01 g0427 ( .a(n7156), .o(n548) );
in01f01 g0428 ( .a(net_6057), .o(n7158) );
in01f01 g0429 ( .a(net_6061), .o(n7159) );
in01f01 g0430 ( .a(net_6056), .o(n7160_1) );
in01f01 g0431 ( .a(net_6058), .o(n7161) );
na04f01 g0432 ( .a(n7161), .b(n7160_1), .c(n7159), .d(n7158), .o(n7162) );
in01f01 g0433 ( .a(net_6060), .o(n7163) );
in01f01 g0434 ( .a(net_6059), .o(n7164_1) );
in01f01 g0435 ( .a(_net_6063), .o(n7165) );
na04f01 g0436 ( .a(n7165), .b(n7164_1), .c(n7163), .d(n6884), .o(n7166) );
oa12f01 g0437 ( .a(_net_392), .b(n7166), .c(n7162), .o(n7167_1) );
in01f01 g0438 ( .a(_net_392), .o(n7168) );
na02f01 g0439 ( .a(n7168), .b(_net_6199), .o(n7169) );
na02f01 g0440 ( .a(n7169), .b(n7167_1), .o(n553) );
in01f01 g0441 ( .a(_net_6293), .o(n7171) );
no02f01 g0442 ( .a(_net_392), .b(n7171), .o(n561) );
in01f01 g0443 ( .a(net_342), .o(n7173) );
no02f01 g0444 ( .a(n6899_1), .b(n7173), .o(n576) );
in01f01 g0445 ( .a(net_361), .o(n7175) );
no02f01 g0446 ( .a(n6867_1), .b(n7175), .o(n595) );
in01f01 g0447 ( .a(_net_7285), .o(n7177_1) );
no02f01 g0448 ( .a(_net_7383), .b(n7026), .o(n7178) );
in01f01 g0449 ( .a(n7178), .o(n7179) );
no02f01 g0450 ( .a(n7179), .b(n6900), .o(n7180) );
na02f01 g0451 ( .a(n6898), .b(net_7237), .o(n7181) );
ao22f01 g0452 ( .a(_net_269), .b(net_331), .c(_net_270), .d(net_329), .o(n7182_1) );
na02f01 g0453 ( .a(n7182_1), .b(n7181), .o(n7183) );
na02f01 g0454 ( .a(n7183), .b(n7180), .o(n7184) );
oa12f01 g0455 ( .a(n7184), .b(n7180), .c(n7177_1), .o(n600) );
in01f01 g0456 ( .a(_net_6209), .o(n7186) );
no02f01 g0457 ( .a(_net_392), .b(n7186), .o(n605) );
in01f01 g0458 ( .a(net_374), .o(n7188) );
no02f01 g0459 ( .a(n6966), .b(n7188), .o(n615) );
in01f01 g0460 ( .a(_net_6004), .o(n7190_1) );
in01f01 g0461 ( .a(_net_5964), .o(n7191) );
oa12f01 g0462 ( .a(n7190_1), .b(n6914), .c(n7191), .o(n620) );
in01f01 g0463 ( .a(_net_7441), .o(n7193) );
in01f01 g0464 ( .a(_net_7533), .o(n7194_1) );
no02f01 g0465 ( .a(n7194_1), .b(_net_7534), .o(n7195) );
in01f01 g0466 ( .a(n7195), .o(n7196) );
no02f01 g0467 ( .a(n7196), .b(n6868), .o(n7197) );
na02f01 g0468 ( .a(n6866), .b(net_7393), .o(n7198) );
ao22f01 g0469 ( .a(net_354), .b(_net_281), .c(net_356), .d(_net_280), .o(n7199_1) );
na02f01 g0470 ( .a(n7199_1), .b(n7198), .o(n7200) );
na02f01 g0471 ( .a(n7200), .b(n7197), .o(n7201) );
oa12f01 g0472 ( .a(n7201), .b(n7197), .c(n7193), .o(n629) );
in01f01 g0473 ( .a(net_356), .o(n7203_1) );
no02f01 g0474 ( .a(n6867_1), .b(n7203_1), .o(n634) );
in01f01 g0475 ( .a(_net_7694), .o(n7205) );
na02f01 g0476 ( .a(_net_6184), .b(x1261), .o(n7206) );
no03f01 g0477 ( .a(n7206), .b(x1286), .c(n6800), .o(n7207_1) );
na02f01 g0478 ( .a(n7207_1), .b(_net_7796), .o(n7208) );
oa12f01 g0479 ( .a(n7208), .b(n7207_1), .c(n7205), .o(n639) );
no02f01 g0480 ( .a(n7010), .b(n6984), .o(n7210) );
na02f01 g0481 ( .a(n7210), .b(n6986_1), .o(n7211) );
in01f01 g0482 ( .a(n7210), .o(n7212_1) );
na02f01 g0483 ( .a(n7212_1), .b(_net_7094), .o(n7213) );
na02f01 g0484 ( .a(n7213), .b(n7211), .o(n7214) );
no04f01 g0485 ( .a(n6978), .b(_net_6031), .c(n6976), .d(_net_6030), .o(n7215) );
na02f01 g0486 ( .a(n7215), .b(n7214), .o(n7216_1) );
na02f01 g0487 ( .a(n6992), .b(n6985), .o(n7217) );
no03f01 g0488 ( .a(n7011), .b(n6978), .c(n6976), .o(n7218) );
in01f01 g0489 ( .a(n6978), .o(n7219) );
no02f01 g0490 ( .a(n7219), .b(n6976), .o(n7220) );
ao22f01 g0491 ( .a(n7220), .b(_net_7094), .c(n7218), .d(n7217), .o(n7221_1) );
na02f01 g0492 ( .a(n7221_1), .b(n7216_1), .o(n644) );
in01f01 g0493 ( .a(net_7529), .o(n7223) );
no02f01 g0494 ( .a(_net_7530), .b(n7223), .o(n7224) );
no02f01 g0495 ( .a(_net_7530), .b(net_7529), .o(n7225) );
ao22f01 g0496 ( .a(n7225), .b(_net_7420), .c(n7224), .d(_net_7452), .o(n7226_1) );
in01f01 g0497 ( .a(_net_7530), .o(n7227) );
no02f01 g0498 ( .a(n7227), .b(net_7529), .o(n7228) );
no02f01 g0499 ( .a(n7227), .b(n7223), .o(n7229) );
ao22f01 g0500 ( .a(n7229), .b(_net_7516), .c(n7228), .d(_net_7484), .o(n7230_1) );
na02f01 g0501 ( .a(n7230_1), .b(n7226_1), .o(n649) );
in01f01 g0502 ( .a(_net_7791), .o(n7232) );
no02f01 g0503 ( .a(n7232), .b(n7164_1), .o(n654) );
ao22f01 g0504 ( .a(n6877), .b(_net_7254), .c(n6876_1), .d(_net_7318), .o(n7234) );
ao22f01 g0505 ( .a(n6881_1), .b(_net_7286), .c(n6880), .d(_net_7350), .o(n7235_1) );
na02f01 g0506 ( .a(n7235_1), .b(n7234), .o(n659) );
in01f01 g0507 ( .a(_net_6207), .o(n7237) );
no02f01 g0508 ( .a(_net_392), .b(n7237), .o(n673) );
in01f01 g0509 ( .a(_net_7330), .o(n7239) );
na02f01 g0510 ( .a(n6898), .b(net_330), .o(n7240_1) );
ao22f01 g0511 ( .a(net_344), .b(_net_269), .c(net_342), .d(_net_270), .o(n7241) );
na02f01 g0512 ( .a(n7241), .b(n7240_1), .o(n7242) );
na02f01 g0513 ( .a(n7242), .b(n7150), .o(n7243) );
oa12f01 g0514 ( .a(n7243), .b(n7150), .c(n7239), .o(n688) );
in01f01 g0515 ( .a(_net_7271), .o(n7245_1) );
in01f01 g0516 ( .a(net_335), .o(n7246) );
no02f01 g0517 ( .a(n6899_1), .b(n7246), .o(n1350) );
na02f01 g0518 ( .a(n1350), .b(n6901), .o(n7248) );
oa12f01 g0519 ( .a(n7248), .b(n6901), .c(n7245_1), .o(n693) );
in01f01 g0520 ( .a(net_383), .o(n7250) );
no02f01 g0521 ( .a(n6966), .b(n7250), .o(n698) );
in01f01 g0522 ( .a(_net_7300), .o(n7252_1) );
in01f01 g0523 ( .a(_net_270), .o(n7253) );
in01f01 g0524 ( .a(net_344), .o(n7254) );
in01f01 g0525 ( .a(net_332), .o(n7255) );
oa22f01 g0526 ( .a(n6899_1), .b(n7255), .c(n7254), .d(n7253), .o(n7256_1) );
na02f01 g0527 ( .a(n7256_1), .b(n7180), .o(n7257) );
oa12f01 g0528 ( .a(n7257), .b(n7180), .c(n7252_1), .o(n708) );
in01f01 g0529 ( .a(_net_6010), .o(n7259) );
no02f01 g0530 ( .a(n7259), .b(_net_6011), .o(n7260_1) );
in01f01 g0531 ( .a(_net_5968), .o(n7261) );
na02f01 g0532 ( .a(_net_6006), .b(_net_6012), .o(n7262) );
ao12f01 g0533 ( .a(n7262), .b(_net_5970), .c(n7261), .o(n7263) );
na02f01 g0534 ( .a(n7263), .b(n7260_1), .o(n7264) );
in01f01 g0535 ( .a(_net_6011), .o(n7265_1) );
in01f01 g0536 ( .a(n7262), .o(n7266) );
na03f01 g0537 ( .a(_net_5970), .b(n7261), .c(_net_5969), .o(n7267) );
na04f01 g0538 ( .a(n7267), .b(n7266), .c(n7259), .d(n7265_1), .o(n7268) );
oa12f01 g0539 ( .a(n7261), .b(_net_5970), .c(_net_5969), .o(n7269) );
na04f01 g0540 ( .a(n7269), .b(n7266), .c(n7259), .d(_net_6011), .o(n7270_1) );
no02f01 g0541 ( .a(n7259), .b(n7265_1), .o(n7271) );
na03f01 g0542 ( .a(n7271), .b(n7266), .c(_net_5968), .o(n7272) );
na04f01 g0543 ( .a(n7272), .b(n7270_1), .c(n7268), .d(n7264), .o(n7273) );
in01f01 g0544 ( .a(n7273), .o(n7274) );
no02f01 g0545 ( .a(n7274), .b(x1006), .o(n713) );
in01f01 g0546 ( .a(net_375), .o(n7276) );
no02f01 g0547 ( .a(n6966), .b(n7276), .o(n718) );
ao22f01 g0548 ( .a(n6738), .b(_net_7558), .c(n6736_1), .d(_net_7622), .o(n7278) );
ao22f01 g0549 ( .a(n6739), .b(_net_7654), .c(n6734), .d(_net_7590), .o(n7279) );
na02f01 g0550 ( .a(n7279), .b(n7278), .o(n727) );
in01f01 g0551 ( .a(x1215), .o(n7281) );
na04f01 g0552 ( .a(x1231), .b(x1286), .c(x1261), .d(n7281), .o(n7282) );
no02f01 g0553 ( .a(x1231), .b(x1261), .o(n7283) );
na04f01 g0554 ( .a(n7283), .b(n6801_1), .c(x1215), .d(n6800), .o(n7284_1) );
na04f01 g0555 ( .a(n7284_1), .b(n7282), .c(x1286), .d(x1322), .o(n7285) );
in01f01 g0556 ( .a(n7285), .o(n7286) );
na04f01 g0557 ( .a(n7284_1), .b(n7282), .c(n6802), .d(n6800), .o(n7287) );
in01f01 g0558 ( .a(n7287), .o(n7288_1) );
ao22f01 g0559 ( .a(n7288_1), .b(_net_6041), .c(n7286), .d(_net_280), .o(n7289) );
na04f01 g0560 ( .a(n7284_1), .b(n7282), .c(x1261), .d(x1322), .o(n7290) );
in01f01 g0561 ( .a(n7290), .o(n7291) );
na02f01 g0562 ( .a(x1286), .b(x1261), .o(n7292_1) );
no02f01 g0563 ( .a(n7282), .b(n6800), .o(n7293) );
in01f01 g0564 ( .a(n7283), .o(n7294) );
na03f01 g0565 ( .a(n6801_1), .b(x1215), .c(n6800), .o(n7295) );
no02f01 g0566 ( .a(n7295), .b(n7294), .o(n7296) );
no02f01 g0567 ( .a(n7282), .b(x1322), .o(n7297_1) );
no04f01 g0568 ( .a(n7297_1), .b(n7296), .c(n7293), .d(n7292_1), .o(n7298) );
ao22f01 g0569 ( .a(n7298), .b(_net_7730), .c(n7291), .d(_net_7701), .o(n7299) );
in01f01 g0570 ( .a(x1261), .o(n7300) );
na04f01 g0571 ( .a(n7284_1), .b(n7282), .c(n6801_1), .d(n6800), .o(n7301) );
no02f01 g0572 ( .a(n7301), .b(n7300), .o(n7302_1) );
na02f01 g0573 ( .a(n7302_1), .b(_net_124), .o(n7303) );
no02f01 g0574 ( .a(x1286), .b(x1261), .o(n7304) );
na04f01 g0575 ( .a(n7304), .b(n7284_1), .c(n7282), .d(x1322), .o(n7305) );
in01f01 g0576 ( .a(n7305), .o(n7306) );
na02f01 g0577 ( .a(x1231), .b(n7281), .o(n7307_1) );
no02f01 g0578 ( .a(n7307_1), .b(n7292_1), .o(n7308) );
na03f01 g0579 ( .a(n7308), .b(net_203), .c(x1322), .o(n7309) );
na02f01 g0580 ( .a(n7296), .b(net_240), .o(n7310) );
na03f01 g0581 ( .a(n7308), .b(net_166), .c(n6800), .o(n7311) );
na03f01 g0582 ( .a(n7311), .b(n7310), .c(n7309), .o(n7312_1) );
ao12f01 g0583 ( .a(n7312_1), .b(n7306), .c(_net_5997), .o(n7313) );
na04f01 g0584 ( .a(n7313), .b(n7303), .c(n7299), .d(n7289), .o(n732) );
in01f01 g0585 ( .a(_net_6037), .o(n7315) );
in01f01 g0586 ( .a(_net_5976), .o(n7316_1) );
oa12f01 g0587 ( .a(n7315), .b(n6978), .c(n7316_1), .o(n736) );
ao22f01 g0588 ( .a(n6738), .b(_net_7557), .c(n6736_1), .d(_net_7621), .o(n7318) );
ao22f01 g0589 ( .a(n6739), .b(_net_7653), .c(n6734), .d(_net_7589), .o(n7319) );
na02f01 g0590 ( .a(n7319), .b(n7318), .o(n746) );
ao22f01 g0591 ( .a(n7000_1), .b(net_6967), .c(n6999), .d(net_7031), .o(n7321_1) );
ao22f01 g0592 ( .a(n7003), .b(net_6999), .c(n7002), .d(net_7063), .o(n7322) );
na02f01 g0593 ( .a(n7322), .b(n7321_1), .o(n7323) );
na02f01 g0594 ( .a(n7323), .b(n6981), .o(n7324) );
ao22f01 g0595 ( .a(n7000_1), .b(net_6965), .c(n6999), .d(net_7029), .o(n7325) );
ao22f01 g0596 ( .a(n7003), .b(net_6997), .c(n7002), .d(net_7061), .o(n7326_1) );
na02f01 g0597 ( .a(n7326_1), .b(n7325), .o(n7327) );
ao22f01 g0598 ( .a(n7327), .b(n6998), .c(n6996), .d(_net_6147), .o(n7328) );
na02f01 g0599 ( .a(n7328), .b(n7324), .o(n756) );
in01f01 g0600 ( .a(_net_7793), .o(n7330_1) );
no02f01 g0601 ( .a(x1286), .b(x1322), .o(n7331) );
na03f01 g0602 ( .a(n7331), .b(_net_6184), .c(n7300), .o(n7332) );
no02f01 g0603 ( .a(n7332), .b(n7330_1), .o(n765) );
in01f01 g0604 ( .a(_net_7732), .o(n7334) );
in01f01 g0605 ( .a(_net_6026), .o(n7335_1) );
in01f01 g0606 ( .a(n7108), .o(n7336) );
in01f01 g0607 ( .a(_net_7688), .o(n7337) );
na03f01 g0608 ( .a(_net_7687), .b(n7337), .c(n7105), .o(n7338) );
no02f01 g0609 ( .a(n7338), .b(n7336), .o(n7339) );
in01f01 g0610 ( .a(n7339), .o(n7340_1) );
in01f01 g0611 ( .a(x1231), .o(n7341) );
na02f01 g0612 ( .a(n7341), .b(n7281), .o(n7342) );
no04f01 g0613 ( .a(n7342), .b(n7340_1), .c(n7292_1), .d(x1322), .o(n7343) );
ao12f01 g0614 ( .a(n7343), .b(n7335_1), .c(n7334), .o(n770) );
in01f01 g0615 ( .a(_net_6012), .o(n7345) );
in01f01 g0616 ( .a(_net_6184), .o(n7346) );
na02f01 g0617 ( .a(n7304), .b(x1322), .o(n7347) );
no02f01 g0618 ( .a(n7347), .b(n7346), .o(n7348) );
na02f01 g0619 ( .a(n7348), .b(_net_7815), .o(n7349_1) );
oa12f01 g0620 ( .a(n7349_1), .b(n7348), .c(n7345), .o(n788) );
in01f01 g0621 ( .a(net_377), .o(n7351) );
no02f01 g0622 ( .a(n6966), .b(n7351), .o(n793) );
in01f01 g0623 ( .a(_net_113), .o(n7353) );
no02f01 g0624 ( .a(_net_7785), .b(_net_7786), .o(n7354_1) );
in01f01 g0625 ( .a(_net_7788), .o(n7355) );
no02f01 g0626 ( .a(n7355), .b(_net_7787), .o(n7356) );
na04f01 g0627 ( .a(n7356), .b(n7354_1), .c(_net_7789), .d(_net_7784), .o(n7357) );
na02f01 g0628 ( .a(n7357), .b(n7353), .o(n7358) );
in01f01 g0629 ( .a(_net_7786), .o(n7359_1) );
na02f01 g0630 ( .a(_net_7784), .b(_net_7785), .o(n7360) );
no02f01 g0631 ( .a(n7360), .b(n7359_1), .o(n7361) );
in01f01 g0632 ( .a(n7360), .o(n7362) );
no02f01 g0633 ( .a(n7362), .b(_net_7786), .o(n7363_1) );
no03f01 g0634 ( .a(n7363_1), .b(n7361), .c(n7358), .o(n806) );
in01f01 g0635 ( .a(_net_121), .o(n7365) );
na02f01 g0636 ( .a(net_317), .b(_net_154), .o(n7366) );
oa12f01 g0637 ( .a(n7366), .b(_net_154), .c(n7365), .o(n820) );
in01f01 g0638 ( .a(_net_120), .o(n7368_1) );
na02f01 g0639 ( .a(net_316), .b(_net_154), .o(n7369) );
oa12f01 g0640 ( .a(n7369), .b(_net_154), .c(n7368_1), .o(n825) );
ao22f01 g0641 ( .a(n7225), .b(_net_7428), .c(n7224), .d(net_7460), .o(n7371) );
ao22f01 g0642 ( .a(n7229), .b(net_7524), .c(n7228), .d(net_7492), .o(n7372_1) );
na02f01 g0643 ( .a(n7372_1), .b(n7371), .o(n834) );
ao22f01 g0644 ( .a(n6877), .b(_net_7265), .c(n6876_1), .d(_net_7329), .o(n7374) );
ao22f01 g0645 ( .a(n6881_1), .b(_net_7297), .c(n6880), .d(_net_7361), .o(n7375) );
na02f01 g0646 ( .a(n7375), .b(n7374), .o(n849) );
na02f01 g0647 ( .a(n6938_1), .b(n6917), .o(n7377) );
ao22f01 g0648 ( .a(n6942), .b(n6935), .c(n6933), .d(_net_6086), .o(n7378) );
na02f01 g0649 ( .a(n7378), .b(n7377), .o(n862) );
no02f01 g0650 ( .a(n6899_1), .b(n7254), .o(n875) );
in01f01 g0651 ( .a(_net_6008), .o(n7381_1) );
na02f01 g0652 ( .a(n7348), .b(_net_7811), .o(n7382) );
oa12f01 g0653 ( .a(n7382), .b(n7348), .c(n7381_1), .o(n885) );
in01f01 g0654 ( .a(_net_7439), .o(n7384) );
na02f01 g0655 ( .a(n6866), .b(net_7391), .o(n7385) );
ao22f01 g0656 ( .a(net_354), .b(_net_280), .c(_net_281), .d(net_352), .o(n7386_1) );
na02f01 g0657 ( .a(n7386_1), .b(n7385), .o(n7387) );
na02f01 g0658 ( .a(n7387), .b(n7197), .o(n7388) );
oa12f01 g0659 ( .a(n7388), .b(n7197), .c(n7384), .o(n903) );
in01f01 g0660 ( .a(_net_7354), .o(n7390) );
na02f01 g0661 ( .a(n6898), .b(net_7242), .o(n7391_1) );
ao22f01 g0662 ( .a(_net_269), .b(net_336), .c(_net_270), .d(net_334), .o(n7392) );
na02f01 g0663 ( .a(n7392), .b(n7391_1), .o(n7393) );
na02f01 g0664 ( .a(n7393), .b(n7030), .o(n7394) );
oa12f01 g0665 ( .a(n7394), .b(n7030), .c(n7390), .o(n925) );
in01f01 g0666 ( .a(_net_7632), .o(n7396) );
in01f01 g0667 ( .a(_net_7685), .o(n7397) );
no02f01 g0668 ( .a(n7397), .b(_net_7684), .o(n7398) );
in01f01 g0669 ( .a(n7398), .o(n7399) );
no02f01 g0670 ( .a(n7399), .b(n6967), .o(n7400_1) );
na02f01 g0671 ( .a(n6965), .b(net_370), .o(n7401) );
ao22f01 g0672 ( .a(net_384), .b(_net_291), .c(_net_292), .d(net_382), .o(n7402) );
na02f01 g0673 ( .a(n7402), .b(n7401), .o(n7403) );
na02f01 g0674 ( .a(n7403), .b(n7400_1), .o(n7404_1) );
oa12f01 g0675 ( .a(n7404_1), .b(n7400_1), .c(n7396), .o(n930) );
in01f01 g0676 ( .a(_net_5851), .o(n7406) );
in01f01 g0677 ( .a(x868), .o(n7407) );
in01f01 g0678 ( .a(_net_282), .o(n7408_1) );
no02f01 g0679 ( .a(_net_283), .b(n7408_1), .o(n7409) );
in01f01 g0680 ( .a(_net_226), .o(n7410) );
na02f01 g0681 ( .a(_net_278), .b(_net_284), .o(n7411) );
ao12f01 g0682 ( .a(n7411), .b(_net_229), .c(n7410), .o(n7412) );
na02f01 g0683 ( .a(n7412), .b(n7409), .o(n7413_1) );
in01f01 g0684 ( .a(n7411), .o(n7414) );
in01f01 g0685 ( .a(_net_283), .o(n7415) );
no02f01 g0686 ( .a(n7415), .b(n7408_1), .o(n7416) );
na03f01 g0687 ( .a(n7416), .b(n7414), .c(_net_226), .o(n7417_1) );
na03f01 g0688 ( .a(_net_228), .b(_net_229), .c(n7410), .o(n7418) );
na04f01 g0689 ( .a(n7418), .b(n7414), .c(n7415), .d(n7408_1), .o(n7419) );
oa12f01 g0690 ( .a(n7410), .b(_net_228), .c(_net_229), .o(n7420) );
na04f01 g0691 ( .a(n7420), .b(n7414), .c(_net_283), .d(n7408_1), .o(n7421) );
na04f01 g0692 ( .a(n7421), .b(n7419), .c(n7417_1), .d(n7413_1), .o(n7422_1) );
na03f01 g0693 ( .a(n7422_1), .b(net_7779), .c(n7407), .o(n7423) );
oa12f01 g0694 ( .a(n7423), .b(n7406), .c(x868), .o(n944) );
in01f01 g0695 ( .a(_net_7629), .o(n7425) );
na02f01 g0696 ( .a(n6965), .b(net_7549), .o(n7426) );
ao22f01 g0697 ( .a(_net_292), .b(net_379), .c(_net_291), .d(net_381), .o(n7427_1) );
na02f01 g0698 ( .a(n7427_1), .b(n7426), .o(n7428) );
na02f01 g0699 ( .a(n7428), .b(n7400_1), .o(n7429) );
oa12f01 g0700 ( .a(n7429), .b(n7400_1), .c(n7425), .o(n961) );
ao22f01 g0701 ( .a(n7225), .b(_net_7412), .c(n7224), .d(_net_7444), .o(n7431) );
ao22f01 g0702 ( .a(n7229), .b(_net_7508), .c(n7228), .d(_net_7476), .o(n7432_1) );
na02f01 g0703 ( .a(n7432_1), .b(n7431), .o(n966) );
in01f01 g0704 ( .a(_net_7296), .o(n7434) );
na02f01 g0705 ( .a(n6898), .b(net_7248), .o(n7435) );
ao22f01 g0706 ( .a(net_342), .b(_net_269), .c(net_340), .d(_net_270), .o(n7436) );
na02f01 g0707 ( .a(n7436), .b(n7435), .o(n7437_1) );
na02f01 g0708 ( .a(n7437_1), .b(n7180), .o(n7438) );
oa12f01 g0709 ( .a(n7438), .b(n7180), .c(n7434), .o(n971) );
no04f01 g0710 ( .a(n7346), .b(n6801_1), .c(x1261), .d(n6800), .o(n7440) );
na02f01 g0711 ( .a(n7440), .b(_net_7805), .o(n7441) );
oa12f01 g0712 ( .a(n7441), .b(n7440), .c(n7408_1), .o(n985) );
in01f01 g0713 ( .a(_net_7653), .o(n7443) );
no02f01 g0714 ( .a(n7397), .b(n6959), .o(n7444) );
in01f01 g0715 ( .a(n7444), .o(n7445) );
no02f01 g0716 ( .a(n7445), .b(n6967), .o(n7446_1) );
na02f01 g0717 ( .a(n6965), .b(net_7541), .o(n7447) );
ao22f01 g0718 ( .a(_net_292), .b(net_371), .c(_net_291), .d(net_373), .o(n7448) );
na02f01 g0719 ( .a(n7448), .b(n7447), .o(n7449) );
na02f01 g0720 ( .a(n7449), .b(n7446_1), .o(n7450_1) );
oa12f01 g0721 ( .a(n7450_1), .b(n7446_1), .c(n7443), .o(n990) );
in01f01 g0722 ( .a(_net_5856), .o(n7452) );
in01f01 g0723 ( .a(x1006), .o(n7453) );
na03f01 g0724 ( .a(n7273), .b(net_7774), .c(n7453), .o(n7454_1) );
oa12f01 g0725 ( .a(n7454_1), .b(n7452), .c(x1006), .o(n995) );
in01f01 g0726 ( .a(_net_7621), .o(n7456) );
na02f01 g0727 ( .a(n7449), .b(n7400_1), .o(n7457) );
oa12f01 g0728 ( .a(n7457), .b(n7400_1), .c(n7456), .o(n1010) );
in01f01 g0729 ( .a(net_6770), .o(n7459_1) );
in01f01 g0730 ( .a(net_6706), .o(n7460) );
oa22f01 g0731 ( .a(n7129), .b(n7460), .c(n7126), .d(n7459_1), .o(n7461) );
in01f01 g0732 ( .a(net_6802), .o(n7462) );
in01f01 g0733 ( .a(net_6738), .o(n7463_1) );
oa22f01 g0734 ( .a(n7134), .b(n7463_1), .c(n7132), .d(n7462), .o(n7464) );
no02f01 g0735 ( .a(n7464), .b(n7461), .o(n7465) );
in01f01 g0736 ( .a(_net_6822), .o(n7466) );
no02f01 g0737 ( .a(_net_6009), .b(_net_6008), .o(n7467) );
na03f01 g0738 ( .a(n7467), .b(n7122), .c(n7466), .o(n7468_1) );
no02f01 g0739 ( .a(n7468_1), .b(n7465), .o(n7469) );
na02f01 g0740 ( .a(n7122), .b(_net_6008), .o(n7470) );
in01f01 g0741 ( .a(net_6708), .o(n7471) );
in01f01 g0742 ( .a(net_6772), .o(n7472) );
oa22f01 g0743 ( .a(n7129), .b(n7471), .c(n7126), .d(n7472), .o(n7473_1) );
in01f01 g0744 ( .a(net_6804), .o(n7474) );
in01f01 g0745 ( .a(net_6740), .o(n7475) );
oa22f01 g0746 ( .a(n7134), .b(n7475), .c(n7132), .d(n7474), .o(n7476) );
no02f01 g0747 ( .a(n7476), .b(n7473_1), .o(n7477) );
no02f01 g0748 ( .a(n7477), .b(n7470), .o(n7478_1) );
in01f01 g0749 ( .a(_net_6120), .o(n7479) );
in01f01 g0750 ( .a(net_6774), .o(n7480) );
in01f01 g0751 ( .a(net_6710), .o(n7481) );
oa22f01 g0752 ( .a(n7129), .b(n7481), .c(n7126), .d(n7480), .o(n7482_1) );
in01f01 g0753 ( .a(net_6806), .o(n7483) );
in01f01 g0754 ( .a(net_6742), .o(n7484) );
oa22f01 g0755 ( .a(n7134), .b(n7484), .c(n7132), .d(n7483), .o(n7485) );
no02f01 g0756 ( .a(n7485), .b(n7482_1), .o(n7486) );
oa22f01 g0757 ( .a(n7486), .b(n7123), .c(n7118), .d(n7479), .o(n7487_1) );
no03f01 g0758 ( .a(n7487_1), .b(n7478_1), .c(n7469), .o(n7488) );
in01f01 g0759 ( .a(net_6754), .o(n7489) );
in01f01 g0760 ( .a(net_6722), .o(n7490) );
na04f01 g0761 ( .a(n7467), .b(n7135), .c(n7122), .d(_net_6822), .o(n7491) );
na04f01 g0762 ( .a(n7467), .b(n7130), .c(n7122), .d(_net_6822), .o(n7492_1) );
oa22f01 g0763 ( .a(n7492_1), .b(n7490), .c(n7491), .d(n7489), .o(n7493) );
in01f01 g0764 ( .a(net_6786), .o(n7494) );
in01f01 g0765 ( .a(net_6818), .o(n7495) );
na04f01 g0766 ( .a(n7467), .b(n7127), .c(n7122), .d(_net_6822), .o(n7496_1) );
na04f01 g0767 ( .a(n7467), .b(n7133_1), .c(n7122), .d(_net_6822), .o(n7497) );
oa22f01 g0768 ( .a(n7497), .b(n7495), .c(n7496_1), .d(n7494), .o(n7498) );
no02f01 g0769 ( .a(n7498), .b(n7493), .o(n7499) );
na02f01 g0770 ( .a(n7499), .b(n7488), .o(n1015) );
in01f01 g0771 ( .a(_net_7447), .o(n7501_1) );
na02f01 g0772 ( .a(n6866), .b(net_7399), .o(n7502) );
ao22f01 g0773 ( .a(_net_281), .b(net_360), .c(_net_280), .d(net_362), .o(n7503) );
na02f01 g0774 ( .a(n7503), .b(n7502), .o(n7504) );
na02f01 g0775 ( .a(n7504), .b(n7197), .o(n7505_1) );
oa12f01 g0776 ( .a(n7505_1), .b(n7197), .c(n7501_1), .o(n1024) );
in01f01 g0777 ( .a(net_334), .o(n7507) );
no02f01 g0778 ( .a(n6899_1), .b(n7507), .o(n1029) );
in01f01 g0779 ( .a(net_343), .o(n7509_1) );
no02f01 g0780 ( .a(n6899_1), .b(n7509_1), .o(n1034) );
in01f01 g0781 ( .a(_net_6259), .o(n7511) );
no02f01 g0782 ( .a(_net_392), .b(n7511), .o(n1039) );
in01f01 g0783 ( .a(_net_7281), .o(n7513_1) );
in01f01 g0784 ( .a(net_345), .o(n7514) );
no02f01 g0785 ( .a(n6899_1), .b(n7514), .o(n6722) );
na02f01 g0786 ( .a(n6722), .b(n6901), .o(n7516) );
oa12f01 g0787 ( .a(n7516), .b(n6901), .c(n7513_1), .o(n1044) );
in01f01 g0788 ( .a(_net_7578), .o(n7518_1) );
no03f01 g0789 ( .a(n6967), .b(_net_7685), .c(_net_7684), .o(n7519) );
in01f01 g0790 ( .a(net_380), .o(n7520) );
no02f01 g0791 ( .a(n6966), .b(n7520), .o(n3546) );
na02f01 g0792 ( .a(n3546), .b(n7519), .o(n7522_1) );
oa12f01 g0793 ( .a(n7522_1), .b(n7519), .c(n7518_1), .o(n1049) );
ao22f01 g0794 ( .a(n7288_1), .b(_net_6034), .c(n7286), .d(_net_273), .o(n7524) );
ao22f01 g0795 ( .a(n7298), .b(_net_7726), .c(n7291), .d(_net_7697), .o(n7525) );
na02f01 g0796 ( .a(n7302_1), .b(_net_120), .o(n7526) );
na03f01 g0797 ( .a(n7308), .b(net_199), .c(x1322), .o(n7527_1) );
na02f01 g0798 ( .a(n7296), .b(net_236), .o(n7528) );
na03f01 g0799 ( .a(n7308), .b(net_162), .c(n6800), .o(n7529) );
na03f01 g0800 ( .a(n7529), .b(n7528), .c(n7527_1), .o(n7530_1) );
ao12f01 g0801 ( .a(n7530_1), .b(n7306), .c(_net_5990), .o(n7531) );
na04f01 g0802 ( .a(n7531), .b(n7526), .c(n7525), .d(n7524), .o(n1058) );
in01f01 g0803 ( .a(_net_5960), .o(n7533) );
oa12f01 g0804 ( .a(n7533), .b(_net_5961), .c(_net_5962), .o(n7534) );
in01f01 g0805 ( .a(_net_5989), .o(n7535_1) );
no03f01 g0806 ( .a(n7535_1), .b(_net_5988), .c(n6759), .o(n7536) );
no02f01 g0807 ( .a(n6759), .b(n7533), .o(n7537) );
in01f01 g0808 ( .a(_net_5988), .o(n7538) );
no02f01 g0809 ( .a(n7535_1), .b(n7538), .o(n7539_1) );
ao22f01 g0810 ( .a(n7539_1), .b(n7537), .c(n7536), .d(n7534), .o(n7540) );
no02f01 g0811 ( .a(_net_5989), .b(n7538), .o(n7541) );
ao12f01 g0812 ( .a(n6759), .b(_net_5962), .c(n7533), .o(n7542) );
na03f01 g0813 ( .a(_net_5961), .b(_net_5962), .c(n7533), .o(n7543_1) );
no03f01 g0814 ( .a(_net_5989), .b(_net_5988), .c(n6759), .o(n7544) );
ao22f01 g0815 ( .a(n7544), .b(n7543_1), .c(n7542), .d(n7541), .o(n7545) );
na02f01 g0816 ( .a(n7545), .b(n7540), .o(n1067) );
in01f01 g0817 ( .a(_net_6285), .o(n7547) );
no02f01 g0818 ( .a(_net_392), .b(n7547), .o(n1072) );
in01f01 g0819 ( .a(_net_7412), .o(n7549) );
no03f01 g0820 ( .a(n6868), .b(_net_7533), .c(_net_7534), .o(n7550) );
na02f01 g0821 ( .a(n6866), .b(net_7396), .o(n7551) );
ao22f01 g0822 ( .a(net_359), .b(_net_280), .c(_net_281), .d(net_357), .o(n7552) );
na02f01 g0823 ( .a(n7552), .b(n7551), .o(n7553_1) );
na02f01 g0824 ( .a(n7553_1), .b(n7550), .o(n7554) );
oa12f01 g0825 ( .a(n7554), .b(n7550), .c(n7549), .o(n1106) );
in01f01 g0826 ( .a(net_7752), .o(n7556) );
na04f01 g0827 ( .a(_net_5995), .b(_net_7791), .c(n7556), .d(net_303), .o(n7557) );
ao12f01 g0828 ( .a(n7557), .b(net_308), .c(_net_5996), .o(n1116) );
in01f01 g0829 ( .a(_net_7274), .o(n7559) );
in01f01 g0830 ( .a(net_338), .o(n7560) );
no02f01 g0831 ( .a(n6899_1), .b(n7560), .o(n4263) );
na02f01 g0832 ( .a(n4263), .b(n6901), .o(n7562) );
oa12f01 g0833 ( .a(n7562), .b(n6901), .c(n7559), .o(n1125) );
in01f01 g0834 ( .a(_net_7299), .o(n7564) );
na02f01 g0835 ( .a(n6898), .b(net_331), .o(n7565) );
ao22f01 g0836 ( .a(_net_269), .b(net_345), .c(net_343), .d(_net_270), .o(n7566) );
na02f01 g0837 ( .a(n7566), .b(n7565), .o(n7567_1) );
na02f01 g0838 ( .a(n7567_1), .b(n7180), .o(n7568) );
oa12f01 g0839 ( .a(n7568), .b(n7180), .c(n7564), .o(n1135) );
in01f01 g0840 ( .a(_net_6039), .o(n7570) );
in01f01 g0841 ( .a(_net_7759), .o(n7571) );
na03f01 g0842 ( .a(net_6056), .b(_net_7791), .c(n7571), .o(n7572_1) );
no02f01 g0843 ( .a(n7572_1), .b(n7570), .o(n7573) );
na02f01 g0844 ( .a(n7573), .b(_net_6042), .o(n7574) );
in01f01 g0845 ( .a(n7574), .o(n7575) );
in01f01 g0846 ( .a(_net_7228), .o(n7576) );
na02f01 g0847 ( .a(n7576), .b(_net_7229), .o(n7577_1) );
in01f01 g0848 ( .a(n7577_1), .o(n7578) );
in01f01 g0849 ( .a(_net_7229), .o(n7579) );
na02f01 g0850 ( .a(n7576), .b(n7579), .o(n7580) );
in01f01 g0851 ( .a(n7580), .o(n7581_1) );
ao22f01 g0852 ( .a(n7581_1), .b(net_7102), .c(n7578), .d(net_7166), .o(n7582) );
na02f01 g0853 ( .a(_net_7228), .b(_net_7229), .o(n7583) );
in01f01 g0854 ( .a(n7583), .o(n7584) );
na02f01 g0855 ( .a(_net_7228), .b(n7579), .o(n7585) );
in01f01 g0856 ( .a(n7585), .o(n7586_1) );
ao22f01 g0857 ( .a(n7586_1), .b(net_7134), .c(n7584), .d(net_7198), .o(n7587) );
na02f01 g0858 ( .a(n7587), .b(n7582), .o(n7588) );
na02f01 g0859 ( .a(n7588), .b(n7575), .o(n7589) );
na02f01 g0860 ( .a(n7572_1), .b(_net_6039), .o(n7590) );
in01f01 g0861 ( .a(n7590), .o(n7591_1) );
na02f01 g0862 ( .a(n7573), .b(_net_6041), .o(n7592) );
in01f01 g0863 ( .a(n7592), .o(n7593) );
ao22f01 g0864 ( .a(n7581_1), .b(net_7100), .c(n7578), .d(net_7164), .o(n7594) );
ao22f01 g0865 ( .a(n7586_1), .b(net_7132), .c(n7584), .d(net_7196), .o(n7595) );
na02f01 g0866 ( .a(n7595), .b(n7594), .o(n7596_1) );
ao22f01 g0867 ( .a(n7596_1), .b(n7593), .c(n7591_1), .d(_net_6167), .o(n7597) );
na02f01 g0868 ( .a(n7597), .b(n7589), .o(n1153) );
in01f01 g0869 ( .a(net_381), .o(n7599_1) );
no02f01 g0870 ( .a(n6966), .b(n7599_1), .o(n1163) );
in01f01 g0871 ( .a(net_360), .o(n7601) );
no02f01 g0872 ( .a(n6867_1), .b(n7601), .o(n1173) );
no02f01 g0873 ( .a(n6833), .b(n6824), .o(n7603) );
no02f01 g0874 ( .a(n6843), .b(n6826_1), .o(n7604_1) );
in01f01 g0875 ( .a(_net_6135), .o(n7605) );
in01f01 g0876 ( .a(net_6904), .o(n7606) );
in01f01 g0877 ( .a(net_6840), .o(n7607) );
oa22f01 g0878 ( .a(n6810), .b(n7607), .c(n6807), .d(n7606), .o(n7608_1) );
in01f01 g0879 ( .a(net_6872), .o(n7609) );
in01f01 g0880 ( .a(net_6936), .o(n7610) );
oa22f01 g0881 ( .a(n6815), .b(n7609), .c(n6813_1), .d(n7610), .o(n7611) );
no02f01 g0882 ( .a(n7611), .b(n7608_1), .o(n7612) );
oa22f01 g0883 ( .a(n7612), .b(n6836_1), .c(n6844), .d(n7605), .o(n7613_1) );
no03f01 g0884 ( .a(n7613_1), .b(n7604_1), .c(n7603), .o(n7614) );
in01f01 g0885 ( .a(net_6852), .o(n7615) );
in01f01 g0886 ( .a(net_6884), .o(n7616) );
oa22f01 g0887 ( .a(n6850_1), .b(n7615), .c(n6849), .d(n7616), .o(n7617) );
in01f01 g0888 ( .a(net_6948), .o(n7618_1) );
in01f01 g0889 ( .a(net_6916), .o(n7619) );
oa22f01 g0890 ( .a(n6855_1), .b(n7618_1), .c(n6854), .d(n7619), .o(n7620) );
no02f01 g0891 ( .a(n7620), .b(n7617), .o(n7621) );
na02f01 g0892 ( .a(n7621), .b(n7614), .o(n1178) );
in01f01 g0893 ( .a(_net_7503), .o(n7623) );
no02f01 g0894 ( .a(n7194_1), .b(n6860_1), .o(n7624) );
in01f01 g0895 ( .a(n7624), .o(n7625) );
no02f01 g0896 ( .a(n7625), .b(n6868), .o(n7626_1) );
na02f01 g0897 ( .a(n7626_1), .b(n7387), .o(n7627) );
oa12f01 g0898 ( .a(n7627), .b(n7626_1), .c(n7623), .o(n1214) );
in01f01 g0899 ( .a(_net_7428), .o(n7629) );
na02f01 g0900 ( .a(n7550), .b(n595), .o(n7630) );
oa12f01 g0901 ( .a(n7630), .b(n7550), .c(n7629), .o(n1219) );
in01f01 g0902 ( .a(_net_7730), .o(n7632) );
in01f01 g0903 ( .a(_net_6016), .o(n7633) );
ao12f01 g0904 ( .a(n7343), .b(n7633), .c(n7632), .o(n1228) );
in01f01 g0905 ( .a(_net_7512), .o(n7635_1) );
na02f01 g0906 ( .a(n6866), .b(net_7400), .o(n7636) );
ao22f01 g0907 ( .a(_net_281), .b(net_361), .c(_net_280), .d(net_363), .o(n7637) );
na02f01 g0908 ( .a(n7637), .b(n7636), .o(n7638) );
na02f01 g0909 ( .a(n7638), .b(n7626_1), .o(n7639) );
oa12f01 g0910 ( .a(n7639), .b(n7626_1), .c(n7635_1), .o(n1253) );
in01f01 g0911 ( .a(_net_7590), .o(n7641) );
na02f01 g0912 ( .a(n6965), .b(net_7542), .o(n7642) );
ao22f01 g0913 ( .a(net_374), .b(_net_291), .c(_net_292), .d(net_372), .o(n7643) );
na02f01 g0914 ( .a(n7643), .b(n7642), .o(n7644_1) );
na02f01 g0915 ( .a(n7644_1), .b(n6968), .o(n7645) );
oa12f01 g0916 ( .a(n7645), .b(n6968), .c(n7641), .o(n1267) );
in01f01 g0917 ( .a(_net_273), .o(n7647) );
na02f01 g0918 ( .a(n7440), .b(net_7799), .o(n7648) );
oa12f01 g0919 ( .a(n7648), .b(n7440), .c(n7647), .o(n1272) );
in01f01 g0920 ( .a(net_354), .o(n7650) );
no02f01 g0921 ( .a(n6867_1), .b(n7650), .o(n1277) );
in01f01 g0922 ( .a(_net_299), .o(n7652) );
in01f01 g0923 ( .a(_net_263), .o(n7653) );
in01f01 g0924 ( .a(n6964_1), .o(n7654_1) );
oa12f01 g0925 ( .a(n7652), .b(n7654_1), .c(n7653), .o(n1282) );
in01f01 g0926 ( .a(_net_7315), .o(n7656) );
na02f01 g0927 ( .a(n6898), .b(net_7235), .o(n7657) );
ao22f01 g0928 ( .a(net_327), .b(_net_270), .c(_net_269), .d(net_329), .o(n7658_1) );
na02f01 g0929 ( .a(n7658_1), .b(n7657), .o(n7659) );
na02f01 g0930 ( .a(n7659), .b(n7150), .o(n7660) );
oa12f01 g0931 ( .a(n7660), .b(n7150), .c(n7656), .o(n1295) );
no02f01 g0932 ( .a(_net_6692), .b(n6921), .o(n7662) );
in01f01 g0933 ( .a(_net_6692), .o(n7663) );
no02f01 g0934 ( .a(n7663), .b(_net_6689), .o(n7664) );
no02f01 g0935 ( .a(n7664), .b(n7662), .o(n7665) );
no02f01 g0936 ( .a(n6918), .b(net_6691), .o(n7666_1) );
no02f01 g0937 ( .a(n7666_1), .b(n7665), .o(n7667) );
no04f01 g0938 ( .a(n7664), .b(n7662), .c(n6918), .d(net_6691), .o(n7668) );
oa12f01 g0939 ( .a(n7156), .b(n7668), .c(n7667), .o(n7669) );
no02f01 g0940 ( .a(n7668), .b(n7667), .o(n7670) );
na02f01 g0941 ( .a(n7670), .b(n548), .o(n7671_1) );
na02f01 g0942 ( .a(n7671_1), .b(n7669), .o(n1309) );
in01f01 g0943 ( .a(_net_6000), .o(n7673) );
na02f01 g0944 ( .a(n7348), .b(_net_7806), .o(n7674) );
oa12f01 g0945 ( .a(n7674), .b(n7348), .c(n7673), .o(n1314) );
in01f01 g0946 ( .a(_net_5991), .o(n7676_1) );
na02f01 g0947 ( .a(n7348), .b(_net_7800), .o(n7677) );
oa12f01 g0948 ( .a(n7677), .b(n7348), .c(n7676_1), .o(n1335) );
in01f01 g0949 ( .a(_net_7707), .o(n7679) );
na02f01 g0950 ( .a(n7207_1), .b(_net_7809), .o(n7680) );
oa12f01 g0951 ( .a(n7680), .b(n7207_1), .c(n7679), .o(n1340) );
in01f01 g0952 ( .a(_net_5975), .o(n7682) );
no02f01 g0953 ( .a(n6819), .b(n7682), .o(n1345) );
ao22f01 g0954 ( .a(n7225), .b(_net_7421), .c(n7224), .d(net_7453), .o(n7684) );
ao22f01 g0955 ( .a(n7229), .b(net_7517), .c(n7228), .d(net_7485), .o(n7685) );
na02f01 g0956 ( .a(n7685), .b(n7684), .o(n1363) );
in01f01 g0957 ( .a(_net_5972), .o(n7687) );
oa12f01 g0958 ( .a(n7687), .b(_net_5973), .c(_net_5974), .o(n7688) );
in01f01 g0959 ( .a(_net_6022), .o(n7689) );
no03f01 g0960 ( .a(n6819), .b(_net_6021), .c(n7689), .o(n7690) );
no02f01 g0961 ( .a(n6819), .b(n7687), .o(n7691_1) );
in01f01 g0962 ( .a(_net_6021), .o(n7692) );
no02f01 g0963 ( .a(n7692), .b(n7689), .o(n7693) );
ao22f01 g0964 ( .a(n7693), .b(n7691_1), .c(n7690), .d(n7688), .o(n7694) );
no02f01 g0965 ( .a(n7692), .b(_net_6022), .o(n7695_1) );
ao12f01 g0966 ( .a(n6819), .b(_net_5974), .c(n7687), .o(n7696) );
na03f01 g0967 ( .a(_net_5973), .b(_net_5974), .c(n7687), .o(n7697) );
no03f01 g0968 ( .a(n6819), .b(_net_6021), .c(_net_6022), .o(n7698) );
ao22f01 g0969 ( .a(n7698), .b(n7697), .c(n7696), .d(n7695_1), .o(n7699) );
na02f01 g0970 ( .a(n7699), .b(n7694), .o(n1368) );
in01f01 g0971 ( .a(_net_5997), .o(n7701) );
na02f01 g0972 ( .a(n7348), .b(_net_7803), .o(n7702) );
oa12f01 g0973 ( .a(n7702), .b(n7348), .c(n7701), .o(n1373) );
in01f01 g0974 ( .a(_net_7658), .o(n7704_1) );
na02f01 g0975 ( .a(n6965), .b(net_7546), .o(n7705) );
ao22f01 g0976 ( .a(_net_292), .b(net_376), .c(_net_291), .d(net_378), .o(n7706) );
na02f01 g0977 ( .a(n7706), .b(n7705), .o(n7707) );
na02f01 g0978 ( .a(n7707), .b(n7446_1), .o(n7708) );
oa12f01 g0979 ( .a(n7708), .b(n7446_1), .c(n7704_1), .o(n1391) );
in01f01 g0980 ( .a(_net_6189), .o(n7710) );
no02f01 g0981 ( .a(_net_392), .b(n7710), .o(n1396) );
in01f01 g0982 ( .a(net_7113), .o(n7712) );
in01f01 g0983 ( .a(net_7177), .o(n7713) );
oa22f01 g0984 ( .a(n7580), .b(n7712), .c(n7577_1), .d(n7713), .o(n7714_1) );
in01f01 g0985 ( .a(net_7145), .o(n7715) );
in01f01 g0986 ( .a(net_7209), .o(n7716) );
oa22f01 g0987 ( .a(n7585), .b(n7715), .c(n7583), .d(n7716), .o(n7717) );
no02f01 g0988 ( .a(n7717), .b(n7714_1), .o(n7718) );
in01f01 g0989 ( .a(_net_7227), .o(n7719_1) );
no02f01 g0990 ( .a(_net_6041), .b(_net_6042), .o(n7720) );
na03f01 g0991 ( .a(n7720), .b(n7573), .c(n7719_1), .o(n7721) );
no02f01 g0992 ( .a(n7721), .b(n7718), .o(n7722) );
in01f01 g0993 ( .a(net_7179), .o(n7723_1) );
in01f01 g0994 ( .a(net_7115), .o(n7724) );
oa22f01 g0995 ( .a(n7580), .b(n7724), .c(n7577_1), .d(n7723_1), .o(n7725) );
in01f01 g0996 ( .a(net_7147), .o(n7726) );
in01f01 g0997 ( .a(net_7211), .o(n7727) );
oa22f01 g0998 ( .a(n7585), .b(n7726), .c(n7583), .d(n7727), .o(n7728_1) );
no02f01 g0999 ( .a(n7728_1), .b(n7725), .o(n7729) );
no02f01 g1000 ( .a(n7729), .b(n7592), .o(n7730) );
ao22f01 g1001 ( .a(n7581_1), .b(net_7117), .c(n7578), .d(net_7181), .o(n7731) );
ao22f01 g1002 ( .a(n7586_1), .b(net_7149), .c(n7584), .d(net_7213), .o(n7732_1) );
ao12f01 g1003 ( .a(n7574), .b(n7732_1), .c(n7731), .o(n7733) );
in01f01 g1004 ( .a(_net_6182), .o(n7734) );
no02f01 g1005 ( .a(n7590), .b(n7734), .o(n7735) );
no04f01 g1006 ( .a(n7735), .b(n7733), .c(n7730), .d(n7722), .o(n7736) );
in01f01 g1007 ( .a(net_7129), .o(n7737_1) );
in01f01 g1008 ( .a(net_7161), .o(n7738) );
na04f01 g1009 ( .a(n7720), .b(n7586_1), .c(n7573), .d(_net_7227), .o(n7739) );
na04f01 g1010 ( .a(n7720), .b(n7581_1), .c(n7573), .d(_net_7227), .o(n7740) );
oa22f01 g1011 ( .a(n7740), .b(n7737_1), .c(n7739), .d(n7738), .o(n7741_1) );
in01f01 g1012 ( .a(net_7225), .o(n7742) );
in01f01 g1013 ( .a(net_7193), .o(n7743) );
na04f01 g1014 ( .a(n7720), .b(n7578), .c(n7573), .d(_net_7227), .o(n7744) );
na04f01 g1015 ( .a(n7720), .b(n7584), .c(n7573), .d(_net_7227), .o(n7745) );
oa22f01 g1016 ( .a(n7745), .b(n7742), .c(n7744), .d(n7743), .o(n7746_1) );
no02f01 g1017 ( .a(n7746_1), .b(n7741_1), .o(n7747) );
na02f01 g1018 ( .a(n7747), .b(n7736), .o(n1405) );
in01f01 g1019 ( .a(_net_6555), .o(n7749) );
no02f01 g1020 ( .a(n6758), .b(n6747), .o(n7750) );
na03f01 g1021 ( .a(n7750), .b(n7749), .c(_net_6554), .o(n7751_1) );
in01f01 g1022 ( .a(n7750), .o(n7752) );
oa12f01 g1023 ( .a(_net_6555), .b(n7752), .c(n6749_1), .o(n7753) );
na02f01 g1024 ( .a(n7753), .b(n7751_1), .o(n7754) );
na02f01 g1025 ( .a(n7754), .b(_net_6558), .o(n7755) );
in01f01 g1026 ( .a(_net_6558), .o(n7756_1) );
na03f01 g1027 ( .a(n7753), .b(n7751_1), .c(n7756_1), .o(n7757) );
na02f01 g1028 ( .a(n6758), .b(_net_6553), .o(n7758) );
na02f01 g1029 ( .a(_net_6552), .b(n6747), .o(n7759) );
na02f01 g1030 ( .a(n7759), .b(n7758), .o(n7760_1) );
na02f01 g1031 ( .a(n7760_1), .b(net_6556), .o(n7761) );
in01f01 g1032 ( .a(net_6556), .o(n7762) );
na03f01 g1033 ( .a(n7759), .b(n7758), .c(n7762), .o(n7763) );
ao22f01 g1034 ( .a(n7763), .b(n7761), .c(n6763), .d(_net_6552), .o(n7764_1) );
in01f01 g1035 ( .a(_net_6557), .o(n7765) );
na02f01 g1036 ( .a(n7750), .b(n6749_1), .o(n7766) );
na02f01 g1037 ( .a(n7752), .b(_net_6554), .o(n7767) );
na02f01 g1038 ( .a(n7767), .b(n7766), .o(n7768_1) );
na02f01 g1039 ( .a(n7768_1), .b(n7765), .o(n7769) );
na03f01 g1040 ( .a(n7767), .b(n7766), .c(_net_6557), .o(n7770) );
na03f01 g1041 ( .a(n7770), .b(n7769), .c(n7764_1), .o(n7771) );
ao12f01 g1042 ( .a(n7771), .b(n7757), .c(n7755), .o(n1410) );
in01f01 g1043 ( .a(_net_7253), .o(n7773_1) );
na02f01 g1044 ( .a(n7183), .b(n6901), .o(n7774) );
oa12f01 g1045 ( .a(n7774), .b(n6901), .c(n7773_1), .o(n1419) );
in01f01 g1046 ( .a(_net_7497), .o(n7776_1) );
na02f01 g1047 ( .a(n6866), .b(net_7385), .o(n7777) );
ao22f01 g1048 ( .a(net_348), .b(_net_280), .c(_net_281), .d(net_346), .o(n7778) );
na02f01 g1049 ( .a(n7778), .b(n7777), .o(n7779_1) );
na02f01 g1050 ( .a(n7779_1), .b(n7626_1), .o(n7780) );
oa12f01 g1051 ( .a(n7780), .b(n7626_1), .c(n7776_1), .o(n1428) );
in01f01 g1052 ( .a(n7331), .o(n7782) );
no02f01 g1053 ( .a(n7782), .b(n7206), .o(n1433) );
in01f01 g1054 ( .a(_net_7565), .o(n7784_1) );
na02f01 g1055 ( .a(n7519), .b(n7428), .o(n7785) );
oa12f01 g1056 ( .a(n7785), .b(n7519), .c(n7784_1), .o(n1442) );
in01f01 g1057 ( .a(_net_7806), .o(n7787) );
na02f01 g1058 ( .a(n6803), .b(_net_6044), .o(n7788_1) );
oa12f01 g1059 ( .a(n7788_1), .b(n6803), .c(n7787), .o(n1451) );
in01f01 g1060 ( .a(_net_7746), .o(n7790) );
in01f01 g1061 ( .a(net_297), .o(n7791) );
ao12f01 g1062 ( .a(n7343), .b(n7791), .c(n7790), .o(n1487) );
in01f01 g1063 ( .a(net_7754), .o(n7793_1) );
na04f01 g1064 ( .a(_net_7791), .b(_net_6006), .c(net_303), .d(n7793_1), .o(n7794) );
ao12f01 g1065 ( .a(n7794), .b(net_307), .c(_net_6007), .o(n1496) );
in01f01 g1066 ( .a(_net_7698), .o(n7796) );
na02f01 g1067 ( .a(n7207_1), .b(_net_7800), .o(n7797) );
oa12f01 g1068 ( .a(n7797), .b(n7207_1), .c(n7796), .o(n1501) );
in01f01 g1069 ( .a(net_6630), .o(n7799) );
in01f01 g1070 ( .a(net_6566), .o(n7800) );
oa22f01 g1071 ( .a(n6922), .b(n7800), .c(n6919_1), .d(n7799), .o(n7801) );
in01f01 g1072 ( .a(net_6598), .o(n7802_1) );
in01f01 g1073 ( .a(net_6662), .o(n7803) );
oa22f01 g1074 ( .a(n6927), .b(n7802_1), .c(n6925), .d(n7803), .o(n7804) );
no02f01 g1075 ( .a(n7804), .b(n7801), .o(n7805) );
no02f01 g1076 ( .a(n7805), .b(n6945), .o(n7806_1) );
in01f01 g1077 ( .a(net_6632), .o(n7807) );
in01f01 g1078 ( .a(net_6568), .o(n7808) );
oa22f01 g1079 ( .a(n6922), .b(n7808), .c(n6919_1), .d(n7807), .o(n7809) );
in01f01 g1080 ( .a(net_6664), .o(n7810_1) );
in01f01 g1081 ( .a(net_6600), .o(n7811) );
oa22f01 g1082 ( .a(n6927), .b(n7811), .c(n6925), .d(n7810_1), .o(n7812) );
no02f01 g1083 ( .a(n7812), .b(n7809), .o(n7813) );
no02f01 g1084 ( .a(n7813), .b(n6934_1), .o(n7814) );
in01f01 g1085 ( .a(_net_6095), .o(n7815_1) );
in01f01 g1086 ( .a(net_6570), .o(n7816) );
in01f01 g1087 ( .a(net_6634), .o(n7817) );
oa22f01 g1088 ( .a(n6922), .b(n7816), .c(n6919_1), .d(n7817), .o(n7818_1) );
in01f01 g1089 ( .a(net_6602), .o(n7819) );
in01f01 g1090 ( .a(net_6666), .o(n7820) );
oa22f01 g1091 ( .a(n6927), .b(n7819), .c(n6925), .d(n7820), .o(n7821) );
no02f01 g1092 ( .a(n7821), .b(n7818_1), .o(n7822_1) );
oa22f01 g1093 ( .a(n7822_1), .b(n6916), .c(n6932), .d(n7815_1), .o(n7823) );
no03f01 g1094 ( .a(n7823), .b(n7814), .c(n7806_1), .o(n7824) );
in01f01 g1095 ( .a(net_6614), .o(n7825) );
in01f01 g1096 ( .a(net_6582), .o(n7826_1) );
oa22f01 g1097 ( .a(n7058_1), .b(n7826_1), .c(n7057), .d(n7825), .o(n7827) );
in01f01 g1098 ( .a(net_6646), .o(n7828) );
in01f01 g1099 ( .a(net_6678), .o(n7829) );
oa22f01 g1100 ( .a(n7063), .b(n7829), .c(n7062_1), .d(n7828), .o(n7830) );
no02f01 g1101 ( .a(n7830), .b(n7827), .o(n7831_1) );
na02f01 g1102 ( .a(n7831_1), .b(n7824), .o(n1519) );
ao22f01 g1103 ( .a(n7225), .b(_net_7411), .c(n7224), .d(_net_7443), .o(n7833) );
ao22f01 g1104 ( .a(n7229), .b(_net_7507), .c(n7228), .d(_net_7475), .o(n7834) );
na02f01 g1105 ( .a(n7834), .b(n7833), .o(n1533) );
na02f01 g1106 ( .a(n7293), .b(net_216), .o(n7836) );
na02f01 g1107 ( .a(n7296), .b(net_253), .o(n7837) );
na02f01 g1108 ( .a(n7297_1), .b(net_179), .o(n7838) );
na03f01 g1109 ( .a(n7838), .b(n7837), .c(n7836), .o(n7839) );
ao12f01 g1110 ( .a(n7839), .b(n7291), .c(net_7714), .o(n7840_1) );
na02f01 g1111 ( .a(n7298), .b(net_7743), .o(n7841) );
ao22f01 g1112 ( .a(n7306), .b(net_6013), .c(n7286), .d(net_296), .o(n7842) );
na03f01 g1113 ( .a(n7842), .b(n7841), .c(n7840_1), .o(n1542) );
na02f01 g1114 ( .a(n6865), .b(_net_278), .o(n7844) );
no02f01 g1115 ( .a(n7844), .b(n6867_1), .o(n7845_1) );
in01f01 g1116 ( .a(_net_7532), .o(n7846) );
oa12f01 g1117 ( .a(n6860_1), .b(n7194_1), .c(n7846), .o(n7847) );
na03f01 g1118 ( .a(_net_7533), .b(_net_7532), .c(_net_7534), .o(n7848_1) );
na03f01 g1119 ( .a(n7848_1), .b(n7847), .c(n7845_1), .o(n7849) );
in01f01 g1120 ( .a(_net_278), .o(n7850) );
in01f01 g1121 ( .a(n6865), .o(n7851) );
no03f01 g1122 ( .a(n6866), .b(n7851), .c(n7850), .o(n7852) );
na02f01 g1123 ( .a(n7196), .b(n6862), .o(n7853_1) );
no02f01 g1124 ( .a(n6865), .b(n7850), .o(n7854) );
ao22f01 g1125 ( .a(n7854), .b(_net_7534), .c(n7853_1), .d(n7852), .o(n7855) );
na02f01 g1126 ( .a(n7855), .b(n7849), .o(n1546) );
in01f01 g1127 ( .a(_net_7406), .o(n7857) );
na02f01 g1128 ( .a(n6866), .b(net_7390), .o(n7858_1) );
ao22f01 g1129 ( .a(_net_281), .b(net_351), .c(_net_280), .d(net_353), .o(n7859) );
na02f01 g1130 ( .a(n7859), .b(n7858_1), .o(n7860) );
na02f01 g1131 ( .a(n7860), .b(n7550), .o(n7861) );
oa12f01 g1132 ( .a(n7861), .b(n7550), .c(n7857), .o(n1555) );
ao22f01 g1133 ( .a(n6736_1), .b(net_7644), .c(n6734), .d(net_7612), .o(n7863_1) );
ao22f01 g1134 ( .a(n6739), .b(net_7676), .c(n6738), .d(_net_7580), .o(n7864) );
na02f01 g1135 ( .a(n7864), .b(n7863_1), .o(n1572) );
na02f01 g1136 ( .a(n7624), .b(_net_7535), .o(n7866) );
in01f01 g1137 ( .a(_net_7535), .o(n7867_1) );
na02f01 g1138 ( .a(n7625), .b(n7867_1), .o(n7868) );
na03f01 g1139 ( .a(n7868), .b(n7866), .c(n7852), .o(n7869) );
na02f01 g1140 ( .a(n7848_1), .b(n7867_1), .o(n7870) );
in01f01 g1141 ( .a(n7848_1), .o(n7871_1) );
na02f01 g1142 ( .a(n7871_1), .b(_net_7535), .o(n7872) );
na03f01 g1143 ( .a(n7872), .b(n7870), .c(n7845_1), .o(n7873) );
na02f01 g1144 ( .a(n7854), .b(_net_7535), .o(n7874) );
na03f01 g1145 ( .a(n7874), .b(n7873), .c(n7869), .o(n1582) );
no02f01 g1146 ( .a(n7160_1), .b(n7232), .o(n1600) );
ao22f01 g1147 ( .a(n6877), .b(_net_7259), .c(n6876_1), .d(_net_7323), .o(n7877) );
ao22f01 g1148 ( .a(n6881_1), .b(_net_7291), .c(n6880), .d(_net_7355), .o(n7878_1) );
na02f01 g1149 ( .a(n7878_1), .b(n7877), .o(n1605) );
in01f01 g1150 ( .a(_net_7498), .o(n7880) );
na02f01 g1151 ( .a(n6866), .b(net_7386), .o(n7881) );
ao22f01 g1152 ( .a(_net_281), .b(net_347), .c(net_349), .d(_net_280), .o(n7882) );
na02f01 g1153 ( .a(n7882), .b(n7881), .o(n7883_1) );
na02f01 g1154 ( .a(n7883_1), .b(n7626_1), .o(n7884) );
oa12f01 g1155 ( .a(n7884), .b(n7626_1), .c(n7880), .o(n1610) );
in01f01 g1156 ( .a(_net_7696), .o(n7886) );
na02f01 g1157 ( .a(n7207_1), .b(_net_7798), .o(n7887) );
oa12f01 g1158 ( .a(n7887), .b(n7207_1), .c(n7886), .o(n1624) );
in01f01 g1159 ( .a(_net_7570), .o(n7889) );
in01f01 g1160 ( .a(net_372), .o(n7890) );
in01f01 g1161 ( .a(net_384), .o(n7891) );
oa22f01 g1162 ( .a(n6966), .b(n7890), .c(n7891), .d(n7143), .o(n7892) );
na02f01 g1163 ( .a(n7892), .b(n7519), .o(n7893_1) );
oa12f01 g1164 ( .a(n7893_1), .b(n7519), .c(n7889), .o(n1634) );
in01f01 g1165 ( .a(net_340), .o(n7895) );
no02f01 g1166 ( .a(n6899_1), .b(n7895), .o(n1639) );
ao22f01 g1167 ( .a(n6736_1), .b(net_7646), .c(n6734), .d(net_7614), .o(n7897_1) );
ao22f01 g1168 ( .a(n6739), .b(net_7678), .c(n6738), .d(_net_7582), .o(n7898) );
na02f01 g1169 ( .a(n7898), .b(n7897_1), .o(n1644) );
ao22f01 g1170 ( .a(n6736_1), .b(_net_7631), .c(n6734), .d(_net_7599), .o(n7900) );
ao22f01 g1171 ( .a(n6739), .b(_net_7663), .c(n6738), .d(_net_7567), .o(n7901) );
na02f01 g1172 ( .a(n7901), .b(n7900), .o(n1658) );
in01f01 g1173 ( .a(_net_7804), .o(n7903) );
na02f01 g1174 ( .a(n6803), .b(_net_6042), .o(n7904) );
oa12f01 g1175 ( .a(n7904), .b(n6803), .c(n7903), .o(n1677) );
ao22f01 g1176 ( .a(n7581_1), .b(net_7103), .c(n7578), .d(net_7167), .o(n7906_1) );
ao22f01 g1177 ( .a(n7586_1), .b(net_7135), .c(n7584), .d(net_7199), .o(n7907) );
na02f01 g1178 ( .a(n7907), .b(n7906_1), .o(n7908) );
na02f01 g1179 ( .a(n7908), .b(n7575), .o(n7909) );
ao22f01 g1180 ( .a(n7581_1), .b(net_7101), .c(n7578), .d(net_7165), .o(n7910) );
ao22f01 g1181 ( .a(n7586_1), .b(net_7133), .c(n7584), .d(net_7197), .o(n7911_1) );
na02f01 g1182 ( .a(n7911_1), .b(n7910), .o(n7912) );
ao22f01 g1183 ( .a(n7912), .b(n7593), .c(n7591_1), .d(_net_6168), .o(n7913) );
in01f01 g1184 ( .a(n7721), .o(n7914) );
ao22f01 g1185 ( .a(n7581_1), .b(net_7099), .c(n7578), .d(net_7163), .o(n7915) );
ao22f01 g1186 ( .a(n7586_1), .b(net_7131), .c(n7584), .d(net_7195), .o(n7916_1) );
na02f01 g1187 ( .a(n7916_1), .b(n7915), .o(n7917) );
na02f01 g1188 ( .a(n7917), .b(n7914), .o(n7918) );
na02f01 g1189 ( .a(n7720), .b(n7573), .o(n7919) );
no02f01 g1190 ( .a(n7919), .b(n7719_1), .o(n7920_1) );
oa12f01 g1191 ( .a(n7920_1), .b(n7728_1), .c(n7725), .o(n7921) );
na04f01 g1192 ( .a(n7921), .b(n7918), .c(n7913), .d(n7909), .o(n1696) );
in01f01 g1193 ( .a(_net_7358), .o(n7923) );
na02f01 g1194 ( .a(n6898), .b(net_7246), .o(n7924_1) );
ao22f01 g1195 ( .a(net_338), .b(_net_270), .c(net_340), .d(_net_269), .o(n7925) );
na02f01 g1196 ( .a(n7925), .b(n7924_1), .o(n7926) );
na02f01 g1197 ( .a(n7926), .b(n7030), .o(n7927) );
oa12f01 g1198 ( .a(n7927), .b(n7030), .c(n7923), .o(n1714) );
in01f01 g1199 ( .a(net_7111), .o(n7929_1) );
in01f01 g1200 ( .a(net_7175), .o(n7930) );
oa22f01 g1201 ( .a(n7580), .b(n7929_1), .c(n7577_1), .d(n7930), .o(n7931) );
in01f01 g1202 ( .a(net_7207), .o(n7932) );
in01f01 g1203 ( .a(net_7143), .o(n7933_1) );
oa22f01 g1204 ( .a(n7585), .b(n7933_1), .c(n7583), .d(n7932), .o(n7934) );
no02f01 g1205 ( .a(n7934), .b(n7931), .o(n7935) );
no02f01 g1206 ( .a(n7935), .b(n7721), .o(n7936) );
no02f01 g1207 ( .a(n7718), .b(n7592), .o(n7937_1) );
in01f01 g1208 ( .a(_net_6180), .o(n7938) );
oa22f01 g1209 ( .a(n7729), .b(n7574), .c(n7590), .d(n7938), .o(n7939) );
no03f01 g1210 ( .a(n7939), .b(n7937_1), .c(n7936), .o(n7940) );
in01f01 g1211 ( .a(net_7159), .o(n7941) );
in01f01 g1212 ( .a(net_7127), .o(n7942_1) );
oa22f01 g1213 ( .a(n7740), .b(n7942_1), .c(n7739), .d(n7941), .o(n7943) );
in01f01 g1214 ( .a(net_7223), .o(n7944) );
in01f01 g1215 ( .a(net_7191), .o(n7945_1) );
oa22f01 g1216 ( .a(n7745), .b(n7944), .c(n7744), .d(n7945_1), .o(n7946) );
no02f01 g1217 ( .a(n7946), .b(n7943), .o(n7947) );
na02f01 g1218 ( .a(n7947), .b(n7940), .o(n1727) );
in01f01 g1219 ( .a(_net_7468), .o(n7949) );
na02f01 g1220 ( .a(n6866), .b(net_7388), .o(n7950_1) );
ao22f01 g1221 ( .a(_net_281), .b(net_349), .c(_net_280), .d(net_351), .o(n7951) );
na02f01 g1222 ( .a(n7951), .b(n7950_1), .o(n7952) );
na02f01 g1223 ( .a(n7952), .b(n6869), .o(n7953) );
oa12f01 g1224 ( .a(n7953), .b(n6869), .c(n7949), .o(n1737) );
in01f01 g1225 ( .a(_net_5996), .o(n7955_1) );
na02f01 g1226 ( .a(n7348), .b(net_7802), .o(n7956) );
oa12f01 g1227 ( .a(n7956), .b(n7348), .c(n7955_1), .o(n1742) );
in01f01 g1228 ( .a(net_6433), .o(n7958_1) );
in01f01 g1229 ( .a(net_6497), .o(n7959) );
oa22f01 g1230 ( .a(n6750), .b(n7958_1), .c(n6748), .d(n7959), .o(n7960) );
in01f01 g1231 ( .a(net_6465), .o(n7961) );
in01f01 g1232 ( .a(net_6529), .o(n7962_1) );
oa22f01 g1233 ( .a(n6755), .b(n7961), .c(n6754), .d(n7962_1), .o(n7963) );
no02f01 g1234 ( .a(n7963), .b(n7960), .o(n7964) );
no02f01 g1235 ( .a(n7964), .b(n6764), .o(n7965) );
no02f01 g1236 ( .a(n7077_1), .b(n6766), .o(n7966) );
in01f01 g1237 ( .a(_net_6077), .o(n7967_1) );
oa22f01 g1238 ( .a(n7085_1), .b(n6775), .c(n6784), .d(n7967_1), .o(n7968) );
no03f01 g1239 ( .a(n7968), .b(n7966), .c(n7965), .o(n7969) );
in01f01 g1240 ( .a(net_6449), .o(n7970_1) );
in01f01 g1241 ( .a(net_6481), .o(n7971) );
oa22f01 g1242 ( .a(n6790), .b(n7970_1), .c(n6789), .d(n7971), .o(n7972) );
in01f01 g1243 ( .a(net_6545), .o(n7973) );
in01f01 g1244 ( .a(net_6513), .o(n7974) );
oa22f01 g1245 ( .a(n6795), .b(n7973), .c(n6794), .d(n7974), .o(n7975_1) );
no02f01 g1246 ( .a(n7975_1), .b(n7972), .o(n7976) );
na02f01 g1247 ( .a(n7976), .b(n7969), .o(n1747) );
in01f01 g1248 ( .a(net_364), .o(n7978) );
no02f01 g1249 ( .a(n6867_1), .b(n7978), .o(n1752) );
in01f01 g1250 ( .a(_net_5985), .o(n7980_1) );
na02f01 g1251 ( .a(n7348), .b(_net_7794), .o(n7981) );
oa12f01 g1252 ( .a(n7981), .b(n7348), .c(n7980_1), .o(n1770) );
in01f01 g1253 ( .a(_net_6295), .o(n7983) );
no02f01 g1254 ( .a(_net_392), .b(n7983), .o(n1787) );
in01f01 g1255 ( .a(n7343), .o(n1792) );
in01f01 g1256 ( .a(_net_6219), .o(n7986) );
no02f01 g1257 ( .a(n7986), .b(_net_392), .o(n1802) );
in01f01 g1258 ( .a(_net_7328), .o(n7988) );
na02f01 g1259 ( .a(n7437_1), .b(n7150), .o(n7989_1) );
oa12f01 g1260 ( .a(n7989_1), .b(n7150), .c(n7988), .o(n1807) );
in01f01 g1261 ( .a(_net_7359), .o(n7991) );
na02f01 g1262 ( .a(n6898), .b(net_7247), .o(n7992) );
ao22f01 g1263 ( .a(net_341), .b(_net_269), .c(_net_270), .d(net_339), .o(n7993) );
na02f01 g1264 ( .a(n7993), .b(n7992), .o(n7994_1) );
na02f01 g1265 ( .a(n7994_1), .b(n7030), .o(n7995) );
oa12f01 g1266 ( .a(n7995), .b(n7030), .c(n7991), .o(n1812) );
in01f01 g1267 ( .a(_net_7650), .o(n7997_1) );
na02f01 g1268 ( .a(n6965), .b(net_7538), .o(n7998) );
ao22f01 g1269 ( .a(net_368), .b(_net_292), .c(net_370), .d(_net_291), .o(n7999) );
na02f01 g1270 ( .a(n7999), .b(n7998), .o(n8000) );
na02f01 g1271 ( .a(n8000), .b(n7446_1), .o(n8001) );
oa12f01 g1272 ( .a(n8001), .b(n7446_1), .c(n7997_1), .o(n1832) );
ao22f01 g1273 ( .a(n6923), .b(net_6562), .c(n6920), .d(net_6626), .o(n8003) );
ao22f01 g1274 ( .a(n6928), .b(net_6594), .c(n6926), .d(net_6658), .o(n8004) );
na02f01 g1275 ( .a(n8004), .b(n8003), .o(n8005_1) );
na02f01 g1276 ( .a(n8005_1), .b(n6917), .o(n8006) );
ao22f01 g1277 ( .a(n6923), .b(net_6560), .c(n6920), .d(net_6624), .o(n8007) );
ao22f01 g1278 ( .a(n6928), .b(net_6592), .c(n6926), .d(net_6656), .o(n8008) );
na02f01 g1279 ( .a(n8008), .b(n8007), .o(n8009) );
ao22f01 g1280 ( .a(n8009), .b(n6935), .c(n6933), .d(_net_6087), .o(n8010_1) );
na02f01 g1281 ( .a(n8010_1), .b(n8006), .o(n1841) );
in01f01 g1282 ( .a(_net_6291), .o(n8012) );
no02f01 g1283 ( .a(_net_392), .b(n8012), .o(n1846) );
in01f01 g1284 ( .a(_net_6222), .o(n8014) );
no02f01 g1285 ( .a(_net_392), .b(n8014), .o(n1851) );
in01f01 g1286 ( .a(_net_7768), .o(n8016) );
in01f01 g1287 ( .a(net_153), .o(n8017) );
no02f01 g1288 ( .a(n8017), .b(n8016), .o(n1860) );
in01f01 g1289 ( .a(_net_7255), .o(n8019_1) );
na02f01 g1290 ( .a(n6898), .b(net_7239), .o(n8020) );
ao22f01 g1291 ( .a(net_333), .b(_net_269), .c(_net_270), .d(net_331), .o(n8021) );
na02f01 g1292 ( .a(n8021), .b(n8020), .o(n8022) );
na02f01 g1293 ( .a(n8022), .b(n6901), .o(n8023) );
oa12f01 g1294 ( .a(n8023), .b(n6901), .c(n8019_1), .o(n1869) );
in01f01 g1295 ( .a(_net_7600), .o(n8025) );
na02f01 g1296 ( .a(n7403), .b(n6968), .o(n8026) );
oa12f01 g1297 ( .a(n8026), .b(n6968), .c(n8025), .o(n1878) );
in01f01 g1298 ( .a(n6775), .o(n8028_1) );
ao22f01 g1299 ( .a(n6777), .b(net_6427), .c(n6776), .d(net_6491), .o(n8029) );
ao22f01 g1300 ( .a(n6780), .b(net_6459), .c(n6779_1), .d(net_6523), .o(n8030) );
na02f01 g1301 ( .a(n8030), .b(n8029), .o(n8031) );
na02f01 g1302 ( .a(n8031), .b(n8028_1), .o(n8032) );
in01f01 g1303 ( .a(n6766), .o(n8033_1) );
in01f01 g1304 ( .a(n6784), .o(n8034) );
ao22f01 g1305 ( .a(n6777), .b(net_6425), .c(n6776), .d(net_6489), .o(n8035) );
ao22f01 g1306 ( .a(n6780), .b(net_6457), .c(n6779_1), .d(net_6521), .o(n8036) );
na02f01 g1307 ( .a(n8036), .b(n8035), .o(n8037) );
ao22f01 g1308 ( .a(n8037), .b(n8033_1), .c(n8034), .d(_net_6067), .o(n8038_1) );
na02f01 g1309 ( .a(n8038_1), .b(n8032), .o(n1883) );
in01f01 g1310 ( .a(_net_7628), .o(n8040) );
na02f01 g1311 ( .a(n6965), .b(net_7548), .o(n8041) );
ao22f01 g1312 ( .a(_net_292), .b(net_378), .c(_net_291), .d(net_380), .o(n8042_1) );
na02f01 g1313 ( .a(n8042_1), .b(n8041), .o(n8043) );
na02f01 g1314 ( .a(n8043), .b(n7400_1), .o(n8044) );
oa12f01 g1315 ( .a(n8044), .b(n7400_1), .c(n8040), .o(n1888) );
in01f01 g1316 ( .a(net_7035), .o(n8046) );
in01f01 g1317 ( .a(net_6971), .o(n8047_1) );
oa22f01 g1318 ( .a(n6987), .b(n8047_1), .c(n6985), .d(n8046), .o(n8048) );
in01f01 g1319 ( .a(net_7067), .o(n8049) );
in01f01 g1320 ( .a(net_7003), .o(n8050) );
oa22f01 g1321 ( .a(n6992), .b(n8050), .c(n6991), .d(n8049), .o(n8051_1) );
no02f01 g1322 ( .a(n8051_1), .b(n8048), .o(n8052) );
no02f01 g1323 ( .a(n8052), .b(n7012), .o(n8053) );
in01f01 g1324 ( .a(net_7037), .o(n8054) );
in01f01 g1325 ( .a(net_6973), .o(n8055) );
oa22f01 g1326 ( .a(n6987), .b(n8055), .c(n6985), .d(n8054), .o(n8056_1) );
in01f01 g1327 ( .a(net_7069), .o(n8057) );
in01f01 g1328 ( .a(net_7005), .o(n8058) );
oa22f01 g1329 ( .a(n6992), .b(n8058), .c(n6991), .d(n8057), .o(n8059_1) );
no02f01 g1330 ( .a(n8059_1), .b(n8056_1), .o(n8060) );
no02f01 g1331 ( .a(n8060), .b(n6997), .o(n8061) );
in01f01 g1332 ( .a(_net_6155), .o(n8062) );
in01f01 g1333 ( .a(net_6975), .o(n8063) );
in01f01 g1334 ( .a(net_7039), .o(n8064_1) );
oa22f01 g1335 ( .a(n6987), .b(n8063), .c(n6985), .d(n8064_1), .o(n8065) );
in01f01 g1336 ( .a(net_7007), .o(n8066) );
in01f01 g1337 ( .a(net_7071), .o(n8067_1) );
oa22f01 g1338 ( .a(n6992), .b(n8066), .c(n6991), .d(n8067_1), .o(n8068) );
no02f01 g1339 ( .a(n8068), .b(n8065), .o(n8069) );
oa22f01 g1340 ( .a(n8069), .b(n6980), .c(n6995_1), .d(n8062), .o(n8070) );
no03f01 g1341 ( .a(n8070), .b(n8061), .c(n8053), .o(n8071) );
in01f01 g1342 ( .a(net_7019), .o(n8072_1) );
in01f01 g1343 ( .a(net_6987), .o(n8073) );
na04f01 g1344 ( .a(n7011), .b(n7003), .c(n6979), .d(_net_7092), .o(n8074) );
na04f01 g1345 ( .a(n7011), .b(n7000_1), .c(n6979), .d(_net_7092), .o(n8075_1) );
oa22f01 g1346 ( .a(n8075_1), .b(n8073), .c(n8074), .d(n8072_1), .o(n8076) );
in01f01 g1347 ( .a(net_7083), .o(n8077) );
in01f01 g1348 ( .a(net_7051), .o(n8078) );
na04f01 g1349 ( .a(n7011), .b(n6999), .c(n6979), .d(_net_7092), .o(n8079) );
na04f01 g1350 ( .a(n7011), .b(n7002), .c(n6979), .d(_net_7092), .o(n8080_1) );
oa22f01 g1351 ( .a(n8080_1), .b(n8077), .c(n8079), .d(n8078), .o(n8081) );
no02f01 g1352 ( .a(n8081), .b(n8076), .o(n8082) );
na02f01 g1353 ( .a(n8082), .b(n8071), .o(n1893) );
in01f01 g1354 ( .a(_net_6411), .o(n8084) );
na04f01 g1355 ( .a(_net_6407), .b(_net_6410), .c(_net_6406), .d(n8084), .o(n8085_1) );
no02f01 g1356 ( .a(_net_6409), .b(_net_6408), .o(n8086) );
in01f01 g1357 ( .a(n8086), .o(n8087) );
in01f01 g1358 ( .a(_net_6404), .o(n8088_1) );
no02f01 g1359 ( .a(_net_6405), .b(n8088_1), .o(n8089) );
in01f01 g1360 ( .a(n8089), .o(n8090) );
no03f01 g1361 ( .a(n8090), .b(n8087), .c(n8085_1), .o(n1898) );
no02f01 g1362 ( .a(n6881_1), .b(n6876_1), .o(n8092_1) );
in01f01 g1363 ( .a(_net_190), .o(n8093) );
in01f01 g1364 ( .a(_net_267), .o(n8094) );
no02f01 g1365 ( .a(n8094), .b(n8093), .o(n3638) );
in01f01 g1366 ( .a(n3638), .o(n8096) );
na02f01 g1367 ( .a(_net_267), .b(n8093), .o(n8097_1) );
oa22f01 g1368 ( .a(n8097_1), .b(n6875), .c(n8096), .d(n8092_1), .o(n1908) );
in01f01 g1369 ( .a(net_6430), .o(n8099) );
in01f01 g1370 ( .a(net_6494), .o(n8100) );
oa22f01 g1371 ( .a(n6750), .b(n8099), .c(n6748), .d(n8100), .o(n8101) );
in01f01 g1372 ( .a(net_6462), .o(n8102_1) );
in01f01 g1373 ( .a(net_6526), .o(n8103) );
oa22f01 g1374 ( .a(n6755), .b(n8102_1), .c(n6754), .d(n8103), .o(n8104) );
oa12f01 g1375 ( .a(n8028_1), .b(n8104), .c(n8101), .o(n8105) );
ao22f01 g1376 ( .a(n6777), .b(net_6428), .c(n6776), .d(net_6492), .o(n8106) );
ao22f01 g1377 ( .a(n6780), .b(net_6460), .c(n6779_1), .d(net_6524), .o(n8107_1) );
na02f01 g1378 ( .a(n8107_1), .b(n8106), .o(n8108) );
ao22f01 g1379 ( .a(n8108), .b(n8033_1), .c(n8034), .d(_net_6070), .o(n8109) );
in01f01 g1380 ( .a(n6764), .o(n8110) );
na02f01 g1381 ( .a(n6781), .b(n6778), .o(n8111) );
na02f01 g1382 ( .a(n6763), .b(n6762), .o(n8112_1) );
no02f01 g1383 ( .a(n8112_1), .b(n6758), .o(n8113) );
ao22f01 g1384 ( .a(n6777), .b(net_6426), .c(n6776), .d(net_6490), .o(n8114) );
ao22f01 g1385 ( .a(n6780), .b(net_6458), .c(n6779_1), .d(net_6522), .o(n8115) );
na02f01 g1386 ( .a(n8115), .b(n8114), .o(n8116_1) );
ao22f01 g1387 ( .a(n8116_1), .b(n8110), .c(n8113), .d(n8111), .o(n8117) );
na03f01 g1388 ( .a(n8117), .b(n8109), .c(n8105), .o(n1922) );
in01f01 g1389 ( .a(_net_6690), .o(n8119) );
no02f01 g1390 ( .a(n6943_1), .b(n6918), .o(n8120) );
na03f01 g1391 ( .a(n8120), .b(_net_6689), .c(n8119), .o(n8121_1) );
in01f01 g1392 ( .a(n8120), .o(n8122) );
oa12f01 g1393 ( .a(_net_6690), .b(n8122), .c(n6921), .o(n8123) );
na02f01 g1394 ( .a(n8123), .b(n8121_1), .o(n8124) );
no04f01 g1395 ( .a(n6914), .b(n6912), .c(_net_5998), .d(_net_5997), .o(n8125_1) );
na02f01 g1396 ( .a(n8125_1), .b(n8124), .o(n8126) );
no03f01 g1397 ( .a(n6944), .b(n6914), .c(n6912), .o(n8127) );
no02f01 g1398 ( .a(n6925), .b(n8119), .o(n8128) );
no02f01 g1399 ( .a(n6926), .b(_net_6690), .o(n8129) );
no02f01 g1400 ( .a(n8129), .b(n8128), .o(n8130_1) );
in01f01 g1401 ( .a(n6914), .o(n8131) );
no02f01 g1402 ( .a(n8131), .b(n6912), .o(n8132) );
ao22f01 g1403 ( .a(n8132), .b(_net_6690), .c(n8130_1), .d(n8127), .o(n8133) );
na02f01 g1404 ( .a(n8133), .b(n8126), .o(n1927) );
ao22f01 g1405 ( .a(n6736_1), .b(_net_7627), .c(n6734), .d(_net_7595), .o(n8135_1) );
ao22f01 g1406 ( .a(n6739), .b(_net_7659), .c(n6738), .d(_net_7563), .o(n8136) );
na02f01 g1407 ( .a(n8136), .b(n8135_1), .o(n1936) );
in01f01 g1408 ( .a(_net_7472), .o(n8138) );
na02f01 g1409 ( .a(n6866), .b(net_7392), .o(n8139) );
ao22f01 g1410 ( .a(_net_281), .b(net_353), .c(net_355), .d(_net_280), .o(n8140_1) );
na02f01 g1411 ( .a(n8140_1), .b(n8139), .o(n8141) );
na02f01 g1412 ( .a(n8141), .b(n6869), .o(n8142) );
oa12f01 g1413 ( .a(n8142), .b(n6869), .c(n8138), .o(n1945) );
in01f01 g1414 ( .a(n7854), .o(n8144_1) );
na02f01 g1415 ( .a(n6867_1), .b(n7846), .o(n8145) );
na02f01 g1416 ( .a(n6866), .b(_net_7532), .o(n8146) );
na02f01 g1417 ( .a(n8146), .b(n8145), .o(n8147_1) );
oa22f01 g1418 ( .a(n8147_1), .b(n7844), .c(n8144_1), .d(n7846), .o(n1950) );
in01f01 g1419 ( .a(_net_129), .o(n8149) );
na02f01 g1420 ( .a(_net_154), .b(net_325), .o(n8150) );
oa12f01 g1421 ( .a(n8150), .b(_net_154), .c(n8149), .o(n1959) );
in01f01 g1422 ( .a(_net_7594), .o(n8152_1) );
na02f01 g1423 ( .a(n7707), .b(n6968), .o(n8153) );
oa12f01 g1424 ( .a(n8153), .b(n6968), .c(n8152_1), .o(n1969) );
ao22f01 g1425 ( .a(n7130), .b(net_6698), .c(n7127), .d(net_6762), .o(n8155) );
ao22f01 g1426 ( .a(n7135), .b(net_6730), .c(n7133_1), .d(net_6794), .o(n8156_1) );
na02f01 g1427 ( .a(n8156_1), .b(n8155), .o(n8157) );
na02f01 g1428 ( .a(n8157), .b(n7124), .o(n8158) );
in01f01 g1429 ( .a(n7470), .o(n8159) );
ao22f01 g1430 ( .a(n7130), .b(net_6696), .c(n7127), .d(net_6760), .o(n8160) );
ao22f01 g1431 ( .a(n7135), .b(net_6728), .c(n7133_1), .d(net_6792), .o(n8161_1) );
na02f01 g1432 ( .a(n8161_1), .b(n8160), .o(n8162) );
ao22f01 g1433 ( .a(n8162), .b(n8159), .c(n7119), .d(_net_6108), .o(n8163) );
in01f01 g1434 ( .a(n7468_1), .o(n8164) );
na02f01 g1435 ( .a(n8164), .b(n7137), .o(n8165) );
na02f01 g1436 ( .a(n7467), .b(n7122), .o(n8166_1) );
no02f01 g1437 ( .a(n8166_1), .b(n7466), .o(n8167) );
oa12f01 g1438 ( .a(n8167), .b(n7485), .c(n7482_1), .o(n8168) );
na04f01 g1439 ( .a(n8168), .b(n8165), .c(n8163), .d(n8158), .o(n1988) );
in01f01 g1440 ( .a(net_357), .o(n8170_1) );
no02f01 g1441 ( .a(n6867_1), .b(n8170_1), .o(n1993) );
in01f01 g1442 ( .a(_net_7426), .o(n8172) );
in01f01 g1443 ( .a(net_359), .o(n8173) );
no02f01 g1444 ( .a(n6867_1), .b(n8173), .o(n2256) );
na02f01 g1445 ( .a(n2256), .b(n7550), .o(n8175) );
oa12f01 g1446 ( .a(n8175), .b(n7550), .c(n8172), .o(n2016) );
no02f01 g1447 ( .a(_net_6410), .b(_net_6411), .o(n8177) );
na02f01 g1448 ( .a(_net_6409), .b(_net_6408), .o(n8178) );
oa12f01 g1449 ( .a(_net_6407), .b(_net_6405), .c(_net_6406), .o(n8179_1) );
oa12f01 g1450 ( .a(n8177), .b(n8179_1), .c(n8178), .o(n2021) );
ao22f01 g1451 ( .a(n7130), .b(net_6697), .c(n7127), .d(net_6761), .o(n8181) );
ao22f01 g1452 ( .a(n7135), .b(net_6729), .c(n7133_1), .d(net_6793), .o(n8182) );
na02f01 g1453 ( .a(n8182), .b(n8181), .o(n8183_1) );
na02f01 g1454 ( .a(n8183_1), .b(n7124), .o(n8184) );
ao22f01 g1455 ( .a(n7130), .b(net_6695), .c(n7127), .d(net_6759), .o(n8185) );
ao22f01 g1456 ( .a(n7135), .b(net_6727), .c(n7133_1), .d(net_6791), .o(n8186) );
na02f01 g1457 ( .a(n8186), .b(n8185), .o(n8187) );
ao22f01 g1458 ( .a(n8187), .b(n8159), .c(n7119), .d(_net_6107), .o(n8188_1) );
na02f01 g1459 ( .a(n8188_1), .b(n8184), .o(n2026) );
in01f01 g1460 ( .a(_net_7483), .o(n8190) );
in01f01 g1461 ( .a(net_352), .o(n8191) );
in01f01 g1462 ( .a(_net_281), .o(n8192_1) );
oa22f01 g1463 ( .a(n6867_1), .b(n8191), .c(n8192_1), .d(n7978), .o(n8193) );
na02f01 g1464 ( .a(n8193), .b(n6869), .o(n8194) );
oa12f01 g1465 ( .a(n8194), .b(n6869), .c(n8190), .o(n2041) );
na02f01 g1466 ( .a(n7218), .b(n6984), .o(n8196) );
na02f01 g1467 ( .a(n7010), .b(_net_7093), .o(n8197_1) );
na02f01 g1468 ( .a(_net_7092), .b(n6984), .o(n8198) );
na02f01 g1469 ( .a(n8198), .b(n8197_1), .o(n8199) );
ao22f01 g1470 ( .a(n8199), .b(n7215), .c(n7220), .d(_net_7093), .o(n8200) );
na02f01 g1471 ( .a(n8200), .b(n8196), .o(n2046) );
in01f01 g1472 ( .a(_net_7465), .o(n8202_1) );
na02f01 g1473 ( .a(n7779_1), .b(n6869), .o(n8203) );
oa12f01 g1474 ( .a(n8203), .b(n6869), .c(n8202_1), .o(n2055) );
in01f01 g1475 ( .a(_net_7352), .o(n8205) );
na02f01 g1476 ( .a(n6898), .b(net_7240), .o(n8206_1) );
ao22f01 g1477 ( .a(net_332), .b(_net_270), .c(_net_269), .d(net_334), .o(n8207) );
na02f01 g1478 ( .a(n8207), .b(n8206_1), .o(n8208) );
na02f01 g1479 ( .a(n8208), .b(n7030), .o(n8209) );
oa12f01 g1480 ( .a(n8209), .b(n7030), .c(n8205), .o(n2060) );
in01f01 g1481 ( .a(n6844), .o(n8211_1) );
na02f01 g1482 ( .a(n8211_1), .b(_net_6125), .o(n8212) );
in01f01 g1483 ( .a(n6836_1), .o(n8213) );
ao22f01 g1484 ( .a(n6811), .b(net_6830), .c(n6808), .d(net_6894), .o(n8214) );
ao22f01 g1485 ( .a(n6816), .b(net_6862), .c(n6814), .d(net_6926), .o(n8215) );
na02f01 g1486 ( .a(n8215), .b(n8214), .o(n8216_1) );
na02f01 g1487 ( .a(n8216_1), .b(n8213), .o(n8217) );
na02f01 g1488 ( .a(n8217), .b(n8212), .o(n2065) );
in01f01 g1489 ( .a(_net_6827), .o(n8219) );
in01f01 g1490 ( .a(net_6826), .o(n8220_1) );
no02f01 g1491 ( .a(n8220_1), .b(_net_6827), .o(n8221) );
no02f01 g1492 ( .a(net_6826), .b(n8219), .o(n8222) );
no02f01 g1493 ( .a(n8222), .b(n8221), .o(n8223) );
in01f01 g1494 ( .a(_net_5971), .o(n8224_1) );
no02f01 g1495 ( .a(n8224_1), .b(n7121), .o(n6427) );
in01f01 g1496 ( .a(n6427), .o(n8226) );
na02f01 g1497 ( .a(n8224_1), .b(_net_6006), .o(n8227) );
oa22f01 g1498 ( .a(n8227), .b(n8219), .c(n8226), .d(n8223), .o(n2070) );
in01f01 g1499 ( .a(net_339), .o(n8229) );
no02f01 g1500 ( .a(n6899_1), .b(n8229), .o(n2084) );
in01f01 g1501 ( .a(_net_7683), .o(n8231) );
na02f01 g1502 ( .a(n6964_1), .b(_net_289), .o(n8232_1) );
na02f01 g1503 ( .a(n6966), .b(n8231), .o(n8233) );
na02f01 g1504 ( .a(n6965), .b(_net_7683), .o(n8234) );
na02f01 g1505 ( .a(n8234), .b(n8233), .o(n8235) );
in01f01 g1506 ( .a(_net_289), .o(n8236) );
no02f01 g1507 ( .a(n6964_1), .b(n8236), .o(n8237_1) );
in01f01 g1508 ( .a(n8237_1), .o(n8238) );
oa22f01 g1509 ( .a(n8238), .b(n8231), .c(n8235), .d(n8232_1), .o(n2140) );
in01f01 g1510 ( .a(_net_7554), .o(n8240) );
na02f01 g1511 ( .a(n8000), .b(n7519), .o(n8241_1) );
oa12f01 g1512 ( .a(n8241_1), .b(n7519), .c(n8240), .o(n2162) );
in01f01 g1513 ( .a(_net_7649), .o(n8243) );
na02f01 g1514 ( .a(n6965), .b(net_7537), .o(n8244) );
ao22f01 g1515 ( .a(_net_292), .b(net_367), .c(_net_291), .d(net_369), .o(n8245_1) );
na02f01 g1516 ( .a(n8245_1), .b(n8244), .o(n8246) );
na02f01 g1517 ( .a(n8246), .b(n7446_1), .o(n8247) );
oa12f01 g1518 ( .a(n8247), .b(n7446_1), .c(n8243), .o(n2167) );
in01f01 g1519 ( .a(_net_6963), .o(n8249_1) );
in01f01 g1520 ( .a(n1345), .o(n8250) );
ao12f01 g1521 ( .a(n8249_1), .b(_net_6962), .c(net_6961), .o(n8251) );
in01f01 g1522 ( .a(net_6961), .o(n8252) );
in01f01 g1523 ( .a(_net_6962), .o(n8253_1) );
no03f01 g1524 ( .a(n8253_1), .b(_net_6963), .c(n8252), .o(n8254) );
no02f01 g1525 ( .a(n8254), .b(n8251), .o(n8255) );
na02f01 g1526 ( .a(_net_6017), .b(n7682), .o(n8256) );
oa22f01 g1527 ( .a(n8256), .b(n8249_1), .c(n8255), .d(n8250), .o(n2172) );
na02f01 g1528 ( .a(n7298), .b(net_7737), .o(n8258_1) );
ao22f01 g1529 ( .a(n7306), .b(_net_6007), .c(n7291), .d(net_7708), .o(n8259) );
na02f01 g1530 ( .a(n7302_1), .b(net_147), .o(n8260) );
na02f01 g1531 ( .a(n7296), .b(net_247), .o(n8261) );
na03f01 g1532 ( .a(n7308), .b(_net_173), .c(n6800), .o(n8262_1) );
na03f01 g1533 ( .a(n7308), .b(_net_210), .c(x1322), .o(n8263) );
na03f01 g1534 ( .a(n8263), .b(n8262_1), .c(n8261), .o(n8264) );
ao12f01 g1535 ( .a(n8264), .b(n7286), .c(_net_290), .o(n8265) );
na04f01 g1536 ( .a(n8265), .b(n8260), .c(n8259), .d(n8258_1), .o(n2177) );
no02f01 g1537 ( .a(n6864), .b(n6863_1), .o(n2181) );
in01f01 g1538 ( .a(net_7108), .o(n8268) );
in01f01 g1539 ( .a(net_7172), .o(n8269) );
oa22f01 g1540 ( .a(n7580), .b(n8268), .c(n7577_1), .d(n8269), .o(n8270) );
in01f01 g1541 ( .a(net_7204), .o(n8271_1) );
in01f01 g1542 ( .a(net_7140), .o(n8272) );
oa22f01 g1543 ( .a(n7585), .b(n8272), .c(n7583), .d(n8271_1), .o(n8273) );
no02f01 g1544 ( .a(n8273), .b(n8270), .o(n8274) );
no02f01 g1545 ( .a(n8274), .b(n7721), .o(n8275) );
in01f01 g1546 ( .a(net_7174), .o(n8276_1) );
in01f01 g1547 ( .a(net_7110), .o(n8277) );
oa22f01 g1548 ( .a(n7580), .b(n8277), .c(n7577_1), .d(n8276_1), .o(n8278) );
in01f01 g1549 ( .a(net_7142), .o(n8279) );
in01f01 g1550 ( .a(net_7206), .o(n8280_1) );
oa22f01 g1551 ( .a(n7585), .b(n8279), .c(n7583), .d(n8280_1), .o(n8281) );
no02f01 g1552 ( .a(n8281), .b(n8278), .o(n8282) );
no02f01 g1553 ( .a(n8282), .b(n7592), .o(n8283) );
in01f01 g1554 ( .a(_net_6177), .o(n8284_1) );
in01f01 g1555 ( .a(net_7176), .o(n8285) );
in01f01 g1556 ( .a(net_7112), .o(n8286) );
oa22f01 g1557 ( .a(n7580), .b(n8286), .c(n7577_1), .d(n8285), .o(n8287) );
in01f01 g1558 ( .a(net_7144), .o(n8288) );
in01f01 g1559 ( .a(net_7208), .o(n8289_1) );
oa22f01 g1560 ( .a(n7585), .b(n8288), .c(n7583), .d(n8289_1), .o(n8290) );
no02f01 g1561 ( .a(n8290), .b(n8287), .o(n8291) );
oa22f01 g1562 ( .a(n8291), .b(n7574), .c(n7590), .d(n8284_1), .o(n8292) );
no03f01 g1563 ( .a(n8292), .b(n8283), .c(n8275), .o(n8293) );
in01f01 g1564 ( .a(net_7124), .o(n8294_1) );
in01f01 g1565 ( .a(net_7156), .o(n8295) );
oa22f01 g1566 ( .a(n7740), .b(n8294_1), .c(n7739), .d(n8295), .o(n8296) );
in01f01 g1567 ( .a(net_7220), .o(n8297) );
in01f01 g1568 ( .a(net_7188), .o(n8298) );
oa22f01 g1569 ( .a(n7745), .b(n8297), .c(n7744), .d(n8298), .o(n8299_1) );
no02f01 g1570 ( .a(n8299_1), .b(n8296), .o(n8300) );
na02f01 g1571 ( .a(n8300), .b(n8293), .o(n2194) );
no02f01 g1572 ( .a(n7576), .b(n7719_1), .o(n8302) );
na02f01 g1573 ( .a(n8302), .b(n7579), .o(n8303_1) );
in01f01 g1574 ( .a(n8302), .o(n8304) );
na02f01 g1575 ( .a(n8304), .b(_net_7229), .o(n8305) );
na02f01 g1576 ( .a(n8305), .b(n8303_1), .o(n8306) );
no04f01 g1577 ( .a(n7572_1), .b(n7570), .c(_net_6041), .d(_net_6042), .o(n8307_1) );
na02f01 g1578 ( .a(n8307_1), .b(n8306), .o(n8308) );
na02f01 g1579 ( .a(n7585), .b(n7577_1), .o(n8309) );
no03f01 g1580 ( .a(n7720), .b(n7572_1), .c(n7570), .o(n8310) );
in01f01 g1581 ( .a(n7572_1), .o(n8311_1) );
no02f01 g1582 ( .a(n8311_1), .b(n7570), .o(n8312) );
ao22f01 g1583 ( .a(n8312), .b(_net_7229), .c(n8310), .d(n8309), .o(n8313) );
na02f01 g1584 ( .a(n8313), .b(n8308), .o(n2199) );
in01f01 g1585 ( .a(n7304), .o(n8315) );
no02f01 g1586 ( .a(n7111_1), .b(n7341), .o(n8316_1) );
na03f01 g1587 ( .a(n8316_1), .b(n7281), .c(n6800), .o(n8317) );
no02f01 g1588 ( .a(n8317), .b(n8315), .o(n2208) );
ao12f01 g1589 ( .a(n8224_1), .b(_net_6828), .c(_net_6825), .o(n8319) );
oa12f01 g1590 ( .a(n8319), .b(_net_6828), .c(_net_6825), .o(n8320_1) );
no02f01 g1591 ( .a(n7128_1), .b(_net_6827), .o(n8321) );
no02f01 g1592 ( .a(_net_6824), .b(n8219), .o(n8322) );
no02f01 g1593 ( .a(n8322), .b(n8321), .o(n8323) );
no02f01 g1594 ( .a(n7125_1), .b(n8220_1), .o(n8324_1) );
no02f01 g1595 ( .a(_net_6823), .b(net_6826), .o(n8325) );
no02f01 g1596 ( .a(n8325), .b(n8324_1), .o(n8326) );
in01f01 g1597 ( .a(n8326), .o(n2948) );
na02f01 g1598 ( .a(n2948), .b(n8323), .o(n8328) );
oa12f01 g1599 ( .a(n7633), .b(n8328), .c(n8320_1), .o(n2213) );
in01f01 g1600 ( .a(_net_5963), .o(n8330) );
no02f01 g1601 ( .a(n6759), .b(n8330), .o(n2222) );
in01f01 g1602 ( .a(_net_6960), .o(n8332) );
no02f01 g1603 ( .a(n6806_1), .b(n6818_1), .o(n8333) );
na03f01 g1604 ( .a(n8333), .b(_net_6959), .c(n8332), .o(n8334_1) );
in01f01 g1605 ( .a(n8333), .o(n8335) );
oa12f01 g1606 ( .a(_net_6960), .b(n8335), .c(n6809_1), .o(n8336) );
na02f01 g1607 ( .a(n8336), .b(n8334_1), .o(n8337_1) );
no04f01 g1608 ( .a(n6821), .b(n6819), .c(_net_6020), .d(_net_6019), .o(n8338) );
na02f01 g1609 ( .a(n8338), .b(n8337_1), .o(n8339) );
no03f01 g1610 ( .a(n6823), .b(n6821), .c(n6819), .o(n8340_1) );
no02f01 g1611 ( .a(n6813_1), .b(n8332), .o(n8341) );
no02f01 g1612 ( .a(n6814), .b(_net_6960), .o(n8342) );
no02f01 g1613 ( .a(n8342), .b(n8341), .o(n8343) );
in01f01 g1614 ( .a(n6821), .o(n8344) );
no02f01 g1615 ( .a(n8344), .b(n6819), .o(n8345_1) );
ao22f01 g1616 ( .a(n8345_1), .b(_net_6960), .c(n8343), .d(n8340_1), .o(n8346) );
na02f01 g1617 ( .a(n8346), .b(n8339), .o(n2227) );
in01f01 g1618 ( .a(_net_7686), .o(n8348) );
in01f01 g1619 ( .a(_net_7682), .o(n8349) );
no02f01 g1620 ( .a(n8349), .b(n8348), .o(n8350_1) );
no02f01 g1621 ( .a(_net_7682), .b(_net_7686), .o(n8351) );
no02f01 g1622 ( .a(n8351), .b(n8350_1), .o(n8352) );
in01f01 g1623 ( .a(n8352), .o(n8353) );
no02f01 g1624 ( .a(n6733), .b(n6959), .o(n8354_1) );
no02f01 g1625 ( .a(net_7680), .b(_net_7684), .o(n8355) );
no02f01 g1626 ( .a(n8355), .b(n8354_1), .o(n8356) );
in01f01 g1627 ( .a(n8356), .o(n4405) );
no02f01 g1628 ( .a(n7397), .b(n6735), .o(n8358) );
no02f01 g1629 ( .a(_net_7685), .b(_net_7681), .o(n8359_1) );
no02f01 g1630 ( .a(n8359_1), .b(n8358), .o(n8360) );
in01f01 g1631 ( .a(n8360), .o(n8361) );
na02f01 g1632 ( .a(n8361), .b(n4405), .o(n8362_1) );
no02f01 g1633 ( .a(n8362_1), .b(n8353), .o(n2232) );
no02f01 g1634 ( .a(n7342), .b(n7111_1), .o(n2237) );
in01f01 g1635 ( .a(_net_7724), .o(n8365) );
in01f01 g1636 ( .a(_net_5994), .o(n8366) );
ao12f01 g1637 ( .a(n7343), .b(n8366), .c(n8365), .o(n2242) );
ao22f01 g1638 ( .a(n7288_1), .b(_net_6044), .c(n7286), .d(_net_283), .o(n8368) );
ao22f01 g1639 ( .a(n7298), .b(_net_7733), .c(n7291), .d(_net_7704), .o(n8369) );
na02f01 g1640 ( .a(n7302_1), .b(_net_127), .o(n8370) );
na03f01 g1641 ( .a(n7308), .b(net_206), .c(x1322), .o(n8371) );
na02f01 g1642 ( .a(n7296), .b(net_243), .o(n8372_1) );
na03f01 g1643 ( .a(n7308), .b(net_169), .c(n6800), .o(n8373) );
na03f01 g1644 ( .a(n8373), .b(n8372_1), .c(n8371), .o(n8374) );
ao12f01 g1645 ( .a(n8374), .b(n7306), .c(_net_6000), .o(n8375) );
na04f01 g1646 ( .a(n8375), .b(n8370), .c(n8369), .d(n8368), .o(n2247) );
in01f01 g1647 ( .a(_net_6402), .o(n8377_1) );
na02f01 g1648 ( .a(n8377_1), .b(net_6403), .o(n8378) );
in01f01 g1649 ( .a(net_6403), .o(n8379) );
na02f01 g1650 ( .a(_net_6402), .b(n8379), .o(n8380) );
na02f01 g1651 ( .a(n8380), .b(n8378), .o(n2251) );
in01f01 g1652 ( .a(_net_7401), .o(n8382_1) );
na02f01 g1653 ( .a(n7779_1), .b(n7550), .o(n8383) );
oa12f01 g1654 ( .a(n8383), .b(n7550), .c(n8382_1), .o(n2265) );
in01f01 g1655 ( .a(net_7096), .o(n8385) );
no02f01 g1656 ( .a(n8385), .b(n6984), .o(n8386) );
no02f01 g1657 ( .a(net_7096), .b(_net_7093), .o(n8387_1) );
no02f01 g1658 ( .a(n8387_1), .b(n8386), .o(n8388) );
in01f01 g1659 ( .a(n8388), .o(n2270) );
no02f01 g1660 ( .a(n7612), .b(n6824), .o(n8390) );
in01f01 g1661 ( .a(net_6906), .o(n8391) );
in01f01 g1662 ( .a(net_6842), .o(n8392_1) );
oa22f01 g1663 ( .a(n6810), .b(n8392_1), .c(n6807), .d(n8391), .o(n8393) );
in01f01 g1664 ( .a(net_6938), .o(n8394) );
in01f01 g1665 ( .a(net_6874), .o(n8395) );
oa22f01 g1666 ( .a(n6815), .b(n8395), .c(n6813_1), .d(n8394), .o(n8396_1) );
no02f01 g1667 ( .a(n8396_1), .b(n8393), .o(n8397) );
no02f01 g1668 ( .a(n8397), .b(n6826_1), .o(n8398) );
in01f01 g1669 ( .a(_net_6139), .o(n8399) );
in01f01 g1670 ( .a(net_6844), .o(n8400) );
in01f01 g1671 ( .a(net_6908), .o(n8401_1) );
oa22f01 g1672 ( .a(n6810), .b(n8400), .c(n6807), .d(n8401_1), .o(n8402) );
in01f01 g1673 ( .a(net_6940), .o(n8403) );
in01f01 g1674 ( .a(net_6876), .o(n8404) );
oa22f01 g1675 ( .a(n6815), .b(n8404), .c(n6813_1), .d(n8403), .o(n8405_1) );
no02f01 g1676 ( .a(n8405_1), .b(n8402), .o(n8406) );
oa22f01 g1677 ( .a(n8406), .b(n6836_1), .c(n6844), .d(n8399), .o(n8407) );
no03f01 g1678 ( .a(n8407), .b(n8398), .c(n8390), .o(n8408) );
in01f01 g1679 ( .a(net_6856), .o(n8409) );
in01f01 g1680 ( .a(net_6888), .o(n8410_1) );
oa22f01 g1681 ( .a(n6850_1), .b(n8409), .c(n6849), .d(n8410_1), .o(n8411) );
in01f01 g1682 ( .a(net_6952), .o(n8412) );
in01f01 g1683 ( .a(net_6920), .o(n8413) );
oa22f01 g1684 ( .a(n6855_1), .b(n8412), .c(n6854), .d(n8413), .o(n8414) );
no02f01 g1685 ( .a(n8414), .b(n8411), .o(n8415_1) );
na02f01 g1686 ( .a(n8415_1), .b(n8408), .o(n2275) );
in01f01 g1687 ( .a(_net_7748), .o(n8417) );
ao12f01 g1688 ( .a(n7343), .b(n8417), .c(n7652), .o(n2280) );
in01f01 g1689 ( .a(_net_6015), .o(n8419) );
oa12f01 g1690 ( .a(n8419), .b(n7117), .c(n7261), .o(n2298) );
in01f01 g1691 ( .a(_net_6186), .o(n8421) );
no02f01 g1692 ( .a(n8421), .b(_net_392), .o(n2303) );
in01f01 g1693 ( .a(_net_7556), .o(n8423) );
na02f01 g1694 ( .a(n6965), .b(net_7540), .o(n8424) );
ao22f01 g1695 ( .a(_net_292), .b(net_370), .c(_net_291), .d(net_372), .o(n8425) );
na02f01 g1696 ( .a(n8425), .b(n8424), .o(n8426_1) );
na02f01 g1697 ( .a(n8426_1), .b(n7519), .o(n8427) );
oa12f01 g1698 ( .a(n8427), .b(n7519), .c(n8423), .o(n2312) );
in01f01 g1699 ( .a(net_6899), .o(n8429) );
in01f01 g1700 ( .a(net_6835), .o(n8430_1) );
oa22f01 g1701 ( .a(n6810), .b(n8430_1), .c(n6807), .d(n8429), .o(n8431) );
in01f01 g1702 ( .a(net_6867), .o(n8432) );
in01f01 g1703 ( .a(net_6931), .o(n8433) );
oa22f01 g1704 ( .a(n6815), .b(n8432), .c(n6813_1), .d(n8433), .o(n8434) );
no02f01 g1705 ( .a(n8434), .b(n8431), .o(n8435_1) );
no02f01 g1706 ( .a(n8435_1), .b(n6824), .o(n8436) );
in01f01 g1707 ( .a(net_6901), .o(n8437) );
in01f01 g1708 ( .a(net_6837), .o(n8438_1) );
oa22f01 g1709 ( .a(n6810), .b(n8438_1), .c(n6807), .d(n8437), .o(n8439) );
in01f01 g1710 ( .a(net_6933), .o(n8440) );
in01f01 g1711 ( .a(net_6869), .o(n8441) );
oa22f01 g1712 ( .a(n6815), .b(n8441), .c(n6813_1), .d(n8440), .o(n8442) );
no02f01 g1713 ( .a(n8442), .b(n8439), .o(n8443_1) );
no02f01 g1714 ( .a(n8443_1), .b(n6826_1), .o(n8444) );
in01f01 g1715 ( .a(_net_6134), .o(n8445) );
in01f01 g1716 ( .a(net_6903), .o(n8446) );
in01f01 g1717 ( .a(net_6839), .o(n8447_1) );
oa22f01 g1718 ( .a(n6810), .b(n8447_1), .c(n6807), .d(n8446), .o(n8448) );
in01f01 g1719 ( .a(net_6935), .o(n8449) );
in01f01 g1720 ( .a(net_6871), .o(n8450) );
oa22f01 g1721 ( .a(n6815), .b(n8450), .c(n6813_1), .d(n8449), .o(n8451_1) );
no02f01 g1722 ( .a(n8451_1), .b(n8448), .o(n8452) );
oa22f01 g1723 ( .a(n8452), .b(n6836_1), .c(n6844), .d(n8445), .o(n8453) );
no03f01 g1724 ( .a(n8453), .b(n8444), .c(n8436), .o(n8454) );
in01f01 g1725 ( .a(net_6883), .o(n8455_1) );
in01f01 g1726 ( .a(net_6851), .o(n8456) );
oa22f01 g1727 ( .a(n6850_1), .b(n8456), .c(n6849), .d(n8455_1), .o(n8457) );
in01f01 g1728 ( .a(net_6915), .o(n8458) );
in01f01 g1729 ( .a(net_6947), .o(n8459_1) );
oa22f01 g1730 ( .a(n6855_1), .b(n8459_1), .c(n6854), .d(n8458), .o(n8460) );
no02f01 g1731 ( .a(n8460), .b(n8457), .o(n8461) );
na02f01 g1732 ( .a(n8461), .b(n8454), .o(n2329) );
in01f01 g1733 ( .a(_net_7747), .o(n8463) );
ao12f01 g1734 ( .a(n7343), .b(n8463), .c(n6907), .o(n2334) );
in01f01 g1735 ( .a(net_6979), .o(n8465) );
in01f01 g1736 ( .a(net_7043), .o(n8466) );
oa22f01 g1737 ( .a(n6987), .b(n8465), .c(n6985), .d(n8466), .o(n8467_1) );
in01f01 g1738 ( .a(net_7075), .o(n8468) );
in01f01 g1739 ( .a(net_7011), .o(n8469) );
oa22f01 g1740 ( .a(n6992), .b(n8469), .c(n6991), .d(n8468), .o(n8470) );
no02f01 g1741 ( .a(n8470), .b(n8467_1), .o(n8471) );
no02f01 g1742 ( .a(n8471), .b(n7012), .o(n8472_1) );
in01f01 g1743 ( .a(net_6981), .o(n8473) );
in01f01 g1744 ( .a(net_7045), .o(n8474) );
oa22f01 g1745 ( .a(n6987), .b(n8473), .c(n6985), .d(n8474), .o(n8475) );
in01f01 g1746 ( .a(net_7013), .o(n8476) );
in01f01 g1747 ( .a(net_7077), .o(n8477_1) );
oa22f01 g1748 ( .a(n6992), .b(n8476), .c(n6991), .d(n8477_1), .o(n8478) );
no02f01 g1749 ( .a(n8478), .b(n8475), .o(n8479) );
no02f01 g1750 ( .a(n8479), .b(n6997), .o(n8480) );
ao22f01 g1751 ( .a(n7000_1), .b(net_6983), .c(n6999), .d(net_7047), .o(n8481_1) );
ao22f01 g1752 ( .a(n7003), .b(net_7015), .c(n7002), .d(net_7079), .o(n8482) );
ao12f01 g1753 ( .a(n6980), .b(n8482), .c(n8481_1), .o(n8483) );
in01f01 g1754 ( .a(_net_6163), .o(n8484) );
no02f01 g1755 ( .a(n6995_1), .b(n8484), .o(n8485) );
no04f01 g1756 ( .a(n8485), .b(n8483), .c(n8480), .d(n8472_1), .o(n8486_1) );
in01f01 g1757 ( .a(net_6995), .o(n8487) );
in01f01 g1758 ( .a(net_7027), .o(n8488) );
oa22f01 g1759 ( .a(n8075_1), .b(n8487), .c(n8074), .d(n8488), .o(n8489) );
in01f01 g1760 ( .a(net_7091), .o(n8490) );
in01f01 g1761 ( .a(net_7059), .o(n8491_1) );
oa22f01 g1762 ( .a(n8080_1), .b(n8490), .c(n8079), .d(n8491_1), .o(n8492) );
no02f01 g1763 ( .a(n8492), .b(n8489), .o(n8493) );
na02f01 g1764 ( .a(n8493), .b(n8486_1), .o(n2365) );
no02f01 g1765 ( .a(_net_154), .b(_net_7720), .o(n8495) );
no02f01 g1766 ( .a(n8495), .b(n7343), .o(n2377) );
ao22f01 g1767 ( .a(n7581_1), .b(net_7104), .c(n7578), .d(net_7168), .o(n8497) );
ao22f01 g1768 ( .a(n7586_1), .b(net_7136), .c(n7584), .d(net_7200), .o(n8498) );
na02f01 g1769 ( .a(n8498), .b(n8497), .o(n8499_1) );
na02f01 g1770 ( .a(n8499_1), .b(n7575), .o(n8500) );
ao22f01 g1771 ( .a(n7593), .b(n7588), .c(n7591_1), .d(_net_6169), .o(n8501) );
na02f01 g1772 ( .a(n7914), .b(n7596_1), .o(n8502) );
in01f01 g1773 ( .a(net_7116), .o(n8503) );
in01f01 g1774 ( .a(net_7180), .o(n8504_1) );
oa22f01 g1775 ( .a(n7580), .b(n8503), .c(n7577_1), .d(n8504_1), .o(n8505) );
in01f01 g1776 ( .a(net_7148), .o(n8506) );
in01f01 g1777 ( .a(net_7212), .o(n8507) );
oa22f01 g1778 ( .a(n7585), .b(n8506), .c(n7583), .d(n8507), .o(n8508_1) );
oa12f01 g1779 ( .a(n7920_1), .b(n8508_1), .c(n8505), .o(n8509) );
na04f01 g1780 ( .a(n8509), .b(n8502), .c(n8501), .d(n8500), .o(n2386) );
ao22f01 g1781 ( .a(n6877), .b(_net_7277), .c(n6876_1), .d(net_7341), .o(n8511) );
ao22f01 g1782 ( .a(n6881_1), .b(net_7309), .c(n6880), .d(net_7373), .o(n8512) );
na02f01 g1783 ( .a(n8512), .b(n8511), .o(n2395) );
in01f01 g1784 ( .a(net_378), .o(n8514) );
no02f01 g1785 ( .a(n6966), .b(n8514), .o(n2404) );
in01f01 g1786 ( .a(_net_7511), .o(n8516) );
na02f01 g1787 ( .a(n7626_1), .b(n7504), .o(n8517_1) );
oa12f01 g1788 ( .a(n8517_1), .b(n7626_1), .c(n8516), .o(n2409) );
ao22f01 g1789 ( .a(n7288_1), .b(_net_6032), .c(n7286), .d(_net_271), .o(n8519) );
ao22f01 g1790 ( .a(n7298), .b(_net_7724), .c(n7291), .d(_net_7695), .o(n8520) );
na02f01 g1791 ( .a(n7302_1), .b(_net_118), .o(n8521) );
na03f01 g1792 ( .a(n7308), .b(net_197), .c(x1322), .o(n8522_1) );
na02f01 g1793 ( .a(n7296), .b(net_234), .o(n8523) );
na03f01 g1794 ( .a(n7308), .b(net_160), .c(n6800), .o(n8524) );
na03f01 g1795 ( .a(n8524), .b(n8523), .c(n8522_1), .o(n8525) );
ao12f01 g1796 ( .a(n8525), .b(n7306), .c(_net_5988), .o(n8526_1) );
na04f01 g1797 ( .a(n8526_1), .b(n8521), .c(n8520), .d(n8519), .o(n2414) );
in01f01 g1798 ( .a(_net_7431), .o(n8528) );
na02f01 g1799 ( .a(n1752), .b(n7550), .o(n8529) );
oa12f01 g1800 ( .a(n8529), .b(n7550), .c(n8528), .o(n2430) );
in01f01 g1801 ( .a(_net_279), .o(n8531_1) );
na02f01 g1802 ( .a(n7440), .b(net_7802), .o(n8532) );
oa12f01 g1803 ( .a(n8532), .b(n7440), .c(n8531_1), .o(n2435) );
na02f01 g1804 ( .a(n8337_1), .b(_net_6963), .o(n8534) );
na03f01 g1805 ( .a(n8336), .b(n8334_1), .c(n8249_1), .o(n8535_1) );
na02f01 g1806 ( .a(_net_6958), .b(n6818_1), .o(n8536) );
na02f01 g1807 ( .a(n6806_1), .b(_net_6957), .o(n8537) );
na02f01 g1808 ( .a(n8537), .b(n8536), .o(n8538) );
na02f01 g1809 ( .a(n8538), .b(net_6961), .o(n8539) );
na03f01 g1810 ( .a(n8537), .b(n8536), .c(n8252), .o(n8540_1) );
ao22f01 g1811 ( .a(n8540_1), .b(n8539), .c(n6823), .d(_net_6957), .o(n8541) );
na02f01 g1812 ( .a(n8333), .b(n6809_1), .o(n8542) );
na02f01 g1813 ( .a(n8335), .b(_net_6959), .o(n8543) );
na02f01 g1814 ( .a(n8543), .b(n8542), .o(n8544_1) );
na02f01 g1815 ( .a(n8544_1), .b(n8253_1), .o(n8545) );
na03f01 g1816 ( .a(n8543), .b(n8542), .c(_net_6962), .o(n8546) );
na03f01 g1817 ( .a(n8546), .b(n8545), .c(n8541), .o(n8547) );
ao12f01 g1818 ( .a(n8547), .b(n8535_1), .c(n8534), .o(n2444) );
na02f01 g1819 ( .a(n7348), .b(_net_7793), .o(n8549_1) );
oa12f01 g1820 ( .a(n8549_1), .b(n7348), .c(n6759), .o(n2457) );
in01f01 g1821 ( .a(net_6704), .o(n8551) );
in01f01 g1822 ( .a(net_6768), .o(n8552_1) );
oa22f01 g1823 ( .a(n7129), .b(n8551), .c(n7126), .d(n8552_1), .o(n8553) );
in01f01 g1824 ( .a(net_6800), .o(n8554) );
in01f01 g1825 ( .a(net_6736), .o(n8555) );
oa22f01 g1826 ( .a(n7134), .b(n8555), .c(n7132), .d(n8554), .o(n8556) );
no02f01 g1827 ( .a(n8556), .b(n8553), .o(n8557_1) );
no02f01 g1828 ( .a(n8557_1), .b(n7468_1), .o(n8558) );
no02f01 g1829 ( .a(n7470), .b(n7465), .o(n8559) );
in01f01 g1830 ( .a(_net_6118), .o(n8560) );
oa22f01 g1831 ( .a(n7477), .b(n7123), .c(n7118), .d(n8560), .o(n8561_1) );
no03f01 g1832 ( .a(n8561_1), .b(n8559), .c(n8558), .o(n8562) );
in01f01 g1833 ( .a(net_6720), .o(n8563) );
in01f01 g1834 ( .a(net_6752), .o(n8564) );
oa22f01 g1835 ( .a(n7492_1), .b(n8563), .c(n7491), .d(n8564), .o(n8565_1) );
in01f01 g1836 ( .a(net_6784), .o(n8566) );
in01f01 g1837 ( .a(net_6816), .o(n8567) );
oa22f01 g1838 ( .a(n7497), .b(n8567), .c(n7496_1), .d(n8566), .o(n8568) );
no02f01 g1839 ( .a(n8568), .b(n8565_1), .o(n8569) );
na02f01 g1840 ( .a(n8569), .b(n8562), .o(n2470) );
in01f01 g1841 ( .a(_net_7294), .o(n8571) );
na02f01 g1842 ( .a(n7926), .b(n7180), .o(n8572) );
oa12f01 g1843 ( .a(n8572), .b(n7180), .c(n8571), .o(n2479) );
ao22f01 g1844 ( .a(n7225), .b(_net_7432), .c(n7224), .d(net_7464), .o(n8574) );
ao22f01 g1845 ( .a(n7229), .b(net_7528), .c(n7228), .d(net_7496), .o(n8575_1) );
na02f01 g1846 ( .a(n8575_1), .b(n8574), .o(n2484) );
in01f01 g1847 ( .a(_net_7704), .o(n8577) );
na02f01 g1848 ( .a(n7207_1), .b(_net_7806), .o(n8578_1) );
oa12f01 g1849 ( .a(n8578_1), .b(n7207_1), .c(n8577), .o(n2505) );
ao22f01 g1850 ( .a(n6736_1), .b(net_7638), .c(n6734), .d(net_7606), .o(n8580) );
ao22f01 g1851 ( .a(n6739), .b(net_7670), .c(n6738), .d(_net_7574), .o(n8581) );
na02f01 g1852 ( .a(n8581), .b(n8580), .o(n2510) );
no03f01 g1853 ( .a(_net_6010), .b(n7121), .c(n7265_1), .o(n8583_1) );
no02f01 g1854 ( .a(n7121), .b(n7261), .o(n8584) );
ao22f01 g1855 ( .a(n8584), .b(n7271), .c(n8583_1), .d(n7269), .o(n8585) );
ao12f01 g1856 ( .a(n7121), .b(_net_5970), .c(n7261), .o(n8586) );
no03f01 g1857 ( .a(_net_6010), .b(n7121), .c(_net_6011), .o(n8587) );
ao22f01 g1858 ( .a(n8587), .b(n7267), .c(n8586), .d(n7260_1), .o(n8588_1) );
na02f01 g1859 ( .a(n8588_1), .b(n8585), .o(n2515) );
ao22f01 g1860 ( .a(n6877), .b(_net_7273), .c(n6876_1), .d(net_7337), .o(n8590) );
ao22f01 g1861 ( .a(n6881_1), .b(net_7305), .c(n6880), .d(net_7369), .o(n8591) );
na02f01 g1862 ( .a(n8591), .b(n8590), .o(n2524) );
in01f01 g1863 ( .a(_net_7419), .o(n8593_1) );
na02f01 g1864 ( .a(n8193), .b(n7550), .o(n8594) );
oa12f01 g1865 ( .a(n8594), .b(n7550), .c(n8593_1), .o(n2529) );
in01f01 g1866 ( .a(net_7040), .o(n8596) );
in01f01 g1867 ( .a(net_6976), .o(n8597) );
oa22f01 g1868 ( .a(n6987), .b(n8597), .c(n6985), .d(n8596), .o(n8598_1) );
in01f01 g1869 ( .a(net_7008), .o(n8599) );
in01f01 g1870 ( .a(net_7072), .o(n8600) );
oa22f01 g1871 ( .a(n6992), .b(n8599), .c(n6991), .d(n8600), .o(n8601) );
no02f01 g1872 ( .a(n8601), .b(n8598_1), .o(n8602_1) );
no02f01 g1873 ( .a(n8602_1), .b(n7012), .o(n8603) );
in01f01 g1874 ( .a(net_7042), .o(n8604) );
in01f01 g1875 ( .a(net_6978), .o(n8605) );
oa22f01 g1876 ( .a(n6987), .b(n8605), .c(n6985), .d(n8604), .o(n8606) );
in01f01 g1877 ( .a(net_7010), .o(n8607_1) );
in01f01 g1878 ( .a(net_7074), .o(n8608) );
oa22f01 g1879 ( .a(n6992), .b(n8607_1), .c(n6991), .d(n8608), .o(n8609) );
no02f01 g1880 ( .a(n8609), .b(n8606), .o(n8610) );
no02f01 g1881 ( .a(n8610), .b(n6997), .o(n8611) );
in01f01 g1882 ( .a(_net_6160), .o(n8612_1) );
in01f01 g1883 ( .a(net_6980), .o(n8613) );
in01f01 g1884 ( .a(net_7044), .o(n8614) );
oa22f01 g1885 ( .a(n6987), .b(n8613), .c(n6985), .d(n8614), .o(n8615) );
in01f01 g1886 ( .a(net_7076), .o(n8616_1) );
in01f01 g1887 ( .a(net_7012), .o(n8617) );
oa22f01 g1888 ( .a(n6992), .b(n8617), .c(n6991), .d(n8616_1), .o(n8618) );
no02f01 g1889 ( .a(n8618), .b(n8615), .o(n8619) );
oa22f01 g1890 ( .a(n8619), .b(n6980), .c(n6995_1), .d(n8612_1), .o(n8620) );
no03f01 g1891 ( .a(n8620), .b(n8611), .c(n8603), .o(n8621_1) );
in01f01 g1892 ( .a(net_7024), .o(n8622) );
in01f01 g1893 ( .a(net_6992), .o(n8623) );
oa22f01 g1894 ( .a(n8075_1), .b(n8623), .c(n8074), .d(n8622), .o(n8624) );
in01f01 g1895 ( .a(net_7056), .o(n8625_1) );
in01f01 g1896 ( .a(net_7088), .o(n8626) );
oa22f01 g1897 ( .a(n8080_1), .b(n8626), .c(n8079), .d(n8625_1), .o(n8627) );
no02f01 g1898 ( .a(n8627), .b(n8624), .o(n8628_1) );
na02f01 g1899 ( .a(n8628_1), .b(n8621_1), .o(n2534) );
in01f01 g1900 ( .a(_net_7445), .o(n8630) );
na02f01 g1901 ( .a(n6866), .b(net_7397), .o(n8631) );
ao22f01 g1902 ( .a(net_358), .b(_net_281), .c(_net_280), .d(net_360), .o(n8632_1) );
na02f01 g1903 ( .a(n8632_1), .b(n8631), .o(n8633) );
na02f01 g1904 ( .a(n8633), .b(n7197), .o(n8634) );
oa12f01 g1905 ( .a(n8634), .b(n7197), .c(n8630), .o(n2552) );
in01f01 g1906 ( .a(_net_7663), .o(n8636) );
na02f01 g1907 ( .a(n6965), .b(net_7551), .o(n8637_1) );
ao22f01 g1908 ( .a(_net_292), .b(net_381), .c(_net_291), .d(net_383), .o(n8638) );
na02f01 g1909 ( .a(n8638), .b(n8637_1), .o(n8639) );
na02f01 g1910 ( .a(n8639), .b(n7446_1), .o(n8640) );
oa12f01 g1911 ( .a(n8640), .b(n7446_1), .c(n8636), .o(n2566) );
ao22f01 g1912 ( .a(n6877), .b(_net_7270), .c(n6876_1), .d(net_7334), .o(n8642) );
ao22f01 g1913 ( .a(n6881_1), .b(net_7302), .c(n6880), .d(net_7366), .o(n8643) );
na02f01 g1914 ( .a(n8643), .b(n8642), .o(n2575) );
ao22f01 g1915 ( .a(n7225), .b(_net_7415), .c(n7224), .d(_net_7447), .o(n8645_1) );
ao22f01 g1916 ( .a(n7229), .b(_net_7511), .c(n7228), .d(_net_7479), .o(n8646) );
na02f01 g1917 ( .a(n8646), .b(n8645_1), .o(n2580) );
in01f01 g1918 ( .a(n7422_1), .o(n8648) );
no02f01 g1919 ( .a(n8648), .b(x868), .o(n2585) );
in01f01 g1920 ( .a(_net_5979), .o(n8650_1) );
no02f01 g1921 ( .a(n6976), .b(n8650_1), .o(n2590) );
no02f01 g1922 ( .a(n6963), .b(n6962), .o(n2632) );
ao22f01 g1923 ( .a(n6736_1), .b(net_7643), .c(n6734), .d(net_7611), .o(n8653) );
ao22f01 g1924 ( .a(n6739), .b(net_7675), .c(n6738), .d(_net_7579), .o(n8654_1) );
na02f01 g1925 ( .a(n8654_1), .b(n8653), .o(n2637) );
ao22f01 g1926 ( .a(n6877), .b(_net_7281), .c(n6876_1), .d(net_7345), .o(n8656) );
ao22f01 g1927 ( .a(n6881_1), .b(net_7313), .c(n6880), .d(net_7377), .o(n8657) );
na02f01 g1928 ( .a(n8657), .b(n8656), .o(n2651) );
in01f01 g1929 ( .a(net_6771), .o(n8659) );
in01f01 g1930 ( .a(net_6707), .o(n8660) );
oa22f01 g1931 ( .a(n7129), .b(n8660), .c(n7126), .d(n8659), .o(n8661) );
in01f01 g1932 ( .a(net_6803), .o(n8662_1) );
in01f01 g1933 ( .a(net_6739), .o(n8663) );
oa22f01 g1934 ( .a(n7134), .b(n8663), .c(n7132), .d(n8662_1), .o(n8664) );
no02f01 g1935 ( .a(n8664), .b(n8661), .o(n8665) );
no02f01 g1936 ( .a(n8665), .b(n7468_1), .o(n8666_1) );
in01f01 g1937 ( .a(net_6773), .o(n8667) );
in01f01 g1938 ( .a(net_6709), .o(n8668) );
oa22f01 g1939 ( .a(n7129), .b(n8668), .c(n7126), .d(n8667), .o(n8669) );
in01f01 g1940 ( .a(net_6741), .o(n8670) );
in01f01 g1941 ( .a(net_6805), .o(n8671_1) );
oa22f01 g1942 ( .a(n7134), .b(n8670), .c(n7132), .d(n8671_1), .o(n8672) );
no02f01 g1943 ( .a(n8672), .b(n8669), .o(n8673) );
no02f01 g1944 ( .a(n8673), .b(n7470), .o(n8674) );
in01f01 g1945 ( .a(_net_6121), .o(n8675) );
in01f01 g1946 ( .a(net_6711), .o(n8676_1) );
in01f01 g1947 ( .a(net_6775), .o(n8677) );
oa22f01 g1948 ( .a(n7129), .b(n8676_1), .c(n7126), .d(n8677), .o(n8678) );
in01f01 g1949 ( .a(net_6743), .o(n8679) );
in01f01 g1950 ( .a(net_6807), .o(n8680) );
oa22f01 g1951 ( .a(n7134), .b(n8679), .c(n7132), .d(n8680), .o(n8681_1) );
no02f01 g1952 ( .a(n8681_1), .b(n8678), .o(n8682) );
oa22f01 g1953 ( .a(n8682), .b(n7123), .c(n7118), .d(n8675), .o(n8683) );
no03f01 g1954 ( .a(n8683), .b(n8674), .c(n8666_1), .o(n8684) );
in01f01 g1955 ( .a(net_6723), .o(n8685_1) );
in01f01 g1956 ( .a(net_6755), .o(n8686) );
oa22f01 g1957 ( .a(n7492_1), .b(n8685_1), .c(n7491), .d(n8686), .o(n8687) );
in01f01 g1958 ( .a(net_6819), .o(n8688) );
in01f01 g1959 ( .a(net_6787), .o(n8689_1) );
oa22f01 g1960 ( .a(n7497), .b(n8688), .c(n7496_1), .d(n8689_1), .o(n8690) );
no02f01 g1961 ( .a(n8690), .b(n8687), .o(n8691) );
na02f01 g1962 ( .a(n8691), .b(n8684), .o(n2665) );
in01f01 g1963 ( .a(_net_6043), .o(n8693) );
no02f01 g1964 ( .a(n8693), .b(_net_6044), .o(n8694_1) );
in01f01 g1965 ( .a(_net_5980), .o(n8695) );
na02f01 g1966 ( .a(_net_6039), .b(_net_6045), .o(n8696) );
ao12f01 g1967 ( .a(n8696), .b(_net_5982), .c(n8695), .o(n8697) );
na02f01 g1968 ( .a(n8697), .b(n8694_1), .o(n8698_1) );
in01f01 g1969 ( .a(_net_6044), .o(n8699) );
in01f01 g1970 ( .a(n8696), .o(n8700) );
na03f01 g1971 ( .a(_net_5982), .b(_net_5981), .c(n8695), .o(n8701) );
na04f01 g1972 ( .a(n8701), .b(n8700), .c(n8693), .d(n8699), .o(n8702) );
oa12f01 g1973 ( .a(n8695), .b(_net_5982), .c(_net_5981), .o(n8703_1) );
na04f01 g1974 ( .a(n8703_1), .b(n8700), .c(n8693), .d(_net_6044), .o(n8704) );
no02f01 g1975 ( .a(n8693), .b(n8699), .o(n8705) );
na03f01 g1976 ( .a(n8705), .b(n8700), .c(_net_5980), .o(n8706) );
na04f01 g1977 ( .a(n8706), .b(n8704), .c(n8702), .d(n8698_1), .o(n8707) );
in01f01 g1978 ( .a(n8707), .o(n8708_1) );
no02f01 g1979 ( .a(n8708_1), .b(x906), .o(n2687) );
in01f01 g1980 ( .a(n7117), .o(n8710) );
na02f01 g1981 ( .a(n8710), .b(_net_6006), .o(n8711_1) );
na03f01 g1982 ( .a(n7467), .b(n8710), .c(_net_6822), .o(n8712) );
na02f01 g1983 ( .a(n7467), .b(n8710), .o(n8713) );
na02f01 g1984 ( .a(n8713), .b(n7466), .o(n8714) );
na02f01 g1985 ( .a(n8714), .b(n8712), .o(n8715_1) );
no02f01 g1986 ( .a(n8710), .b(n7121), .o(n8716) );
na02f01 g1987 ( .a(n8716), .b(_net_6822), .o(n8717) );
oa12f01 g1988 ( .a(n8717), .b(n8715_1), .c(n8711_1), .o(n2696) );
in01f01 g1989 ( .a(_net_126), .o(n8719) );
na02f01 g1990 ( .a(_net_154), .b(net_322), .o(n8720_1) );
oa12f01 g1991 ( .a(n8720_1), .b(_net_154), .c(n8719), .o(n2713) );
ao22f01 g1992 ( .a(n6736_1), .b(_net_7624), .c(n6734), .d(_net_7592), .o(n8722) );
ao22f01 g1993 ( .a(n6739), .b(_net_7656), .c(n6738), .d(_net_7560), .o(n8723) );
na02f01 g1994 ( .a(n8723), .b(n8722), .o(n2718) );
in01f01 g1995 ( .a(_net_280), .o(n8725_1) );
na02f01 g1996 ( .a(n7440), .b(_net_7803), .o(n8726) );
oa12f01 g1997 ( .a(n8726), .b(n7440), .c(n8725_1), .o(n2723) );
in01f01 g1998 ( .a(_net_7314), .o(n8728) );
na02f01 g1999 ( .a(n6898), .b(net_7234), .o(n8729) );
ao22f01 g2000 ( .a(net_328), .b(_net_269), .c(_net_270), .d(net_326), .o(n8730_1) );
na02f01 g2001 ( .a(n8730_1), .b(n8729), .o(n8731) );
na02f01 g2002 ( .a(n8731), .b(n7150), .o(n8732) );
oa12f01 g2003 ( .a(n8732), .b(n7150), .c(n8728), .o(n2732) );
ao22f01 g2004 ( .a(n6877), .b(_net_7257), .c(n6876_1), .d(_net_7321), .o(n8734_1) );
ao22f01 g2005 ( .a(n6881_1), .b(_net_7289), .c(n6880), .d(_net_7353), .o(n8735) );
na02f01 g2006 ( .a(n8735), .b(n8734_1), .o(n2753) );
no02f01 g2007 ( .a(n7813), .b(n6945), .o(n8737) );
no02f01 g2008 ( .a(n7822_1), .b(n6934_1), .o(n8738) );
in01f01 g2009 ( .a(_net_6097), .o(n8739_1) );
in01f01 g2010 ( .a(net_6636), .o(n8740) );
in01f01 g2011 ( .a(net_6572), .o(n8741) );
oa22f01 g2012 ( .a(n6922), .b(n8741), .c(n6919_1), .d(n8740), .o(n8742) );
in01f01 g2013 ( .a(net_6668), .o(n8743_1) );
in01f01 g2014 ( .a(net_6604), .o(n8744) );
oa22f01 g2015 ( .a(n6927), .b(n8744), .c(n6925), .d(n8743_1), .o(n8745) );
no02f01 g2016 ( .a(n8745), .b(n8742), .o(n8746) );
oa22f01 g2017 ( .a(n8746), .b(n6916), .c(n6932), .d(n8739_1), .o(n8747) );
no03f01 g2018 ( .a(n8747), .b(n8738), .c(n8737), .o(n8748_1) );
in01f01 g2019 ( .a(net_6616), .o(n8749) );
in01f01 g2020 ( .a(net_6584), .o(n8750) );
oa22f01 g2021 ( .a(n7058_1), .b(n8750), .c(n7057), .d(n8749), .o(n8751) );
in01f01 g2022 ( .a(net_6680), .o(n8752) );
in01f01 g2023 ( .a(net_6648), .o(n8753_1) );
oa22f01 g2024 ( .a(n7063), .b(n8752), .c(n7062_1), .d(n8753_1), .o(n8754) );
no02f01 g2025 ( .a(n8754), .b(n8751), .o(n8755) );
na02f01 g2026 ( .a(n8755), .b(n8748_1), .o(n2758) );
na02f01 g2027 ( .a(n7348), .b(_net_7822), .o(n8757_1) );
oa12f01 g2028 ( .a(n8757_1), .b(n7348), .c(n7689), .o(n2771) );
no02f01 g2029 ( .a(_net_7097), .b(n6986_1), .o(n8759) );
in01f01 g2030 ( .a(_net_7097), .o(n8760) );
no02f01 g2031 ( .a(n8760), .b(_net_7094), .o(n8761) );
no02f01 g2032 ( .a(n8761), .b(n8759), .o(n8762_1) );
no02f01 g2033 ( .a(net_7096), .b(n6984), .o(n8763) );
no02f01 g2034 ( .a(n8763), .b(n8762_1), .o(n8764) );
no04f01 g2035 ( .a(n8761), .b(n8759), .c(net_7096), .d(n6984), .o(n8765) );
oa12f01 g2036 ( .a(n8388), .b(n8765), .c(n8764), .o(n8766) );
no02f01 g2037 ( .a(n8765), .b(n8764), .o(n8767_1) );
na02f01 g2038 ( .a(n8767_1), .b(n2270), .o(n8768) );
na02f01 g2039 ( .a(n8768), .b(n8766), .o(n2776) );
ao22f01 g2040 ( .a(n6738), .b(_net_7554), .c(n6736_1), .d(_net_7618), .o(n8770) );
ao22f01 g2041 ( .a(n6739), .b(_net_7650), .c(n6734), .d(_net_7586), .o(n8771_1) );
na02f01 g2042 ( .a(n8771_1), .b(n8770), .o(n2797) );
ao22f01 g2043 ( .a(n7225), .b(_net_7422), .c(n7224), .d(net_7454), .o(n8773) );
ao22f01 g2044 ( .a(n7229), .b(net_7518), .c(n7228), .d(net_7486), .o(n8774) );
na02f01 g2045 ( .a(n8774), .b(n8773), .o(n2810) );
in01f01 g2046 ( .a(net_7036), .o(n8776) );
in01f01 g2047 ( .a(net_6972), .o(n8777) );
oa22f01 g2048 ( .a(n6987), .b(n8777), .c(n6985), .d(n8776), .o(n8778) );
in01f01 g2049 ( .a(net_7004), .o(n8779) );
in01f01 g2050 ( .a(net_7068), .o(n8780_1) );
oa22f01 g2051 ( .a(n6992), .b(n8779), .c(n6991), .d(n8780_1), .o(n8781) );
no02f01 g2052 ( .a(n8781), .b(n8778), .o(n8782) );
no02f01 g2053 ( .a(n8782), .b(n7012), .o(n8783) );
in01f01 g2054 ( .a(net_6974), .o(n8784_1) );
in01f01 g2055 ( .a(net_7038), .o(n8785) );
oa22f01 g2056 ( .a(n6987), .b(n8784_1), .c(n6985), .d(n8785), .o(n8786) );
in01f01 g2057 ( .a(net_7070), .o(n8787) );
in01f01 g2058 ( .a(net_7006), .o(n8788_1) );
oa22f01 g2059 ( .a(n6992), .b(n8788_1), .c(n6991), .d(n8787), .o(n8789) );
no02f01 g2060 ( .a(n8789), .b(n8786), .o(n8790) );
no02f01 g2061 ( .a(n8790), .b(n6997), .o(n8791) );
in01f01 g2062 ( .a(_net_6156), .o(n8792) );
oa22f01 g2063 ( .a(n8602_1), .b(n6980), .c(n6995_1), .d(n8792), .o(n8793_1) );
no03f01 g2064 ( .a(n8793_1), .b(n8791), .c(n8783), .o(n8794) );
in01f01 g2065 ( .a(net_6988), .o(n8795) );
in01f01 g2066 ( .a(net_7020), .o(n8796) );
oa22f01 g2067 ( .a(n8075_1), .b(n8795), .c(n8074), .d(n8796), .o(n8797_1) );
in01f01 g2068 ( .a(net_7052), .o(n8798) );
in01f01 g2069 ( .a(net_7084), .o(n8799) );
oa22f01 g2070 ( .a(n8080_1), .b(n8799), .c(n8079), .d(n8798), .o(n8800_1) );
no02f01 g2071 ( .a(n8800_1), .b(n8797_1), .o(n8801) );
na02f01 g2072 ( .a(n8801), .b(n8794), .o(n2831) );
in01f01 g2073 ( .a(_net_7794), .o(n8803) );
na02f01 g2074 ( .a(n6803), .b(_net_6029), .o(n8804) );
oa12f01 g2075 ( .a(n8804), .b(n6803), .c(n8803), .o(n2836) );
in01f01 g2076 ( .a(_net_7261), .o(n8806) );
na02f01 g2077 ( .a(n6898), .b(net_7245), .o(n8807) );
ao22f01 g2078 ( .a(_net_269), .b(net_339), .c(_net_270), .d(net_337), .o(n8808) );
na02f01 g2079 ( .a(n8808), .b(n8807), .o(n8809_1) );
na02f01 g2080 ( .a(n8809_1), .b(n6901), .o(n8810) );
oa12f01 g2081 ( .a(n8810), .b(n6901), .c(n8806), .o(n2845) );
in01f01 g2082 ( .a(net_376), .o(n8812) );
no02f01 g2083 ( .a(n6966), .b(n8812), .o(n2850) );
in01f01 g2084 ( .a(_net_7501), .o(n8814) );
na02f01 g2085 ( .a(n6866), .b(net_7389), .o(n8815) );
ao22f01 g2086 ( .a(net_350), .b(_net_281), .c(_net_280), .d(net_352), .o(n8816) );
na02f01 g2087 ( .a(n8816), .b(n8815), .o(n8817) );
na02f01 g2088 ( .a(n8817), .b(n7626_1), .o(n8818_1) );
oa12f01 g2089 ( .a(n8818_1), .b(n7626_1), .c(n8814), .o(n2855) );
in01f01 g2090 ( .a(_net_7572), .o(n8820) );
na02f01 g2091 ( .a(n7519), .b(n615), .o(n8821) );
oa12f01 g2092 ( .a(n8821), .b(n7519), .c(n8820), .o(n2890) );
in01f01 g2093 ( .a(net_5992), .o(n8823_1) );
in01f01 g2094 ( .a(_net_7722), .o(n8824) );
ao12f01 g2095 ( .a(n7343), .b(n8824), .c(n8823_1), .o(n2900) );
in01f01 g2096 ( .a(net_336), .o(n8826_1) );
no02f01 g2097 ( .a(n6899_1), .b(n8826_1), .o(n2913) );
na02f01 g2098 ( .a(n7298), .b(net_7742), .o(n8828) );
ao22f01 g2099 ( .a(n7306), .b(_net_6012), .c(n7291), .d(net_7713), .o(n8829) );
na02f01 g2100 ( .a(n7302_1), .b(net_152), .o(n8830) );
na02f01 g2101 ( .a(n7296), .b(net_252), .o(n8831_1) );
na03f01 g2102 ( .a(n7308), .b(_net_178), .c(n6800), .o(n8832) );
na03f01 g2103 ( .a(n7308), .b(_net_215), .c(x1322), .o(n8833) );
na03f01 g2104 ( .a(n8833), .b(n8832), .c(n8831_1), .o(n8834) );
ao12f01 g2105 ( .a(n8834), .b(n7286), .c(_net_295), .o(n8835_1) );
na04f01 g2106 ( .a(n8835_1), .b(n8830), .c(n8829), .d(n8828), .o(n2918) );
in01f01 g2107 ( .a(_net_6220), .o(n8837) );
no02f01 g2108 ( .a(_net_392), .b(n8837), .o(n2930) );
in01f01 g2109 ( .a(_net_7552), .o(n8839) );
na02f01 g2110 ( .a(n6965), .b(net_7536), .o(n8840_1) );
ao22f01 g2111 ( .a(net_366), .b(_net_292), .c(net_368), .d(_net_291), .o(n8841) );
na02f01 g2112 ( .a(n8841), .b(n8840_1), .o(n8842) );
na02f01 g2113 ( .a(n8842), .b(n7519), .o(n8843) );
oa12f01 g2114 ( .a(n8843), .b(n7519), .c(n8839), .o(n2953) );
in01f01 g2115 ( .a(net_358), .o(n8845_1) );
no02f01 g2116 ( .a(n6867_1), .b(n8845_1), .o(n2958) );
no02f01 g2117 ( .a(net_7680), .b(n6959), .o(n8847) );
in01f01 g2118 ( .a(n8847), .o(n8848) );
no02f01 g2119 ( .a(n8848), .b(n8360), .o(n8849) );
no02f01 g2120 ( .a(n8847), .b(n8361), .o(n8850_1) );
oa12f01 g2121 ( .a(n8356), .b(n8850_1), .c(n8849), .o(n8851) );
no02f01 g2122 ( .a(n8850_1), .b(n8849), .o(n8852) );
na02f01 g2123 ( .a(n8852), .b(n4405), .o(n8853) );
na02f01 g2124 ( .a(n8853), .b(n8851), .o(n2976) );
in01f01 g2125 ( .a(n6761_1), .o(n8855_1) );
na02f01 g2126 ( .a(n6763), .b(n8855_1), .o(n8856) );
in01f01 g2127 ( .a(n8856), .o(n8857) );
na02f01 g2128 ( .a(n8855_1), .b(_net_5984), .o(n8858) );
no02f01 g2129 ( .a(n8858), .b(n8857), .o(n8859) );
na02f01 g2130 ( .a(n8859), .b(n6747), .o(n8860_1) );
no02f01 g2131 ( .a(n8858), .b(n8856), .o(n8861) );
no02f01 g2132 ( .a(n8855_1), .b(n6759), .o(n8862) );
ao22f01 g2133 ( .a(n8862), .b(_net_6553), .c(n8861), .d(n7760_1), .o(n8863) );
na02f01 g2134 ( .a(n8863), .b(n8860_1), .o(n2981) );
oa12f01 g2135 ( .a(n6886_1), .b(_net_7791), .c(n7165), .o(n2986) );
in01f01 g2136 ( .a(_net_7531), .o(n8866) );
no02f01 g2137 ( .a(n7229), .b(n8866), .o(n8867) );
no03f01 g2138 ( .a(n7227), .b(n7223), .c(_net_7531), .o(n8868) );
no02f01 g2139 ( .a(n8868), .b(n8867), .o(n8869_1) );
in01f01 g2140 ( .a(_net_227), .o(n8870) );
no02f01 g2141 ( .a(n7850), .b(n8870), .o(n5792) );
in01f01 g2142 ( .a(n5792), .o(n8872) );
na02f01 g2143 ( .a(_net_278), .b(n8870), .o(n8873_1) );
oa22f01 g2144 ( .a(n8873_1), .b(n8866), .c(n8872), .d(n8869_1), .o(n2991) );
in01f01 g2145 ( .a(_net_6038), .o(n8875) );
ao12f01 g2146 ( .a(n8650_1), .b(_net_7098), .c(_net_7095), .o(n8876) );
oa12f01 g2147 ( .a(n8876), .b(_net_7098), .c(_net_7095), .o(n8877_1) );
na02f01 g2148 ( .a(n8762_1), .b(n2270), .o(n8878) );
oa12f01 g2149 ( .a(n8875), .b(n8878), .c(n8877_1), .o(n3000) );
in01f01 g2150 ( .a(net_6629), .o(n8880) );
in01f01 g2151 ( .a(net_6565), .o(n8881) );
oa22f01 g2152 ( .a(n6922), .b(n8881), .c(n6919_1), .d(n8880), .o(n8882_1) );
in01f01 g2153 ( .a(net_6661), .o(n8883) );
in01f01 g2154 ( .a(net_6597), .o(n8884) );
oa22f01 g2155 ( .a(n6927), .b(n8884), .c(n6925), .d(n8883), .o(n8885) );
oa12f01 g2156 ( .a(n6917), .b(n8885), .c(n8882_1), .o(n8886_1) );
ao22f01 g2157 ( .a(n6935), .b(n6930), .c(n6933), .d(_net_6090), .o(n8887) );
in01f01 g2158 ( .a(net_6641), .o(n8888) );
in01f01 g2159 ( .a(net_6577), .o(n8889) );
oa22f01 g2160 ( .a(n6922), .b(n8889), .c(n6919_1), .d(n8888), .o(n8890) );
in01f01 g2161 ( .a(net_6609), .o(n8891_1) );
in01f01 g2162 ( .a(net_6673), .o(n8892) );
oa22f01 g2163 ( .a(n6927), .b(n8891_1), .c(n6925), .d(n8892), .o(n8893) );
no02f01 g2164 ( .a(n8893), .b(n8890), .o(n8894) );
no03f01 g2165 ( .a(n8894), .b(n6947_1), .c(n6943_1), .o(n8895_1) );
ao12f01 g2166 ( .a(n8895_1), .b(n6946), .c(n6938_1), .o(n8896) );
na03f01 g2167 ( .a(n8896), .b(n8887), .c(n8886_1), .o(n3005) );
no02f01 g2168 ( .a(n7232), .b(n7163), .o(n3010) );
in01f01 g2169 ( .a(net_379), .o(n8899_1) );
no02f01 g2170 ( .a(n6966), .b(n8899_1), .o(n3015) );
in01f01 g2171 ( .a(_net_7320), .o(n8901) );
na02f01 g2172 ( .a(n8208), .b(n7150), .o(n8902) );
oa12f01 g2173 ( .a(n8902), .b(n7150), .c(n8901), .o(n3020) );
ao22f01 g2174 ( .a(n6877), .b(_net_7267), .c(n6876_1), .d(_net_7331), .o(n8904) );
ao22f01 g2175 ( .a(n6881_1), .b(_net_7299), .c(n6880), .d(_net_7363), .o(n8905) );
na02f01 g2176 ( .a(n8905), .b(n8904), .o(n3025) );
in01f01 g2177 ( .a(_net_6023), .o(n8907) );
na02f01 g2178 ( .a(n7348), .b(_net_7823), .o(n8908_1) );
oa12f01 g2179 ( .a(n8908_1), .b(n7348), .c(n8907), .o(n3042) );
in01f01 g2180 ( .a(_net_7667), .o(n8910) );
na02f01 g2181 ( .a(n7446_1), .b(n7144), .o(n8911) );
oa12f01 g2182 ( .a(n8911), .b(n7446_1), .c(n8910), .o(n3047) );
no02f01 g2183 ( .a(n8866), .b(n7867_1), .o(n8913) );
no02f01 g2184 ( .a(_net_7531), .b(_net_7535), .o(n8914) );
no02f01 g2185 ( .a(n8914), .b(n8913), .o(n8915) );
in01f01 g2186 ( .a(n8915), .o(n8916) );
no02f01 g2187 ( .a(n7194_1), .b(n7223), .o(n8917_1) );
no02f01 g2188 ( .a(_net_7533), .b(net_7529), .o(n8918) );
no02f01 g2189 ( .a(n8918), .b(n8917_1), .o(n8919) );
in01f01 g2190 ( .a(n8919), .o(n8850) );
no02f01 g2191 ( .a(n7227), .b(n6860_1), .o(n8921) );
no02f01 g2192 ( .a(_net_7530), .b(_net_7534), .o(n8922_1) );
no02f01 g2193 ( .a(n8922_1), .b(n8921), .o(n8923) );
in01f01 g2194 ( .a(n8923), .o(n8924) );
na02f01 g2195 ( .a(n8924), .b(n8850), .o(n8925) );
no02f01 g2196 ( .a(n8925), .b(n8916), .o(n3056) );
ao22f01 g2197 ( .a(n6877), .b(_net_7278), .c(n6876_1), .d(net_7342), .o(n8927) );
ao22f01 g2198 ( .a(n6881_1), .b(net_7310), .c(n6880), .d(net_7374), .o(n8928) );
na02f01 g2199 ( .a(n8928), .b(n8927), .o(n3065) );
ao22f01 g2200 ( .a(n6738), .b(_net_7555), .c(n6736_1), .d(_net_7619), .o(n8930) );
ao22f01 g2201 ( .a(n6739), .b(_net_7651), .c(n6734), .d(_net_7587), .o(n8931_1) );
na02f01 g2202 ( .a(n8931_1), .b(n8930), .o(n3078) );
na02f01 g2203 ( .a(n8127), .b(n6918), .o(n8933) );
na02f01 g2204 ( .a(n6943_1), .b(_net_6688), .o(n8934_1) );
na02f01 g2205 ( .a(_net_6687), .b(n6918), .o(n8935) );
na02f01 g2206 ( .a(n8935), .b(n8934_1), .o(n8936) );
ao22f01 g2207 ( .a(n8936), .b(n8125_1), .c(n8132), .d(_net_6688), .o(n8937) );
na02f01 g2208 ( .a(n8937), .b(n8933), .o(n3087) );
in01f01 g2209 ( .a(_net_6280), .o(n8939_1) );
no02f01 g2210 ( .a(n8939_1), .b(_net_392), .o(n3092) );
in01f01 g2211 ( .a(_net_128), .o(n8941) );
na02f01 g2212 ( .a(net_324), .b(_net_154), .o(n8942) );
oa12f01 g2213 ( .a(n8942), .b(_net_154), .c(n8941), .o(n3097) );
in01f01 g2214 ( .a(_net_7410), .o(n8944) );
na02f01 g2215 ( .a(n7550), .b(n6891), .o(n8945) );
oa12f01 g2216 ( .a(n8945), .b(n7550), .c(n8944), .o(n3130) );
in01f01 g2217 ( .a(_net_7557), .o(n8947) );
na02f01 g2218 ( .a(n7519), .b(n7449), .o(n8948_1) );
oa12f01 g2219 ( .a(n8948_1), .b(n7519), .c(n8947), .o(n3139) );
in01f01 g2220 ( .a(_net_7449), .o(n8950) );
na02f01 g2221 ( .a(n7197), .b(n6872_1), .o(n8951) );
oa12f01 g2222 ( .a(n8951), .b(n7197), .c(n8950), .o(n3148) );
no03f01 g2223 ( .a(n7336), .b(n7109), .c(n7105), .o(n3157) );
in01f01 g2224 ( .a(_net_7470), .o(n8954) );
na02f01 g2225 ( .a(n7860), .b(n6869), .o(n8955) );
oa12f01 g2226 ( .a(n8955), .b(n6869), .c(n8954), .o(n3170) );
in01f01 g2227 ( .a(_net_7350), .o(n8957) );
na02f01 g2228 ( .a(n6898), .b(net_7238), .o(n8958_1) );
ao22f01 g2229 ( .a(net_332), .b(_net_269), .c(net_330), .d(_net_270), .o(n8959) );
na02f01 g2230 ( .a(n8959), .b(n8958_1), .o(n8960) );
na02f01 g2231 ( .a(n8960), .b(n7030), .o(n8961) );
oa12f01 g2232 ( .a(n8961), .b(n7030), .c(n8957), .o(n3182) );
in01f01 g2233 ( .a(_net_7277), .o(n8963_1) );
in01f01 g2234 ( .a(net_341), .o(n8964) );
no02f01 g2235 ( .a(n6899_1), .b(n8964), .o(n6376) );
na02f01 g2236 ( .a(n6376), .b(n6901), .o(n8966) );
oa12f01 g2237 ( .a(n8966), .b(n6901), .c(n8963_1), .o(n3194) );
ao22f01 g2238 ( .a(n6877), .b(_net_7272), .c(n6876_1), .d(net_7336), .o(n8968) );
ao22f01 g2239 ( .a(n6881_1), .b(net_7304), .c(n6880), .d(net_7368), .o(n8969) );
na02f01 g2240 ( .a(n8969), .b(n8968), .o(n3203) );
in01f01 g2241 ( .a(_net_7326), .o(n8971_1) );
na02f01 g2242 ( .a(n7926), .b(n7150), .o(n8972) );
oa12f01 g2243 ( .a(n8972), .b(n7150), .c(n8971_1), .o(n3212) );
in01f01 g2244 ( .a(net_6764), .o(n8974) );
in01f01 g2245 ( .a(net_6700), .o(n8975) );
oa22f01 g2246 ( .a(n7129), .b(n8975), .c(n7126), .d(n8974), .o(n8976_1) );
in01f01 g2247 ( .a(net_6732), .o(n8977) );
in01f01 g2248 ( .a(net_6796), .o(n8978) );
oa22f01 g2249 ( .a(n7134), .b(n8977), .c(n7132), .d(n8978), .o(n8979) );
oa12f01 g2250 ( .a(n7124), .b(n8979), .c(n8976_1), .o(n8980) );
ao22f01 g2251 ( .a(n8157), .b(n8159), .c(n7119), .d(_net_6110), .o(n8981_1) );
na02f01 g2252 ( .a(n8162), .b(n8164), .o(n8982) );
in01f01 g2253 ( .a(net_6776), .o(n8983) );
in01f01 g2254 ( .a(net_6712), .o(n8984) );
oa22f01 g2255 ( .a(n7129), .b(n8984), .c(n7126), .d(n8983), .o(n8985) );
in01f01 g2256 ( .a(net_6808), .o(n8986_1) );
in01f01 g2257 ( .a(net_6744), .o(n8987) );
oa22f01 g2258 ( .a(n7134), .b(n8987), .c(n7132), .d(n8986_1), .o(n8988) );
oa12f01 g2259 ( .a(n8167), .b(n8988), .c(n8985), .o(n8989) );
na04f01 g2260 ( .a(n8989), .b(n8982), .c(n8981_1), .d(n8980), .o(n3217) );
in01f01 g2261 ( .a(_net_7478), .o(n8991) );
na02f01 g2262 ( .a(n6866), .b(net_7398), .o(n8992) );
ao22f01 g2263 ( .a(net_359), .b(_net_281), .c(_net_280), .d(net_361), .o(n8993) );
na02f01 g2264 ( .a(n8993), .b(n8992), .o(n8994) );
na02f01 g2265 ( .a(n8994), .b(n6869), .o(n8995_1) );
oa12f01 g2266 ( .a(n8995_1), .b(n6869), .c(n8991), .o(n3222) );
in01f01 g2267 ( .a(net_7770), .o(n8997) );
no03f01 g2268 ( .a(n7232), .b(n8997), .c(net_7771), .o(n3231) );
in01f01 g2269 ( .a(net_7106), .o(n8999) );
in01f01 g2270 ( .a(net_7170), .o(n9000_1) );
oa22f01 g2271 ( .a(n7580), .b(n8999), .c(n7577_1), .d(n9000_1), .o(n9001) );
in01f01 g2272 ( .a(net_7202), .o(n9002) );
in01f01 g2273 ( .a(net_7138), .o(n9003) );
oa22f01 g2274 ( .a(n7585), .b(n9003), .c(n7583), .d(n9002), .o(n9004) );
no02f01 g2275 ( .a(n9004), .b(n9001), .o(n9005_1) );
no02f01 g2276 ( .a(n9005_1), .b(n7721), .o(n9006) );
no02f01 g2277 ( .a(n8274), .b(n7592), .o(n9007) );
in01f01 g2278 ( .a(_net_6175), .o(n9008) );
oa22f01 g2279 ( .a(n8282), .b(n7574), .c(n7590), .d(n9008), .o(n9009) );
no03f01 g2280 ( .a(n9009), .b(n9007), .c(n9006), .o(n9010_1) );
in01f01 g2281 ( .a(net_7154), .o(n9011) );
in01f01 g2282 ( .a(net_7122), .o(n9012) );
oa22f01 g2283 ( .a(n7740), .b(n9012), .c(n7739), .d(n9011), .o(n9013) );
in01f01 g2284 ( .a(net_7186), .o(n9014_1) );
in01f01 g2285 ( .a(net_7218), .o(n9015) );
oa22f01 g2286 ( .a(n7745), .b(n9015), .c(n7744), .d(n9014_1), .o(n9016) );
no02f01 g2287 ( .a(n9016), .b(n9013), .o(n9017_1) );
na02f01 g2288 ( .a(n9017_1), .b(n9010_1), .o(n3240) );
in01f01 g2289 ( .a(_net_272), .o(n9019) );
na02f01 g2290 ( .a(n7440), .b(_net_7798), .o(n9020) );
oa12f01 g2291 ( .a(n9020), .b(n7440), .c(n9019), .o(n3254) );
in01f01 g2292 ( .a(_net_116), .o(n9022_1) );
na02f01 g2293 ( .a(net_312), .b(_net_154), .o(n9023) );
oa12f01 g2294 ( .a(n9023), .b(n9022_1), .c(_net_154), .o(n3263) );
no02f01 g2295 ( .a(n7050), .b(n6945), .o(n9025_1) );
no02f01 g2296 ( .a(n6954), .b(n6934_1), .o(n9026) );
in01f01 g2297 ( .a(_net_6102), .o(n9027) );
oa22f01 g2298 ( .a(n8894), .b(n6916), .c(n6932), .d(n9027), .o(n9028) );
no03f01 g2299 ( .a(n9028), .b(n9026), .c(n9025_1), .o(n9029) );
in01f01 g2300 ( .a(net_6589), .o(n9030_1) );
in01f01 g2301 ( .a(net_6621), .o(n9031) );
oa22f01 g2302 ( .a(n7058_1), .b(n9030_1), .c(n7057), .d(n9031), .o(n9032) );
in01f01 g2303 ( .a(net_6653), .o(n9033) );
in01f01 g2304 ( .a(net_6685), .o(n9034_1) );
oa22f01 g2305 ( .a(n7063), .b(n9034_1), .c(n7062_1), .d(n9033), .o(n9035) );
no02f01 g2306 ( .a(n9035), .b(n9032), .o(n9036) );
na02f01 g2307 ( .a(n9036), .b(n9029), .o(n3268) );
in01f01 g2308 ( .a(_net_6203), .o(n9038) );
no02f01 g2309 ( .a(n9038), .b(_net_392), .o(n3285) );
no02f01 g2310 ( .a(n7094), .b(n6764), .o(n9040) );
in01f01 g2311 ( .a(net_6505), .o(n9041) );
in01f01 g2312 ( .a(net_6441), .o(n9042_1) );
oa22f01 g2313 ( .a(n6750), .b(n9042_1), .c(n6748), .d(n9041), .o(n9043) );
in01f01 g2314 ( .a(net_6537), .o(n9044) );
in01f01 g2315 ( .a(net_6473), .o(n9045) );
oa22f01 g2316 ( .a(n6755), .b(n9045), .c(n6754), .d(n9044), .o(n9046) );
no02f01 g2317 ( .a(n9046), .b(n9043), .o(n9047_1) );
no02f01 g2318 ( .a(n9047_1), .b(n6766), .o(n9048) );
ao22f01 g2319 ( .a(n6777), .b(net_6443), .c(n6776), .d(net_6507), .o(n9049) );
ao22f01 g2320 ( .a(n6780), .b(net_6475), .c(n6779_1), .d(net_6539), .o(n9050) );
ao12f01 g2321 ( .a(n6775), .b(n9050), .c(n9049), .o(n9051) );
in01f01 g2322 ( .a(_net_6083), .o(n9052_1) );
no02f01 g2323 ( .a(n6784), .b(n9052_1), .o(n9053) );
no04f01 g2324 ( .a(n9053), .b(n9051), .c(n9048), .d(n9040), .o(n9054) );
in01f01 g2325 ( .a(net_6487), .o(n9055) );
in01f01 g2326 ( .a(net_6455), .o(n9056) );
oa22f01 g2327 ( .a(n6790), .b(n9056), .c(n6789), .d(n9055), .o(n9057_1) );
in01f01 g2328 ( .a(net_6551), .o(n9058) );
in01f01 g2329 ( .a(net_6519), .o(n9059) );
oa22f01 g2330 ( .a(n6795), .b(n9058), .c(n6794), .d(n9059), .o(n9060_1) );
no02f01 g2331 ( .a(n9060_1), .b(n9057_1), .o(n9061) );
na02f01 g2332 ( .a(n9061), .b(n9054), .o(n3294) );
in01f01 g2333 ( .a(_net_7266), .o(n9063) );
na02f01 g2334 ( .a(n7242), .b(n6901), .o(n9064) );
oa12f01 g2335 ( .a(n9064), .b(n6901), .c(n9063), .o(n3308) );
oa12f01 g2336 ( .a(n7575), .b(n9004), .c(n9001), .o(n9066) );
ao22f01 g2337 ( .a(n8499_1), .b(n7593), .c(n7591_1), .d(_net_6171), .o(n9067) );
na02f01 g2338 ( .a(n7914), .b(n7588), .o(n9068) );
in01f01 g2339 ( .a(net_7182), .o(n9069_1) );
in01f01 g2340 ( .a(net_7118), .o(n9070) );
oa22f01 g2341 ( .a(n7580), .b(n9070), .c(n7577_1), .d(n9069_1), .o(n9071) );
in01f01 g2342 ( .a(net_7150), .o(n9072) );
in01f01 g2343 ( .a(net_7214), .o(n9073) );
oa22f01 g2344 ( .a(n7585), .b(n9072), .c(n7583), .d(n9073), .o(n9074_1) );
oa12f01 g2345 ( .a(n7920_1), .b(n9074_1), .c(n9071), .o(n9075) );
na04f01 g2346 ( .a(n9075), .b(n9068), .c(n9067), .d(n9066), .o(n3313) );
ao22f01 g2347 ( .a(n7288_1), .b(net_6046), .c(n7286), .d(net_285), .o(n9077) );
ao22f01 g2348 ( .a(n7298), .b(_net_7735), .c(n7291), .d(_net_7706), .o(n9078) );
na02f01 g2349 ( .a(n7302_1), .b(_net_129), .o(n9079_1) );
na03f01 g2350 ( .a(n7308), .b(net_208), .c(x1322), .o(n9080) );
na02f01 g2351 ( .a(n7296), .b(net_245), .o(n9081) );
na03f01 g2352 ( .a(n7308), .b(net_171), .c(n6800), .o(n9082_1) );
na03f01 g2353 ( .a(n9082_1), .b(n9081), .c(n9080), .o(n9083) );
ao12f01 g2354 ( .a(n9083), .b(n7306), .c(_net_6002), .o(n9084) );
na04f01 g2355 ( .a(n9084), .b(n9079_1), .c(n9078), .d(n9077), .o(n3322) );
in01f01 g2356 ( .a(_net_7803), .o(n9086_1) );
na02f01 g2357 ( .a(n6803), .b(_net_6041), .o(n9087) );
oa12f01 g2358 ( .a(n9087), .b(n6803), .c(n9086_1), .o(n3338) );
ao22f01 g2359 ( .a(n7288_1), .b(_net_6040), .c(n7286), .d(_net_279), .o(n9089) );
ao22f01 g2360 ( .a(n7298), .b(_net_7729), .c(n7291), .d(_net_7700), .o(n9090) );
na02f01 g2361 ( .a(n7302_1), .b(_net_123), .o(n9091_1) );
na03f01 g2362 ( .a(n7308), .b(net_202), .c(x1322), .o(n9092) );
na02f01 g2363 ( .a(n7296), .b(net_239), .o(n9093) );
na03f01 g2364 ( .a(n7308), .b(net_165), .c(n6800), .o(n9094) );
na03f01 g2365 ( .a(n9094), .b(n9093), .c(n9092), .o(n9095) );
ao12f01 g2366 ( .a(n9095), .b(n7306), .c(_net_5996), .o(n9096_1) );
na04f01 g2367 ( .a(n9096_1), .b(n9091_1), .c(n9090), .d(n9089), .o(n3352) );
in01f01 g2368 ( .a(_net_7583), .o(n9098) );
no02f01 g2369 ( .a(n6966), .b(n7142_1), .o(n5628) );
na02f01 g2370 ( .a(n5628), .b(n7519), .o(n9100) );
oa12f01 g2371 ( .a(n9100), .b(n7519), .c(n9098), .o(n3356) );
in01f01 g2372 ( .a(_net_7230), .o(n9102) );
na03f01 g2373 ( .a(n8302), .b(n9102), .c(_net_7229), .o(n9103) );
oa12f01 g2374 ( .a(_net_7230), .b(n8304), .c(n7579), .o(n9104) );
na02f01 g2375 ( .a(n9104), .b(n9103), .o(n9105) );
na02f01 g2376 ( .a(n9105), .b(_net_7233), .o(n9106_1) );
in01f01 g2377 ( .a(_net_7233), .o(n9107) );
na03f01 g2378 ( .a(n9104), .b(n9103), .c(n9107), .o(n9108) );
na02f01 g2379 ( .a(_net_7228), .b(n7719_1), .o(n9109) );
na02f01 g2380 ( .a(n7576), .b(_net_7227), .o(n9110_1) );
na02f01 g2381 ( .a(n9110_1), .b(n9109), .o(n9111) );
na02f01 g2382 ( .a(n9111), .b(net_7231), .o(n9112) );
in01f01 g2383 ( .a(net_7231), .o(n9113) );
na03f01 g2384 ( .a(n9110_1), .b(n9109), .c(n9113), .o(n9114) );
ao22f01 g2385 ( .a(n9114), .b(n9112), .c(n7720), .d(_net_7227), .o(n9115_1) );
in01f01 g2386 ( .a(_net_7232), .o(n9116) );
na02f01 g2387 ( .a(n8306), .b(n9116), .o(n9117) );
na03f01 g2388 ( .a(n8305), .b(n8303_1), .c(_net_7232), .o(n9118) );
na03f01 g2389 ( .a(n9118), .b(n9117), .c(n9115_1), .o(n9119) );
ao12f01 g2390 ( .a(n9119), .b(n9108), .c(n9106_1), .o(n3370) );
in01f01 g2391 ( .a(net_6907), .o(n9121) );
in01f01 g2392 ( .a(net_6843), .o(n9122) );
oa22f01 g2393 ( .a(n6810), .b(n9122), .c(n6807), .d(n9121), .o(n9123) );
in01f01 g2394 ( .a(net_6939), .o(n9124_1) );
in01f01 g2395 ( .a(net_6875), .o(n9125) );
oa22f01 g2396 ( .a(n6815), .b(n9125), .c(n6813_1), .d(n9124_1), .o(n9126) );
no02f01 g2397 ( .a(n9126), .b(n9123), .o(n9127) );
no02f01 g2398 ( .a(n9127), .b(n6824), .o(n9128) );
in01f01 g2399 ( .a(net_6845), .o(n9129_1) );
in01f01 g2400 ( .a(net_6909), .o(n9130) );
oa22f01 g2401 ( .a(n6810), .b(n9129_1), .c(n6807), .d(n9130), .o(n9131) );
in01f01 g2402 ( .a(net_6877), .o(n9132) );
in01f01 g2403 ( .a(net_6941), .o(n9133) );
oa22f01 g2404 ( .a(n6815), .b(n9132), .c(n6813_1), .d(n9133), .o(n9134_1) );
no02f01 g2405 ( .a(n9134_1), .b(n9131), .o(n9135) );
no02f01 g2406 ( .a(n9135), .b(n6826_1), .o(n9136) );
ao22f01 g2407 ( .a(n6811), .b(net_6847), .c(n6808), .d(net_6911), .o(n9137) );
ao22f01 g2408 ( .a(n6816), .b(net_6879), .c(n6814), .d(net_6943), .o(n9138_1) );
ao12f01 g2409 ( .a(n6836_1), .b(n9138_1), .c(n9137), .o(n9139) );
in01f01 g2410 ( .a(_net_6142), .o(n9140) );
no02f01 g2411 ( .a(n6844), .b(n9140), .o(n9141) );
no04f01 g2412 ( .a(n9141), .b(n9139), .c(n9136), .d(n9128), .o(n9142) );
in01f01 g2413 ( .a(net_6859), .o(n9143_1) );
in01f01 g2414 ( .a(net_6891), .o(n9144) );
oa22f01 g2415 ( .a(n6850_1), .b(n9143_1), .c(n6849), .d(n9144), .o(n9145) );
in01f01 g2416 ( .a(net_6955), .o(n9146_1) );
in01f01 g2417 ( .a(net_6923), .o(n9147) );
oa22f01 g2418 ( .a(n6855_1), .b(n9146_1), .c(n6854), .d(n9147), .o(n9148) );
no02f01 g2419 ( .a(n9148), .b(n9145), .o(n9149) );
na02f01 g2420 ( .a(n9149), .b(n9142), .o(n3395) );
in01f01 g2421 ( .a(_net_7619), .o(n9151_1) );
na02f01 g2422 ( .a(n6965), .b(net_7539), .o(n9152) );
ao22f01 g2423 ( .a(_net_292), .b(net_369), .c(_net_291), .d(net_371), .o(n9153) );
na02f01 g2424 ( .a(n9153), .b(n9152), .o(n9154) );
na02f01 g2425 ( .a(n9154), .b(n7400_1), .o(n9155) );
oa12f01 g2426 ( .a(n9155), .b(n7400_1), .c(n9151_1), .o(n3400) );
ao22f01 g2427 ( .a(n7225), .b(_net_7405), .c(n7224), .d(_net_7437), .o(n9157) );
ao22f01 g2428 ( .a(n7229), .b(_net_7501), .c(n7228), .d(_net_7469), .o(n9158) );
na02f01 g2429 ( .a(n9158), .b(n9157), .o(n3422) );
in01f01 g2430 ( .a(_net_7618), .o(n9160_1) );
na02f01 g2431 ( .a(n8000), .b(n7400_1), .o(n9161) );
oa12f01 g2432 ( .a(n9161), .b(n7400_1), .c(n9160_1), .o(n3427) );
ao22f01 g2433 ( .a(n7225), .b(_net_7419), .c(n7224), .d(_net_7451), .o(n9163) );
ao22f01 g2434 ( .a(n7229), .b(_net_7515), .c(n7228), .d(_net_7483), .o(n9164_1) );
na02f01 g2435 ( .a(n9164_1), .b(n9163), .o(n3440) );
ao22f01 g2436 ( .a(n7306), .b(_net_5984), .c(n7298), .d(_net_7720), .o(n9166) );
ao22f01 g2437 ( .a(n7288_1), .b(_net_6028), .c(n7286), .d(_net_267), .o(n9167) );
na02f01 g2438 ( .a(n7302_1), .b(_net_114), .o(n9168) );
na03f01 g2439 ( .a(n7308), .b(_net_193), .c(x1322), .o(n9169_1) );
na02f01 g2440 ( .a(n7296), .b(net_230), .o(n9170) );
na03f01 g2441 ( .a(n7308), .b(net_156), .c(n6800), .o(n9171) );
na03f01 g2442 ( .a(n9171), .b(n9170), .c(n9169_1), .o(n9172) );
ao12f01 g2443 ( .a(n9172), .b(n7291), .c(net_7691), .o(n9173_1) );
na04f01 g2444 ( .a(n9173_1), .b(n9168), .c(n9167), .d(n9166), .o(n3455) );
in01f01 g2445 ( .a(net_6431), .o(n9175) );
in01f01 g2446 ( .a(net_6495), .o(n9176) );
oa22f01 g2447 ( .a(n6750), .b(n9175), .c(n6748), .d(n9176), .o(n9177) );
in01f01 g2448 ( .a(net_6463), .o(n9178_1) );
in01f01 g2449 ( .a(net_6527), .o(n9179) );
oa22f01 g2450 ( .a(n6755), .b(n9178_1), .c(n6754), .d(n9179), .o(n9180) );
no02f01 g2451 ( .a(n9180), .b(n9177), .o(n9181) );
no02f01 g2452 ( .a(n9181), .b(n6764), .o(n9182_1) );
no02f01 g2453 ( .a(n7964), .b(n6766), .o(n9183) );
in01f01 g2454 ( .a(_net_6075), .o(n9184) );
oa22f01 g2455 ( .a(n7077_1), .b(n6775), .c(n6784), .d(n9184), .o(n9185) );
no03f01 g2456 ( .a(n9185), .b(n9183), .c(n9182_1), .o(n9186) );
in01f01 g2457 ( .a(net_6447), .o(n9187_1) );
in01f01 g2458 ( .a(net_6479), .o(n9188) );
oa22f01 g2459 ( .a(n6790), .b(n9187_1), .c(n6789), .d(n9188), .o(n9189) );
in01f01 g2460 ( .a(net_6543), .o(n9190) );
in01f01 g2461 ( .a(net_6511), .o(n9191) );
oa22f01 g2462 ( .a(n6795), .b(n9190), .c(n6794), .d(n9191), .o(n9192_1) );
no02f01 g2463 ( .a(n9192_1), .b(n9189), .o(n9193) );
na02f01 g2464 ( .a(n9193), .b(n9186), .o(n3459) );
no02f01 g2465 ( .a(n7026), .b(n6879), .o(n9195) );
no02f01 g2466 ( .a(_net_7382), .b(net_7378), .o(n9196_1) );
no02f01 g2467 ( .a(n9196_1), .b(n9195), .o(n9197) );
in01f01 g2468 ( .a(n9197), .o(n3464) );
oa12f01 g2469 ( .a(n8213), .b(n8434), .c(n8431), .o(n9199) );
in01f01 g2470 ( .a(n6826_1), .o(n9200) );
ao22f01 g2471 ( .a(n6811), .b(net_6833), .c(n6808), .d(net_6897), .o(n9201_1) );
ao22f01 g2472 ( .a(n6816), .b(net_6865), .c(n6814), .d(net_6929), .o(n9202) );
na02f01 g2473 ( .a(n9202), .b(n9201_1), .o(n9203) );
ao22f01 g2474 ( .a(n9203), .b(n9200), .c(n8211_1), .d(_net_6130), .o(n9204) );
in01f01 g2475 ( .a(n6824), .o(n9205) );
na02f01 g2476 ( .a(n6823), .b(n6822_1), .o(n9206_1) );
no02f01 g2477 ( .a(n9206_1), .b(n6818_1), .o(n9207) );
na02f01 g2478 ( .a(n9138_1), .b(n9137), .o(n9208) );
ao22f01 g2479 ( .a(n6811), .b(net_6831), .c(n6808), .d(net_6895), .o(n9209) );
ao22f01 g2480 ( .a(n6816), .b(net_6863), .c(n6814), .d(net_6927), .o(n9210) );
na02f01 g2481 ( .a(n9210), .b(n9209), .o(n9211_1) );
ao22f01 g2482 ( .a(n9211_1), .b(n9205), .c(n9208), .d(n9207), .o(n9212) );
na03f01 g2483 ( .a(n9212), .b(n9204), .c(n9199), .o(n3474) );
in01f01 g2484 ( .a(_net_6289), .o(n9214) );
no02f01 g2485 ( .a(n9214), .b(_net_392), .o(n3484) );
in01f01 g2486 ( .a(_net_7362), .o(n9216) );
na02f01 g2487 ( .a(n7242), .b(n7030), .o(n9217) );
oa12f01 g2488 ( .a(n9217), .b(n7030), .c(n9216), .o(n3489) );
in01f01 g2489 ( .a(net_6434), .o(n9219) );
in01f01 g2490 ( .a(net_6498), .o(n9220_1) );
oa22f01 g2491 ( .a(n6750), .b(n9219), .c(n6748), .d(n9220_1), .o(n9221) );
in01f01 g2492 ( .a(net_6530), .o(n9222) );
in01f01 g2493 ( .a(net_6466), .o(n9223) );
oa22f01 g2494 ( .a(n6755), .b(n9223), .c(n6754), .d(n9222), .o(n9224) );
no02f01 g2495 ( .a(n9224), .b(n9221), .o(n9225_1) );
no02f01 g2496 ( .a(n9225_1), .b(n6764), .o(n9226) );
in01f01 g2497 ( .a(net_6500), .o(n9227) );
in01f01 g2498 ( .a(net_6436), .o(n9228_1) );
oa22f01 g2499 ( .a(n6750), .b(n9228_1), .c(n6748), .d(n9227), .o(n9229) );
in01f01 g2500 ( .a(net_6468), .o(n9230) );
in01f01 g2501 ( .a(net_6532), .o(n9231) );
oa22f01 g2502 ( .a(n6755), .b(n9230), .c(n6754), .d(n9231), .o(n9232) );
no02f01 g2503 ( .a(n9232), .b(n9229), .o(n9233_1) );
no02f01 g2504 ( .a(n9233_1), .b(n6766), .o(n9234) );
in01f01 g2505 ( .a(_net_6078), .o(n9235) );
oa22f01 g2506 ( .a(n6784), .b(n9235), .c(n6775), .d(n6757), .o(n9236) );
no03f01 g2507 ( .a(n9236), .b(n9234), .c(n9226), .o(n9237) );
in01f01 g2508 ( .a(net_6482), .o(n9238_1) );
in01f01 g2509 ( .a(net_6450), .o(n9239) );
oa22f01 g2510 ( .a(n6790), .b(n9239), .c(n6789), .d(n9238_1), .o(n9240) );
in01f01 g2511 ( .a(net_6514), .o(n9241) );
in01f01 g2512 ( .a(net_6546), .o(n9242_1) );
oa22f01 g2513 ( .a(n6795), .b(n9242_1), .c(n6794), .d(n9241), .o(n9243) );
no02f01 g2514 ( .a(n9243), .b(n9240), .o(n9244) );
na02f01 g2515 ( .a(n9244), .b(n9237), .o(n3507) );
no02f01 g2516 ( .a(n6914), .b(n6912), .o(n9246) );
na03f01 g2517 ( .a(n6944), .b(n8131), .c(_net_6687), .o(n9247) );
na02f01 g2518 ( .a(n6944), .b(n8131), .o(n9248) );
na02f01 g2519 ( .a(n9248), .b(n6943_1), .o(n9249) );
na03f01 g2520 ( .a(n9249), .b(n9247), .c(n9246), .o(n9250_1) );
na02f01 g2521 ( .a(n8132), .b(_net_6687), .o(n9251) );
na02f01 g2522 ( .a(n9251), .b(n9250_1), .o(n3516) );
in01f01 g2523 ( .a(_net_5983), .o(n9253) );
no02f01 g2524 ( .a(n9253), .b(n7570), .o(n3551) );
in01f01 g2525 ( .a(_net_7703), .o(n9255) );
na02f01 g2526 ( .a(n7207_1), .b(_net_7805), .o(n9256) );
oa12f01 g2527 ( .a(n9256), .b(n7207_1), .c(n9255), .o(n3572) );
in01f01 g2528 ( .a(_net_6406), .o(n9258_1) );
na02f01 g2529 ( .a(_net_6405), .b(_net_6404), .o(n9259) );
no02f01 g2530 ( .a(n9259), .b(n9258_1), .o(n9260) );
na02f01 g2531 ( .a(n9260), .b(_net_6407), .o(n9261) );
ao12f01 g2532 ( .a(x38), .b(n9261), .c(_net_6408), .o(n9262) );
oa12f01 g2533 ( .a(n9262), .b(n9261), .c(_net_6408), .o(n3577) );
ao22f01 g2534 ( .a(n6736_1), .b(net_7641), .c(n6734), .d(net_7609), .o(n9264) );
ao22f01 g2535 ( .a(n6739), .b(net_7673), .c(n6738), .d(_net_7577), .o(n9265) );
na02f01 g2536 ( .a(n9265), .b(n9264), .o(n3582) );
no02f01 g2537 ( .a(_net_6557), .b(n6749_1), .o(n9267_1) );
no02f01 g2538 ( .a(n7765), .b(_net_6554), .o(n9268) );
no02f01 g2539 ( .a(n9268), .b(n9267_1), .o(n9269) );
no02f01 g2540 ( .a(n6747), .b(net_6556), .o(n9270) );
no02f01 g2541 ( .a(n9270), .b(n9269), .o(n9271) );
no04f01 g2542 ( .a(n9268), .b(n9267_1), .c(n6747), .d(net_6556), .o(n9272_1) );
no02f01 g2543 ( .a(n6747), .b(n7762), .o(n9273) );
no02f01 g2544 ( .a(_net_6553), .b(net_6556), .o(n9274) );
no02f01 g2545 ( .a(n9274), .b(n9273), .o(n9275) );
oa12f01 g2546 ( .a(n9275), .b(n9272_1), .c(n9271), .o(n9276) );
no02f01 g2547 ( .a(n9272_1), .b(n9271), .o(n9277_1) );
in01f01 g2548 ( .a(n9275), .o(n8472) );
na02f01 g2549 ( .a(n8472), .b(n9277_1), .o(n9279) );
na02f01 g2550 ( .a(n9279), .b(n9276), .o(n3595) );
no02f01 g2551 ( .a(n6966), .b(n7891), .o(n3604) );
ao12f01 g2552 ( .a(n6945), .b(n6929_1), .c(n6924_1), .o(n9282_1) );
no02f01 g2553 ( .a(n8885), .b(n8882_1), .o(n9283) );
no02f01 g2554 ( .a(n9283), .b(n6934_1), .o(n9284) );
in01f01 g2555 ( .a(_net_6092), .o(n9285) );
in01f01 g2556 ( .a(net_6631), .o(n9286) );
in01f01 g2557 ( .a(net_6567), .o(n9287_1) );
oa22f01 g2558 ( .a(n6922), .b(n9287_1), .c(n6919_1), .d(n9286), .o(n9288) );
in01f01 g2559 ( .a(net_6599), .o(n9289) );
in01f01 g2560 ( .a(net_6663), .o(n9290_1) );
oa22f01 g2561 ( .a(n6927), .b(n9289), .c(n6925), .d(n9290_1), .o(n9291) );
no02f01 g2562 ( .a(n9291), .b(n9288), .o(n9292) );
oa22f01 g2563 ( .a(n9292), .b(n6916), .c(n6932), .d(n9285), .o(n9293) );
no03f01 g2564 ( .a(n9293), .b(n9284), .c(n9282_1), .o(n9294_1) );
in01f01 g2565 ( .a(net_6579), .o(n9295) );
in01f01 g2566 ( .a(net_6611), .o(n9296) );
oa22f01 g2567 ( .a(n7058_1), .b(n9295), .c(n7057), .d(n9296), .o(n9297) );
in01f01 g2568 ( .a(net_6643), .o(n9298_1) );
in01f01 g2569 ( .a(net_6675), .o(n9299) );
oa22f01 g2570 ( .a(n7063), .b(n9299), .c(n7062_1), .d(n9298_1), .o(n9300) );
no02f01 g2571 ( .a(n9300), .b(n9297), .o(n9301) );
na02f01 g2572 ( .a(n9301), .b(n9294_1), .o(n3609) );
na02f01 g2573 ( .a(n7348), .b(_net_7797), .o(n9303) );
oa12f01 g2574 ( .a(n9303), .b(n7348), .c(n7538), .o(n3614) );
in01f01 g2575 ( .a(n7357), .o(n9305) );
in01f01 g2576 ( .a(_net_7783), .o(n9306) );
in01f01 g2577 ( .a(_net_7781), .o(n9307_1) );
in01f01 g2578 ( .a(_net_7782), .o(n9308) );
na02f01 g2579 ( .a(n9308), .b(n9307_1), .o(n9309) );
no02f01 g2580 ( .a(n9309), .b(n9306), .o(n9310) );
no02f01 g2581 ( .a(n9310), .b(_net_113), .o(n9311) );
ao12f01 g2582 ( .a(_net_7781), .b(n9311), .c(n9305), .o(n9312_1) );
oa12f01 g2583 ( .a(n7353), .b(n9310), .c(n7357), .o(n9313) );
ao12f01 g2584 ( .a(n9312_1), .b(n9313), .c(_net_7781), .o(n3628) );
in01f01 g2585 ( .a(_net_7665), .o(n9315) );
na02f01 g2586 ( .a(n6965), .b(net_371), .o(n9316_1) );
ao22f01 g2587 ( .a(_net_292), .b(net_383), .c(_net_291), .d(net_385), .o(n9317) );
na02f01 g2588 ( .a(n9317), .b(n9316_1), .o(n9318) );
na02f01 g2589 ( .a(n9318), .b(n7446_1), .o(n9319) );
oa12f01 g2590 ( .a(n9319), .b(n7446_1), .c(n9315), .o(n3633) );
na02f01 g2591 ( .a(n7306), .b(_net_6020), .o(n9321_1) );
na02f01 g2592 ( .a(n7293), .b(net_220), .o(n9322) );
ao22f01 g2593 ( .a(n7297_1), .b(net_183), .c(n7296), .d(net_257), .o(n9323) );
ao22f01 g2594 ( .a(n7298), .b(_net_7747), .c(n7291), .d(_net_7718), .o(n9324) );
na04f01 g2595 ( .a(n9324), .b(n9323), .c(n9322), .d(n9321_1), .o(n3647) );
in01f01 g2596 ( .a(_net_7424), .o(n9326_1) );
na02f01 g2597 ( .a(n1993), .b(n7550), .o(n9327) );
oa12f01 g2598 ( .a(n9327), .b(n7550), .c(n9326_1), .o(n3666) );
in01f01 g2599 ( .a(net_6014), .o(n9329) );
in01f01 g2600 ( .a(_net_7728), .o(n9330_1) );
ao12f01 g2601 ( .a(n7343), .b(n9330_1), .c(n9329), .o(n3675) );
in01f01 g2602 ( .a(_net_5854), .o(n9332) );
in01f01 g2603 ( .a(x940), .o(n9333) );
in01f01 g2604 ( .a(_net_6032), .o(n9334) );
no02f01 g2605 ( .a(_net_6033), .b(n9334), .o(n9335_1) );
na02f01 g2606 ( .a(_net_6028), .b(_net_6034), .o(n9336) );
ao12f01 g2607 ( .a(n9336), .b(n7316_1), .c(_net_5978), .o(n9337) );
na02f01 g2608 ( .a(n9337), .b(n9335_1), .o(n9338) );
in01f01 g2609 ( .a(_net_6033), .o(n9339_1) );
in01f01 g2610 ( .a(n9336), .o(n9340) );
na03f01 g2611 ( .a(n7316_1), .b(_net_5978), .c(_net_5977), .o(n9341) );
na04f01 g2612 ( .a(n9341), .b(n9340), .c(n9339_1), .d(n9334), .o(n9342) );
oa12f01 g2613 ( .a(n7316_1), .b(_net_5978), .c(_net_5977), .o(n9343_1) );
na04f01 g2614 ( .a(n9343_1), .b(n9340), .c(_net_6033), .d(n9334), .o(n9344) );
no02f01 g2615 ( .a(n9339_1), .b(n9334), .o(n9345) );
na03f01 g2616 ( .a(n9345), .b(n9340), .c(_net_5976), .o(n9346) );
na04f01 g2617 ( .a(n9346), .b(n9344), .c(n9342), .d(n9338), .o(n9347) );
na03f01 g2618 ( .a(n9347), .b(net_7776), .c(n9333), .o(n9348_1) );
oa12f01 g2619 ( .a(n9348_1), .b(n9332), .c(x940), .o(n3684) );
in01f01 g2620 ( .a(_net_7250), .o(n9350) );
na02f01 g2621 ( .a(n8731), .b(n6901), .o(n9351) );
oa12f01 g2622 ( .a(n9351), .b(n6901), .c(n9350), .o(n3693) );
in01f01 g2623 ( .a(_net_5853), .o(n9353) );
in01f01 g2624 ( .a(x906), .o(n9354) );
na03f01 g2625 ( .a(n8707), .b(net_7777), .c(n9354), .o(n9355) );
oa12f01 g2626 ( .a(n9355), .b(n9353), .c(x906), .o(n3698) );
na02f01 g2627 ( .a(_net_6017), .b(_net_6023), .o(n9357) );
ao12f01 g2628 ( .a(n9357), .b(_net_5974), .c(n7687), .o(n9358) );
na02f01 g2629 ( .a(n9358), .b(n7695_1), .o(n9359) );
in01f01 g2630 ( .a(n9357), .o(n9360) );
na04f01 g2631 ( .a(n9360), .b(n7697), .c(n7692), .d(n7689), .o(n9361_1) );
na04f01 g2632 ( .a(n9360), .b(n7688), .c(n7692), .d(_net_6022), .o(n9362) );
na03f01 g2633 ( .a(n9360), .b(n7693), .c(_net_5972), .o(n9363) );
na04f01 g2634 ( .a(n9363), .b(n9362), .c(n9361_1), .d(n9359), .o(n9364) );
in01f01 g2635 ( .a(n9364), .o(n9365_1) );
no02f01 g2636 ( .a(n9365_1), .b(x977), .o(n3711) );
in01f01 g2637 ( .a(_net_7444), .o(n9367) );
na02f01 g2638 ( .a(n7553_1), .b(n7197), .o(n9368) );
oa12f01 g2639 ( .a(n9368), .b(n7197), .c(n9367), .o(n3737) );
in01f01 g2640 ( .a(_net_7598), .o(n9370_1) );
na02f01 g2641 ( .a(n6965), .b(net_7550), .o(n9371) );
ao22f01 g2642 ( .a(_net_292), .b(net_380), .c(_net_291), .d(net_382), .o(n9372) );
na02f01 g2643 ( .a(n9372), .b(n9371), .o(n9373_1) );
na02f01 g2644 ( .a(n9373_1), .b(n6968), .o(n9374) );
oa12f01 g2645 ( .a(n9374), .b(n6968), .c(n9370_1), .o(n3742) );
in01f01 g2646 ( .a(_net_290), .o(n9376) );
na02f01 g2647 ( .a(n7440), .b(_net_7810), .o(n9377_1) );
oa12f01 g2648 ( .a(n9377_1), .b(n7440), .c(n9376), .o(n3765) );
in01f01 g2649 ( .a(_net_7626), .o(n9379) );
na02f01 g2650 ( .a(n7707), .b(n7400_1), .o(n9380) );
oa12f01 g2651 ( .a(n9380), .b(n7400_1), .c(n9379), .o(n3782) );
no02f01 g2652 ( .a(n6978), .b(n6976), .o(n9382) );
na03f01 g2653 ( .a(n7011), .b(n7219), .c(_net_7092), .o(n9383) );
na02f01 g2654 ( .a(n7011), .b(n7219), .o(n9384) );
na02f01 g2655 ( .a(n9384), .b(n7010), .o(n9385_1) );
na03f01 g2656 ( .a(n9385_1), .b(n9383), .c(n9382), .o(n9386) );
na02f01 g2657 ( .a(n7220), .b(_net_7092), .o(n9387) );
na02f01 g2658 ( .a(n9387), .b(n9386), .o(n3787) );
no02f01 g2659 ( .a(_net_7784), .b(_net_7785), .o(n9389) );
no03f01 g2660 ( .a(n9389), .b(n7362), .c(n7358), .o(n3796) );
ao22f01 g2661 ( .a(n6877), .b(_net_7276), .c(n6876_1), .d(net_7340), .o(n9391) );
ao22f01 g2662 ( .a(n6881_1), .b(net_7308), .c(n6880), .d(net_7372), .o(n9392) );
na02f01 g2663 ( .a(n9392), .b(n9391), .o(n3813) );
no03f01 g2664 ( .a(n7850), .b(n7415), .c(_net_282), .o(n9394) );
no02f01 g2665 ( .a(n7850), .b(n7410), .o(n9395) );
ao22f01 g2666 ( .a(n9395), .b(n7416), .c(n9394), .d(n7420), .o(n9396) );
ao12f01 g2667 ( .a(n7850), .b(_net_229), .c(n7410), .o(n9397) );
no03f01 g2668 ( .a(n7850), .b(_net_283), .c(_net_282), .o(n9398_1) );
ao22f01 g2669 ( .a(n9398_1), .b(n7418), .c(n9397), .d(n7409), .o(n9399) );
na02f01 g2670 ( .a(n9399), .b(n9396), .o(n3827) );
in01f01 g2671 ( .a(_net_6419), .o(n9401) );
in01f01 g2672 ( .a(_net_6401), .o(n9402_1) );
in01f01 g2673 ( .a(_net_6422), .o(n9403) );
in01f01 g2674 ( .a(_net_6423), .o(n9404) );
in01f01 g2675 ( .a(_net_6418), .o(n9405_1) );
no04f01 g2676 ( .a(_net_6421), .b(n9405_1), .c(n9404), .d(_net_6420), .o(n9406) );
na03f01 g2677 ( .a(n9406), .b(n9403), .c(n9401), .o(n9407) );
in01f01 g2678 ( .a(n9407), .o(n7691) );
na02f01 g2679 ( .a(n7691), .b(n9402_1), .o(n9409) );
no02f01 g2680 ( .a(n7691), .b(_net_6401), .o(n9410_1) );
in01f01 g2681 ( .a(n9410_1), .o(n9411) );
na02f01 g2682 ( .a(_net_6418), .b(_net_6419), .o(n9412) );
na02f01 g2683 ( .a(n9405_1), .b(n9401), .o(n9413) );
na02f01 g2684 ( .a(n9413), .b(n9412), .o(n9414) );
oa22f01 g2685 ( .a(n9414), .b(n9411), .c(n9409), .d(n9401), .o(n3836) );
in01f01 g2686 ( .a(_net_7652), .o(n9416) );
na02f01 g2687 ( .a(n8426_1), .b(n7446_1), .o(n9417) );
oa12f01 g2688 ( .a(n9417), .b(n7446_1), .c(n9416), .o(n3841) );
no02f01 g2689 ( .a(n8790), .b(n7012), .o(n9419) );
no02f01 g2690 ( .a(n8602_1), .b(n6997), .o(n9420_1) );
in01f01 g2691 ( .a(_net_6158), .o(n9421) );
oa22f01 g2692 ( .a(n8610), .b(n6980), .c(n6995_1), .d(n9421), .o(n9422) );
no03f01 g2693 ( .a(n9422), .b(n9420_1), .c(n9419), .o(n9423) );
in01f01 g2694 ( .a(net_7022), .o(n9424) );
in01f01 g2695 ( .a(net_6990), .o(n9425_1) );
oa22f01 g2696 ( .a(n8075_1), .b(n9425_1), .c(n8074), .d(n9424), .o(n9426) );
in01f01 g2697 ( .a(net_7054), .o(n9427) );
in01f01 g2698 ( .a(net_7086), .o(n9428_1) );
oa22f01 g2699 ( .a(n8080_1), .b(n9428_1), .c(n8079), .d(n9427), .o(n9429) );
no02f01 g2700 ( .a(n9429), .b(n9426), .o(n9430) );
na02f01 g2701 ( .a(n9430), .b(n9423), .o(n3846) );
in01f01 g2702 ( .a(_net_7290), .o(n9432) );
na02f01 g2703 ( .a(n7393), .b(n7180), .o(n9433) );
oa12f01 g2704 ( .a(n9433), .b(n7180), .c(n9432), .o(n3859) );
no02f01 g2705 ( .a(n7027_1), .b(n6875), .o(n9435) );
no02f01 g2706 ( .a(_net_7383), .b(_net_7379), .o(n9436_1) );
no02f01 g2707 ( .a(n9436_1), .b(n9435), .o(n9437) );
in01f01 g2708 ( .a(n9437), .o(n9438) );
na02f01 g2709 ( .a(n9438), .b(n3464), .o(n9439) );
in01f01 g2710 ( .a(_net_7380), .o(n9440) );
in01f01 g2711 ( .a(_net_7384), .o(n9441_1) );
no02f01 g2712 ( .a(n9441_1), .b(n9440), .o(n9442) );
no02f01 g2713 ( .a(_net_7384), .b(_net_7380), .o(n9443) );
no02f01 g2714 ( .a(n9443), .b(n9442), .o(n9444) );
no04f01 g2715 ( .a(n9444), .b(n9439), .c(n6899_1), .d(_net_7381), .o(n3872) );
na02f01 g2716 ( .a(n8034), .b(_net_6065), .o(n9446) );
na02f01 g2717 ( .a(n8037), .b(n8028_1), .o(n9447) );
na02f01 g2718 ( .a(n9447), .b(n9446), .o(n3877) );
in01f01 g2719 ( .a(_net_7574), .o(n9449_1) );
na02f01 g2720 ( .a(n2850), .b(n7519), .o(n9450) );
oa12f01 g2721 ( .a(n9450), .b(n7519), .c(n9449_1), .o(n3886) );
in01f01 g2722 ( .a(_net_123), .o(n9452) );
na02f01 g2723 ( .a(_net_154), .b(net_319), .o(n9453) );
oa12f01 g2724 ( .a(n9453), .b(n9452), .c(_net_154), .o(n3891) );
ao22f01 g2725 ( .a(n7225), .b(_net_7431), .c(n7224), .d(net_7463), .o(n9455) );
ao22f01 g2726 ( .a(n7229), .b(net_7527), .c(n7228), .d(net_7495), .o(n9456) );
na02f01 g2727 ( .a(n9456), .b(n9455), .o(n3908) );
in01f01 g2728 ( .a(_net_7270), .o(n9458) );
na02f01 g2729 ( .a(n1029), .b(n6901), .o(n9459_1) );
oa12f01 g2730 ( .a(n9459_1), .b(n6901), .c(n9458), .o(n3913) );
in01f01 g2731 ( .a(net_6766), .o(n9461) );
in01f01 g2732 ( .a(net_6702), .o(n9462_1) );
oa22f01 g2733 ( .a(n7129), .b(n9462_1), .c(n7126), .d(n9461), .o(n9463) );
in01f01 g2734 ( .a(net_6734), .o(n9464) );
in01f01 g2735 ( .a(net_6798), .o(n9465) );
oa22f01 g2736 ( .a(n7134), .b(n9464), .c(n7132), .d(n9465), .o(n9466) );
no02f01 g2737 ( .a(n9466), .b(n9463), .o(n9467_1) );
no02f01 g2738 ( .a(n9467_1), .b(n7468_1), .o(n9468) );
no02f01 g2739 ( .a(n8557_1), .b(n7470), .o(n9469) );
in01f01 g2740 ( .a(_net_6116), .o(n9470_1) );
oa22f01 g2741 ( .a(n7465), .b(n7123), .c(n7118), .d(n9470_1), .o(n9471) );
no03f01 g2742 ( .a(n9471), .b(n9469), .c(n9468), .o(n9472) );
in01f01 g2743 ( .a(net_6718), .o(n9473) );
in01f01 g2744 ( .a(net_6750), .o(n9474) );
oa22f01 g2745 ( .a(n7492_1), .b(n9473), .c(n7491), .d(n9474), .o(n9475_1) );
in01f01 g2746 ( .a(net_6814), .o(n9476) );
in01f01 g2747 ( .a(net_6782), .o(n9477) );
oa22f01 g2748 ( .a(n7497), .b(n9476), .c(n7496_1), .d(n9477), .o(n9478_1) );
no02f01 g2749 ( .a(n9478_1), .b(n9475_1), .o(n9479) );
na02f01 g2750 ( .a(n9479), .b(n9472), .o(n3922) );
in01f01 g2751 ( .a(_net_7563), .o(n9481) );
na02f01 g2752 ( .a(n7519), .b(n6971), .o(n9482) );
oa12f01 g2753 ( .a(n9482), .b(n7519), .c(n9481), .o(n3927) );
in01f01 g2754 ( .a(_net_7418), .o(n9484) );
na02f01 g2755 ( .a(n6866), .b(net_351), .o(n9485) );
ao22f01 g2756 ( .a(_net_281), .b(net_363), .c(_net_280), .d(net_365), .o(n9486) );
na02f01 g2757 ( .a(n9486), .b(n9485), .o(n9487_1) );
na02f01 g2758 ( .a(n9487_1), .b(n7550), .o(n9488) );
oa12f01 g2759 ( .a(n9488), .b(n7550), .c(n9484), .o(n3932) );
in01f01 g2760 ( .a(_net_7591), .o(n9490) );
na02f01 g2761 ( .a(n6965), .b(net_7543), .o(n9491) );
ao22f01 g2762 ( .a(_net_292), .b(net_373), .c(_net_291), .d(net_375), .o(n9492_1) );
na02f01 g2763 ( .a(n9492_1), .b(n9491), .o(n9493) );
na02f01 g2764 ( .a(n9493), .b(n6968), .o(n9494) );
oa12f01 g2765 ( .a(n9494), .b(n6968), .c(n9490), .o(n3941) );
in01f01 g2766 ( .a(_net_7510), .o(n9496) );
na02f01 g2767 ( .a(n8994), .b(n7626_1), .o(n9497_1) );
oa12f01 g2768 ( .a(n9497_1), .b(n7626_1), .c(n9496), .o(n3967) );
in01f01 g2769 ( .a(_net_6201), .o(n9499) );
no02f01 g2770 ( .a(n9499), .b(_net_392), .o(n3976) );
ao12f01 g2771 ( .a(n7468_1), .b(n8156_1), .c(n8155), .o(n9501) );
no02f01 g2772 ( .a(n8979), .b(n8976_1), .o(n9502_1) );
no02f01 g2773 ( .a(n9502_1), .b(n7470), .o(n9503) );
in01f01 g2774 ( .a(_net_6112), .o(n9504) );
oa22f01 g2775 ( .a(n9467_1), .b(n7123), .c(n7118), .d(n9504), .o(n9505) );
no03f01 g2776 ( .a(n9505), .b(n9503), .c(n9501), .o(n9506) );
in01f01 g2777 ( .a(net_6746), .o(n9507_1) );
in01f01 g2778 ( .a(net_6714), .o(n9508) );
oa22f01 g2779 ( .a(n7492_1), .b(n9508), .c(n7491), .d(n9507_1), .o(n9509) );
in01f01 g2780 ( .a(net_6810), .o(n9510) );
in01f01 g2781 ( .a(net_6778), .o(n9511) );
oa22f01 g2782 ( .a(n7497), .b(n9510), .c(n7496_1), .d(n9511), .o(n9512_1) );
no02f01 g2783 ( .a(n9512_1), .b(n9509), .o(n9513) );
na02f01 g2784 ( .a(n9513), .b(n9506), .o(n3981) );
in01f01 g2785 ( .a(_net_7095), .o(n9515) );
na03f01 g2786 ( .a(n7210), .b(n9515), .c(_net_7094), .o(n9516) );
oa12f01 g2787 ( .a(_net_7095), .b(n7212_1), .c(n6986_1), .o(n9517_1) );
na02f01 g2788 ( .a(n9517_1), .b(n9516), .o(n9518) );
na02f01 g2789 ( .a(n9518), .b(n7215), .o(n9519) );
no02f01 g2790 ( .a(n6991), .b(n9515), .o(n9520_1) );
no02f01 g2791 ( .a(n7002), .b(_net_7095), .o(n9521) );
no02f01 g2792 ( .a(n9521), .b(n9520_1), .o(n9522) );
ao22f01 g2793 ( .a(n9522), .b(n7218), .c(n7220), .d(_net_7095), .o(n9523) );
na02f01 g2794 ( .a(n9523), .b(n9519), .o(n3998) );
in01f01 g2795 ( .a(_net_7733), .o(n9525_1) );
in01f01 g2796 ( .a(_net_6027), .o(n9526) );
ao12f01 g2797 ( .a(n7343), .b(n9526), .c(n9525_1), .o(n4016) );
in01f01 g2798 ( .a(_net_7601), .o(n9528_1) );
na02f01 g2799 ( .a(n9318), .b(n6968), .o(n9529) );
oa12f01 g2800 ( .a(n9529), .b(n6968), .c(n9528_1), .o(n4029) );
in01f01 g2801 ( .a(_net_7633), .o(n9531) );
na02f01 g2802 ( .a(n9318), .b(n7400_1), .o(n9532) );
oa12f01 g2803 ( .a(n9532), .b(n7400_1), .c(n9531), .o(n4042) );
in01f01 g2804 ( .a(_net_7329), .o(n9534) );
na02f01 g2805 ( .a(n6898), .b(net_7249), .o(n9535) );
ao22f01 g2806 ( .a(net_341), .b(_net_270), .c(_net_269), .d(net_343), .o(n9536) );
na02f01 g2807 ( .a(n9536), .b(n9535), .o(n9537_1) );
na02f01 g2808 ( .a(n9537_1), .b(n7150), .o(n9538) );
oa12f01 g2809 ( .a(n9538), .b(n7150), .c(n9534), .o(n4063) );
in01f01 g2810 ( .a(_net_294), .o(n9540) );
na02f01 g2811 ( .a(n7440), .b(_net_7814), .o(n9541_1) );
oa12f01 g2812 ( .a(n9541_1), .b(n7440), .c(n9540), .o(n4084) );
no02f01 g2813 ( .a(n9261), .b(n8178), .o(n9543) );
na03f01 g2814 ( .a(n9543), .b(_net_6410), .c(n8084), .o(n9544) );
in01f01 g2815 ( .a(_net_6410), .o(n9545) );
in01f01 g2816 ( .a(n9543), .o(n9546_1) );
oa12f01 g2817 ( .a(_net_6411), .b(n9546_1), .c(n9545), .o(n9547) );
na03f01 g2818 ( .a(n9547), .b(n9544), .c(n6910_1), .o(n4089) );
in01f01 g2819 ( .a(_net_7404), .o(n9549_1) );
na02f01 g2820 ( .a(n7952), .b(n7550), .o(n9550) );
oa12f01 g2821 ( .a(n9550), .b(n7550), .c(n9549_1), .o(n4094) );
in01f01 g2822 ( .a(_net_7719), .o(n9552) );
na02f01 g2823 ( .a(n7207_1), .b(_net_7821), .o(n9553) );
oa12f01 g2824 ( .a(n9553), .b(n7207_1), .c(n9552), .o(n4107) );
in01f01 g2825 ( .a(_net_7364), .o(n9555) );
na02f01 g2826 ( .a(n7256_1), .b(n7030), .o(n9556) );
oa12f01 g2827 ( .a(n9556), .b(n7030), .c(n9555), .o(n4116) );
in01f01 g2828 ( .a(_net_276), .o(n9558) );
na02f01 g2829 ( .a(_net_190), .b(_net_188), .o(n9559_1) );
na02f01 g2830 ( .a(n9559_1), .b(n9558), .o(n4121) );
no02f01 g2831 ( .a(n7572_1), .b(n7570), .o(n9561) );
na03f01 g2832 ( .a(n7720), .b(n8311_1), .c(_net_7227), .o(n9562) );
na02f01 g2833 ( .a(n7720), .b(n8311_1), .o(n9563) );
na02f01 g2834 ( .a(n9563), .b(n7719_1), .o(n9564_1) );
na03f01 g2835 ( .a(n9564_1), .b(n9562), .c(n9561), .o(n9565) );
na02f01 g2836 ( .a(n8312), .b(_net_7227), .o(n9566) );
na02f01 g2837 ( .a(n9566), .b(n9565), .o(n4126) );
in01f01 g2838 ( .a(n3551), .o(n9568) );
no02f01 g2839 ( .a(_net_7232), .b(n9113), .o(n9569_1) );
no02f01 g2840 ( .a(n9116), .b(net_7231), .o(n9570) );
no02f01 g2841 ( .a(n9570), .b(n9569_1), .o(n9571) );
na02f01 g2842 ( .a(n9253), .b(_net_6039), .o(n9572) );
oa22f01 g2843 ( .a(n9572), .b(n9116), .c(n9571), .d(n9568), .o(n4135) );
in01f01 g2844 ( .a(_net_7347), .o(n9574_1) );
na02f01 g2845 ( .a(n7659), .b(n7030), .o(n9575) );
oa12f01 g2846 ( .a(n9575), .b(n7030), .c(n9574_1), .o(n4140) );
in01f01 g2847 ( .a(_net_7437), .o(n9577) );
na02f01 g2848 ( .a(n8817), .b(n7197), .o(n9578) );
oa12f01 g2849 ( .a(n9578), .b(n7197), .c(n9577), .o(n4166) );
no02f01 g2850 ( .a(_net_7784), .b(_net_113), .o(n4171) );
ao22f01 g2851 ( .a(n6738), .b(_net_7556), .c(n6736_1), .d(_net_7620), .o(n9581) );
ao22f01 g2852 ( .a(n6739), .b(_net_7652), .c(n6734), .d(_net_7588), .o(n9582) );
na02f01 g2853 ( .a(n9582), .b(n9581), .o(n4181) );
in01f01 g2854 ( .a(_net_7321), .o(n9584) );
na02f01 g2855 ( .a(n6898), .b(net_7241), .o(n9585) );
ao22f01 g2856 ( .a(net_333), .b(_net_270), .c(net_335), .d(_net_269), .o(n9586) );
na02f01 g2857 ( .a(n9586), .b(n9585), .o(n9587) );
na02f01 g2858 ( .a(n9587), .b(n7150), .o(n9588_1) );
oa12f01 g2859 ( .a(n9588_1), .b(n7150), .c(n9584), .o(n4186) );
in01f01 g2860 ( .a(_net_277), .o(n9590) );
in01f01 g2861 ( .a(_net_189), .o(n9591) );
in01f01 g2862 ( .a(n6897), .o(n9592_1) );
oa12f01 g2863 ( .a(n9590), .b(n9592_1), .c(n9591), .o(n4203) );
ao22f01 g2864 ( .a(n7225), .b(_net_7414), .c(n7224), .d(_net_7446), .o(n9594) );
ao22f01 g2865 ( .a(n7229), .b(_net_7510), .c(n7228), .d(_net_7478), .o(n9595) );
na02f01 g2866 ( .a(n9595), .b(n9594), .o(n4212) );
in01f01 g2867 ( .a(_net_7630), .o(n9597_1) );
na02f01 g2868 ( .a(n9373_1), .b(n7400_1), .o(n9598) );
oa12f01 g2869 ( .a(n9598), .b(n7400_1), .c(n9597_1), .o(n4217) );
in01f01 g2870 ( .a(_net_6825), .o(n9600) );
no02f01 g2871 ( .a(n7125_1), .b(n7466), .o(n9601) );
na03f01 g2872 ( .a(n9601), .b(_net_6824), .c(n9600), .o(n9602_1) );
in01f01 g2873 ( .a(n9601), .o(n9603) );
oa12f01 g2874 ( .a(_net_6825), .b(n9603), .c(n7128_1), .o(n9604) );
na02f01 g2875 ( .a(n9604), .b(n9602_1), .o(n9605) );
na02f01 g2876 ( .a(n9605), .b(_net_6828), .o(n9606_1) );
in01f01 g2877 ( .a(_net_6828), .o(n9607) );
na03f01 g2878 ( .a(n9604), .b(n9602_1), .c(n9607), .o(n9608) );
na02f01 g2879 ( .a(_net_6823), .b(n7466), .o(n9609) );
na02f01 g2880 ( .a(n7125_1), .b(_net_6822), .o(n9610) );
na02f01 g2881 ( .a(n9610), .b(n9609), .o(n9611_1) );
na02f01 g2882 ( .a(n9611_1), .b(net_6826), .o(n9612) );
na03f01 g2883 ( .a(n9610), .b(n9609), .c(n8220_1), .o(n9613) );
ao22f01 g2884 ( .a(n9613), .b(n9612), .c(n7467), .d(_net_6822), .o(n9614) );
na02f01 g2885 ( .a(n9601), .b(n7128_1), .o(n9615) );
na02f01 g2886 ( .a(n9603), .b(_net_6824), .o(n9616_1) );
na02f01 g2887 ( .a(n9616_1), .b(n9615), .o(n9617) );
na02f01 g2888 ( .a(n9617), .b(n8219), .o(n9618) );
na03f01 g2889 ( .a(n9616_1), .b(n9615), .c(_net_6827), .o(n9619) );
na03f01 g2890 ( .a(n9619), .b(n9618), .c(n9614), .o(n9620_1) );
ao12f01 g2891 ( .a(n9620_1), .b(n9608), .c(n9606_1), .o(n4226) );
in01f01 g2892 ( .a(_net_7635), .o(n9622) );
na02f01 g2893 ( .a(n7400_1), .b(n7144), .o(n9623) );
oa12f01 g2894 ( .a(n9623), .b(n7400_1), .c(n9622), .o(n4240) );
ao12f01 g2895 ( .a(n7012), .b(n7004), .c(n7001), .o(n9625) );
no02f01 g2896 ( .a(n6993), .b(n6988), .o(n9626) );
no02f01 g2897 ( .a(n6997), .b(n9626), .o(n9627) );
in01f01 g2898 ( .a(_net_6152), .o(n9628_1) );
oa22f01 g2899 ( .a(n8782), .b(n6980), .c(n6995_1), .d(n9628_1), .o(n9629) );
no03f01 g2900 ( .a(n9629), .b(n9627), .c(n9625), .o(n9630) );
in01f01 g2901 ( .a(net_7016), .o(n9631) );
in01f01 g2902 ( .a(net_6984), .o(n9632) );
oa22f01 g2903 ( .a(n8075_1), .b(n9632), .c(n8074), .d(n9631), .o(n9633_1) );
in01f01 g2904 ( .a(net_7048), .o(n9634) );
in01f01 g2905 ( .a(net_7080), .o(n9635) );
oa22f01 g2906 ( .a(n8080_1), .b(n9635), .c(n8079), .d(n9634), .o(n9636) );
no02f01 g2907 ( .a(n9636), .b(n9633_1), .o(n9637) );
na02f01 g2908 ( .a(n9637), .b(n9630), .o(n4249) );
no02f01 g2909 ( .a(n7576), .b(n9113), .o(n9639) );
no02f01 g2910 ( .a(_net_7228), .b(net_7231), .o(n9640) );
no02f01 g2911 ( .a(n9640), .b(n9639), .o(n9641) );
in01f01 g2912 ( .a(n9641), .o(n4276) );
no02f01 g2913 ( .a(n7194_1), .b(net_7529), .o(n9643) );
in01f01 g2914 ( .a(n9643), .o(n9644) );
no02f01 g2915 ( .a(n9644), .b(n8923), .o(n9645) );
no02f01 g2916 ( .a(n9643), .b(n8924), .o(n9646) );
oa12f01 g2917 ( .a(n8919), .b(n9646), .c(n9645), .o(n9647_1) );
no02f01 g2918 ( .a(n9646), .b(n9645), .o(n9648) );
na02f01 g2919 ( .a(n9648), .b(n8850), .o(n9649) );
na02f01 g2920 ( .a(n9649), .b(n9647_1), .o(n4289) );
in01f01 g2921 ( .a(_net_7318), .o(n9651_1) );
na02f01 g2922 ( .a(n8960), .b(n7150), .o(n9652) );
oa12f01 g2923 ( .a(n9652), .b(n7150), .c(n9651_1), .o(n4294) );
na02f01 g2924 ( .a(n9203), .b(n8213), .o(n9654) );
ao22f01 g2925 ( .a(n9211_1), .b(n9200), .c(n8211_1), .d(_net_6128), .o(n9655_1) );
ao22f01 g2926 ( .a(n6811), .b(net_6829), .c(n6808), .d(net_6893), .o(n9656) );
ao22f01 g2927 ( .a(n6816), .b(net_6861), .c(n6814), .d(net_6925), .o(n9657) );
na02f01 g2928 ( .a(n9657), .b(n9656), .o(n9658) );
na02f01 g2929 ( .a(n9658), .b(n9205), .o(n9659) );
oa12f01 g2930 ( .a(n9207), .b(n9134_1), .c(n9131), .o(n9660_1) );
na04f01 g2931 ( .a(n9660_1), .b(n9659), .c(n9655_1), .d(n9654), .o(n4299) );
no04f01 g2932 ( .a(n7338), .b(n7107_1), .c(n7106), .d(x1155), .o(n4304) );
in01f01 g2933 ( .a(_net_6421), .o(n9663) );
na03f01 g2934 ( .a(_net_6418), .b(_net_6420), .c(_net_6419), .o(n9664_1) );
no02f01 g2935 ( .a(n9664_1), .b(n9663), .o(n9665) );
no02f01 g2936 ( .a(n9665), .b(_net_6422), .o(n9666) );
na02f01 g2937 ( .a(n9665), .b(_net_6422), .o(n9667) );
na02f01 g2938 ( .a(n9667), .b(n9410_1), .o(n9668_1) );
oa22f01 g2939 ( .a(n9668_1), .b(n9666), .c(n9409), .d(n9403), .o(n4313) );
na03f01 g2940 ( .a(n8089), .b(n8084), .c(_net_6408), .o(n9670) );
in01f01 g2941 ( .a(_net_6409), .o(n9671) );
na02f01 g2942 ( .a(n9671), .b(n9545), .o(n9672) );
no04f01 g2943 ( .a(n9672), .b(n9670), .c(_net_6407), .d(_net_6406), .o(n4322) );
in01f01 g2944 ( .a(_net_7505), .o(n9674) );
na02f01 g2945 ( .a(n7626_1), .b(n7200), .o(n9675) );
oa12f01 g2946 ( .a(n9675), .b(n7626_1), .c(n9674), .o(n4348) );
in01f01 g2947 ( .a(_net_6009), .o(n9677) );
na02f01 g2948 ( .a(n7348), .b(_net_7812), .o(n9678_1) );
oa12f01 g2949 ( .a(n9678_1), .b(n7348), .c(n9677), .o(n4357) );
in01f01 g2950 ( .a(_net_7278), .o(n9680) );
na02f01 g2951 ( .a(n576), .b(n6901), .o(n9681) );
oa12f01 g2952 ( .a(n9681), .b(n6901), .c(n9680), .o(n4379) );
in01f01 g2953 ( .a(_net_7301), .o(n9683_1) );
in01f01 g2954 ( .a(net_333), .o(n9684) );
oa22f01 g2955 ( .a(n6899_1), .b(n9684), .c(n7253), .d(n7514), .o(n9685) );
na02f01 g2956 ( .a(n9685), .b(n7180), .o(n9686) );
oa12f01 g2957 ( .a(n9686), .b(n7180), .c(n9683_1), .o(n4392) );
in01f01 g2958 ( .a(_net_7718), .o(n9688) );
na02f01 g2959 ( .a(n7207_1), .b(_net_7820), .o(n9689) );
oa12f01 g2960 ( .a(n9689), .b(n7207_1), .c(n9688), .o(n4414) );
in01f01 g2961 ( .a(net_7807), .o(n9691) );
na02f01 g2962 ( .a(n6803), .b(_net_6045), .o(n9692_1) );
oa12f01 g2963 ( .a(n9692_1), .b(n6803), .c(n9691), .o(n4424) );
in01f01 g2964 ( .a(_net_7332), .o(n9694) );
na02f01 g2965 ( .a(n7256_1), .b(n7150), .o(n9695_1) );
oa12f01 g2966 ( .a(n9695_1), .b(n7150), .c(n9694), .o(n4433) );
in01f01 g2967 ( .a(_net_7403), .o(n9697) );
na02f01 g2968 ( .a(n6866), .b(net_7387), .o(n9698) );
ao22f01 g2969 ( .a(net_350), .b(_net_280), .c(net_348), .d(_net_281), .o(n9699) );
na02f01 g2970 ( .a(n9699), .b(n9698), .o(n9700_1) );
na02f01 g2971 ( .a(n9700_1), .b(n7550), .o(n9701) );
oa12f01 g2972 ( .a(n9701), .b(n7550), .c(n9697), .o(n4438) );
in01f01 g2973 ( .a(_net_6205), .o(n9703) );
no02f01 g2974 ( .a(_net_392), .b(n9703), .o(n4443) );
oa12f01 g2975 ( .a(n7284_1), .b(n7282), .c(x1322), .o(n9705) );
no02f01 g2976 ( .a(n9705), .b(n7293), .o(n9706) );
in01f01 g2977 ( .a(n7347), .o(n9707) );
na03f01 g2978 ( .a(n9707), .b(n9706), .c(_net_6023), .o(n9708) );
na02f01 g2979 ( .a(n7293), .b(net_223), .o(n9709_1) );
ao22f01 g2980 ( .a(n7297_1), .b(net_186), .c(n7296), .d(net_260), .o(n9710) );
na03f01 g2981 ( .a(n9710), .b(n9709_1), .c(n9708), .o(n4456) );
in01f01 g2982 ( .a(_net_7323), .o(n9712) );
na02f01 g2983 ( .a(n7150), .b(n7033), .o(n9713) );
oa12f01 g2984 ( .a(n9713), .b(n7150), .c(n9712), .o(n4464) );
na02f01 g2985 ( .a(n7005_1), .b(n6981), .o(n9715) );
ao22f01 g2986 ( .a(n7009_1), .b(n6998), .c(n6996), .d(_net_6148), .o(n9716) );
ao22f01 g2987 ( .a(n7000_1), .b(net_6964), .c(n6999), .d(net_7028), .o(n9717) );
ao22f01 g2988 ( .a(n7003), .b(net_6996), .c(n7002), .d(net_7060), .o(n9718) );
na02f01 g2989 ( .a(n9718), .b(n9717), .o(n9719_1) );
na02f01 g2990 ( .a(n9719_1), .b(n7013_1), .o(n9720) );
oa12f01 g2991 ( .a(n7022), .b(n8618), .c(n8615), .o(n9721) );
na04f01 g2992 ( .a(n9721), .b(n9720), .c(n9716), .d(n9715), .o(n4482) );
in01f01 g2993 ( .a(_net_6018), .o(n9723) );
na02f01 g2994 ( .a(n7348), .b(_net_7818), .o(n9724_1) );
oa12f01 g2995 ( .a(n9724_1), .b(n7348), .c(n9723), .o(n4491) );
no02f01 g2996 ( .a(net_153), .b(n8016), .o(n4501) );
in01f01 g2997 ( .a(_net_7469), .o(n9727) );
na02f01 g2998 ( .a(n8817), .b(n6869), .o(n9728) );
oa12f01 g2999 ( .a(n9728), .b(n6869), .c(n9727), .o(n4510) );
ao12f01 g3000 ( .a(n7721), .b(n8498), .c(n8497), .o(n9730) );
no02f01 g3001 ( .a(n9005_1), .b(n7592), .o(n9731) );
in01f01 g3002 ( .a(_net_6173), .o(n9732) );
oa22f01 g3003 ( .a(n8274), .b(n7574), .c(n7590), .d(n9732), .o(n9733_1) );
no03f01 g3004 ( .a(n9733_1), .b(n9731), .c(n9730), .o(n9734) );
in01f01 g3005 ( .a(net_7120), .o(n9735) );
in01f01 g3006 ( .a(net_7152), .o(n9736) );
oa22f01 g3007 ( .a(n7740), .b(n9735), .c(n7739), .d(n9736), .o(n9737_1) );
in01f01 g3008 ( .a(net_7184), .o(n9738) );
in01f01 g3009 ( .a(net_7216), .o(n9739) );
oa22f01 g3010 ( .a(n7745), .b(n9739), .c(n7744), .d(n9738), .o(n9740) );
no02f01 g3011 ( .a(n9740), .b(n9737_1), .o(n9741) );
na02f01 g3012 ( .a(n9741), .b(n9734), .o(n4515) );
ao22f01 g3013 ( .a(n6736_1), .b(_net_7632), .c(n6734), .d(_net_7600), .o(n9743) );
ao22f01 g3014 ( .a(n6739), .b(_net_7664), .c(n6738), .d(_net_7568), .o(n9744) );
na02f01 g3015 ( .a(n9744), .b(n9743), .o(n4520) );
in01f01 g3016 ( .a(_net_6188), .o(n9746_1) );
no02f01 g3017 ( .a(n9746_1), .b(_net_392), .o(n4529) );
in01f01 g3018 ( .a(_net_6194), .o(n9748) );
no02f01 g3019 ( .a(_net_392), .b(n9748), .o(n4534) );
ao12f01 g3020 ( .a(n7721), .b(n7907), .c(n7906_1), .o(n9750_1) );
in01f01 g3021 ( .a(net_7105), .o(n9751) );
in01f01 g3022 ( .a(net_7169), .o(n9752) );
oa22f01 g3023 ( .a(n7580), .b(n9751), .c(n7577_1), .d(n9752), .o(n9753) );
in01f01 g3024 ( .a(net_7201), .o(n9754_1) );
in01f01 g3025 ( .a(net_7137), .o(n9755) );
oa22f01 g3026 ( .a(n7585), .b(n9755), .c(n7583), .d(n9754_1), .o(n9756) );
no02f01 g3027 ( .a(n9756), .b(n9753), .o(n9757) );
no02f01 g3028 ( .a(n9757), .b(n7592), .o(n9758_1) );
in01f01 g3029 ( .a(_net_6172), .o(n9759) );
in01f01 g3030 ( .a(net_7171), .o(n9760) );
in01f01 g3031 ( .a(net_7107), .o(n9761) );
oa22f01 g3032 ( .a(n7580), .b(n9761), .c(n7577_1), .d(n9760), .o(n9762) );
in01f01 g3033 ( .a(net_7203), .o(n9763_1) );
in01f01 g3034 ( .a(net_7139), .o(n9764) );
oa22f01 g3035 ( .a(n7585), .b(n9764), .c(n7583), .d(n9763_1), .o(n9765) );
no02f01 g3036 ( .a(n9765), .b(n9762), .o(n9766) );
oa22f01 g3037 ( .a(n9766), .b(n7574), .c(n7590), .d(n9759), .o(n9767) );
no03f01 g3038 ( .a(n9767), .b(n9758_1), .c(n9750_1), .o(n9768_1) );
in01f01 g3039 ( .a(net_7119), .o(n9769) );
in01f01 g3040 ( .a(net_7151), .o(n9770) );
oa22f01 g3041 ( .a(n7740), .b(n9769), .c(n7739), .d(n9770), .o(n9771) );
in01f01 g3042 ( .a(net_7215), .o(n9772) );
in01f01 g3043 ( .a(net_7183), .o(n9773_1) );
oa22f01 g3044 ( .a(n7745), .b(n9772), .c(n7744), .d(n9773_1), .o(n9774) );
no02f01 g3045 ( .a(n9774), .b(n9771), .o(n9775) );
na02f01 g3046 ( .a(n9775), .b(n9768_1), .o(n4539) );
in01f01 g3047 ( .a(_net_7480), .o(n9777) );
na02f01 g3048 ( .a(n7638), .b(n6869), .o(n9778_1) );
oa12f01 g3049 ( .a(n9778_1), .b(n6869), .c(n9777), .o(n4544) );
na02f01 g3050 ( .a(n7591_1), .b(_net_6165), .o(n9780) );
na02f01 g3051 ( .a(n7596_1), .b(n7575), .o(n9781) );
na02f01 g3052 ( .a(n9781), .b(n9780), .o(n4553) );
in01f01 g3053 ( .a(_net_7475), .o(n9783_1) );
na02f01 g3054 ( .a(n6866), .b(net_7395), .o(n9784) );
ao22f01 g3055 ( .a(net_358), .b(_net_280), .c(_net_281), .d(net_356), .o(n9785) );
na02f01 g3056 ( .a(n9785), .b(n9784), .o(n9786) );
na02f01 g3057 ( .a(n9786), .b(n6869), .o(n9787_1) );
oa12f01 g3058 ( .a(n9787_1), .b(n6869), .c(n9783_1), .o(n4572) );
in01f01 g3059 ( .a(_net_6296), .o(n9789) );
no02f01 g3060 ( .a(_net_392), .b(n9789), .o(n4586) );
ao12f01 g3061 ( .a(n9107), .b(_net_7232), .c(net_7231), .o(n9791) );
no03f01 g3062 ( .a(_net_7233), .b(n9116), .c(n9113), .o(n9792_1) );
no02f01 g3063 ( .a(n9792_1), .b(n9791), .o(n9793) );
oa22f01 g3064 ( .a(n9793), .b(n9568), .c(n9572), .d(n9107), .o(n4591) );
in01f01 g3065 ( .a(_net_7413), .o(n9795) );
na02f01 g3066 ( .a(n8633), .b(n7550), .o(n9796_1) );
oa12f01 g3067 ( .a(n9796_1), .b(n7550), .c(n9795), .o(n4596) );
in01f01 g3068 ( .a(_net_7586), .o(n9798) );
na02f01 g3069 ( .a(n8000), .b(n6968), .o(n9799) );
oa12f01 g3070 ( .a(n9799), .b(n6968), .c(n9798), .o(n4609) );
in01f01 g3071 ( .a(_net_7346), .o(n9801_1) );
na02f01 g3072 ( .a(n8731), .b(n7030), .o(n9802) );
oa12f01 g3073 ( .a(n9802), .b(n7030), .c(n9801_1), .o(n4627) );
ao22f01 g3074 ( .a(n6736_1), .b(net_7639), .c(n6734), .d(net_7607), .o(n9804) );
ao22f01 g3075 ( .a(n6739), .b(net_7671), .c(n6738), .d(_net_7575), .o(n9805_1) );
na02f01 g3076 ( .a(n9805_1), .b(n9804), .o(n4636) );
na02f01 g3077 ( .a(n8034), .b(_net_6064), .o(n9807) );
ao22f01 g3078 ( .a(n6777), .b(net_6424), .c(n6776), .d(net_6488), .o(n9808) );
ao22f01 g3079 ( .a(n6780), .b(net_6456), .c(n6779_1), .d(net_6520), .o(n9809_1) );
na02f01 g3080 ( .a(n9809_1), .b(n9808), .o(n9810) );
na02f01 g3081 ( .a(n9810), .b(n8028_1), .o(n9811) );
na02f01 g3082 ( .a(n9811), .b(n9807), .o(n4641) );
in01f01 g3083 ( .a(_net_7269), .o(n9813) );
na02f01 g3084 ( .a(n9685), .b(n6901), .o(n9814_1) );
oa12f01 g3085 ( .a(n9814_1), .b(n6901), .c(n9813), .o(n4646) );
in01f01 g3086 ( .a(_net_7288), .o(n9816) );
na02f01 g3087 ( .a(n8208), .b(n7180), .o(n9817) );
oa12f01 g3088 ( .a(n9817), .b(n7180), .c(n9816), .o(n4656) );
na03f01 g3089 ( .a(n8089), .b(_net_6407), .c(n9258_1), .o(n9819_1) );
no04f01 g3090 ( .a(n9819_1), .b(n9672), .c(n8084), .d(_net_6408), .o(n4673) );
ao22f01 g3091 ( .a(n7288_1), .b(_net_6030), .c(n7286), .d(_net_269), .o(n9821) );
ao22f01 g3092 ( .a(n7298), .b(_net_7722), .c(n7291), .d(_net_7693), .o(n9822) );
na02f01 g3093 ( .a(n7302_1), .b(_net_116), .o(n9823) );
na03f01 g3094 ( .a(n7308), .b(net_195), .c(x1322), .o(n9824_1) );
na02f01 g3095 ( .a(n7296), .b(net_232), .o(n9825) );
na03f01 g3096 ( .a(n7308), .b(net_158), .c(n6800), .o(n9826) );
na03f01 g3097 ( .a(n9826), .b(n9825), .c(n9824_1), .o(n9827) );
ao12f01 g3098 ( .a(n9827), .b(n7306), .c(_net_5986), .o(n9828_1) );
na04f01 g3099 ( .a(n9828_1), .b(n9823), .c(n9822), .d(n9821), .o(n4678) );
no02f01 g3100 ( .a(n7232), .b(n7159), .o(n4703) );
ao22f01 g3101 ( .a(n6777), .b(net_6429), .c(n6776), .d(net_6493), .o(n9831) );
ao22f01 g3102 ( .a(n6780), .b(net_6461), .c(n6779_1), .d(net_6525), .o(n9832) );
ao12f01 g3103 ( .a(n6764), .b(n9832), .c(n9831), .o(n9833_1) );
no02f01 g3104 ( .a(n9181), .b(n6766), .o(n9834) );
in01f01 g3105 ( .a(_net_6073), .o(n9835) );
oa22f01 g3106 ( .a(n7964), .b(n6775), .c(n6784), .d(n9835), .o(n9836) );
no03f01 g3107 ( .a(n9836), .b(n9834), .c(n9833_1), .o(n9837_1) );
in01f01 g3108 ( .a(net_6477), .o(n9838) );
in01f01 g3109 ( .a(net_6445), .o(n9839) );
oa22f01 g3110 ( .a(n6790), .b(n9839), .c(n6789), .d(n9838), .o(n9840_1) );
in01f01 g3111 ( .a(net_6541), .o(n9841) );
in01f01 g3112 ( .a(net_6509), .o(n9842) );
oa22f01 g3113 ( .a(n6795), .b(n9841), .c(n6794), .d(n9842), .o(n9843) );
no02f01 g3114 ( .a(n9843), .b(n9840_1), .o(n9844_1) );
na02f01 g3115 ( .a(n9844_1), .b(n9837_1), .o(n4708) );
in01f01 g3116 ( .a(_net_7692), .o(n9846) );
na02f01 g3117 ( .a(n7207_1), .b(_net_7794), .o(n9847) );
oa12f01 g3118 ( .a(n9847), .b(n7207_1), .c(n9846), .o(n4727) );
in01f01 g3119 ( .a(_net_7286), .o(n9849_1) );
na02f01 g3120 ( .a(n8960), .b(n7180), .o(n9850) );
oa12f01 g3121 ( .a(n9850), .b(n7180), .c(n9849_1), .o(n4732) );
no03f01 g3122 ( .a(n6898), .b(n9592_1), .c(n8094), .o(n9852) );
na02f01 g3123 ( .a(n9852), .b(n7026), .o(n9853_1) );
in01f01 g3124 ( .a(_net_7381), .o(n9854) );
no02f01 g3125 ( .a(n9854), .b(_net_7382), .o(n9855) );
no02f01 g3126 ( .a(_net_7381), .b(n7026), .o(n9856) );
na02f01 g3127 ( .a(n6897), .b(_net_267), .o(n9857) );
no02f01 g3128 ( .a(n9857), .b(n6899_1), .o(n9858_1) );
oa12f01 g3129 ( .a(n9858_1), .b(n9856), .c(n9855), .o(n9859) );
no02f01 g3130 ( .a(n6897), .b(n8094), .o(n9860) );
na02f01 g3131 ( .a(n9860), .b(_net_7382), .o(n9861) );
na03f01 g3132 ( .a(n9861), .b(n9859), .c(n9853_1), .o(n4737) );
in01f01 g3133 ( .a(_net_7706), .o(n9863_1) );
na02f01 g3134 ( .a(n7207_1), .b(_net_7808), .o(n9864) );
oa12f01 g3135 ( .a(n9864), .b(n7207_1), .c(n9863_1), .o(n4760) );
in01f01 g3136 ( .a(_net_7559), .o(n9866) );
na02f01 g3137 ( .a(n9493), .b(n7519), .o(n9867_1) );
oa12f01 g3138 ( .a(n9867_1), .b(n7519), .c(n9866), .o(n4787) );
in01f01 g3139 ( .a(_net_7452), .o(n9869) );
in01f01 g3140 ( .a(net_365), .o(n9870) );
in01f01 g3141 ( .a(net_353), .o(n9871_1) );
oa22f01 g3142 ( .a(n6867_1), .b(n9871_1), .c(n8192_1), .d(n9870), .o(n9872) );
na02f01 g3143 ( .a(n9872), .b(n7197), .o(n9873) );
oa12f01 g3144 ( .a(n9873), .b(n7197), .c(n9869), .o(n4800) );
in01f01 g3145 ( .a(_net_7655), .o(n9875_1) );
na02f01 g3146 ( .a(n9493), .b(n7446_1), .o(n9876) );
oa12f01 g3147 ( .a(n9876), .b(n7446_1), .c(n9875_1), .o(n4809) );
in01f01 g3148 ( .a(_net_7624), .o(n9878) );
na02f01 g3149 ( .a(n6965), .b(net_7544), .o(n9879) );
ao22f01 g3150 ( .a(net_374), .b(_net_292), .c(_net_291), .d(net_376), .o(n9880_1) );
na02f01 g3151 ( .a(n9880_1), .b(n9879), .o(n9881) );
na02f01 g3152 ( .a(n9881), .b(n7400_1), .o(n9882) );
oa12f01 g3153 ( .a(n9882), .b(n7400_1), .c(n9878), .o(n4818) );
na02f01 g3154 ( .a(n7306), .b(_net_6019), .o(n9884) );
na02f01 g3155 ( .a(n7293), .b(net_219), .o(n9885_1) );
ao22f01 g3156 ( .a(n7297_1), .b(net_182), .c(n7296), .d(net_256), .o(n9886) );
ao22f01 g3157 ( .a(n7298), .b(_net_7746), .c(n7291), .d(_net_7717), .o(n9887) );
na04f01 g3158 ( .a(n9887), .b(n9886), .c(n9885_1), .d(n9884), .o(n4831) );
in01f01 g3159 ( .a(_net_6019), .o(n9889_1) );
na02f01 g3160 ( .a(n7348), .b(_net_7819), .o(n9890) );
oa12f01 g3161 ( .a(n9890), .b(n7348), .c(n9889_1), .o(n4843) );
in01f01 g3162 ( .a(n6802), .o(n9892) );
na03f01 g3163 ( .a(n8316_1), .b(n7281), .c(x1322), .o(n9893) );
no02f01 g3164 ( .a(n9893), .b(n9892), .o(n4857) );
in01f01 g3165 ( .a(_net_284), .o(n9895) );
na02f01 g3166 ( .a(n7440), .b(net_7807), .o(n9896) );
oa12f01 g3167 ( .a(n9896), .b(n7440), .c(n9895), .o(n4872) );
ao12f01 g3168 ( .a(x38), .b(n9259), .c(_net_6406), .o(n9898) );
oa12f01 g3169 ( .a(n9898), .b(n9259), .c(_net_6406), .o(n4877) );
ao22f01 g3170 ( .a(n7225), .b(_net_7410), .c(n7224), .d(_net_7442), .o(n9900) );
ao22f01 g3171 ( .a(n7229), .b(_net_7506), .c(n7228), .d(_net_7474), .o(n9901) );
na02f01 g3172 ( .a(n9901), .b(n9900), .o(n4886) );
no02f01 g3173 ( .a(n9893), .b(n8315), .o(n4908) );
na02f01 g3174 ( .a(n7348), .b(_net_7814), .o(n9904) );
oa12f01 g3175 ( .a(n9904), .b(n7348), .c(n7265_1), .o(n4917) );
no02f01 g3176 ( .a(n7125_1), .b(net_6826), .o(n9906) );
no02f01 g3177 ( .a(n9906), .b(n8323), .o(n9907_1) );
no04f01 g3178 ( .a(n8322), .b(n8321), .c(n7125_1), .d(net_6826), .o(n9908) );
oa12f01 g3179 ( .a(n8326), .b(n9908), .c(n9907_1), .o(n9909) );
no02f01 g3180 ( .a(n9908), .b(n9907_1), .o(n9910) );
na02f01 g3181 ( .a(n9910), .b(n2948), .o(n9911_1) );
na02f01 g3182 ( .a(n9911_1), .b(n9909), .o(n4922) );
na02f01 g3183 ( .a(n9311), .b(n9305), .o(n9913) );
no02f01 g3184 ( .a(n9308), .b(n9307_1), .o(n9914_1) );
in01f01 g3185 ( .a(n9914_1), .o(n9915) );
na02f01 g3186 ( .a(n9915), .b(n9309), .o(n9916) );
oa22f01 g3187 ( .a(n9916), .b(n9913), .c(n9313), .d(n9308), .o(n4927) );
in01f01 g3188 ( .a(_net_7659), .o(n9918_1) );
na02f01 g3189 ( .a(n7446_1), .b(n6971), .o(n9919) );
oa12f01 g3190 ( .a(n9919), .b(n7446_1), .c(n9918_1), .o(n4936) );
in01f01 g3191 ( .a(_net_295), .o(n9921) );
na02f01 g3192 ( .a(n7440), .b(_net_7815), .o(n9922) );
oa12f01 g3193 ( .a(n9922), .b(n7440), .c(n9921), .o(n4952) );
in01f01 g3194 ( .a(_net_7651), .o(n9924) );
na02f01 g3195 ( .a(n9154), .b(n7446_1), .o(n9925) );
oa12f01 g3196 ( .a(n9925), .b(n7446_1), .c(n9924), .o(n4961) );
no02f01 g3197 ( .a(n8060), .b(n7012), .o(n9927) );
in01f01 g3198 ( .a(net_6977), .o(n9928) );
in01f01 g3199 ( .a(net_7041), .o(n9929) );
oa22f01 g3200 ( .a(n6987), .b(n9928), .c(n6985), .d(n9929), .o(n9930_1) );
in01f01 g3201 ( .a(net_7073), .o(n9931) );
in01f01 g3202 ( .a(net_7009), .o(n9932) );
oa22f01 g3203 ( .a(n6992), .b(n9932), .c(n6991), .d(n9931), .o(n9933) );
no02f01 g3204 ( .a(n9933), .b(n9930_1), .o(n9934) );
no02f01 g3205 ( .a(n9934), .b(n6980), .o(n9935_1) );
in01f01 g3206 ( .a(_net_6157), .o(n9936) );
oa22f01 g3207 ( .a(n8069), .b(n6997), .c(n6995_1), .d(n9936), .o(n9937) );
no03f01 g3208 ( .a(n9937), .b(n9935_1), .c(n9927), .o(n9938) );
in01f01 g3209 ( .a(net_6989), .o(n9939_1) );
in01f01 g3210 ( .a(net_7021), .o(n9940) );
oa22f01 g3211 ( .a(n8075_1), .b(n9939_1), .c(n8074), .d(n9940), .o(n9941) );
in01f01 g3212 ( .a(net_7085), .o(n9942) );
in01f01 g3213 ( .a(net_7053), .o(n9943) );
oa22f01 g3214 ( .a(n8080_1), .b(n9942), .c(n8079), .d(n9943), .o(n9944_1) );
no02f01 g3215 ( .a(n9944_1), .b(n9941), .o(n9945) );
na02f01 g3216 ( .a(n9945), .b(n9938), .o(n4974) );
in01f01 g3217 ( .a(_net_7571), .o(n9947) );
na02f01 g3218 ( .a(n7519), .b(n7144), .o(n9948) );
oa12f01 g3219 ( .a(n9948), .b(n7519), .c(n9947), .o(n4987) );
in01f01 g3220 ( .a(_net_6029), .o(n9950) );
no02f01 g3221 ( .a(n7287), .b(n9950), .o(n9951) );
in01f01 g3222 ( .a(_net_7721), .o(n9952) );
no04f01 g3223 ( .a(n9705), .b(n7293), .c(n7292_1), .d(n9952), .o(n9953_1) );
na02f01 g3224 ( .a(x38), .b(n7300), .o(n9954) );
no02f01 g3225 ( .a(n9954), .b(n7301), .o(n9955) );
no03f01 g3226 ( .a(n9955), .b(n9953_1), .c(n9951), .o(n9956) );
na02f01 g3227 ( .a(n7302_1), .b(_net_115), .o(n9957_1) );
in01f01 g3228 ( .a(net_157), .o(n9958) );
no04f01 g3229 ( .a(n7307_1), .b(n7292_1), .c(n9958), .d(x1322), .o(n9959) );
in01f01 g3230 ( .a(net_231), .o(n9960) );
no03f01 g3231 ( .a(n7295), .b(n7294), .c(n9960), .o(n9961_1) );
in01f01 g3232 ( .a(net_194), .o(n9962) );
no04f01 g3233 ( .a(n7307_1), .b(n7292_1), .c(n9962), .d(n6800), .o(n9963) );
no03f01 g3234 ( .a(n9963), .b(n9961_1), .c(n9959), .o(n9964) );
oa12f01 g3235 ( .a(n9964), .b(n7305), .c(n7980_1), .o(n9965) );
in01f01 g3236 ( .a(_net_268), .o(n9966_1) );
oa22f01 g3237 ( .a(n7290), .b(n9846), .c(n7285), .d(n9966_1), .o(n9967) );
no02f01 g3238 ( .a(n9967), .b(n9965), .o(n9968) );
na03f01 g3239 ( .a(n9968), .b(n9957_1), .c(n9956), .o(n4992) );
in01f01 g3240 ( .a(_net_7727), .o(n9970) );
in01f01 g3241 ( .a(_net_6005), .o(n9971_1) );
ao12f01 g3242 ( .a(n7343), .b(n9971_1), .c(n9970), .o(n5013) );
in01f01 g3243 ( .a(_net_6693), .o(n9973) );
in01f01 g3244 ( .a(n513), .o(n9974) );
ao12f01 g3245 ( .a(n9973), .b(_net_6692), .c(net_6691), .o(n9975) );
no03f01 g3246 ( .a(n7663), .b(_net_6693), .c(n7153), .o(n9976_1) );
no02f01 g3247 ( .a(n9976_1), .b(n9975), .o(n9977) );
na02f01 g3248 ( .a(_net_5995), .b(n7067_1), .o(n9978) );
oa22f01 g3249 ( .a(n9978), .b(n9973), .c(n9977), .d(n9974), .o(n5018) );
in01f01 g3250 ( .a(net_355), .o(n9980) );
no02f01 g3251 ( .a(n6867_1), .b(n9980), .o(n5027) );
in01f01 g3252 ( .a(net_7799), .o(n9982) );
na02f01 g3253 ( .a(n6803), .b(_net_6034), .o(n9983) );
oa12f01 g3254 ( .a(n9983), .b(n6803), .c(n9982), .o(n5040) );
in01f01 g3255 ( .a(_net_7507), .o(n9985_1) );
na02f01 g3256 ( .a(n9786), .b(n7626_1), .o(n9986) );
oa12f01 g3257 ( .a(n9986), .b(n7626_1), .c(n9985_1), .o(n5061) );
in01f01 g3258 ( .a(_net_7508), .o(n9988_1) );
na02f01 g3259 ( .a(n7626_1), .b(n7553_1), .o(n9989) );
oa12f01 g3260 ( .a(n9989), .b(n7626_1), .c(n9988_1), .o(n5075) );
in01f01 g3261 ( .a(_net_7514), .o(n9991) );
na02f01 g3262 ( .a(n9487_1), .b(n7626_1), .o(n9992_1) );
oa12f01 g3263 ( .a(n9992_1), .b(n7626_1), .c(n9991), .o(n5080) );
in01f01 g3264 ( .a(net_7758), .o(n9994) );
na04f01 g3265 ( .a(_net_6028), .b(_net_7791), .c(net_303), .d(n9994), .o(n9995) );
ao12f01 g3266 ( .a(n9995), .b(net_305), .c(_net_6029), .o(n5085) );
in01f01 g3267 ( .a(_net_7433), .o(n9997_1) );
na02f01 g3268 ( .a(n7779_1), .b(n7197), .o(n9998) );
oa12f01 g3269 ( .a(n9998), .b(n7197), .c(n9997_1), .o(n5094) );
na02f01 g3270 ( .a(n7298), .b(net_7739), .o(n10000) );
ao22f01 g3271 ( .a(n7306), .b(_net_6009), .c(n7291), .d(net_7710), .o(n10001_1) );
na02f01 g3272 ( .a(n7302_1), .b(net_149), .o(n10002) );
na02f01 g3273 ( .a(n7296), .b(net_249), .o(n10003) );
na03f01 g3274 ( .a(n7308), .b(_net_175), .c(n6800), .o(n10004) );
na03f01 g3275 ( .a(n7308), .b(_net_212), .c(x1322), .o(n10005) );
na03f01 g3276 ( .a(n10005), .b(n10004), .c(n10003), .o(n10006_1) );
ao12f01 g3277 ( .a(n10006_1), .b(n7286), .c(_net_292), .o(n10007) );
na04f01 g3278 ( .a(n10007), .b(n10002), .c(n10001_1), .d(n10000), .o(n5103) );
ao22f01 g3279 ( .a(n7225), .b(_net_7416), .c(n7224), .d(_net_7448), .o(n10009) );
ao22f01 g3280 ( .a(n7229), .b(_net_7512), .c(n7228), .d(_net_7480), .o(n10010_1) );
na02f01 g3281 ( .a(n10010_1), .b(n10009), .o(n5107) );
in01f01 g3282 ( .a(_net_6415), .o(n10012) );
na02f01 g3283 ( .a(n7357), .b(net_6417), .o(n10013) );
na02f01 g3284 ( .a(n9305), .b(net_6417), .o(n10014_1) );
in01f01 g3285 ( .a(net_6412), .o(n10015) );
in01f01 g3286 ( .a(_net_6413), .o(n10016) );
no02f01 g3287 ( .a(n10016), .b(n10015), .o(n10017) );
na03f01 g3288 ( .a(n10017), .b(_net_6414), .c(_net_6415), .o(n10018) );
in01f01 g3289 ( .a(_net_6414), .o(n10019_1) );
in01f01 g3290 ( .a(n10017), .o(n10020) );
oa12f01 g3291 ( .a(n10012), .b(n10020), .c(n10019_1), .o(n10021) );
na02f01 g3292 ( .a(n10021), .b(n10018), .o(n10022) );
oa22f01 g3293 ( .a(n10022), .b(n10014_1), .c(n10013), .d(n10012), .o(n5112) );
na02f01 g3294 ( .a(n7339), .b(x1231), .o(n10024) );
no04f01 g3295 ( .a(n10024), .b(n7292_1), .c(x1215), .d(n6800), .o(n5117) );
no02f01 g3296 ( .a(n7339), .b(n7112), .o(n10026) );
no03f01 g3297 ( .a(n10026), .b(n7336), .c(x149), .o(n5130) );
ao22f01 g3298 ( .a(n7225), .b(_net_7426), .c(n7224), .d(net_7458), .o(n10028_1) );
ao22f01 g3299 ( .a(n7229), .b(net_7522), .c(n7228), .d(net_7490), .o(n10029) );
na02f01 g3300 ( .a(n10029), .b(n10028_1), .o(n5134) );
in01f01 g3301 ( .a(_net_7272), .o(n10031) );
na02f01 g3302 ( .a(n2913), .b(n6901), .o(n10032_1) );
oa12f01 g3303 ( .a(n10032_1), .b(n6901), .c(n10031), .o(n5143) );
in01f01 g3304 ( .a(_net_271), .o(n10034) );
na02f01 g3305 ( .a(n7440), .b(_net_7797), .o(n10035) );
oa12f01 g3306 ( .a(n10035), .b(n7440), .c(n10034), .o(n5164) );
in01f01 g3307 ( .a(_net_7435), .o(n10037_1) );
na02f01 g3308 ( .a(n9700_1), .b(n7197), .o(n10038) );
oa12f01 g3309 ( .a(n10038), .b(n7197), .c(n10037_1), .o(n5169) );
na02f01 g3310 ( .a(n6933), .b(_net_6084), .o(n10040) );
na02f01 g3311 ( .a(n6942), .b(n6917), .o(n10041) );
na02f01 g3312 ( .a(n10041), .b(n10040), .o(n5198) );
no03f01 g3313 ( .a(n6965), .b(n7654_1), .c(n8236), .o(n10043) );
na02f01 g3314 ( .a(n7444), .b(_net_7686), .o(n10044) );
na02f01 g3315 ( .a(n7445), .b(n8348), .o(n10045) );
na03f01 g3316 ( .a(n10045), .b(n10044), .c(n10043), .o(n10046) );
no02f01 g3317 ( .a(n8232_1), .b(n6966), .o(n10047_1) );
na03f01 g3318 ( .a(_net_7685), .b(_net_7684), .c(_net_7683), .o(n10048) );
na02f01 g3319 ( .a(n10048), .b(n8348), .o(n10049) );
in01f01 g3320 ( .a(n10048), .o(n10050) );
na02f01 g3321 ( .a(n10050), .b(_net_7686), .o(n10051) );
na03f01 g3322 ( .a(n10051), .b(n10049), .c(n10047_1), .o(n10052_1) );
na02f01 g3323 ( .a(n8237_1), .b(_net_7686), .o(n10053) );
na03f01 g3324 ( .a(n10053), .b(n10052_1), .c(n10046), .o(n5207) );
no02f01 g3325 ( .a(n9502_1), .b(n7468_1), .o(n10055) );
no02f01 g3326 ( .a(n9467_1), .b(n7470), .o(n10056_1) );
in01f01 g3327 ( .a(_net_6114), .o(n10057) );
oa22f01 g3328 ( .a(n8557_1), .b(n7123), .c(n7118), .d(n10057), .o(n10058) );
no03f01 g3329 ( .a(n10058), .b(n10056_1), .c(n10055), .o(n10059) );
in01f01 g3330 ( .a(net_6716), .o(n10060) );
in01f01 g3331 ( .a(net_6748), .o(n10061_1) );
oa22f01 g3332 ( .a(n7492_1), .b(n10060), .c(n7491), .d(n10061_1), .o(n10062) );
in01f01 g3333 ( .a(net_6812), .o(n10063) );
in01f01 g3334 ( .a(net_6780), .o(n10064) );
oa22f01 g3335 ( .a(n7497), .b(n10063), .c(n7496_1), .d(n10064), .o(n10065) );
no02f01 g3336 ( .a(n10065), .b(n10062), .o(n10066_1) );
na02f01 g3337 ( .a(n10066_1), .b(n10059), .o(n5212) );
in01f01 g3338 ( .a(_net_7593), .o(n10068) );
na02f01 g3339 ( .a(n6965), .b(net_7545), .o(n10069) );
ao22f01 g3340 ( .a(_net_292), .b(net_375), .c(_net_291), .d(net_377), .o(n10070_1) );
na02f01 g3341 ( .a(n10070_1), .b(n10069), .o(n10071) );
na02f01 g3342 ( .a(n10071), .b(n6968), .o(n10072) );
oa12f01 g3343 ( .a(n10072), .b(n6968), .c(n10068), .o(n5225) );
in01f01 g3344 ( .a(_net_7422), .o(n10074_1) );
na02f01 g3345 ( .a(n5027), .b(n7550), .o(n10075) );
oa12f01 g3346 ( .a(n10075), .b(n7550), .c(n10074_1), .o(n5230) );
in01f01 g3347 ( .a(_net_7297), .o(n10077) );
na02f01 g3348 ( .a(n9537_1), .b(n7180), .o(n10078) );
oa12f01 g3349 ( .a(n10078), .b(n7180), .c(n10077), .o(n5251) );
in01f01 g3350 ( .a(_net_7567), .o(n10080) );
na02f01 g3351 ( .a(n8639), .b(n7519), .o(n10081) );
oa12f01 g3352 ( .a(n10081), .b(n7519), .c(n10080), .o(n5256) );
in01f01 g3353 ( .a(_net_7416), .o(n10083) );
na02f01 g3354 ( .a(n7638), .b(n7550), .o(n10084_1) );
oa12f01 g3355 ( .a(n10084_1), .b(n7550), .c(n10083), .o(n5265) );
in01f01 g3356 ( .a(_net_7292), .o(n10086) );
na02f01 g3357 ( .a(n6898), .b(net_7244), .o(n10087) );
ao22f01 g3358 ( .a(net_338), .b(_net_269), .c(_net_270), .d(net_336), .o(n10088) );
na02f01 g3359 ( .a(n10088), .b(n10087), .o(n10089_1) );
na02f01 g3360 ( .a(n10089_1), .b(n7180), .o(n10090) );
oa12f01 g3361 ( .a(n10090), .b(n7180), .c(n10086), .o(n5274) );
in01f01 g3362 ( .a(net_6025), .o(n10092) );
in01f01 g3363 ( .a(_net_7731), .o(n10093) );
ao12f01 g3364 ( .a(n7343), .b(n10093), .c(n10092), .o(n5279) );
in01f01 g3365 ( .a(_net_6283), .o(n10095) );
no02f01 g3366 ( .a(_net_392), .b(n10095), .o(n5284) );
in01f01 g3367 ( .a(_net_7599), .o(n10097) );
na02f01 g3368 ( .a(n8639), .b(n6968), .o(n10098) );
oa12f01 g3369 ( .a(n10098), .b(n6968), .c(n10097), .o(n5293) );
in01f01 g3370 ( .a(_net_7411), .o(n10100) );
na02f01 g3371 ( .a(n9786), .b(n7550), .o(n10101) );
oa12f01 g3372 ( .a(n10101), .b(n7550), .c(n10100), .o(n5307) );
in01f01 g3373 ( .a(net_7750), .o(n10103_1) );
na04f01 g3374 ( .a(_net_7791), .b(net_303), .c(_net_5984), .d(n10103_1), .o(n10104) );
ao12f01 g3375 ( .a(n10104), .b(net_309), .c(_net_5985), .o(n5316) );
na02f01 g3376 ( .a(n10043), .b(n6959), .o(n10106) );
no02f01 g3377 ( .a(_net_7684), .b(n8231), .o(n10107_1) );
no02f01 g3378 ( .a(n6959), .b(_net_7683), .o(n10108) );
oa12f01 g3379 ( .a(n10047_1), .b(n10108), .c(n10107_1), .o(n10109) );
na02f01 g3380 ( .a(n8237_1), .b(_net_7684), .o(n10110) );
na03f01 g3381 ( .a(n10110), .b(n10109), .c(n10106), .o(n5321) );
in01f01 g3382 ( .a(_net_7662), .o(n10112_1) );
na02f01 g3383 ( .a(n9373_1), .b(n7446_1), .o(n10113) );
oa12f01 g3384 ( .a(n10113), .b(n7446_1), .c(n10112_1), .o(n5330) );
in01f01 g3385 ( .a(_net_6420), .o(n10115) );
na02f01 g3386 ( .a(n9412), .b(n10115), .o(n10116_1) );
na02f01 g3387 ( .a(n10116_1), .b(n9664_1), .o(n10117) );
oa22f01 g3388 ( .a(n10117), .b(n9411), .c(n9409), .d(n10115), .o(n5344) );
in01f01 g3389 ( .a(_net_7280), .o(n10119) );
na02f01 g3390 ( .a(n875), .b(n6901), .o(n10120_1) );
oa12f01 g3391 ( .a(n10120_1), .b(n6901), .c(n10119), .o(n5353) );
in01f01 g3392 ( .a(_net_7657), .o(n10122) );
na02f01 g3393 ( .a(n10071), .b(n7446_1), .o(n10123) );
oa12f01 g3394 ( .a(n10123), .b(n7446_1), .c(n10122), .o(n5370) );
no02f01 g3395 ( .a(n9292), .b(n6945), .o(n10125) );
in01f01 g3396 ( .a(net_6633), .o(n10126) );
in01f01 g3397 ( .a(net_6569), .o(n10127) );
oa22f01 g3398 ( .a(n6922), .b(n10127), .c(n6919_1), .d(n10126), .o(n10128_1) );
in01f01 g3399 ( .a(net_6665), .o(n10129) );
in01f01 g3400 ( .a(net_6601), .o(n10130) );
oa22f01 g3401 ( .a(n6927), .b(n10130), .c(n6925), .d(n10129), .o(n10131) );
no02f01 g3402 ( .a(n10131), .b(n10128_1), .o(n10132_1) );
no02f01 g3403 ( .a(n10132_1), .b(n6934_1), .o(n10133) );
in01f01 g3404 ( .a(_net_6096), .o(n10134) );
oa22f01 g3405 ( .a(n7042), .b(n6916), .c(n6932), .d(n10134), .o(n10135) );
no03f01 g3406 ( .a(n10135), .b(n10133), .c(n10125), .o(n10136) );
in01f01 g3407 ( .a(net_6583), .o(n10137_1) );
in01f01 g3408 ( .a(net_6615), .o(n10138) );
oa22f01 g3409 ( .a(n7058_1), .b(n10137_1), .c(n7057), .d(n10138), .o(n10139) );
in01f01 g3410 ( .a(net_6679), .o(n10140) );
in01f01 g3411 ( .a(net_6647), .o(n10141_1) );
oa22f01 g3412 ( .a(n7063), .b(n10140), .c(n7062_1), .d(n10141_1), .o(n10142) );
no02f01 g3413 ( .a(n10142), .b(n10139), .o(n10143) );
na02f01 g3414 ( .a(n10143), .b(n10136), .o(n5388) );
ao22f01 g3415 ( .a(n6877), .b(_net_7253), .c(n6876_1), .d(_net_7317), .o(n10145_1) );
ao22f01 g3416 ( .a(n6881_1), .b(_net_7285), .c(n6880), .d(_net_7349), .o(n10146) );
na02f01 g3417 ( .a(n10146), .b(n10145_1), .o(n5397) );
in01f01 g3418 ( .a(_net_7429), .o(n10148) );
na02f01 g3419 ( .a(n7550), .b(n420), .o(n10149) );
oa12f01 g3420 ( .a(n10149), .b(n7550), .c(n10148), .o(n5406) );
in01f01 g3421 ( .a(_net_7631), .o(n10151) );
na02f01 g3422 ( .a(n8639), .b(n7400_1), .o(n10152) );
oa12f01 g3423 ( .a(n10152), .b(n7400_1), .c(n10151), .o(n5411) );
in01f01 g3424 ( .a(_net_7295), .o(n10154_1) );
na02f01 g3425 ( .a(n7994_1), .b(n7180), .o(n10155) );
oa12f01 g3426 ( .a(n10155), .b(n7180), .c(n10154_1), .o(n5420) );
in01f01 g3427 ( .a(_net_7795), .o(n10157) );
na02f01 g3428 ( .a(n6803), .b(_net_6030), .o(n10158_1) );
oa12f01 g3429 ( .a(n10158_1), .b(n6803), .c(n10157), .o(n5429) );
in01f01 g3430 ( .a(_net_119), .o(n10160) );
na02f01 g3431 ( .a(net_315), .b(_net_154), .o(n10161) );
oa12f01 g3432 ( .a(n10161), .b(n10160), .c(_net_154), .o(n5446) );
in01f01 g3433 ( .a(_net_5987), .o(n10163) );
na02f01 g3434 ( .a(n7348), .b(_net_7796), .o(n10164) );
oa12f01 g3435 ( .a(n10164), .b(n7348), .c(n10163), .o(n5455) );
in01f01 g3436 ( .a(_net_7587), .o(n10166) );
na02f01 g3437 ( .a(n9154), .b(n6968), .o(n10167) );
oa12f01 g3438 ( .a(n10167), .b(n6968), .c(n10166), .o(n5477) );
in01f01 g3439 ( .a(_net_7513), .o(n10169) );
na02f01 g3440 ( .a(n7626_1), .b(n6872_1), .o(n10170) );
oa12f01 g3441 ( .a(n10170), .b(n7626_1), .c(n10169), .o(n5490) );
na02f01 g3442 ( .a(n7440), .b(_net_7796), .o(n10172) );
oa12f01 g3443 ( .a(n10172), .b(n7440), .c(n7253), .o(n5495) );
in01f01 g3444 ( .a(_net_7467), .o(n10174) );
na02f01 g3445 ( .a(n9700_1), .b(n6869), .o(n10175) );
oa12f01 g3446 ( .a(n10175), .b(n6869), .c(n10174), .o(n5508) );
na02f01 g3447 ( .a(n7298), .b(net_7738), .o(n10177) );
ao22f01 g3448 ( .a(n7306), .b(_net_6008), .c(n7291), .d(net_7709), .o(n10178) );
na02f01 g3449 ( .a(n7302_1), .b(net_148), .o(n10179) );
na02f01 g3450 ( .a(n7296), .b(net_248), .o(n10180) );
na03f01 g3451 ( .a(n7308), .b(_net_174), .c(n6800), .o(n10181) );
na03f01 g3452 ( .a(n7308), .b(_net_211), .c(x1322), .o(n10182) );
na03f01 g3453 ( .a(n10182), .b(n10181), .c(n10180), .o(n10183) );
ao12f01 g3454 ( .a(n10183), .b(n7286), .c(_net_291), .o(n10184) );
na04f01 g3455 ( .a(n10184), .b(n10179), .c(n10178), .d(n10177), .o(n5517) );
na02f01 g3456 ( .a(n7302_1), .b(net_153), .o(n10186) );
na02f01 g3457 ( .a(n7306), .b(net_6024), .o(n10187) );
na02f01 g3458 ( .a(n7296), .b(net_261), .o(n10188) );
ao22f01 g3459 ( .a(n7297_1), .b(net_187), .c(n7293), .d(net_224), .o(n10189) );
na04f01 g3460 ( .a(n10189), .b(n10188), .c(n10187), .d(n10186), .o(n5525) );
in01f01 g3461 ( .a(_net_293), .o(n10191) );
no02f01 g3462 ( .a(n10191), .b(_net_294), .o(n10192) );
na02f01 g3463 ( .a(_net_289), .b(_net_295), .o(n10193) );
ao12f01 g3464 ( .a(n10193), .b(_net_266), .c(n7653), .o(n10194) );
na02f01 g3465 ( .a(n10194), .b(n10192), .o(n10195) );
in01f01 g3466 ( .a(n10193), .o(n10196) );
no02f01 g3467 ( .a(n10191), .b(n9540), .o(n10197) );
na03f01 g3468 ( .a(n10197), .b(n10196), .c(_net_263), .o(n10198) );
na03f01 g3469 ( .a(_net_265), .b(_net_266), .c(n7653), .o(n10199) );
na04f01 g3470 ( .a(n10199), .b(n10196), .c(n10191), .d(n9540), .o(n10200) );
oa12f01 g3471 ( .a(n7653), .b(_net_265), .c(_net_266), .o(n10201) );
na04f01 g3472 ( .a(n10201), .b(n10196), .c(n10191), .d(_net_294), .o(n10202) );
na04f01 g3473 ( .a(n10202), .b(n10200), .c(n10198), .d(n10195), .o(n10203) );
in01f01 g3474 ( .a(n10203), .o(n10204) );
no02f01 g3475 ( .a(n10204), .b(x837), .o(n5529) );
na02f01 g3476 ( .a(n7232), .b(net_7771), .o(n10206) );
no02f01 g3477 ( .a(n10206), .b(n6885), .o(n10207) );
no02f01 g3478 ( .a(n10207), .b(_net_7721), .o(n10208) );
no02f01 g3479 ( .a(n10208), .b(n7343), .o(n5534) );
in01f01 g3480 ( .a(_net_7577), .o(n10210) );
na02f01 g3481 ( .a(n3015), .b(n7519), .o(n10211) );
oa12f01 g3482 ( .a(n10211), .b(n7519), .c(n10210), .o(n5543) );
no02f01 g3483 ( .a(n6867_1), .b(n9870), .o(n5552) );
in01f01 g3484 ( .a(_net_7430), .o(n10214) );
in01f01 g3485 ( .a(net_363), .o(n10215) );
no02f01 g3486 ( .a(n6867_1), .b(n10215), .o(n6437) );
na02f01 g3487 ( .a(n6437), .b(n7550), .o(n10217) );
oa12f01 g3488 ( .a(n10217), .b(n7550), .c(n10214), .o(n5565) );
in01f01 g3489 ( .a(_net_7502), .o(n10219) );
na02f01 g3490 ( .a(n7860), .b(n7626_1), .o(n10220) );
oa12f01 g3491 ( .a(n10220), .b(n7626_1), .c(n10219), .o(n5570) );
in01f01 g3492 ( .a(_net_7622), .o(n10222) );
na02f01 g3493 ( .a(n7644_1), .b(n7400_1), .o(n10223) );
oa12f01 g3494 ( .a(n10223), .b(n7400_1), .c(n10222), .o(n5579) );
no02f01 g3495 ( .a(n8610), .b(n7012), .o(n10225) );
no02f01 g3496 ( .a(n8619), .b(n6997), .o(n10226) );
in01f01 g3497 ( .a(_net_6162), .o(n10227) );
no02f01 g3498 ( .a(n7020), .b(n7017), .o(n10228) );
oa22f01 g3499 ( .a(n10228), .b(n6980), .c(n6995_1), .d(n10227), .o(n10229) );
no03f01 g3500 ( .a(n10229), .b(n10226), .c(n10225), .o(n10230) );
in01f01 g3501 ( .a(net_7026), .o(n10231) );
in01f01 g3502 ( .a(net_6994), .o(n10232) );
oa22f01 g3503 ( .a(n8075_1), .b(n10232), .c(n8074), .d(n10231), .o(n10233) );
in01f01 g3504 ( .a(net_7058), .o(n10234) );
in01f01 g3505 ( .a(net_7090), .o(n10235) );
oa22f01 g3506 ( .a(n8080_1), .b(n10235), .c(n8079), .d(n10234), .o(n10236) );
no02f01 g3507 ( .a(n10236), .b(n10233), .o(n10237) );
na02f01 g3508 ( .a(n10237), .b(n10230), .o(n5596) );
in01f01 g3509 ( .a(_net_7420), .o(n10239) );
na02f01 g3510 ( .a(n9872), .b(n7550), .o(n10240) );
oa12f01 g3511 ( .a(n10240), .b(n7550), .c(n10239), .o(n5601) );
no02f01 g3512 ( .a(n8452), .b(n6824), .o(n10242) );
in01f01 g3513 ( .a(net_6841), .o(n10243) );
in01f01 g3514 ( .a(net_6905), .o(n10244) );
oa22f01 g3515 ( .a(n6810), .b(n10243), .c(n6807), .d(n10244), .o(n10245) );
in01f01 g3516 ( .a(net_6873), .o(n10246) );
in01f01 g3517 ( .a(net_6937), .o(n10247) );
oa22f01 g3518 ( .a(n6815), .b(n10246), .c(n6813_1), .d(n10247), .o(n10248) );
no02f01 g3519 ( .a(n10248), .b(n10245), .o(n10249) );
no02f01 g3520 ( .a(n10249), .b(n6826_1), .o(n10250) );
in01f01 g3521 ( .a(_net_6138), .o(n10251) );
oa22f01 g3522 ( .a(n9127), .b(n6836_1), .c(n6844), .d(n10251), .o(n10252) );
no03f01 g3523 ( .a(n10252), .b(n10250), .c(n10242), .o(n10253) );
in01f01 g3524 ( .a(net_6855), .o(n10254) );
in01f01 g3525 ( .a(net_6887), .o(n10255) );
oa22f01 g3526 ( .a(n6850_1), .b(n10254), .c(n6849), .d(n10255), .o(n10256) );
in01f01 g3527 ( .a(net_6951), .o(n10257) );
in01f01 g3528 ( .a(net_6919), .o(n10258) );
oa22f01 g3529 ( .a(n6855_1), .b(n10257), .c(n6854), .d(n10258), .o(n10259) );
no02f01 g3530 ( .a(n10259), .b(n10256), .o(n10260) );
na02f01 g3531 ( .a(n10260), .b(n10253), .o(n5623) );
in01f01 g3532 ( .a(_net_7736), .o(n10262) );
ao12f01 g3533 ( .a(n7343), .b(n10262), .c(n8875), .o(n5633) );
in01f01 g3534 ( .a(_net_6204), .o(n10264) );
no02f01 g3535 ( .a(_net_392), .b(n10264), .o(n5638) );
in01f01 g3536 ( .a(_net_7634), .o(n10266) );
na02f01 g3537 ( .a(n7892), .b(n7400_1), .o(n10267) );
oa12f01 g3538 ( .a(n10267), .b(n7400_1), .c(n10266), .o(n5643) );
no02f01 g3539 ( .a(n7332), .b(n8803), .o(n5660) );
no02f01 g3540 ( .a(n6880), .b(n9440), .o(n10270) );
no03f01 g3541 ( .a(_net_7380), .b(n6879), .c(n6875), .o(n10271) );
no02f01 g3542 ( .a(n10271), .b(n10270), .o(n10272) );
oa22f01 g3543 ( .a(n10272), .b(n8096), .c(n8097_1), .d(n9440), .o(n5669) );
in01f01 g3544 ( .a(_net_7564), .o(n10274) );
na02f01 g3545 ( .a(n8043), .b(n7519), .o(n10275) );
oa12f01 g3546 ( .a(n10275), .b(n7519), .c(n10274), .o(n5674) );
in01f01 g3547 ( .a(_net_6282), .o(n10277) );
no02f01 g3548 ( .a(n10277), .b(_net_392), .o(n5691) );
ao22f01 g3549 ( .a(n6877), .b(_net_7263), .c(n6876_1), .d(_net_7327), .o(n10279) );
ao22f01 g3550 ( .a(n6881_1), .b(_net_7295), .c(n6880), .d(_net_7359), .o(n10280) );
na02f01 g3551 ( .a(n10280), .b(n10279), .o(n5700) );
in01f01 g3552 ( .a(n10014_1), .o(n5709) );
in01f01 g3553 ( .a(_net_269), .o(n10283) );
na02f01 g3554 ( .a(n7440), .b(_net_7795), .o(n10284) );
oa12f01 g3555 ( .a(n10284), .b(n7440), .c(n10283), .o(n5722) );
in01f01 g3556 ( .a(_net_5998), .o(n10286) );
na02f01 g3557 ( .a(n7348), .b(_net_7804), .o(n10287) );
oa12f01 g3558 ( .a(n10287), .b(n7348), .c(n10286), .o(n5739) );
no02f01 g3559 ( .a(n8711_1), .b(n8713), .o(n10289) );
na02f01 g3560 ( .a(n10289), .b(n9605), .o(n10290) );
no03f01 g3561 ( .a(n7467), .b(n7117), .c(n7121), .o(n10291) );
no02f01 g3562 ( .a(n7132), .b(n9600), .o(n10292) );
no02f01 g3563 ( .a(n7133_1), .b(_net_6825), .o(n10293) );
no02f01 g3564 ( .a(n10293), .b(n10292), .o(n10294) );
ao22f01 g3565 ( .a(n10294), .b(n10291), .c(n8716), .d(_net_6825), .o(n10295) );
na02f01 g3566 ( .a(n10295), .b(n10290), .o(n5748) );
no02f01 g3567 ( .a(n10017), .b(n10019_1), .o(n10297) );
no02f01 g3568 ( .a(n10020), .b(_net_6414), .o(n10298) );
no02f01 g3569 ( .a(n10298), .b(n10297), .o(n10299) );
oa22f01 g3570 ( .a(n10299), .b(n10014_1), .c(n10013), .d(n10019_1), .o(n5753) );
no02f01 g3571 ( .a(n7012), .b(n9626), .o(n10301) );
no02f01 g3572 ( .a(n8782), .b(n6997), .o(n10302) );
in01f01 g3573 ( .a(_net_6154), .o(n10303) );
oa22f01 g3574 ( .a(n8790), .b(n6980), .c(n6995_1), .d(n10303), .o(n10304) );
no03f01 g3575 ( .a(n10304), .b(n10302), .c(n10301), .o(n10305) );
in01f01 g3576 ( .a(net_6986), .o(n10306) );
in01f01 g3577 ( .a(net_7018), .o(n10307) );
oa22f01 g3578 ( .a(n8075_1), .b(n10306), .c(n8074), .d(n10307), .o(n10308) );
in01f01 g3579 ( .a(net_7082), .o(n10309) );
in01f01 g3580 ( .a(net_7050), .o(n10310) );
oa22f01 g3581 ( .a(n8080_1), .b(n10309), .c(n8079), .d(n10310), .o(n10311) );
no02f01 g3582 ( .a(n10311), .b(n10308), .o(n10312) );
na02f01 g3583 ( .a(n10312), .b(n10305), .o(n5775) );
in01f01 g3584 ( .a(_net_7561), .o(n10314) );
na02f01 g3585 ( .a(n10071), .b(n7519), .o(n10315) );
oa12f01 g3586 ( .a(n10315), .b(n7519), .c(n10314), .o(n5809) );
in01f01 g3587 ( .a(net_382), .o(n10317) );
no02f01 g3588 ( .a(n6966), .b(n10317), .o(n5814) );
ao22f01 g3589 ( .a(n6736_1), .b(_net_7633), .c(n6734), .d(_net_7601), .o(n10319) );
ao22f01 g3590 ( .a(n6739), .b(_net_7665), .c(n6738), .d(_net_7569), .o(n10320) );
na02f01 g3591 ( .a(n10320), .b(n10319), .o(n5819) );
ao22f01 g3592 ( .a(n6877), .b(_net_7258), .c(n6876_1), .d(_net_7322), .o(n10322) );
ao22f01 g3593 ( .a(n6881_1), .b(_net_7290), .c(n6880), .d(_net_7354), .o(n10323) );
na02f01 g3594 ( .a(n10323), .b(n10322), .o(n5828) );
ao22f01 g3595 ( .a(n6736_1), .b(net_7645), .c(n6734), .d(net_7613), .o(n10325) );
ao22f01 g3596 ( .a(n6739), .b(net_7677), .c(n6738), .d(_net_7581), .o(n10326) );
na02f01 g3597 ( .a(n10326), .b(n10325), .o(n5845) );
in01f01 g3598 ( .a(_net_7734), .o(n10328) );
in01f01 g3599 ( .a(net_6036), .o(n10329) );
ao12f01 g3600 ( .a(n7343), .b(n10329), .c(n10328), .o(n5850) );
na02f01 g3601 ( .a(n8177), .b(n8086), .o(n10331) );
no03f01 g3602 ( .a(_net_6407), .b(_net_6405), .c(_net_6406), .o(n10332) );
na02f01 g3603 ( .a(n10332), .b(n8088_1), .o(n10333) );
no04f01 g3604 ( .a(_net_6407), .b(_net_6405), .c(_net_6406), .d(_net_6404), .o(n10334) );
ao12f01 g3605 ( .a(n10331), .b(n10334), .c(n10333), .o(n5855) );
no02f01 g3606 ( .a(_net_7232), .b(n7579), .o(n10336) );
no02f01 g3607 ( .a(n9116), .b(_net_7229), .o(n10337) );
no02f01 g3608 ( .a(n10337), .b(n10336), .o(n10338) );
no02f01 g3609 ( .a(n7576), .b(net_7231), .o(n10339) );
no02f01 g3610 ( .a(n10339), .b(n10338), .o(n10340) );
no04f01 g3611 ( .a(n10337), .b(n10336), .c(n7576), .d(net_7231), .o(n10341) );
oa12f01 g3612 ( .a(n9641), .b(n10341), .c(n10340), .o(n10342) );
no02f01 g3613 ( .a(n10341), .b(n10340), .o(n10343) );
na02f01 g3614 ( .a(n10343), .b(n4276), .o(n10344) );
na02f01 g3615 ( .a(n10344), .b(n10342), .o(n5885) );
na02f01 g3616 ( .a(n7440), .b(_net_7806), .o(n10346) );
oa12f01 g3617 ( .a(n10346), .b(n7440), .c(n7415), .o(n5890) );
in01f01 g3618 ( .a(_net_7407), .o(n10348) );
na02f01 g3619 ( .a(n7550), .b(n7387), .o(n10349) );
oa12f01 g3620 ( .a(n10349), .b(n7550), .c(n10348), .o(n5899) );
in01f01 g3621 ( .a(net_7802), .o(n10351) );
na02f01 g3622 ( .a(n6803), .b(_net_6040), .o(n10352) );
oa12f01 g3623 ( .a(n10352), .b(n6803), .c(n10351), .o(n5925) );
in01f01 g3624 ( .a(_net_7553), .o(n10354) );
na02f01 g3625 ( .a(n8246), .b(n7519), .o(n10355) );
oa12f01 g3626 ( .a(n10355), .b(n7519), .c(n10354), .o(n5938) );
na02f01 g3627 ( .a(n7348), .b(_net_7809), .o(n10357) );
oa12f01 g3628 ( .a(n10357), .b(n7348), .c(n7121), .o(n5960) );
in01f01 g3629 ( .a(_net_7360), .o(n10359) );
na02f01 g3630 ( .a(n7437_1), .b(n7030), .o(n10360) );
oa12f01 g3631 ( .a(n10360), .b(n7030), .c(n10359), .o(n5973) );
na02f01 g3632 ( .a(n8120), .b(n6921), .o(n10362) );
na02f01 g3633 ( .a(n8122), .b(_net_6689), .o(n10363) );
na02f01 g3634 ( .a(n10363), .b(n10362), .o(n10364) );
na02f01 g3635 ( .a(n10364), .b(n8125_1), .o(n10365) );
na02f01 g3636 ( .a(n6927), .b(n6919_1), .o(n10366) );
ao22f01 g3637 ( .a(n10366), .b(n8127), .c(n8132), .d(_net_6689), .o(n10367) );
na02f01 g3638 ( .a(n10367), .b(n10365), .o(n5982) );
ao12f01 g3639 ( .a(x38), .b(n9546_1), .c(_net_6410), .o(n10369) );
oa12f01 g3640 ( .a(n10369), .b(n9546_1), .c(_net_6410), .o(n5987) );
in01f01 g3641 ( .a(_net_7357), .o(n10371) );
na02f01 g3642 ( .a(n8809_1), .b(n7030), .o(n10372) );
oa12f01 g3643 ( .a(n10372), .b(n7030), .c(n10371), .o(n5992) );
na02f01 g3644 ( .a(n8116_1), .b(n8028_1), .o(n10374) );
ao22f01 g3645 ( .a(n9810), .b(n8033_1), .c(n8034), .d(_net_6066), .o(n10375) );
na02f01 g3646 ( .a(n10375), .b(n10374), .o(n5997) );
in01f01 g3647 ( .a(_net_7596), .o(n10377) );
na02f01 g3648 ( .a(n8043), .b(n6968), .o(n10378) );
oa12f01 g3649 ( .a(n10378), .b(n6968), .c(n10377), .o(n6024) );
no02f01 g3650 ( .a(n7085_1), .b(n6764), .o(n10380) );
no02f01 g3651 ( .a(n7094), .b(n6766), .o(n10381) );
in01f01 g3652 ( .a(_net_6081), .o(n10382) );
oa22f01 g3653 ( .a(n9047_1), .b(n6775), .c(n6784), .d(n10382), .o(n10383) );
no03f01 g3654 ( .a(n10383), .b(n10381), .c(n10380), .o(n10384) );
in01f01 g3655 ( .a(net_6453), .o(n10385) );
in01f01 g3656 ( .a(net_6485), .o(n10386) );
oa22f01 g3657 ( .a(n6790), .b(n10385), .c(n6789), .d(n10386), .o(n10387) );
in01f01 g3658 ( .a(net_6517), .o(n10388) );
in01f01 g3659 ( .a(net_6549), .o(n10389) );
oa22f01 g3660 ( .a(n6795), .b(n10389), .c(n6794), .d(n10388), .o(n10390) );
no02f01 g3661 ( .a(n10390), .b(n10387), .o(n10391) );
na02f01 g3662 ( .a(n10391), .b(n10384), .o(n6029) );
ao22f01 g3663 ( .a(n6736_1), .b(net_7637), .c(n6734), .d(net_7605), .o(n10393) );
ao22f01 g3664 ( .a(n6739), .b(net_7669), .c(n6738), .d(_net_7573), .o(n10394) );
na02f01 g3665 ( .a(n10394), .b(n10393), .o(n6038) );
ao12f01 g3666 ( .a(n6824), .b(n9202), .c(n9201_1), .o(n10396) );
no02f01 g3667 ( .a(n8435_1), .b(n6826_1), .o(n10397) );
in01f01 g3668 ( .a(_net_6132), .o(n10398) );
oa22f01 g3669 ( .a(n8443_1), .b(n6836_1), .c(n6844), .d(n10398), .o(n10399) );
no03f01 g3670 ( .a(n10399), .b(n10397), .c(n10396), .o(n10400) );
in01f01 g3671 ( .a(net_6849), .o(n10401) );
in01f01 g3672 ( .a(net_6881), .o(n10402) );
oa22f01 g3673 ( .a(n6850_1), .b(n10401), .c(n6849), .d(n10402), .o(n10403) );
in01f01 g3674 ( .a(net_6913), .o(n10404) );
in01f01 g3675 ( .a(net_6945), .o(n10405) );
oa22f01 g3676 ( .a(n6855_1), .b(n10405), .c(n6854), .d(n10404), .o(n10406) );
no02f01 g3677 ( .a(n10406), .b(n10403), .o(n10407) );
na02f01 g3678 ( .a(n10407), .b(n10400), .o(n6052) );
in01f01 g3679 ( .a(_net_7482), .o(n10409) );
na02f01 g3680 ( .a(n9487_1), .b(n6869), .o(n10410) );
oa12f01 g3681 ( .a(n10410), .b(n6869), .c(n10409), .o(n6061) );
in01f01 g3682 ( .a(n2222), .o(n10412) );
ao12f01 g3683 ( .a(n7756_1), .b(_net_6557), .c(net_6556), .o(n10413) );
no03f01 g3684 ( .a(n7765), .b(_net_6558), .c(n7762), .o(n10414) );
no02f01 g3685 ( .a(n10414), .b(n10413), .o(n10415) );
na02f01 g3686 ( .a(_net_5984), .b(n8330), .o(n10416) );
oa22f01 g3687 ( .a(n10416), .b(n7756_1), .c(n10415), .d(n10412), .o(n6074) );
ao22f01 g3688 ( .a(n6736_1), .b(net_7647), .c(n6734), .d(net_7615), .o(n10418) );
ao22f01 g3689 ( .a(n6739), .b(net_7679), .c(n6738), .d(_net_7583), .o(n10419) );
na02f01 g3690 ( .a(n10419), .b(n10418), .o(n6083) );
in01f01 g3691 ( .a(_net_6407), .o(n10421) );
na04f01 g3692 ( .a(n10421), .b(_net_6410), .c(n9258_1), .d(n8084), .o(n10422) );
in01f01 g3693 ( .a(_net_6408), .o(n10423) );
na02f01 g3694 ( .a(_net_6409), .b(n10423), .o(n10424) );
no03f01 g3695 ( .a(n10424), .b(n10422), .c(n8090), .o(n6088) );
in01f01 g3696 ( .a(_net_7405), .o(n10426) );
na02f01 g3697 ( .a(n8817), .b(n7550), .o(n10427) );
oa12f01 g3698 ( .a(n10427), .b(n7550), .c(n10426), .o(n6093) );
no02f01 g3699 ( .a(n8291), .b(n7721), .o(n10429) );
in01f01 g3700 ( .a(net_7114), .o(n10430) );
in01f01 g3701 ( .a(net_7178), .o(n10431) );
oa22f01 g3702 ( .a(n7580), .b(n10430), .c(n7577_1), .d(n10431), .o(n10432) );
in01f01 g3703 ( .a(net_7146), .o(n10433) );
in01f01 g3704 ( .a(net_7210), .o(n10434) );
oa22f01 g3705 ( .a(n7585), .b(n10433), .c(n7583), .d(n10434), .o(n10435) );
no02f01 g3706 ( .a(n10435), .b(n10432), .o(n10436) );
no02f01 g3707 ( .a(n10436), .b(n7592), .o(n10437) );
in01f01 g3708 ( .a(_net_6181), .o(n10438) );
no02f01 g3709 ( .a(n8508_1), .b(n8505), .o(n10439) );
oa22f01 g3710 ( .a(n10439), .b(n7574), .c(n7590), .d(n10438), .o(n10440) );
no03f01 g3711 ( .a(n10440), .b(n10437), .c(n10429), .o(n10441) );
in01f01 g3712 ( .a(net_7128), .o(n10442) );
in01f01 g3713 ( .a(net_7160), .o(n10443) );
oa22f01 g3714 ( .a(n7740), .b(n10442), .c(n7739), .d(n10443), .o(n10444) );
in01f01 g3715 ( .a(net_7224), .o(n10445) );
in01f01 g3716 ( .a(net_7192), .o(n10446) );
oa22f01 g3717 ( .a(n7745), .b(n10445), .c(n7744), .d(n10446), .o(n10447) );
no02f01 g3718 ( .a(n10447), .b(n10444), .o(n10448) );
na02f01 g3719 ( .a(n10448), .b(n10441), .o(n6119) );
in01f01 g3720 ( .a(_net_7729), .o(n10450) );
ao12f01 g3721 ( .a(n7343), .b(n10450), .c(n8419), .o(n6124) );
no02f01 g3722 ( .a(n6736_1), .b(n6734), .o(n10452) );
in01f01 g3723 ( .a(_net_264), .o(n10453) );
no02f01 g3724 ( .a(n8236), .b(n10453), .o(n8038) );
in01f01 g3725 ( .a(n8038), .o(n10455) );
na02f01 g3726 ( .a(_net_289), .b(n10453), .o(n10456) );
oa22f01 g3727 ( .a(n10456), .b(n6735), .c(n10455), .d(n10452), .o(n6140) );
in01f01 g3728 ( .a(_net_6292), .o(n10458) );
no02f01 g3729 ( .a(_net_392), .b(n10458), .o(n6153) );
in01f01 g3730 ( .a(_net_6208), .o(n10460) );
no02f01 g3731 ( .a(_net_392), .b(n10460), .o(n6166) );
oa12f01 g3732 ( .a(n8028_1), .b(n9180), .c(n9177), .o(n10462) );
na02f01 g3733 ( .a(n9832), .b(n9831), .o(n10463) );
ao22f01 g3734 ( .a(n10463), .b(n8033_1), .c(n8034), .d(_net_6071), .o(n10464) );
na02f01 g3735 ( .a(n9050), .b(n9049), .o(n10465) );
ao22f01 g3736 ( .a(n10465), .b(n8113), .c(n8031), .d(n8110), .o(n10466) );
na03f01 g3737 ( .a(n10466), .b(n10464), .c(n10462), .o(n6171) );
na02f01 g3738 ( .a(n8211_1), .b(_net_6124), .o(n10468) );
na02f01 g3739 ( .a(n9658), .b(n8213), .o(n10469) );
na02f01 g3740 ( .a(n10469), .b(n10468), .o(n6186) );
ao22f01 g3741 ( .a(n7000_1), .b(net_6969), .c(n6999), .d(net_7033), .o(n10471) );
ao22f01 g3742 ( .a(n7003), .b(net_7001), .c(n7002), .d(net_7065), .o(n10472) );
na02f01 g3743 ( .a(n10472), .b(n10471), .o(n10473) );
na02f01 g3744 ( .a(n10473), .b(n6981), .o(n10474) );
ao22f01 g3745 ( .a(n7323), .b(n6998), .c(n6996), .d(_net_6149), .o(n10475) );
na02f01 g3746 ( .a(n7327), .b(n7013_1), .o(n10476) );
oa12f01 g3747 ( .a(n7022), .b(n8478), .c(n8475), .o(n10477) );
na04f01 g3748 ( .a(n10477), .b(n10476), .c(n10475), .d(n10474), .o(n6191) );
in01f01 g3749 ( .a(_net_7693), .o(n10479) );
na02f01 g3750 ( .a(n7207_1), .b(_net_7795), .o(n10480) );
oa12f01 g3751 ( .a(n10480), .b(n7207_1), .c(n10479), .o(n6200) );
in01f01 g3752 ( .a(_net_7254), .o(n10482) );
na02f01 g3753 ( .a(n8960), .b(n6901), .o(n10483) );
oa12f01 g3754 ( .a(n10483), .b(n6901), .c(n10482), .o(n6209) );
no02f01 g3755 ( .a(n7822_1), .b(n6945), .o(n10485) );
no02f01 g3756 ( .a(n8746), .b(n6934_1), .o(n10486) );
in01f01 g3757 ( .a(_net_6099), .o(n10487) );
in01f01 g3758 ( .a(net_6574), .o(n10488) );
in01f01 g3759 ( .a(net_6638), .o(n10489) );
oa22f01 g3760 ( .a(n6922), .b(n10488), .c(n6919_1), .d(n10489), .o(n10490) );
in01f01 g3761 ( .a(net_6606), .o(n10491) );
in01f01 g3762 ( .a(net_6670), .o(n10492) );
oa22f01 g3763 ( .a(n6927), .b(n10491), .c(n6925), .d(n10492), .o(n10493) );
no02f01 g3764 ( .a(n10493), .b(n10490), .o(n10494) );
oa22f01 g3765 ( .a(n10494), .b(n6916), .c(n6932), .d(n10487), .o(n10495) );
no03f01 g3766 ( .a(n10495), .b(n10486), .c(n10485), .o(n10496) );
in01f01 g3767 ( .a(net_6586), .o(n10497) );
in01f01 g3768 ( .a(net_6618), .o(n10498) );
oa22f01 g3769 ( .a(n7058_1), .b(n10497), .c(n7057), .d(n10498), .o(n10499) );
in01f01 g3770 ( .a(net_6650), .o(n10500) );
in01f01 g3771 ( .a(net_6682), .o(n10501) );
oa22f01 g3772 ( .a(n7063), .b(n10501), .c(n7062_1), .d(n10500), .o(n10502) );
no02f01 g3773 ( .a(n10502), .b(n10499), .o(n10503) );
na02f01 g3774 ( .a(n10503), .b(n10496), .o(n6218) );
ao22f01 g3775 ( .a(n6877), .b(_net_7280), .c(n6876_1), .d(net_7344), .o(n10505) );
ao22f01 g3776 ( .a(n6881_1), .b(net_7312), .c(n6880), .d(net_7376), .o(n10506) );
na02f01 g3777 ( .a(n10506), .b(n10505), .o(n6227) );
ao22f01 g3778 ( .a(n7225), .b(_net_7418), .c(n7224), .d(_net_7450), .o(n10508) );
ao22f01 g3779 ( .a(n7229), .b(_net_7514), .c(n7228), .d(_net_7482), .o(n10509) );
na02f01 g3780 ( .a(n10509), .b(n10508), .o(n6244) );
ao22f01 g3781 ( .a(n7225), .b(_net_7409), .c(n7224), .d(_net_7441), .o(n10511) );
ao22f01 g3782 ( .a(n7229), .b(_net_7505), .c(n7228), .d(_net_7473), .o(n10512) );
na02f01 g3783 ( .a(n10512), .b(n10511), .o(n6249) );
in01f01 g3784 ( .a(_net_7434), .o(n10514) );
na02f01 g3785 ( .a(n7883_1), .b(n7197), .o(n10515) );
oa12f01 g3786 ( .a(n10515), .b(n7197), .c(n10514), .o(n6266) );
ao22f01 g3787 ( .a(n6877), .b(_net_7261), .c(n6876_1), .d(_net_7325), .o(n10517) );
ao22f01 g3788 ( .a(n6881_1), .b(_net_7293), .c(n6880), .d(_net_7357), .o(n10518) );
na02f01 g3789 ( .a(n10518), .b(n10517), .o(n6271) );
ao22f01 g3790 ( .a(n6877), .b(_net_7268), .c(n6876_1), .d(_net_7332), .o(n10520) );
ao22f01 g3791 ( .a(n6881_1), .b(_net_7300), .c(n6880), .d(_net_7364), .o(n10521) );
na02f01 g3792 ( .a(n10521), .b(n10520), .o(n6281) );
ao22f01 g3793 ( .a(n7298), .b(_net_7723), .c(n7288_1), .d(_net_6031), .o(n10523) );
ao22f01 g3794 ( .a(n7306), .b(_net_5987), .c(n7286), .d(_net_270), .o(n10524) );
na02f01 g3795 ( .a(n7302_1), .b(_net_117), .o(n10525) );
na03f01 g3796 ( .a(n7308), .b(net_159), .c(n6800), .o(n10526) );
na03f01 g3797 ( .a(n7308), .b(net_196), .c(x1322), .o(n10527) );
na02f01 g3798 ( .a(n7296), .b(net_233), .o(n10528) );
na03f01 g3799 ( .a(n10528), .b(n10527), .c(n10526), .o(n10529) );
ao12f01 g3800 ( .a(n10529), .b(n7291), .c(_net_7694), .o(n10530) );
na04f01 g3801 ( .a(n10530), .b(n10525), .c(n10524), .d(n10523), .o(n6290) );
in01f01 g3802 ( .a(_net_7787), .o(n10532) );
no04f01 g3803 ( .a(n7360), .b(n7355), .c(n10532), .d(n7359_1), .o(n10533) );
no02f01 g3804 ( .a(n10533), .b(_net_7789), .o(n10534) );
in01f01 g3805 ( .a(_net_7789), .o(n10535) );
in01f01 g3806 ( .a(n10533), .o(n10536) );
no02f01 g3807 ( .a(n10536), .b(n10535), .o(n10537) );
no03f01 g3808 ( .a(n10537), .b(n10534), .c(n7358), .o(n6294) );
ao12f01 g3809 ( .a(n8330), .b(_net_6555), .c(_net_6558), .o(n10539) );
oa12f01 g3810 ( .a(n10539), .b(_net_6555), .c(_net_6558), .o(n10540) );
na02f01 g3811 ( .a(n8472), .b(n9269), .o(n10541) );
oa12f01 g3812 ( .a(n8366), .b(n10541), .c(n10540), .o(n6311) );
in01f01 g3813 ( .a(_net_6001), .o(n10543) );
na02f01 g3814 ( .a(n7348), .b(net_7807), .o(n10544) );
oa12f01 g3815 ( .a(n10544), .b(n7348), .c(n10543), .o(n6324) );
no02f01 g3816 ( .a(n8104), .b(n8101), .o(n10546) );
no02f01 g3817 ( .a(n10546), .b(n6764), .o(n10547) );
in01f01 g3818 ( .a(net_6432), .o(n10548) );
in01f01 g3819 ( .a(net_6496), .o(n10549) );
oa22f01 g3820 ( .a(n6750), .b(n10548), .c(n6748), .d(n10549), .o(n10550) );
in01f01 g3821 ( .a(net_6528), .o(n10551) );
in01f01 g3822 ( .a(net_6464), .o(n10552) );
oa22f01 g3823 ( .a(n6755), .b(n10552), .c(n6754), .d(n10551), .o(n10553) );
no02f01 g3824 ( .a(n10553), .b(n10550), .o(n10554) );
no02f01 g3825 ( .a(n10554), .b(n6766), .o(n10555) );
in01f01 g3826 ( .a(_net_6074), .o(n10556) );
oa22f01 g3827 ( .a(n9225_1), .b(n6775), .c(n6784), .d(n10556), .o(n10557) );
no03f01 g3828 ( .a(n10557), .b(n10555), .c(n10547), .o(n10558) );
in01f01 g3829 ( .a(net_6478), .o(n10559) );
in01f01 g3830 ( .a(net_6446), .o(n10560) );
oa22f01 g3831 ( .a(n6790), .b(n10560), .c(n6789), .d(n10559), .o(n10561) );
in01f01 g3832 ( .a(net_6510), .o(n10562) );
in01f01 g3833 ( .a(net_6542), .o(n10563) );
oa22f01 g3834 ( .a(n6795), .b(n10563), .c(n6794), .d(n10562), .o(n10564) );
no02f01 g3835 ( .a(n10564), .b(n10561), .o(n10565) );
na02f01 g3836 ( .a(n10565), .b(n10558), .o(n6337) );
in01f01 g3837 ( .a(_net_7353), .o(n10567) );
na02f01 g3838 ( .a(n9587), .b(n7030), .o(n10568) );
oa12f01 g3839 ( .a(n10568), .b(n7030), .c(n10567), .o(n6346) );
in01f01 g3840 ( .a(_net_7440), .o(n10570) );
na02f01 g3841 ( .a(n8141), .b(n7197), .o(n10571) );
oa12f01 g3842 ( .a(n10571), .b(n7197), .c(n10570), .o(n6362) );
in01f01 g3843 ( .a(_net_7098), .o(n10573) );
in01f01 g3844 ( .a(n2590), .o(n10574) );
ao12f01 g3845 ( .a(n10573), .b(_net_7097), .c(net_7096), .o(n10575) );
no03f01 g3846 ( .a(n8760), .b(_net_7098), .c(n8385), .o(n10576) );
no02f01 g3847 ( .a(n10576), .b(n10575), .o(n10577) );
na02f01 g3848 ( .a(_net_6028), .b(n8650_1), .o(n10578) );
oa22f01 g3849 ( .a(n10578), .b(n10573), .c(n10577), .d(n10574), .o(n6371) );
in01f01 g3850 ( .a(_net_7661), .o(n10580) );
na02f01 g3851 ( .a(n7446_1), .b(n7428), .o(n10581) );
oa12f01 g3852 ( .a(n10581), .b(n7446_1), .c(n10580), .o(n6381) );
no02f01 g3853 ( .a(n8746), .b(n6945), .o(n10583) );
no02f01 g3854 ( .a(n10494), .b(n6934_1), .o(n10584) );
in01f01 g3855 ( .a(_net_6101), .o(n10585) );
in01f01 g3856 ( .a(net_6576), .o(n10586) );
in01f01 g3857 ( .a(net_6640), .o(n10587) );
oa22f01 g3858 ( .a(n6922), .b(n10586), .c(n6919_1), .d(n10587), .o(n10588) );
in01f01 g3859 ( .a(net_6608), .o(n10589) );
in01f01 g3860 ( .a(net_6672), .o(n10590) );
oa22f01 g3861 ( .a(n6927), .b(n10589), .c(n6925), .d(n10590), .o(n10591) );
no02f01 g3862 ( .a(n10591), .b(n10588), .o(n10592) );
oa22f01 g3863 ( .a(n10592), .b(n6916), .c(n6932), .d(n10585), .o(n10593) );
no03f01 g3864 ( .a(n10593), .b(n10584), .c(n10583), .o(n10594) );
in01f01 g3865 ( .a(net_6588), .o(n10595) );
in01f01 g3866 ( .a(net_6620), .o(n10596) );
oa22f01 g3867 ( .a(n7058_1), .b(n10595), .c(n7057), .d(n10596), .o(n10597) );
in01f01 g3868 ( .a(net_6652), .o(n10598) );
in01f01 g3869 ( .a(net_6684), .o(n10599) );
oa22f01 g3870 ( .a(n7063), .b(n10599), .c(n7062_1), .d(n10598), .o(n10600) );
no02f01 g3871 ( .a(n10600), .b(n10597), .o(n10601) );
na02f01 g3872 ( .a(n10601), .b(n10594), .o(n6395) );
in01f01 g3873 ( .a(_net_7438), .o(n10603) );
na02f01 g3874 ( .a(n7860), .b(n7197), .o(n10604) );
oa12f01 g3875 ( .a(n10604), .b(n7197), .c(n10603), .o(n6411) );
ao22f01 g3876 ( .a(n6877), .b(_net_7250), .c(n6876_1), .d(_net_7314), .o(n10606) );
ao22f01 g3877 ( .a(n6881_1), .b(_net_7282), .c(n6880), .d(_net_7346), .o(n10607) );
na02f01 g3878 ( .a(n10607), .b(n10606), .o(n6432) );
no02f01 g3879 ( .a(_net_6692), .b(n7153), .o(n10609) );
no02f01 g3880 ( .a(n7663), .b(net_6691), .o(n10610) );
no02f01 g3881 ( .a(n10610), .b(n10609), .o(n10611) );
oa22f01 g3882 ( .a(n10611), .b(n9974), .c(n9978), .d(n7663), .o(n6450) );
in01f01 g3883 ( .a(_net_7257), .o(n10613) );
na02f01 g3884 ( .a(n9587), .b(n6901), .o(n10614) );
oa12f01 g3885 ( .a(n10614), .b(n6901), .c(n10613), .o(n6455) );
ao22f01 g3886 ( .a(n7225), .b(_net_7413), .c(n7224), .d(_net_7445), .o(n10616) );
ao22f01 g3887 ( .a(n7229), .b(_net_7509), .c(n7228), .d(_net_7477), .o(n10617) );
na02f01 g3888 ( .a(n10617), .b(n10616), .o(n6493) );
in01f01 g3889 ( .a(_net_5857), .o(n10619) );
in01f01 g3890 ( .a(x1034), .o(n10620) );
in01f01 g3891 ( .a(_net_5999), .o(n10621) );
no02f01 g3892 ( .a(n10621), .b(_net_6000), .o(n10622) );
na02f01 g3893 ( .a(_net_5995), .b(_net_6001), .o(n10623) );
ao12f01 g3894 ( .a(n10623), .b(n7191), .c(_net_5966), .o(n10624) );
na02f01 g3895 ( .a(n10624), .b(n10622), .o(n10625) );
in01f01 g3896 ( .a(n10623), .o(n10626) );
na03f01 g3897 ( .a(n7191), .b(_net_5966), .c(_net_5965), .o(n10627) );
na04f01 g3898 ( .a(n10627), .b(n10626), .c(n10621), .d(n7673), .o(n10628) );
oa12f01 g3899 ( .a(n7191), .b(_net_5966), .c(_net_5965), .o(n10629) );
na04f01 g3900 ( .a(n10629), .b(n10626), .c(n10621), .d(_net_6000), .o(n10630) );
no02f01 g3901 ( .a(n10621), .b(n7673), .o(n10631) );
na03f01 g3902 ( .a(n10631), .b(n10626), .c(_net_5964), .o(n10632) );
na04f01 g3903 ( .a(n10632), .b(n10630), .c(n10628), .d(n10625), .o(n10633) );
na03f01 g3904 ( .a(n10633), .b(net_7773), .c(n10620), .o(n10634) );
oa12f01 g3905 ( .a(n10634), .b(n10619), .c(x1034), .o(n6527) );
na02f01 g3906 ( .a(n9211_1), .b(n8213), .o(n10636) );
ao22f01 g3907 ( .a(n9658), .b(n9200), .c(n8211_1), .d(_net_6126), .o(n10637) );
na02f01 g3908 ( .a(n10637), .b(n10636), .o(n6540) );
in01f01 g3909 ( .a(_net_118), .o(n10639) );
na02f01 g3910 ( .a(net_314), .b(_net_154), .o(n10640) );
oa12f01 g3911 ( .a(n10640), .b(n10639), .c(_net_154), .o(n6545) );
in01f01 g3912 ( .a(_net_7654), .o(n10642) );
na02f01 g3913 ( .a(n7644_1), .b(n7446_1), .o(n10643) );
oa12f01 g3914 ( .a(n10643), .b(n7446_1), .c(n10642), .o(n6558) );
na02f01 g3915 ( .a(n7009_1), .b(n6981), .o(n10645) );
ao22f01 g3916 ( .a(n9719_1), .b(n6998), .c(n6996), .d(_net_6146), .o(n10646) );
na02f01 g3917 ( .a(n10646), .b(n10645), .o(n6570) );
na03f01 g3918 ( .a(_net_6407), .b(_net_6405), .c(_net_6406), .o(n10648) );
no02f01 g3919 ( .a(n8087), .b(_net_6411), .o(n10649) );
ao12f01 g3920 ( .a(n8177), .b(n10649), .c(n10648), .o(n6583) );
ao22f01 g3921 ( .a(n6877), .b(_net_7251), .c(n6876_1), .d(_net_7315), .o(n10651) );
ao22f01 g3922 ( .a(n6881_1), .b(_net_7283), .c(n6880), .d(_net_7347), .o(n10652) );
na02f01 g3923 ( .a(n10652), .b(n10651), .o(n6591) );
in01f01 g3924 ( .a(net_6769), .o(n10654) );
in01f01 g3925 ( .a(net_6705), .o(n10655) );
oa22f01 g3926 ( .a(n7129), .b(n10655), .c(n7126), .d(n10654), .o(n10656) );
in01f01 g3927 ( .a(net_6737), .o(n10657) );
in01f01 g3928 ( .a(net_6801), .o(n10658) );
oa22f01 g3929 ( .a(n7134), .b(n10657), .c(n7132), .d(n10658), .o(n10659) );
no02f01 g3930 ( .a(n10659), .b(n10656), .o(n10660) );
no02f01 g3931 ( .a(n10660), .b(n7468_1), .o(n10661) );
no02f01 g3932 ( .a(n8665), .b(n7470), .o(n10662) );
in01f01 g3933 ( .a(_net_6119), .o(n10663) );
oa22f01 g3934 ( .a(n8673), .b(n7123), .c(n7118), .d(n10663), .o(n10664) );
no03f01 g3935 ( .a(n10664), .b(n10662), .c(n10661), .o(n10665) );
in01f01 g3936 ( .a(net_6721), .o(n10666) );
in01f01 g3937 ( .a(net_6753), .o(n10667) );
oa22f01 g3938 ( .a(n7492_1), .b(n10666), .c(n7491), .d(n10667), .o(n10668) );
in01f01 g3939 ( .a(net_6817), .o(n10669) );
in01f01 g3940 ( .a(net_6785), .o(n10670) );
oa22f01 g3941 ( .a(n7497), .b(n10669), .c(n7496_1), .d(n10670), .o(n10671) );
no02f01 g3942 ( .a(n10671), .b(n10668), .o(n10672) );
na02f01 g3943 ( .a(n10672), .b(n10665), .o(n6596) );
in01f01 g3944 ( .a(_net_7448), .o(n10674) );
na02f01 g3945 ( .a(n7638), .b(n7197), .o(n10675) );
oa12f01 g3946 ( .a(n10675), .b(n7197), .c(n10674), .o(n6601) );
na02f01 g3947 ( .a(n9518), .b(_net_7098), .o(n10677) );
na03f01 g3948 ( .a(n9517_1), .b(n9516), .c(n10573), .o(n10678) );
na02f01 g3949 ( .a(n8199), .b(net_7096), .o(n10679) );
na03f01 g3950 ( .a(n8198), .b(n8197_1), .c(n8385), .o(n10680) );
ao22f01 g3951 ( .a(n10680), .b(n10679), .c(n7011), .d(_net_7092), .o(n10681) );
na02f01 g3952 ( .a(n7214), .b(n8760), .o(n10682) );
na03f01 g3953 ( .a(n7213), .b(n7211), .c(_net_7097), .o(n10683) );
na03f01 g3954 ( .a(n10683), .b(n10682), .c(n10681), .o(n10684) );
ao12f01 g3955 ( .a(n10684), .b(n10678), .c(n10677), .o(n6606) );
ao22f01 g3956 ( .a(n6877), .b(_net_7262), .c(n6876_1), .d(_net_7326), .o(n10686) );
ao22f01 g3957 ( .a(n6881_1), .b(_net_7294), .c(n6880), .d(_net_7358), .o(n10687) );
na02f01 g3958 ( .a(n10687), .b(n10686), .o(n6624) );
oa12f01 g3959 ( .a(n7575), .b(n9756), .c(n9753), .o(n10689) );
ao22f01 g3960 ( .a(n7908), .b(n7593), .c(n7591_1), .d(_net_6170), .o(n10690) );
na02f01 g3961 ( .a(n7732_1), .b(n7731), .o(n10691) );
ao22f01 g3962 ( .a(n7912), .b(n7914), .c(n7920_1), .d(n10691), .o(n10692) );
na03f01 g3963 ( .a(n10692), .b(n10690), .c(n10689), .o(n6634) );
no03f01 g3964 ( .a(n6912), .b(_net_5999), .c(n7673), .o(n10694) );
no02f01 g3965 ( .a(n7191), .b(n6912), .o(n10695) );
ao22f01 g3966 ( .a(n10695), .b(n10631), .c(n10694), .d(n10629), .o(n10696) );
ao12f01 g3967 ( .a(n6912), .b(n7191), .c(_net_5966), .o(n10697) );
no03f01 g3968 ( .a(n6912), .b(_net_5999), .c(_net_6000), .o(n10698) );
ao22f01 g3969 ( .a(n10698), .b(n10627), .c(n10697), .d(n10622), .o(n10699) );
na02f01 g3970 ( .a(n10699), .b(n10696), .o(n6643) );
in01f01 g3971 ( .a(_net_124), .o(n10701) );
na02f01 g3972 ( .a(net_320), .b(_net_154), .o(n10702) );
oa12f01 g3973 ( .a(n10702), .b(n10701), .c(_net_154), .o(n6652) );
na02f01 g3974 ( .a(n6817), .b(n6812), .o(n10704) );
na02f01 g3975 ( .a(n8213), .b(n10704), .o(n10705) );
ao22f01 g3976 ( .a(n6811), .b(net_6832), .c(n6808), .d(net_6896), .o(n10706) );
ao22f01 g3977 ( .a(n6816), .b(net_6864), .c(n6814), .d(net_6928), .o(n10707) );
na02f01 g3978 ( .a(n10707), .b(n10706), .o(n10708) );
ao22f01 g3979 ( .a(n10708), .b(n9200), .c(n8211_1), .d(_net_6129), .o(n10709) );
na02f01 g3980 ( .a(n8216_1), .b(n9205), .o(n10710) );
in01f01 g3981 ( .a(net_6846), .o(n10711) );
in01f01 g3982 ( .a(net_6910), .o(n10712) );
oa22f01 g3983 ( .a(n6810), .b(n10711), .c(n6807), .d(n10712), .o(n10713) );
in01f01 g3984 ( .a(net_6942), .o(n10714) );
in01f01 g3985 ( .a(net_6878), .o(n10715) );
oa22f01 g3986 ( .a(n6815), .b(n10715), .c(n6813_1), .d(n10714), .o(n10716) );
oa12f01 g3987 ( .a(n9207), .b(n10716), .c(n10713), .o(n10717) );
na04f01 g3988 ( .a(n10717), .b(n10710), .c(n10709), .d(n10705), .o(n6665) );
na02f01 g3989 ( .a(n7440), .b(_net_7801), .o(n10719) );
oa12f01 g3990 ( .a(n10719), .b(n7440), .c(n7850), .o(n6682) );
ao22f01 g3991 ( .a(n7288_1), .b(_net_6033), .c(n7286), .d(_net_272), .o(n10721) );
ao22f01 g3992 ( .a(n7298), .b(_net_7725), .c(n7291), .d(_net_7696), .o(n10722) );
na02f01 g3993 ( .a(n7302_1), .b(_net_119), .o(n10723) );
na03f01 g3994 ( .a(n7308), .b(net_198), .c(x1322), .o(n10724) );
na02f01 g3995 ( .a(n7296), .b(net_235), .o(n10725) );
na03f01 g3996 ( .a(n7308), .b(net_161), .c(n6800), .o(n10726) );
na03f01 g3997 ( .a(n10726), .b(n10725), .c(n10724), .o(n10727) );
ao12f01 g3998 ( .a(n10727), .b(n7306), .c(_net_5989), .o(n10728) );
na04f01 g3999 ( .a(n10728), .b(n10723), .c(n10722), .d(n10721), .o(n6691) );
in01f01 g4000 ( .a(_net_7623), .o(n10730) );
na02f01 g4001 ( .a(n9493), .b(n7400_1), .o(n10731) );
oa12f01 g4002 ( .a(n10731), .b(n7400_1), .c(n10730), .o(n6695) );
in01f01 g4003 ( .a(_net_7279), .o(n10733) );
na02f01 g4004 ( .a(n1034), .b(n6901), .o(n10734) );
oa12f01 g4005 ( .a(n10734), .b(n6901), .c(n10733), .o(n6709) );
ao22f01 g4006 ( .a(n7130), .b(net_6699), .c(n7127), .d(net_6763), .o(n10736) );
ao22f01 g4007 ( .a(n7135), .b(net_6731), .c(n7133_1), .d(net_6795), .o(n10737) );
ao12f01 g4008 ( .a(n7468_1), .b(n10737), .c(n10736), .o(n10738) );
in01f01 g4009 ( .a(net_6765), .o(n10739) );
in01f01 g4010 ( .a(net_6701), .o(n10740) );
oa22f01 g4011 ( .a(n7129), .b(n10740), .c(n7126), .d(n10739), .o(n10741) );
in01f01 g4012 ( .a(net_6733), .o(n10742) );
in01f01 g4013 ( .a(net_6797), .o(n10743) );
oa22f01 g4014 ( .a(n7134), .b(n10742), .c(n7132), .d(n10743), .o(n10744) );
no02f01 g4015 ( .a(n10744), .b(n10741), .o(n10745) );
no02f01 g4016 ( .a(n10745), .b(n7470), .o(n10746) );
in01f01 g4017 ( .a(_net_6113), .o(n10747) );
in01f01 g4018 ( .a(net_6767), .o(n10748) );
in01f01 g4019 ( .a(net_6703), .o(n10749) );
oa22f01 g4020 ( .a(n7129), .b(n10749), .c(n7126), .d(n10748), .o(n10750) );
in01f01 g4021 ( .a(net_6799), .o(n10751) );
in01f01 g4022 ( .a(net_6735), .o(n10752) );
oa22f01 g4023 ( .a(n7134), .b(n10752), .c(n7132), .d(n10751), .o(n10753) );
no02f01 g4024 ( .a(n10753), .b(n10750), .o(n10754) );
oa22f01 g4025 ( .a(n10754), .b(n7123), .c(n7118), .d(n10747), .o(n10755) );
no03f01 g4026 ( .a(n10755), .b(n10746), .c(n10738), .o(n10756) );
in01f01 g4027 ( .a(net_6747), .o(n10757) );
in01f01 g4028 ( .a(net_6715), .o(n10758) );
oa22f01 g4029 ( .a(n7492_1), .b(n10758), .c(n7491), .d(n10757), .o(n10759) );
in01f01 g4030 ( .a(net_6779), .o(n10760) );
in01f01 g4031 ( .a(net_6811), .o(n10761) );
oa22f01 g4032 ( .a(n7497), .b(n10761), .c(n7496_1), .d(n10760), .o(n10762) );
no02f01 g4033 ( .a(n10762), .b(n10759), .o(n10763) );
na02f01 g4034 ( .a(n10763), .b(n10756), .o(n6727) );
in01f01 g4035 ( .a(_net_7620), .o(n10765) );
na02f01 g4036 ( .a(n8426_1), .b(n7400_1), .o(n10766) );
oa12f01 g4037 ( .a(n10766), .b(n7400_1), .c(n10765), .o(n6741) );
no02f01 g4038 ( .a(n8443_1), .b(n6824), .o(n10768) );
no02f01 g4039 ( .a(n8452), .b(n6826_1), .o(n10769) );
in01f01 g4040 ( .a(_net_6136), .o(n10770) );
oa22f01 g4041 ( .a(n10249), .b(n6836_1), .c(n6844), .d(n10770), .o(n10771) );
no03f01 g4042 ( .a(n10771), .b(n10769), .c(n10768), .o(n10772) );
in01f01 g4043 ( .a(net_6885), .o(n10773) );
in01f01 g4044 ( .a(net_6853), .o(n10774) );
oa22f01 g4045 ( .a(n6850_1), .b(n10774), .c(n6849), .d(n10773), .o(n10775) );
in01f01 g4046 ( .a(net_6949), .o(n10776) );
in01f01 g4047 ( .a(net_6917), .o(n10777) );
oa22f01 g4048 ( .a(n6855_1), .b(n10776), .c(n6854), .d(n10777), .o(n10778) );
no02f01 g4049 ( .a(n10778), .b(n10775), .o(n10779) );
na02f01 g4050 ( .a(n10779), .b(n10772), .o(n6765) );
no02f01 g4051 ( .a(n10754), .b(n7468_1), .o(n10781) );
no02f01 g4052 ( .a(n10660), .b(n7470), .o(n10782) );
in01f01 g4053 ( .a(_net_6117), .o(n10783) );
oa22f01 g4054 ( .a(n8665), .b(n7123), .c(n7118), .d(n10783), .o(n10784) );
no03f01 g4055 ( .a(n10784), .b(n10782), .c(n10781), .o(n10785) );
in01f01 g4056 ( .a(net_6751), .o(n10786) );
in01f01 g4057 ( .a(net_6719), .o(n10787) );
oa22f01 g4058 ( .a(n7492_1), .b(n10787), .c(n7491), .d(n10786), .o(n10788) );
in01f01 g4059 ( .a(net_6783), .o(n10789) );
in01f01 g4060 ( .a(net_6815), .o(n10790) );
oa22f01 g4061 ( .a(n7497), .b(n10790), .c(n7496_1), .d(n10789), .o(n10791) );
no02f01 g4062 ( .a(n10791), .b(n10788), .o(n10792) );
na02f01 g4063 ( .a(n10792), .b(n10785), .o(n6774) );
in01f01 g4064 ( .a(_net_7723), .o(n10794) );
in01f01 g4065 ( .a(_net_5993), .o(n10795) );
ao12f01 g4066 ( .a(n7343), .b(n10795), .c(n10794), .o(n6779) );
in01f01 g4067 ( .a(_net_7446), .o(n10797) );
na02f01 g4068 ( .a(n8994), .b(n7197), .o(n10798) );
oa12f01 g4069 ( .a(n10798), .b(n7197), .c(n10797), .o(n6788) );
in01f01 g4070 ( .a(_net_7258), .o(n10800) );
na02f01 g4071 ( .a(n7393), .b(n6901), .o(n10801) );
oa12f01 g4072 ( .a(n10801), .b(n6901), .c(n10800), .o(n6801) );
in01f01 g4073 ( .a(_net_7700), .o(n10803) );
na02f01 g4074 ( .a(n7207_1), .b(net_7802), .o(n10804) );
oa12f01 g4075 ( .a(n10804), .b(n7207_1), .c(n10803), .o(n6818) );
in01f01 g4076 ( .a(_net_7584), .o(n10806) );
na02f01 g4077 ( .a(n8842), .b(n6968), .o(n10807) );
oa12f01 g4078 ( .a(n10807), .b(n6968), .c(n10806), .o(n6831) );
oa12f01 g4079 ( .a(n10795), .b(n6761_1), .c(n7533), .o(n6840) );
in01f01 g4080 ( .a(_net_7325), .o(n10810) );
na02f01 g4081 ( .a(n8809_1), .b(n7150), .o(n10811) );
oa12f01 g4082 ( .a(n10811), .b(n7150), .c(n10810), .o(n6845) );
ao22f01 g4083 ( .a(n6736_1), .b(_net_7626), .c(n6734), .d(_net_7594), .o(n10813) );
ao22f01 g4084 ( .a(n6739), .b(_net_7658), .c(n6738), .d(_net_7562), .o(n10814) );
na02f01 g4085 ( .a(n10814), .b(n10813), .o(n6850) );
in01f01 g4086 ( .a(_net_5990), .o(n10816) );
na02f01 g4087 ( .a(n7348), .b(net_7799), .o(n10817) );
oa12f01 g4088 ( .a(n10817), .b(n7348), .c(n10816), .o(n6855) );
ao22f01 g4089 ( .a(n7225), .b(_net_7424), .c(n7224), .d(net_7456), .o(n10819) );
ao22f01 g4090 ( .a(n7229), .b(net_7520), .c(n7228), .d(net_7488), .o(n10820) );
na02f01 g4091 ( .a(n10820), .b(n10819), .o(n6872) );
no02f01 g4092 ( .a(n9934), .b(n7012), .o(n10822) );
no02f01 g4093 ( .a(n8471), .b(n6997), .o(n10823) );
in01f01 g4094 ( .a(_net_6161), .o(n10824) );
oa22f01 g4095 ( .a(n8479), .b(n6980), .c(n6995_1), .d(n10824), .o(n10825) );
no03f01 g4096 ( .a(n10825), .b(n10823), .c(n10822), .o(n10826) );
in01f01 g4097 ( .a(net_6993), .o(n10827) );
in01f01 g4098 ( .a(net_7025), .o(n10828) );
oa22f01 g4099 ( .a(n8075_1), .b(n10827), .c(n8074), .d(n10828), .o(n10829) );
in01f01 g4100 ( .a(net_7089), .o(n10830) );
in01f01 g4101 ( .a(net_7057), .o(n10831) );
oa22f01 g4102 ( .a(n8080_1), .b(n10830), .c(n8079), .d(n10831), .o(n10832) );
no02f01 g4103 ( .a(n10832), .b(n10829), .o(n10833) );
na02f01 g4104 ( .a(n10833), .b(n10826), .o(n6881) );
in01f01 g4105 ( .a(_net_7427), .o(n10835) );
na02f01 g4106 ( .a(n1173), .b(n7550), .o(n10836) );
oa12f01 g4107 ( .a(n10836), .b(n7550), .c(n10835), .o(n6890) );
ao22f01 g4108 ( .a(n7225), .b(_net_7423), .c(n7224), .d(net_7455), .o(n10838) );
ao22f01 g4109 ( .a(n7229), .b(net_7519), .c(n7228), .d(net_7487), .o(n10839) );
na02f01 g4110 ( .a(n10839), .b(n10838), .o(n6915) );
in01f01 g4111 ( .a(_net_7443), .o(n10841) );
na02f01 g4112 ( .a(n9786), .b(n7197), .o(n10842) );
oa12f01 g4113 ( .a(n10842), .b(n7197), .c(n10841), .o(n6924) );
ao22f01 g4114 ( .a(n6736_1), .b(_net_7630), .c(n6734), .d(_net_7598), .o(n10844) );
ao22f01 g4115 ( .a(n6739), .b(_net_7662), .c(n6738), .d(_net_7566), .o(n10845) );
na02f01 g4116 ( .a(n10845), .b(n10844), .o(n6929) );
in01f01 g4117 ( .a(_net_114), .o(n10847) );
na02f01 g4118 ( .a(net_310), .b(_net_154), .o(n10848) );
oa12f01 g4119 ( .a(n10848), .b(n10847), .c(_net_154), .o(n6938) );
in01f01 g4120 ( .a(_net_7589), .o(n10850) );
na02f01 g4121 ( .a(n7449), .b(n6968), .o(n10851) );
oa12f01 g4122 ( .a(n10851), .b(n6968), .c(n10850), .o(n6943) );
in01f01 g4123 ( .a(_net_7500), .o(n10853) );
na02f01 g4124 ( .a(n7952), .b(n7626_1), .o(n10854) );
oa12f01 g4125 ( .a(n10854), .b(n7626_1), .c(n10853), .o(n6952) );
no02f01 g4126 ( .a(n10132_1), .b(n6945), .o(n10856) );
no02f01 g4127 ( .a(n7042), .b(n6934_1), .o(n10857) );
in01f01 g4128 ( .a(_net_6098), .o(n10858) );
oa22f01 g4129 ( .a(n7050), .b(n6916), .c(n6932), .d(n10858), .o(n10859) );
no03f01 g4130 ( .a(n10859), .b(n10857), .c(n10856), .o(n10860) );
in01f01 g4131 ( .a(net_6617), .o(n10861) );
in01f01 g4132 ( .a(net_6585), .o(n10862) );
oa22f01 g4133 ( .a(n7058_1), .b(n10862), .c(n7057), .d(n10861), .o(n10863) );
in01f01 g4134 ( .a(net_6681), .o(n10864) );
in01f01 g4135 ( .a(net_6649), .o(n10865) );
oa22f01 g4136 ( .a(n7063), .b(n10864), .c(n7062_1), .d(n10865), .o(n10866) );
no02f01 g4137 ( .a(n10866), .b(n10863), .o(n10867) );
na02f01 g4138 ( .a(n10867), .b(n10860), .o(n6964) );
ao22f01 g4139 ( .a(n7225), .b(_net_7402), .c(n7224), .d(_net_7434), .o(n10869) );
ao22f01 g4140 ( .a(n7229), .b(_net_7498), .c(n7228), .d(_net_7466), .o(n10870) );
na02f01 g4141 ( .a(n10870), .b(n10869), .o(n6969) );
in01f01 g4142 ( .a(_net_7256), .o(n10872) );
na02f01 g4143 ( .a(n8208), .b(n6901), .o(n10873) );
oa12f01 g4144 ( .a(n10873), .b(n6901), .c(n10872), .o(n6995) );
na02f01 g4145 ( .a(n7440), .b(_net_7804), .o(n10875) );
oa12f01 g4146 ( .a(n10875), .b(n7440), .c(n8192_1), .o(n7000) );
in01f01 g4147 ( .a(_net_7408), .o(n10877) );
na02f01 g4148 ( .a(n8141), .b(n7550), .o(n10878) );
oa12f01 g4149 ( .a(n10878), .b(n7550), .c(n10877), .o(n7013) );
no02f01 g4150 ( .a(n10249), .b(n6824), .o(n10880) );
no02f01 g4151 ( .a(n9127), .b(n6826_1), .o(n10881) );
in01f01 g4152 ( .a(_net_6140), .o(n10882) );
oa22f01 g4153 ( .a(n9135), .b(n6836_1), .c(n6844), .d(n10882), .o(n10883) );
no03f01 g4154 ( .a(n10883), .b(n10881), .c(n10880), .o(n10884) );
in01f01 g4155 ( .a(net_6857), .o(n10885) );
in01f01 g4156 ( .a(net_6889), .o(n10886) );
oa22f01 g4157 ( .a(n6850_1), .b(n10885), .c(n6849), .d(n10886), .o(n10887) );
in01f01 g4158 ( .a(net_6953), .o(n10888) );
in01f01 g4159 ( .a(net_6921), .o(n10889) );
oa22f01 g4160 ( .a(n6855_1), .b(n10888), .c(n6854), .d(n10889), .o(n10890) );
no02f01 g4161 ( .a(n10890), .b(n10887), .o(n10891) );
na02f01 g4162 ( .a(n10891), .b(n10884), .o(n7018) );
ao22f01 g4163 ( .a(n7225), .b(_net_7430), .c(n7224), .d(net_7462), .o(n10893) );
ao22f01 g4164 ( .a(n7229), .b(net_7526), .c(n7228), .d(net_7494), .o(n10894) );
na02f01 g4165 ( .a(n10894), .b(n10893), .o(n7023) );
in01f01 g4166 ( .a(_net_7298), .o(n10896) );
na02f01 g4167 ( .a(n7242), .b(n7180), .o(n10897) );
oa12f01 g4168 ( .a(n10897), .b(n7180), .c(n10896), .o(n7032) );
in01f01 g4169 ( .a(_net_7579), .o(n10899) );
na02f01 g4170 ( .a(n1163), .b(n7519), .o(n10900) );
oa12f01 g4171 ( .a(n10900), .b(n7519), .c(n10899), .o(n7053) );
in01f01 g4172 ( .a(_net_7268), .o(n10902) );
na02f01 g4173 ( .a(n7256_1), .b(n6901), .o(n10903) );
oa12f01 g4174 ( .a(n10903), .b(n6901), .c(n10902), .o(n7058) );
no02f01 g4175 ( .a(n7477), .b(n7468_1), .o(n10905) );
no02f01 g4176 ( .a(n7486), .b(n7470), .o(n10906) );
in01f01 g4177 ( .a(_net_6122), .o(n10907) );
no02f01 g4178 ( .a(n8988), .b(n8985), .o(n10908) );
oa22f01 g4179 ( .a(n10908), .b(n7123), .c(n7118), .d(n10907), .o(n10909) );
no03f01 g4180 ( .a(n10909), .b(n10906), .c(n10905), .o(n10910) );
in01f01 g4181 ( .a(net_6724), .o(n10911) );
in01f01 g4182 ( .a(net_6756), .o(n10912) );
oa22f01 g4183 ( .a(n7492_1), .b(n10911), .c(n7491), .d(n10912), .o(n10913) );
in01f01 g4184 ( .a(net_6788), .o(n10914) );
in01f01 g4185 ( .a(net_6820), .o(n10915) );
oa22f01 g4186 ( .a(n7497), .b(n10915), .c(n7496_1), .d(n10914), .o(n10916) );
no02f01 g4187 ( .a(n10916), .b(n10913), .o(n10917) );
na02f01 g4188 ( .a(n10917), .b(n10910), .o(n7067) );
no02f01 g4189 ( .a(n6896), .b(n6895_1), .o(n7072) );
in01f01 g4190 ( .a(_net_6284), .o(n10920) );
no02f01 g4191 ( .a(_net_392), .b(n10920), .o(n7077) );
ao22f01 g4192 ( .a(n7225), .b(_net_7401), .c(n7224), .d(_net_7433), .o(n10922) );
ao22f01 g4193 ( .a(n7229), .b(_net_7497), .c(n7228), .d(_net_7465), .o(n10923) );
na02f01 g4194 ( .a(n10923), .b(n10922), .o(n7102) );
in01f01 g4195 ( .a(net_7767), .o(n10925) );
na02f01 g4196 ( .a(net_7769), .b(n8997), .o(n10926) );
oa12f01 g4197 ( .a(n10926), .b(n10206), .c(n10925), .o(n7107) );
in01f01 g4198 ( .a(_net_7705), .o(n10928) );
na02f01 g4199 ( .a(n7207_1), .b(net_7807), .o(n10929) );
oa12f01 g4200 ( .a(n10929), .b(n7207_1), .c(n10928), .o(n7133) );
in01f01 g4201 ( .a(_net_5848), .o(n10931) );
ao12f01 g4202 ( .a(n10925), .b(n10206), .c(n10931), .o(n7138) );
na02f01 g4203 ( .a(n7291), .b(_net_7719), .o(n10933) );
na02f01 g4204 ( .a(n7293), .b(_net_221), .o(n10934) );
ao22f01 g4205 ( .a(n7297_1), .b(_net_184), .c(n7296), .d(net_258), .o(n10935) );
ao22f01 g4206 ( .a(n7306), .b(_net_6021), .c(n7298), .d(_net_7748), .o(n10936) );
na04f01 g4207 ( .a(n10936), .b(n10935), .c(n10934), .d(n10933), .o(n7164) );
na02f01 g4208 ( .a(n6801_1), .b(x1261), .o(n10938) );
no02f01 g4209 ( .a(n10938), .b(n8317), .o(n7172) );
ao22f01 g4210 ( .a(n6877), .b(_net_7255), .c(n6876_1), .d(_net_7319), .o(n10940) );
ao22f01 g4211 ( .a(n6881_1), .b(_net_7287), .c(n6880), .d(_net_7351), .o(n10941) );
na02f01 g4212 ( .a(n10941), .b(n10940), .o(n7177) );
na02f01 g4213 ( .a(n8861), .b(n7768_1), .o(n10943) );
na02f01 g4214 ( .a(n6755), .b(n6748), .o(n10944) );
ao22f01 g4215 ( .a(n10944), .b(n8859), .c(n8862), .d(_net_6554), .o(n10945) );
na02f01 g4216 ( .a(n10945), .b(n10943), .o(n7194) );
no02f01 g4217 ( .a(n9233_1), .b(n6764), .o(n10947) );
no02f01 g4218 ( .a(n6766), .b(n6757), .o(n10948) );
in01f01 g4219 ( .a(_net_6080), .o(n10949) );
oa22f01 g4220 ( .a(n6784), .b(n10949), .c(n6775), .d(n6773), .o(n10950) );
no03f01 g4221 ( .a(n10950), .b(n10948), .c(n10947), .o(n10951) );
in01f01 g4222 ( .a(net_6452), .o(n10952) );
in01f01 g4223 ( .a(net_6484), .o(n10953) );
oa22f01 g4224 ( .a(n6790), .b(n10952), .c(n6789), .d(n10953), .o(n10954) );
in01f01 g4225 ( .a(net_6548), .o(n10955) );
in01f01 g4226 ( .a(net_6516), .o(n10956) );
oa22f01 g4227 ( .a(n6795), .b(n10955), .c(n6794), .d(n10956), .o(n10957) );
no02f01 g4228 ( .a(n10957), .b(n10954), .o(n10958) );
na02f01 g4229 ( .a(n10958), .b(n10951), .o(n7207) );
in01f01 g4230 ( .a(_net_7361), .o(n10960) );
na02f01 g4231 ( .a(n9537_1), .b(n7030), .o(n10961) );
oa12f01 g4232 ( .a(n10961), .b(n7030), .c(n10960), .o(n7216) );
in01f01 g4233 ( .a(_net_6210), .o(n10963) );
no02f01 g4234 ( .a(_net_392), .b(n10963), .o(n7221) );
in01f01 g4235 ( .a(_net_6239), .o(n10965) );
no02f01 g4236 ( .a(_net_392), .b(n10965), .o(n7226) );
in01f01 g4237 ( .a(_net_6294), .o(n10967) );
no02f01 g4238 ( .a(_net_392), .b(n10967), .o(n7235) );
na02f01 g4239 ( .a(n6996), .b(_net_6145), .o(n10969) );
na02f01 g4240 ( .a(n7327), .b(n6981), .o(n10970) );
na02f01 g4241 ( .a(n10970), .b(n10969), .o(n7240) );
na02f01 g4242 ( .a(n9667), .b(n9404), .o(n10972) );
na03f01 g4243 ( .a(n9665), .b(_net_6423), .c(_net_6422), .o(n10973) );
na03f01 g4244 ( .a(n10973), .b(n10972), .c(n9410_1), .o(n10974) );
oa12f01 g4245 ( .a(n10974), .b(n9409), .c(n9404), .o(n7245) );
oa12f01 g4246 ( .a(n6981), .b(n8051_1), .c(n8048), .o(n10977) );
ao22f01 g4247 ( .a(n10473), .b(n6998), .c(n6996), .d(_net_6151), .o(n10978) );
na02f01 g4248 ( .a(n8482), .b(n8481_1), .o(n10979) );
ao22f01 g4249 ( .a(n10979), .b(n7022), .c(n7323), .d(n7013_1), .o(n10980) );
na03f01 g4250 ( .a(n10980), .b(n10978), .c(n10977), .o(n7270) );
in01f01 g4251 ( .a(_net_6290), .o(n10982) );
no02f01 g4252 ( .a(_net_392), .b(n10982), .o(n7275) );
oa12f01 g4253 ( .a(n7335_1), .b(n6821), .c(n7687), .o(n7280) );
na02f01 g4254 ( .a(n6803), .b(_net_6028), .o(n10985) );
oa12f01 g4255 ( .a(n10985), .b(n6803), .c(n7330_1), .o(n7297) );
in01f01 g4256 ( .a(_net_6287), .o(n10987) );
no02f01 g4257 ( .a(n10987), .b(_net_392), .o(n7302) );
in01f01 g4258 ( .a(_net_7697), .o(n10989) );
na02f01 g4259 ( .a(n7207_1), .b(net_7799), .o(n10990) );
oa12f01 g4260 ( .a(n10990), .b(n7207_1), .c(n10989), .o(n7307) );
in01f01 g4261 ( .a(_net_7365), .o(n10992) );
na02f01 g4262 ( .a(n9685), .b(n7030), .o(n10993) );
oa12f01 g4263 ( .a(n10993), .b(n7030), .c(n10992), .o(n7321) );
no02f01 g4264 ( .a(n8282), .b(n7721), .o(n10995) );
no02f01 g4265 ( .a(n8291), .b(n7592), .o(n10996) );
in01f01 g4266 ( .a(_net_6179), .o(n10997) );
oa22f01 g4267 ( .a(n10436), .b(n7574), .c(n7590), .d(n10997), .o(n10998) );
no03f01 g4268 ( .a(n10998), .b(n10996), .c(n10995), .o(n10999) );
in01f01 g4269 ( .a(net_7126), .o(n11000) );
in01f01 g4270 ( .a(net_7158), .o(n11001) );
oa22f01 g4271 ( .a(n7740), .b(n11000), .c(n7739), .d(n11001), .o(n11002) );
in01f01 g4272 ( .a(net_7222), .o(n11003) );
in01f01 g4273 ( .a(net_7190), .o(n11004) );
oa22f01 g4274 ( .a(n7745), .b(n11003), .c(n7744), .d(n11004), .o(n11005) );
no02f01 g4275 ( .a(n11005), .b(n11002), .o(n11006) );
na02f01 g4276 ( .a(n11006), .b(n10999), .o(n7340) );
ao22f01 g4277 ( .a(n6736_1), .b(net_7636), .c(n6734), .d(net_7604), .o(n11008) );
ao22f01 g4278 ( .a(n6739), .b(net_7668), .c(n6738), .d(_net_7572), .o(n11009) );
na02f01 g4279 ( .a(n11009), .b(n11008), .o(n7354) );
ao22f01 g4280 ( .a(n6877), .b(_net_7279), .c(n6876_1), .d(net_7343), .o(n11011) );
ao22f01 g4281 ( .a(n6881_1), .b(net_7311), .c(n6880), .d(net_7375), .o(n11012) );
na02f01 g4282 ( .a(n11012), .b(n11011), .o(n7363) );
in01f01 g4283 ( .a(_net_7666), .o(n11014) );
na02f01 g4284 ( .a(n7892), .b(n7446_1), .o(n11015) );
oa12f01 g4285 ( .a(n11015), .b(n7446_1), .c(n11014), .o(n7381) );
na02f01 g4286 ( .a(n7119), .b(_net_6105), .o(n11017) );
na02f01 g4287 ( .a(n8187), .b(n7124), .o(n11018) );
na02f01 g4288 ( .a(n11018), .b(n11017), .o(n7386) );
in01f01 g4289 ( .a(_net_117), .o(n11020) );
na02f01 g4290 ( .a(net_313), .b(_net_154), .o(n11021) );
oa12f01 g4291 ( .a(n11021), .b(n11020), .c(_net_154), .o(n7395) );
in01f01 g4292 ( .a(_net_7473), .o(n11023) );
na02f01 g4293 ( .a(n7200), .b(n6869), .o(n11024) );
oa12f01 g4294 ( .a(n11024), .b(n6869), .c(n11023), .o(n7400) );
no02f01 g4295 ( .a(n6821), .b(n6819), .o(n11026) );
na03f01 g4296 ( .a(n6823), .b(n8344), .c(_net_6957), .o(n11027) );
na02f01 g4297 ( .a(n6823), .b(n8344), .o(n11028) );
na02f01 g4298 ( .a(n11028), .b(n6818_1), .o(n11029) );
na03f01 g4299 ( .a(n11029), .b(n11027), .c(n11026), .o(n11030) );
na02f01 g4300 ( .a(n8345_1), .b(_net_6957), .o(n11031) );
na02f01 g4301 ( .a(n11031), .b(n11030), .o(n7422) );
no02f01 g4302 ( .a(n7232), .b(n7158), .o(n7432) );
na02f01 g4303 ( .a(n10463), .b(n8028_1), .o(n11034) );
ao22f01 g4304 ( .a(n8031), .b(n8033_1), .c(n8034), .d(_net_6069), .o(n11035) );
na02f01 g4305 ( .a(n8037), .b(n8110), .o(n11036) );
oa12f01 g4306 ( .a(n8113), .b(n9046), .c(n9043), .o(n11037) );
na04f01 g4307 ( .a(n11037), .b(n11036), .c(n11035), .d(n11034), .o(n7437) );
in01f01 g4308 ( .a(_net_6007), .o(n11039) );
na02f01 g4309 ( .a(n7348), .b(_net_7810), .o(n11040) );
oa12f01 g4310 ( .a(n11040), .b(n7348), .c(n11039), .o(n7454) );
in01f01 g4311 ( .a(_net_7263), .o(n11042) );
na02f01 g4312 ( .a(n7994_1), .b(n6901), .o(n11043) );
oa12f01 g4313 ( .a(n11043), .b(n6901), .c(n11042), .o(n7459) );
in01f01 g4314 ( .a(_net_6221), .o(n11045) );
no02f01 g4315 ( .a(_net_392), .b(n11045), .o(n7473) );
in01f01 g4316 ( .a(_net_7351), .o(n11047) );
na02f01 g4317 ( .a(n8022), .b(n7030), .o(n11048) );
oa12f01 g4318 ( .a(n11048), .b(n7030), .c(n11047), .o(n7478) );
no02f01 g4319 ( .a(_net_6962), .b(n8252), .o(n11050) );
no02f01 g4320 ( .a(n8253_1), .b(net_6961), .o(n11051) );
no02f01 g4321 ( .a(n11051), .b(n11050), .o(n11052) );
oa22f01 g4322 ( .a(n11052), .b(n8250), .c(n8256), .d(n8253_1), .o(n7487) );
na02f01 g4323 ( .a(n8108), .b(n8028_1), .o(n11054) );
ao22f01 g4324 ( .a(n8116_1), .b(n8033_1), .c(n8034), .d(_net_6068), .o(n11055) );
na02f01 g4325 ( .a(n9810), .b(n8110), .o(n11056) );
oa12f01 g4326 ( .a(n8113), .b(n6772), .c(n6769), .o(n11057) );
na04f01 g4327 ( .a(n11057), .b(n11056), .c(n11055), .d(n11054), .o(n7496) );
no04f01 g4328 ( .a(n7340_1), .b(n7782), .c(n7294), .d(n7281), .o(n7501) );
in01f01 g4329 ( .a(_net_7471), .o(n11060) );
na02f01 g4330 ( .a(n7387), .b(n6869), .o(n11061) );
oa12f01 g4331 ( .a(n11061), .b(n6869), .c(n11060), .o(n7518) );
ao22f01 g4332 ( .a(n7288_1), .b(_net_6045), .c(n7286), .d(_net_284), .o(n11063) );
ao22f01 g4333 ( .a(n7298), .b(_net_7734), .c(n7291), .d(_net_7705), .o(n11064) );
na02f01 g4334 ( .a(n7302_1), .b(_net_128), .o(n11065) );
na03f01 g4335 ( .a(n7308), .b(net_207), .c(x1322), .o(n11066) );
na02f01 g4336 ( .a(n7296), .b(net_244), .o(n11067) );
na03f01 g4337 ( .a(n7308), .b(net_170), .c(n6800), .o(n11068) );
na03f01 g4338 ( .a(n11068), .b(n11067), .c(n11066), .o(n11069) );
ao12f01 g4339 ( .a(n11069), .b(n7306), .c(_net_6001), .o(n11070) );
na04f01 g4340 ( .a(n11070), .b(n11065), .c(n11064), .d(n11063), .o(n7539) );
ao22f01 g4341 ( .a(n6877), .b(_net_7271), .c(n6876_1), .d(net_7335), .o(n11072) );
ao22f01 g4342 ( .a(n6881_1), .b(net_7303), .c(n6880), .d(net_7367), .o(n11073) );
na02f01 g4343 ( .a(n11073), .b(n11072), .o(n7543) );
ao22f01 g4344 ( .a(n6736_1), .b(_net_7629), .c(n6734), .d(_net_7597), .o(n11075) );
ao22f01 g4345 ( .a(n6739), .b(_net_7661), .c(n6738), .d(_net_7565), .o(n11076) );
na02f01 g4346 ( .a(n11076), .b(n11075), .o(n7548) );
in01f01 g4347 ( .a(n9860), .o(n11078) );
na02f01 g4348 ( .a(n6899_1), .b(n9854), .o(n11079) );
na02f01 g4349 ( .a(n6898), .b(_net_7381), .o(n11080) );
na02f01 g4350 ( .a(n11080), .b(n11079), .o(n11081) );
oa22f01 g4351 ( .a(n11081), .b(n9857), .c(n11078), .d(n9854), .o(n7558) );
in01f01 g4352 ( .a(_net_7293), .o(n11083) );
na02f01 g4353 ( .a(n8809_1), .b(n7180), .o(n11084) );
oa12f01 g4354 ( .a(n11084), .b(n7180), .c(n11083), .o(n7563) );
na02f01 g4355 ( .a(n10708), .b(n8213), .o(n11086) );
ao22f01 g4356 ( .a(n8216_1), .b(n9200), .c(n8211_1), .d(_net_6127), .o(n11087) );
na02f01 g4357 ( .a(n11087), .b(n11086), .o(n7572) );
in01f01 g4358 ( .a(_net_7798), .o(n11089) );
na02f01 g4359 ( .a(n6803), .b(_net_6033), .o(n11090) );
oa12f01 g4360 ( .a(n11090), .b(n6803), .c(n11089), .o(n7586) );
in01f01 g4361 ( .a(_net_127), .o(n11092) );
na02f01 g4362 ( .a(_net_154), .b(net_323), .o(n11093) );
oa12f01 g4363 ( .a(n11093), .b(n11092), .c(_net_154), .o(n7591) );
na03f01 g4364 ( .a(n9707), .b(n9706), .c(_net_6022), .o(n11095) );
na02f01 g4365 ( .a(n7293), .b(net_222), .o(n11096) );
ao22f01 g4366 ( .a(n7297_1), .b(net_185), .c(n7296), .d(net_259), .o(n11097) );
na03f01 g4367 ( .a(n11097), .b(n11096), .c(n11095), .o(n7596) );
na02f01 g4368 ( .a(n8544_1), .b(n8338), .o(n11099) );
na02f01 g4369 ( .a(n6815), .b(n6807), .o(n11100) );
ao22f01 g4370 ( .a(n11100), .b(n8340_1), .c(n8345_1), .d(_net_6959), .o(n11101) );
na02f01 g4371 ( .a(n11101), .b(n11099), .o(n7608) );
ao22f01 g4372 ( .a(n7225), .b(_net_7407), .c(n7224), .d(_net_7439), .o(n11103) );
ao22f01 g4373 ( .a(n7229), .b(_net_7503), .c(n7228), .d(_net_7471), .o(n11104) );
na02f01 g4374 ( .a(n11104), .b(n11103), .o(n7613) );
in01f01 g4375 ( .a(_net_6206), .o(n11106) );
no02f01 g4376 ( .a(_net_392), .b(n11106), .o(n7622) );
in01f01 g4377 ( .a(_net_7331), .o(n11108) );
na02f01 g4378 ( .a(n7567_1), .b(n7150), .o(n11109) );
oa12f01 g4379 ( .a(n11109), .b(n7150), .c(n11108), .o(n7631) );
na02f01 g4380 ( .a(n7348), .b(_net_7805), .o(n11111) );
oa12f01 g4381 ( .a(n11111), .b(n7348), .c(n10621), .o(n7640) );
in01f01 g4382 ( .a(_net_6298), .o(n11113) );
no02f01 g4383 ( .a(n11113), .b(_net_392), .o(n7649) );
na02f01 g4384 ( .a(n8310), .b(n7576), .o(n11115) );
ao22f01 g4385 ( .a(n9111), .b(n8307_1), .c(n8312), .d(_net_7228), .o(n11116) );
na02f01 g4386 ( .a(n11116), .b(n11115), .o(n7666) );
oa12f01 g4387 ( .a(n6917), .b(n7804), .c(n7801), .o(n11118) );
ao22f01 g4388 ( .a(n6923), .b(net_6564), .c(n6920), .d(net_6628), .o(n11119) );
ao22f01 g4389 ( .a(n6928), .b(net_6596), .c(n6926), .d(net_6660), .o(n11120) );
na02f01 g4390 ( .a(n11120), .b(n11119), .o(n11121) );
ao22f01 g4391 ( .a(n11121), .b(n6935), .c(n6933), .d(_net_6091), .o(n11122) );
in01f01 g4392 ( .a(net_6578), .o(n11123) );
in01f01 g4393 ( .a(net_6642), .o(n11124) );
oa22f01 g4394 ( .a(n6922), .b(n11123), .c(n6919_1), .d(n11124), .o(n11125) );
in01f01 g4395 ( .a(net_6674), .o(n11126) );
in01f01 g4396 ( .a(net_6610), .o(n11127) );
oa22f01 g4397 ( .a(n6927), .b(n11127), .c(n6925), .d(n11126), .o(n11128) );
no02f01 g4398 ( .a(n11128), .b(n11125), .o(n11129) );
no03f01 g4399 ( .a(n11129), .b(n6947_1), .c(n6943_1), .o(n11130) );
ao12f01 g4400 ( .a(n11130), .b(n8005_1), .c(n6946), .o(n11131) );
na03f01 g4401 ( .a(n11131), .b(n11122), .c(n11118), .o(n7671) );
no02f01 g4402 ( .a(n10494), .b(n6945), .o(n11133) );
no02f01 g4403 ( .a(n10592), .b(n6934_1), .o(n11134) );
in01f01 g4404 ( .a(_net_6103), .o(n11135) );
oa22f01 g4405 ( .a(n11129), .b(n6916), .c(n6932), .d(n11135), .o(n11136) );
no03f01 g4406 ( .a(n11136), .b(n11134), .c(n11133), .o(n11137) );
in01f01 g4407 ( .a(net_6590), .o(n11138) );
in01f01 g4408 ( .a(net_6622), .o(n11139) );
oa22f01 g4409 ( .a(n7058_1), .b(n11138), .c(n7057), .d(n11139), .o(n11140) );
in01f01 g4410 ( .a(net_6654), .o(n11141) );
in01f01 g4411 ( .a(net_6686), .o(n11142) );
oa22f01 g4412 ( .a(n7063), .b(n11142), .c(n7062_1), .d(n11141), .o(n11143) );
no02f01 g4413 ( .a(n11143), .b(n11140), .o(n11144) );
na02f01 g4414 ( .a(n11144), .b(n11137), .o(n7676) );
in01f01 g4415 ( .a(_net_125), .o(n11146) );
na02f01 g4416 ( .a(net_321), .b(_net_154), .o(n11147) );
oa12f01 g4417 ( .a(n11147), .b(n11146), .c(_net_154), .o(n7681) );
ao22f01 g4418 ( .a(n6738), .b(_net_7553), .c(n6736_1), .d(_net_7617), .o(n11149) );
ao22f01 g4419 ( .a(n6739), .b(_net_7649), .c(n6734), .d(_net_7585), .o(n11150) );
na02f01 g4420 ( .a(n11150), .b(n11149), .o(n7686) );
na02f01 g4421 ( .a(n7348), .b(_net_7801), .o(n11152) );
oa12f01 g4422 ( .a(n11152), .b(n7348), .c(n6912), .o(n7695) );
no03f01 g4423 ( .a(_net_6043), .b(n7570), .c(n8699), .o(n11154) );
no02f01 g4424 ( .a(n7570), .b(n8695), .o(n11155) );
ao22f01 g4425 ( .a(n11155), .b(n8705), .c(n11154), .d(n8703_1), .o(n11156) );
ao12f01 g4426 ( .a(n7570), .b(_net_5982), .c(n8695), .o(n11157) );
no03f01 g4427 ( .a(_net_6043), .b(n7570), .c(_net_6044), .o(n11158) );
ao22f01 g4428 ( .a(n11158), .b(n8701), .c(n11157), .d(n8694_1), .o(n11159) );
na02f01 g4429 ( .a(n11159), .b(n11156), .o(n7709) );
in01f01 g4430 ( .a(_net_7273), .o(n11161) );
na02f01 g4431 ( .a(n518), .b(n6901), .o(n11162) );
oa12f01 g4432 ( .a(n11162), .b(n6901), .c(n11161), .o(n7723) );
in01f01 g4433 ( .a(_net_7289), .o(n11164) );
na02f01 g4434 ( .a(n9587), .b(n7180), .o(n11165) );
oa12f01 g4435 ( .a(n11165), .b(n7180), .c(n11164), .o(n7728) );
ao22f01 g4436 ( .a(n7288_1), .b(_net_6043), .c(n7286), .d(_net_282), .o(n11167) );
ao22f01 g4437 ( .a(n7298), .b(_net_7732), .c(n7291), .d(_net_7703), .o(n11168) );
na02f01 g4438 ( .a(n7302_1), .b(_net_126), .o(n11169) );
na03f01 g4439 ( .a(n7308), .b(net_205), .c(x1322), .o(n11170) );
na02f01 g4440 ( .a(n7296), .b(net_242), .o(n11171) );
na03f01 g4441 ( .a(n7308), .b(net_168), .c(n6800), .o(n11172) );
na03f01 g4442 ( .a(n11172), .b(n11171), .c(n11170), .o(n11173) );
ao12f01 g4443 ( .a(n11173), .b(n7306), .c(_net_5999), .o(n11174) );
na04f01 g4444 ( .a(n11174), .b(n11169), .c(n11168), .d(n11167), .o(n7737) );
no02f01 g4445 ( .a(n10333), .b(n10331), .o(n7741) );
ao12f01 g4446 ( .a(n9607), .b(net_6826), .c(_net_6827), .o(n11177) );
no03f01 g4447 ( .a(_net_6828), .b(n8220_1), .c(n8219), .o(n11178) );
no02f01 g4448 ( .a(n11178), .b(n11177), .o(n11179) );
oa22f01 g4449 ( .a(n11179), .b(n8226), .c(n8227), .d(n9607), .o(n7746) );
in01f01 g4450 ( .a(_net_7555), .o(n11181) );
na02f01 g4451 ( .a(n9154), .b(n7519), .o(n11182) );
oa12f01 g4452 ( .a(n11182), .b(n7519), .c(n11181), .o(n7751) );
in01f01 g4453 ( .a(_net_7699), .o(n11184) );
na02f01 g4454 ( .a(n7207_1), .b(_net_7801), .o(n11185) );
oa12f01 g4455 ( .a(n11185), .b(n7207_1), .c(n11184), .o(n7768) );
na02f01 g4456 ( .a(n7298), .b(_net_7736), .o(n11187) );
ao22f01 g4457 ( .a(n7306), .b(_net_6006), .c(n7291), .d(_net_7707), .o(n11188) );
na02f01 g4458 ( .a(n7302_1), .b(net_146), .o(n11189) );
na02f01 g4459 ( .a(n7296), .b(net_246), .o(n11190) );
na03f01 g4460 ( .a(n7308), .b(_net_172), .c(n6800), .o(n11191) );
na03f01 g4461 ( .a(n7308), .b(_net_209), .c(x1322), .o(n11192) );
na03f01 g4462 ( .a(n11192), .b(n11191), .c(n11190), .o(n11193) );
ao12f01 g4463 ( .a(n11193), .b(n7286), .c(_net_289), .o(n11194) );
na04f01 g4464 ( .a(n11194), .b(n11189), .c(n11188), .d(n11187), .o(n7773) );
ao12f01 g4465 ( .a(n6945), .b(n11120), .c(n11119), .o(n11196) );
no02f01 g4466 ( .a(n7805), .b(n6934_1), .o(n11197) );
in01f01 g4467 ( .a(_net_6093), .o(n11198) );
oa22f01 g4468 ( .a(n7813), .b(n6916), .c(n6932), .d(n11198), .o(n11199) );
no03f01 g4469 ( .a(n11199), .b(n11197), .c(n11196), .o(n11200) );
in01f01 g4470 ( .a(net_6612), .o(n11201) );
in01f01 g4471 ( .a(net_6580), .o(n11202) );
oa22f01 g4472 ( .a(n7058_1), .b(n11202), .c(n7057), .d(n11201), .o(n11203) );
in01f01 g4473 ( .a(net_6676), .o(n11204) );
in01f01 g4474 ( .a(net_6644), .o(n11205) );
oa22f01 g4475 ( .a(n7063), .b(n11204), .c(n7062_1), .d(n11205), .o(n11206) );
no02f01 g4476 ( .a(n11206), .b(n11203), .o(n11207) );
na02f01 g4477 ( .a(n11207), .b(n11200), .o(n7788) );
in01f01 g4478 ( .a(_net_6049), .o(n11209) );
ao12f01 g4479 ( .a(n9253), .b(_net_7230), .c(_net_7233), .o(n11210) );
oa12f01 g4480 ( .a(n11210), .b(_net_7230), .c(_net_7233), .o(n11211) );
na02f01 g4481 ( .a(n10338), .b(n4276), .o(n11212) );
oa12f01 g4482 ( .a(n11209), .b(n11212), .c(n11211), .o(n7793) );
in01f01 g4483 ( .a(_net_7442), .o(n11214) );
na02f01 g4484 ( .a(n7197), .b(n6891), .o(n11215) );
oa12f01 g4485 ( .a(n11215), .b(n7197), .c(n11214), .o(n7798) );
no02f01 g4486 ( .a(n6809_1), .b(_net_6962), .o(n11217) );
no02f01 g4487 ( .a(_net_6959), .b(n8253_1), .o(n11218) );
no02f01 g4488 ( .a(n11218), .b(n11217), .o(n11219) );
no02f01 g4489 ( .a(n6806_1), .b(net_6961), .o(n11220) );
no02f01 g4490 ( .a(n11220), .b(n11219), .o(n11221) );
no04f01 g4491 ( .a(n11218), .b(n11217), .c(n6806_1), .d(net_6961), .o(n11222) );
no02f01 g4492 ( .a(n6806_1), .b(n8252), .o(n11223) );
no02f01 g4493 ( .a(_net_6958), .b(net_6961), .o(n11224) );
no02f01 g4494 ( .a(n11224), .b(n11223), .o(n11225) );
oa12f01 g4495 ( .a(n11225), .b(n11222), .c(n11221), .o(n11226) );
no02f01 g4496 ( .a(n11222), .b(n11221), .o(n11227) );
in01f01 g4497 ( .a(n11225), .o(n9778) );
na02f01 g4498 ( .a(n9778), .b(n11227), .o(n11229) );
na02f01 g4499 ( .a(n11229), .b(n11226), .o(n7822) );
in01f01 g4500 ( .a(_net_7276), .o(n11231) );
na02f01 g4501 ( .a(n1639), .b(n6901), .o(n11232) );
oa12f01 g4502 ( .a(n11232), .b(n6901), .c(n11231), .o(n7835) );
na02f01 g4503 ( .a(n7291), .b(net_7715), .o(n11234) );
na02f01 g4504 ( .a(n7293), .b(_net_217), .o(n11235) );
ao22f01 g4505 ( .a(n7297_1), .b(_net_180), .c(n7296), .d(net_254), .o(n11236) );
ao22f01 g4506 ( .a(n7306), .b(_net_6017), .c(n7298), .d(net_7744), .o(n11237) );
na04f01 g4507 ( .a(n11237), .b(n11236), .c(n11235), .d(n11234), .o(n7845) );
ao22f01 g4508 ( .a(n7225), .b(_net_7408), .c(n7224), .d(_net_7440), .o(n11239) );
ao22f01 g4509 ( .a(n7229), .b(_net_7504), .c(n7228), .d(_net_7472), .o(n11240) );
na02f01 g4510 ( .a(n11240), .b(n11239), .o(n7853) );
no02f01 g4511 ( .a(n8317), .b(n9892), .o(n7858) );
na03f01 g4512 ( .a(n9260), .b(_net_6407), .c(_net_6408), .o(n11243) );
ao12f01 g4513 ( .a(x38), .b(n11243), .c(_net_6409), .o(n11244) );
oa12f01 g4514 ( .a(n11244), .b(n11243), .c(_net_6409), .o(n7863) );
in01f01 g4515 ( .a(_net_7484), .o(n11246) );
na02f01 g4516 ( .a(n9872), .b(n6869), .o(n11247) );
oa12f01 g4517 ( .a(n11247), .b(n6869), .c(n11246), .o(n7888) );
in01f01 g4518 ( .a(_net_5850), .o(n11249) );
in01f01 g4519 ( .a(x837), .o(n11250) );
na03f01 g4520 ( .a(n10203), .b(net_7780), .c(n11250), .o(n11251) );
oa12f01 g4521 ( .a(n11251), .b(n11249), .c(x837), .o(n7897) );
in01f01 g4522 ( .a(_net_7796), .o(n11253) );
na02f01 g4523 ( .a(n6803), .b(_net_6031), .o(n11254) );
oa12f01 g4524 ( .a(n11254), .b(n6803), .c(n11253), .o(n7902) );
na02f01 g4525 ( .a(n8857), .b(_net_6552), .o(n11256) );
na02f01 g4526 ( .a(n8856), .b(n6758), .o(n11257) );
na02f01 g4527 ( .a(n11257), .b(n11256), .o(n11258) );
na02f01 g4528 ( .a(n8862), .b(_net_6552), .o(n11259) );
oa12f01 g4529 ( .a(n11259), .b(n11258), .c(n8858), .o(n7911) );
ao22f01 g4530 ( .a(n6736_1), .b(_net_7623), .c(n6734), .d(_net_7591), .o(n11261) );
ao22f01 g4531 ( .a(n6739), .b(_net_7655), .c(n6738), .d(_net_7559), .o(n11262) );
na02f01 g4532 ( .a(n11262), .b(n11261), .o(n7933) );
in01f01 g4533 ( .a(net_7760), .o(n11264) );
na04f01 g4534 ( .a(_net_6039), .b(_net_7791), .c(net_303), .d(n11264), .o(n11265) );
ao12f01 g4535 ( .a(n11265), .b(net_304), .c(_net_6040), .o(n7950) );
in01f01 g4536 ( .a(_net_5855), .o(n11267) );
in01f01 g4537 ( .a(x977), .o(n11268) );
na03f01 g4538 ( .a(n9364), .b(net_7775), .c(n11268), .o(n11269) );
oa12f01 g4539 ( .a(n11269), .b(n11267), .c(x977), .o(n7975) );
ao22f01 g4540 ( .a(n6877), .b(_net_7252), .c(n6876_1), .d(_net_7316), .o(n11271) );
ao22f01 g4541 ( .a(n6881_1), .b(_net_7284), .c(n6880), .d(_net_7348), .o(n11272) );
na02f01 g4542 ( .a(n11272), .b(n11271), .o(n7980) );
in01f01 g4543 ( .a(_net_7425), .o(n11274) );
na02f01 g4544 ( .a(n2958), .b(n7550), .o(n11275) );
oa12f01 g4545 ( .a(n11275), .b(n7550), .c(n11274), .o(n7985) );
in01f01 g4546 ( .a(_net_5852), .o(n11277) );
in01f01 g4547 ( .a(x889), .o(n11278) );
no02f01 g4548 ( .a(n10034), .b(_net_272), .o(n11279) );
na02f01 g4549 ( .a(_net_267), .b(_net_273), .o(n11280) );
ao12f01 g4550 ( .a(n11280), .b(_net_192), .c(n9591), .o(n11281) );
na02f01 g4551 ( .a(n11281), .b(n11279), .o(n11282) );
in01f01 g4552 ( .a(n11280), .o(n11283) );
no02f01 g4553 ( .a(n10034), .b(n9019), .o(n11284) );
na03f01 g4554 ( .a(n11284), .b(n11283), .c(_net_189), .o(n11285) );
na03f01 g4555 ( .a(_net_192), .b(n9591), .c(_net_191), .o(n11286) );
na04f01 g4556 ( .a(n11286), .b(n11283), .c(n10034), .d(n9019), .o(n11287) );
oa12f01 g4557 ( .a(n9591), .b(_net_192), .c(_net_191), .o(n11288) );
na04f01 g4558 ( .a(n11288), .b(n11283), .c(n10034), .d(_net_272), .o(n11289) );
na04f01 g4559 ( .a(n11289), .b(n11287), .c(n11285), .d(n11282), .o(n11290) );
na03f01 g4560 ( .a(n11290), .b(net_7778), .c(n11278), .o(n11291) );
oa12f01 g4561 ( .a(n11291), .b(n11277), .c(x889), .o(n8010) );
in01f01 g4562 ( .a(_net_291), .o(n11293) );
na02f01 g4563 ( .a(n7440), .b(_net_7811), .o(n11294) );
oa12f01 g4564 ( .a(n11294), .b(n7440), .c(n11293), .o(n8019) );
in01f01 g4565 ( .a(_net_6286), .o(n11296) );
no02f01 g4566 ( .a(_net_392), .b(n11296), .o(n8024) );
ao12f01 g4567 ( .a(n6764), .b(n8107_1), .c(n8106), .o(n11298) );
no02f01 g4568 ( .a(n10546), .b(n6766), .o(n11299) );
in01f01 g4569 ( .a(_net_6072), .o(n11300) );
oa22f01 g4570 ( .a(n10554), .b(n6775), .c(n6784), .d(n11300), .o(n11301) );
no03f01 g4571 ( .a(n11301), .b(n11299), .c(n11298), .o(n11302) );
in01f01 g4572 ( .a(net_6476), .o(n11303) );
in01f01 g4573 ( .a(net_6444), .o(n11304) );
oa22f01 g4574 ( .a(n6790), .b(n11304), .c(n6789), .d(n11303), .o(n11305) );
in01f01 g4575 ( .a(net_6540), .o(n11306) );
in01f01 g4576 ( .a(net_6508), .o(n11307) );
oa22f01 g4577 ( .a(n6795), .b(n11306), .c(n6794), .d(n11307), .o(n11308) );
no02f01 g4578 ( .a(n11308), .b(n11305), .o(n11309) );
na02f01 g4579 ( .a(n11309), .b(n11302), .o(n8033) );
in01f01 g4580 ( .a(_net_7262), .o(n11311) );
na02f01 g4581 ( .a(n7926), .b(n6901), .o(n11312) );
oa12f01 g4582 ( .a(n11312), .b(n6901), .c(n11311), .o(n8080) );
in01f01 g4583 ( .a(_net_7573), .o(n11314) );
na02f01 g4584 ( .a(n7519), .b(n718), .o(n11315) );
oa12f01 g4585 ( .a(n11315), .b(n7519), .c(n11314), .o(n8097) );
in01f01 g4586 ( .a(_net_7499), .o(n11317) );
na02f01 g4587 ( .a(n9700_1), .b(n7626_1), .o(n11318) );
oa12f01 g4588 ( .a(n11318), .b(n7626_1), .c(n11317), .o(n8102) );
in01f01 g4589 ( .a(_net_7417), .o(n11320) );
na02f01 g4590 ( .a(n7550), .b(n6872_1), .o(n11321) );
oa12f01 g4591 ( .a(n11321), .b(n7550), .c(n11320), .o(n8107) );
no02f01 g4592 ( .a(n10745), .b(n7468_1), .o(n11323) );
no02f01 g4593 ( .a(n10754), .b(n7470), .o(n11324) );
in01f01 g4594 ( .a(_net_6115), .o(n11325) );
oa22f01 g4595 ( .a(n10660), .b(n7123), .c(n7118), .d(n11325), .o(n11326) );
no03f01 g4596 ( .a(n11326), .b(n11324), .c(n11323), .o(n11327) );
in01f01 g4597 ( .a(net_6717), .o(n11328) );
in01f01 g4598 ( .a(net_6749), .o(n11329) );
oa22f01 g4599 ( .a(n7492_1), .b(n11328), .c(n7491), .d(n11329), .o(n11330) );
in01f01 g4600 ( .a(net_6813), .o(n11331) );
in01f01 g4601 ( .a(net_6781), .o(n11332) );
oa22f01 g4602 ( .a(n7497), .b(n11331), .c(n7496_1), .d(n11332), .o(n11333) );
no02f01 g4603 ( .a(n11333), .b(n11330), .o(n11334) );
na02f01 g4604 ( .a(n11334), .b(n11327), .o(n8112) );
in01f01 g4605 ( .a(_net_7562), .o(n11336) );
na02f01 g4606 ( .a(n7707), .b(n7519), .o(n11337) );
oa12f01 g4607 ( .a(n11337), .b(n7519), .c(n11336), .o(n8121) );
in01f01 g4608 ( .a(_net_7291), .o(n11339) );
na02f01 g4609 ( .a(n7180), .b(n7033), .o(n11340) );
oa12f01 g4610 ( .a(n11340), .b(n7180), .c(n11339), .o(n8130) );
in01f01 g4611 ( .a(_net_7592), .o(n11342) );
na02f01 g4612 ( .a(n9881), .b(n6968), .o(n11343) );
oa12f01 g4613 ( .a(n11343), .b(n6968), .c(n11342), .o(n8135) );
no04f01 g4614 ( .a(n8362_1), .b(n8352), .c(n6966), .d(_net_7683), .o(n8152) );
ao22f01 g4615 ( .a(n6736_1), .b(_net_7628), .c(n6734), .d(_net_7596), .o(n11346) );
ao22f01 g4616 ( .a(n6739), .b(_net_7660), .c(n6738), .d(_net_7564), .o(n11347) );
na02f01 g4617 ( .a(n11347), .b(n11346), .o(n8161) );
ao22f01 g4618 ( .a(n7225), .b(_net_7429), .c(n7224), .d(net_7461), .o(n11349) );
ao22f01 g4619 ( .a(n7229), .b(net_7525), .c(n7228), .d(net_7493), .o(n11350) );
na02f01 g4620 ( .a(n11350), .b(n11349), .o(n8170) );
ao22f01 g4621 ( .a(n6877), .b(_net_7274), .c(n6876_1), .d(net_7338), .o(n11352) );
ao22f01 g4622 ( .a(n6881_1), .b(net_7306), .c(n6880), .d(net_7370), .o(n11353) );
na02f01 g4623 ( .a(n11353), .b(n11352), .o(n8179) );
in01f01 g4624 ( .a(_net_7275), .o(n11355) );
na02f01 g4625 ( .a(n2084), .b(n6901), .o(n11356) );
oa12f01 g4626 ( .a(n11356), .b(n6901), .c(n11355), .o(n8192) );
no03f01 g4627 ( .a(n8094), .b(_net_271), .c(n9019), .o(n11358) );
no02f01 g4628 ( .a(n8094), .b(n9591), .o(n11359) );
ao22f01 g4629 ( .a(n11359), .b(n11284), .c(n11358), .d(n11288), .o(n11360) );
ao12f01 g4630 ( .a(n8094), .b(_net_192), .c(n9591), .o(n11361) );
no03f01 g4631 ( .a(n8094), .b(_net_271), .c(_net_272), .o(n11362) );
ao22f01 g4632 ( .a(n11362), .b(n11286), .c(n11361), .d(n11279), .o(n11363) );
na02f01 g4633 ( .a(n11363), .b(n11360), .o(n8197) );
no02f01 g4634 ( .a(n8069), .b(n7012), .o(n11365) );
no02f01 g4635 ( .a(n9934), .b(n6997), .o(n11366) );
in01f01 g4636 ( .a(_net_6159), .o(n11367) );
oa22f01 g4637 ( .a(n8471), .b(n6980), .c(n6995_1), .d(n11367), .o(n11368) );
no03f01 g4638 ( .a(n11368), .b(n11366), .c(n11365), .o(n11369) );
in01f01 g4639 ( .a(net_6991), .o(n11370) );
in01f01 g4640 ( .a(net_7023), .o(n11371) );
oa22f01 g4641 ( .a(n8075_1), .b(n11370), .c(n8074), .d(n11371), .o(n11372) );
in01f01 g4642 ( .a(net_7055), .o(n11373) );
in01f01 g4643 ( .a(net_7087), .o(n11374) );
oa22f01 g4644 ( .a(n8080_1), .b(n11374), .c(n8079), .d(n11373), .o(n11375) );
no02f01 g4645 ( .a(n11375), .b(n11372), .o(n11376) );
na02f01 g4646 ( .a(n11376), .b(n11369), .o(n8202) );
na02f01 g4647 ( .a(_net_5990), .b(_net_5984), .o(n11378) );
ao12f01 g4648 ( .a(n11378), .b(_net_5962), .c(n7533), .o(n11379) );
na02f01 g4649 ( .a(n11379), .b(n7541), .o(n11380) );
in01f01 g4650 ( .a(n11378), .o(n11381) );
na04f01 g4651 ( .a(n11381), .b(n7543_1), .c(n7535_1), .d(n7538), .o(n11382) );
na04f01 g4652 ( .a(n11381), .b(n7534), .c(_net_5989), .d(n7538), .o(n11383) );
na03f01 g4653 ( .a(n11381), .b(n7539_1), .c(_net_5960), .o(n11384) );
na04f01 g4654 ( .a(n11384), .b(n11383), .c(n11382), .d(n11380), .o(n11385) );
in01f01 g4655 ( .a(n11385), .o(n11386) );
no02f01 g4656 ( .a(n11386), .b(x1062), .o(n8211) );
in01f01 g4657 ( .a(_net_7702), .o(n11388) );
na02f01 g4658 ( .a(n7207_1), .b(_net_7804), .o(n11389) );
oa12f01 g4659 ( .a(n11389), .b(n7207_1), .c(n11388), .o(n8216) );
no02f01 g4660 ( .a(n7161), .b(n7232), .o(n8224) );
in01f01 g4661 ( .a(_net_7580), .o(n11392) );
na02f01 g4662 ( .a(n5814), .b(n7519), .o(n11393) );
oa12f01 g4663 ( .a(n11393), .b(n7519), .c(n11392), .o(n8237) );
in01f01 g4664 ( .a(_net_7432), .o(n11395) );
na02f01 g4665 ( .a(n5552), .b(n7550), .o(n11396) );
oa12f01 g4666 ( .a(n11396), .b(n7550), .c(n11395), .o(n8253) );
ao22f01 g4667 ( .a(n7225), .b(_net_7404), .c(n7224), .d(_net_7436), .o(n11398) );
ao22f01 g4668 ( .a(n7229), .b(_net_7500), .c(n7228), .d(_net_7468), .o(n11399) );
na02f01 g4669 ( .a(n11399), .b(n11398), .o(n8258) );
na02f01 g4670 ( .a(n10016), .b(n10015), .o(n11401) );
na02f01 g4671 ( .a(n11401), .b(n10020), .o(n11402) );
oa22f01 g4672 ( .a(n11402), .b(n10014_1), .c(n10013), .d(n10016), .o(n8284) );
in01f01 g4673 ( .a(_net_7648), .o(n11404) );
na02f01 g4674 ( .a(n8842), .b(n7446_1), .o(n11405) );
oa12f01 g4675 ( .a(n11405), .b(n7446_1), .c(n11404), .o(n8294) );
in01f01 g4676 ( .a(_net_6020), .o(n11407) );
na02f01 g4677 ( .a(n7348), .b(_net_7820), .o(n11408) );
oa12f01 g4678 ( .a(n11408), .b(n7348), .c(n11407), .o(n8299) );
in01f01 g4679 ( .a(_net_6200), .o(n11410) );
no02f01 g4680 ( .a(_net_392), .b(n11410), .o(n8324) );
no02f01 g4681 ( .a(n8673), .b(n7468_1), .o(n11412) );
no02f01 g4682 ( .a(n8682), .b(n7470), .o(n11413) );
ao22f01 g4683 ( .a(n7130), .b(net_6713), .c(n7127), .d(net_6777), .o(n11414) );
ao22f01 g4684 ( .a(n7135), .b(net_6745), .c(n7133_1), .d(net_6809), .o(n11415) );
ao12f01 g4685 ( .a(n7123), .b(n11415), .c(n11414), .o(n11416) );
in01f01 g4686 ( .a(_net_6123), .o(n11417) );
no02f01 g4687 ( .a(n7118), .b(n11417), .o(n11418) );
no04f01 g4688 ( .a(n11418), .b(n11416), .c(n11413), .d(n11412), .o(n11419) );
in01f01 g4689 ( .a(net_6725), .o(n11420) );
in01f01 g4690 ( .a(net_6757), .o(n11421) );
oa22f01 g4691 ( .a(n7492_1), .b(n11420), .c(n7491), .d(n11421), .o(n11422) );
in01f01 g4692 ( .a(net_6821), .o(n11423) );
in01f01 g4693 ( .a(net_6789), .o(n11424) );
oa22f01 g4694 ( .a(n7497), .b(n11423), .c(n7496_1), .d(n11424), .o(n11425) );
no02f01 g4695 ( .a(n11425), .b(n11422), .o(n11426) );
na02f01 g4696 ( .a(n11426), .b(n11419), .o(n8345) );
na02f01 g4697 ( .a(n10291), .b(n7125_1), .o(n11428) );
ao22f01 g4698 ( .a(n10289), .b(n9611_1), .c(n8716), .d(_net_6823), .o(n11429) );
na02f01 g4699 ( .a(n11429), .b(n11428), .o(n8354) );
in01f01 g4700 ( .a(n9444), .o(n11431) );
no02f01 g4701 ( .a(n11431), .b(n9439), .o(n8367) );
oa12f01 g4702 ( .a(n7397), .b(n6959), .c(n8231), .o(n11433) );
na03f01 g4703 ( .a(n11433), .b(n10048), .c(n10047_1), .o(n11434) );
na02f01 g4704 ( .a(n7399), .b(n6961), .o(n11435) );
ao22f01 g4705 ( .a(n11435), .b(n10043), .c(n8237_1), .d(_net_7685), .o(n11436) );
na02f01 g4706 ( .a(n11436), .b(n11434), .o(n8372) );
in01f01 g4707 ( .a(_net_7735), .o(n11438) );
ao12f01 g4708 ( .a(n7343), .b(n11438), .c(n7315), .o(n8377) );
in01f01 g4709 ( .a(_net_7602), .o(n11440) );
na02f01 g4710 ( .a(n7892), .b(n6968), .o(n11441) );
oa12f01 g4711 ( .a(n11441), .b(n6968), .c(n11440), .o(n8382) );
ao12f01 g4712 ( .a(n7682), .b(_net_6960), .c(_net_6963), .o(n11443) );
oa12f01 g4713 ( .a(n11443), .b(_net_6960), .c(_net_6963), .o(n11444) );
na02f01 g4714 ( .a(n9778), .b(n11219), .o(n11445) );
oa12f01 g4715 ( .a(n9526), .b(n11445), .c(n11444), .o(n8387) );
in01f01 g4716 ( .a(_net_7568), .o(n11447) );
na02f01 g4717 ( .a(n7519), .b(n7403), .o(n11448) );
oa12f01 g4718 ( .a(n11448), .b(n7519), .c(n11447), .o(n8396) );
na02f01 g4719 ( .a(n8340_1), .b(n6806_1), .o(n11450) );
ao22f01 g4720 ( .a(n8538), .b(n8338), .c(n8345_1), .d(_net_6958), .o(n11451) );
na02f01 g4721 ( .a(n11451), .b(n11450), .o(n8405) );
in01f01 g4722 ( .a(_net_7333), .o(n11453) );
na02f01 g4723 ( .a(n9685), .b(n7150), .o(n11454) );
oa12f01 g4724 ( .a(n11454), .b(n7150), .c(n11453), .o(n8410) );
na02f01 g4725 ( .a(n11121), .b(n6917), .o(n11456) );
ao22f01 g4726 ( .a(n8005_1), .b(n6935), .c(n6933), .d(_net_6089), .o(n11457) );
no03f01 g4727 ( .a(n10592), .b(n6947_1), .c(n6943_1), .o(n11458) );
ao12f01 g4728 ( .a(n11458), .b(n8009), .c(n6946), .o(n11459) );
na03f01 g4729 ( .a(n11459), .b(n11457), .c(n11456), .o(n8426) );
na02f01 g4730 ( .a(n7298), .b(net_7741), .o(n11461) );
ao22f01 g4731 ( .a(n7306), .b(_net_6011), .c(n7291), .d(net_7712), .o(n11462) );
na02f01 g4732 ( .a(n7302_1), .b(net_151), .o(n11463) );
na02f01 g4733 ( .a(n7296), .b(net_251), .o(n11464) );
na03f01 g4734 ( .a(n7308), .b(_net_177), .c(n6800), .o(n11465) );
na03f01 g4735 ( .a(n7308), .b(_net_214), .c(x1322), .o(n11466) );
na03f01 g4736 ( .a(n11466), .b(n11465), .c(n11464), .o(n11467) );
ao12f01 g4737 ( .a(n11467), .b(n7286), .c(_net_294), .o(n11468) );
na04f01 g4738 ( .a(n11468), .b(n11463), .c(n11462), .d(n11461), .o(n8435) );
no03f01 g4739 ( .a(n7114), .b(_net_7688), .c(x1155), .o(n8443) );
in01f01 g4740 ( .a(_net_7450), .o(n11471) );
na02f01 g4741 ( .a(n9487_1), .b(n7197), .o(n11472) );
oa12f01 g4742 ( .a(n11472), .b(n7197), .c(n11471), .o(n8481) );
in01f01 g4743 ( .a(net_7173), .o(n11474) );
in01f01 g4744 ( .a(net_7109), .o(n11475) );
oa22f01 g4745 ( .a(n7580), .b(n11475), .c(n7577_1), .d(n11474), .o(n11476) );
in01f01 g4746 ( .a(net_7141), .o(n11477) );
in01f01 g4747 ( .a(net_7205), .o(n11478) );
oa22f01 g4748 ( .a(n7585), .b(n11477), .c(n7583), .d(n11478), .o(n11479) );
no02f01 g4749 ( .a(n11479), .b(n11476), .o(n11480) );
no02f01 g4750 ( .a(n11480), .b(n7721), .o(n11481) );
no02f01 g4751 ( .a(n7935), .b(n7592), .o(n11482) );
in01f01 g4752 ( .a(_net_6178), .o(n11483) );
oa22f01 g4753 ( .a(n7718), .b(n7574), .c(n7590), .d(n11483), .o(n11484) );
no03f01 g4754 ( .a(n11484), .b(n11482), .c(n11481), .o(n11485) );
in01f01 g4755 ( .a(net_7157), .o(n11486) );
in01f01 g4756 ( .a(net_7125), .o(n11487) );
oa22f01 g4757 ( .a(n7740), .b(n11487), .c(n7739), .d(n11486), .o(n11488) );
in01f01 g4758 ( .a(net_7189), .o(n11489) );
in01f01 g4759 ( .a(net_7221), .o(n11490) );
oa22f01 g4760 ( .a(n7745), .b(n11490), .c(n7744), .d(n11489), .o(n11491) );
no02f01 g4761 ( .a(n11491), .b(n11488), .o(n11492) );
na02f01 g4762 ( .a(n11492), .b(n11485), .o(n8486) );
in01f01 g4763 ( .a(_net_7801), .o(n11494) );
na02f01 g4764 ( .a(n6803), .b(_net_6039), .o(n11495) );
oa12f01 g4765 ( .a(n11495), .b(n6803), .c(n11494), .o(n8499) );
no02f01 g4766 ( .a(_net_6557), .b(n7762), .o(n11497) );
no02f01 g4767 ( .a(n7765), .b(net_6556), .o(n11498) );
no02f01 g4768 ( .a(n11498), .b(n11497), .o(n11499) );
oa22f01 g4769 ( .a(n11499), .b(n10412), .c(n10416), .d(n7765), .o(n8508) );
in01f01 g4770 ( .a(_net_7575), .o(n11501) );
na02f01 g4771 ( .a(n7519), .b(n793), .o(n11502) );
oa12f01 g4772 ( .a(n11502), .b(n7519), .c(n11501), .o(n8517) );
in01f01 g4773 ( .a(_net_7349), .o(n11504) );
na02f01 g4774 ( .a(n7183), .b(n7030), .o(n11505) );
oa12f01 g4775 ( .a(n11505), .b(n7030), .c(n11504), .o(n8526) );
in01f01 g4776 ( .a(_net_7284), .o(n11507) );
na02f01 g4777 ( .a(n7180), .b(n6904), .o(n11508) );
oa12f01 g4778 ( .a(n11508), .b(n7180), .c(n11507), .o(n8531) );
ao22f01 g4779 ( .a(n6736_1), .b(_net_7625), .c(n6734), .d(_net_7593), .o(n11510) );
ao22f01 g4780 ( .a(n6739), .b(_net_7657), .c(n6738), .d(_net_7561), .o(n11511) );
na02f01 g4781 ( .a(n11511), .b(n11510), .o(n8540) );
ao22f01 g4782 ( .a(n6877), .b(_net_7260), .c(n6876_1), .d(_net_7324), .o(n11513) );
ao22f01 g4783 ( .a(n6881_1), .b(_net_7292), .c(n6880), .d(_net_7356), .o(n11514) );
na02f01 g4784 ( .a(n11514), .b(n11513), .o(n8557) );
in01f01 g4785 ( .a(_net_122), .o(n11516) );
na02f01 g4786 ( .a(net_318), .b(_net_154), .o(n11517) );
oa12f01 g4787 ( .a(n11517), .b(n11516), .c(_net_154), .o(n8570) );
in01f01 g4788 ( .a(_net_6281), .o(n11519) );
no02f01 g4789 ( .a(_net_392), .b(n11519), .o(n8583) );
in01f01 g4790 ( .a(n11290), .o(n11521) );
no02f01 g4791 ( .a(n11521), .b(x889), .o(n8588) );
in01f01 g4792 ( .a(_net_7695), .o(n11523) );
na02f01 g4793 ( .a(n7207_1), .b(_net_7797), .o(n11524) );
oa12f01 g4794 ( .a(n11524), .b(n7207_1), .c(n11523), .o(n8593) );
in01f01 g4795 ( .a(_net_7319), .o(n11526) );
na02f01 g4796 ( .a(n8022), .b(n7150), .o(n11527) );
oa12f01 g4797 ( .a(n11527), .b(n7150), .c(n11526), .o(n8602) );
ao22f01 g4798 ( .a(n6877), .b(_net_7275), .c(n6876_1), .d(net_7339), .o(n11529) );
ao22f01 g4799 ( .a(n6881_1), .b(net_7307), .c(n6880), .d(net_7371), .o(n11530) );
na02f01 g4800 ( .a(n11530), .b(n11529), .o(n8607) );
in01f01 g4801 ( .a(_net_6164), .o(n11532) );
no02f01 g4802 ( .a(n11532), .b(n7168), .o(n8616) );
no02f01 g4803 ( .a(n8087), .b(_net_6410), .o(n11534) );
ao12f01 g4804 ( .a(n8084), .b(n11534), .c(n8179_1), .o(n8625) );
no02f01 g4805 ( .a(n8397), .b(n6824), .o(n11536) );
no02f01 g4806 ( .a(n8406), .b(n6826_1), .o(n11537) );
in01f01 g4807 ( .a(_net_6141), .o(n11538) );
no02f01 g4808 ( .a(n10716), .b(n10713), .o(n11539) );
oa22f01 g4809 ( .a(n11539), .b(n6836_1), .c(n6844), .d(n11538), .o(n11540) );
no03f01 g4810 ( .a(n11540), .b(n11537), .c(n11536), .o(n11541) );
in01f01 g4811 ( .a(net_6890), .o(n11542) );
in01f01 g4812 ( .a(net_6858), .o(n11543) );
oa22f01 g4813 ( .a(n6850_1), .b(n11543), .c(n6849), .d(n11542), .o(n11544) );
in01f01 g4814 ( .a(net_6922), .o(n11545) );
in01f01 g4815 ( .a(net_6954), .o(n11546) );
oa22f01 g4816 ( .a(n6855_1), .b(n11546), .c(n6854), .d(n11545), .o(n11547) );
no02f01 g4817 ( .a(n11547), .b(n11544), .o(n11548) );
na02f01 g4818 ( .a(n11548), .b(n11541), .o(n8645) );
ao22f01 g4819 ( .a(n7225), .b(_net_7406), .c(n7224), .d(_net_7438), .o(n11550) );
ao22f01 g4820 ( .a(n7229), .b(_net_7502), .c(n7228), .d(_net_7470), .o(n11551) );
na02f01 g4821 ( .a(n11551), .b(n11550), .o(n8662) );
in01f01 g4822 ( .a(_net_7267), .o(n11553) );
na02f01 g4823 ( .a(n7567_1), .b(n6901), .o(n11554) );
oa12f01 g4824 ( .a(n11554), .b(n6901), .c(n11553), .o(n8671) );
na02f01 g4825 ( .a(n9410_1), .b(n9405_1), .o(n11556) );
oa12f01 g4826 ( .a(n11556), .b(n9409), .c(n9405_1), .o(n8676) );
in01f01 g4827 ( .a(_net_7627), .o(n11558) );
na02f01 g4828 ( .a(n7400_1), .b(n6971), .o(n11559) );
oa12f01 g4829 ( .a(n11559), .b(n7400_1), .c(n11558), .o(n8689) );
na02f01 g4830 ( .a(n6996), .b(_net_6144), .o(n11561) );
na02f01 g4831 ( .a(n9719_1), .b(n6981), .o(n11562) );
na02f01 g4832 ( .a(n11562), .b(n11561), .o(n8694) );
na02f01 g4833 ( .a(n7348), .b(_net_7813), .o(n11564) );
oa12f01 g4834 ( .a(n11564), .b(n7348), .c(n7259), .o(n8703) );
ao22f01 g4835 ( .a(n7298), .b(_net_7731), .c(n7288_1), .d(_net_6042), .o(n11566) );
ao22f01 g4836 ( .a(n7306), .b(_net_5998), .c(n7286), .d(_net_281), .o(n11567) );
na02f01 g4837 ( .a(n7302_1), .b(_net_125), .o(n11568) );
na03f01 g4838 ( .a(n7308), .b(net_167), .c(n6800), .o(n11569) );
na03f01 g4839 ( .a(n7308), .b(net_204), .c(x1322), .o(n11570) );
na02f01 g4840 ( .a(n7296), .b(net_241), .o(n11571) );
na03f01 g4841 ( .a(n11571), .b(n11570), .c(n11569), .o(n11572) );
ao12f01 g4842 ( .a(n11572), .b(n7291), .c(_net_7702), .o(n11573) );
na04f01 g4843 ( .a(n11573), .b(n11568), .c(n11567), .d(n11566), .o(n8708) );
in01f01 g4844 ( .a(_net_7477), .o(n11575) );
na02f01 g4845 ( .a(n8633), .b(n6869), .o(n11576) );
oa12f01 g4846 ( .a(n11576), .b(n6869), .c(n11575), .o(n8720) );
na02f01 g4847 ( .a(n10289), .b(n9617), .o(n11578) );
na02f01 g4848 ( .a(n7134), .b(n7126), .o(n11579) );
ao22f01 g4849 ( .a(n11579), .b(n10291), .c(n8716), .d(_net_6824), .o(n11580) );
na02f01 g4850 ( .a(n11580), .b(n11578), .o(n8725) );
na02f01 g4851 ( .a(n10737), .b(n10736), .o(n11582) );
na02f01 g4852 ( .a(n11582), .b(n7124), .o(n11583) );
ao22f01 g4853 ( .a(n8183_1), .b(n8159), .c(n7119), .d(_net_6109), .o(n11584) );
na02f01 g4854 ( .a(n8187), .b(n8164), .o(n11585) );
oa12f01 g4855 ( .a(n8167), .b(n8681_1), .c(n8678), .o(n11586) );
na04f01 g4856 ( .a(n11586), .b(n11585), .c(n11584), .d(n11583), .o(n8730) );
in01f01 g4857 ( .a(_net_7805), .o(n11588) );
na02f01 g4858 ( .a(n6803), .b(_net_6043), .o(n11589) );
oa12f01 g4859 ( .a(n11589), .b(n6803), .c(n11588), .o(n8743) );
in01f01 g4860 ( .a(_net_7476), .o(n11591) );
na02f01 g4861 ( .a(n7553_1), .b(n6869), .o(n11592) );
oa12f01 g4862 ( .a(n11592), .b(n6869), .c(n11591), .o(n8748) );
in01f01 g4863 ( .a(_net_7585), .o(n11594) );
na02f01 g4864 ( .a(n8246), .b(n6968), .o(n11595) );
oa12f01 g4865 ( .a(n11595), .b(n6968), .c(n11594), .o(n8753) );
in01f01 g4866 ( .a(_net_6288), .o(n11597) );
no02f01 g4867 ( .a(_net_392), .b(n11597), .o(n8762) );
ao12f01 g4868 ( .a(n9671), .b(n10332), .c(n10423), .o(n11599) );
no02f01 g4869 ( .a(n11599), .b(_net_6411), .o(n11600) );
no02f01 g4870 ( .a(n11600), .b(n8177), .o(n8771) );
na02f01 g4871 ( .a(n9105), .b(n8307_1), .o(n11602) );
no02f01 g4872 ( .a(n7583), .b(n9102), .o(n11603) );
no02f01 g4873 ( .a(n7584), .b(_net_7230), .o(n11604) );
no02f01 g4874 ( .a(n11604), .b(n11603), .o(n11605) );
ao22f01 g4875 ( .a(n11605), .b(n8310), .c(n8312), .d(_net_7230), .o(n11606) );
na02f01 g4876 ( .a(n11606), .b(n11602), .o(n8775) );
in01f01 g4877 ( .a(_net_7265), .o(n11608) );
na02f01 g4878 ( .a(n9537_1), .b(n6901), .o(n11609) );
oa12f01 g4879 ( .a(n11609), .b(n6901), .c(n11608), .o(n8780) );
na04f01 g4880 ( .a(n10016), .b(_net_6414), .c(net_6412), .d(n10012), .o(n8809) );
in01f01 g4881 ( .a(_net_7409), .o(n11612) );
na02f01 g4882 ( .a(n7550), .b(n7200), .o(n11613) );
oa12f01 g4883 ( .a(n11613), .b(n7550), .c(n11612), .o(n8818) );
ao22f01 g4884 ( .a(n7225), .b(_net_7403), .c(n7224), .d(_net_7435), .o(n11615) );
ao22f01 g4885 ( .a(n7229), .b(_net_7499), .c(n7228), .d(_net_7467), .o(n11616) );
na02f01 g4886 ( .a(n11616), .b(n11615), .o(n8831) );
in01f01 g4887 ( .a(_net_7664), .o(n11618) );
na02f01 g4888 ( .a(n7446_1), .b(n7403), .o(n11619) );
oa12f01 g4889 ( .a(n11619), .b(n7446_1), .c(n11618), .o(n8840) );
in01f01 g4890 ( .a(_net_6048), .o(n11621) );
oa12f01 g4891 ( .a(n11621), .b(n7572_1), .c(n8695), .o(n8845) );
in01f01 g4892 ( .a(_net_7363), .o(n11623) );
na02f01 g4893 ( .a(n7567_1), .b(n7030), .o(n11624) );
oa12f01 g4894 ( .a(n11624), .b(n7030), .c(n11623), .o(n8855) );
in01f01 g4895 ( .a(_net_7625), .o(n11626) );
na02f01 g4896 ( .a(n10071), .b(n7400_1), .o(n11627) );
oa12f01 g4897 ( .a(n11627), .b(n7400_1), .c(n11626), .o(n8860) );
in01f01 g4898 ( .a(_net_6185), .o(n11629) );
no02f01 g4899 ( .a(_net_392), .b(n11629), .o(n8869) );
in01f01 g4900 ( .a(_net_6297), .o(n11631) );
no02f01 g4901 ( .a(_net_392), .b(n11631), .o(n8895) );
na02f01 g4902 ( .a(n7912), .b(n7575), .o(n11633) );
ao22f01 g4903 ( .a(n7917), .b(n7593), .c(n7591_1), .d(_net_6166), .o(n11634) );
na02f01 g4904 ( .a(n11634), .b(n11633), .o(n8917) );
no03f01 g4905 ( .a(n7360), .b(n10532), .c(n7359_1), .o(n11636) );
no02f01 g4906 ( .a(n7361), .b(_net_7787), .o(n11637) );
no03f01 g4907 ( .a(n11637), .b(n11636), .c(n7358), .o(n8922) );
in01f01 g4908 ( .a(_net_7322), .o(n11639) );
na02f01 g4909 ( .a(n7393), .b(n7150), .o(n11640) );
oa12f01 g4910 ( .a(n11640), .b(n7150), .c(n11639), .o(n8948) );
in01f01 g4911 ( .a(_net_7451), .o(n11642) );
na02f01 g4912 ( .a(n8193), .b(n7197), .o(n11643) );
oa12f01 g4913 ( .a(n11643), .b(n7197), .c(n11642), .o(n8953) );
ao22f01 g4914 ( .a(n7225), .b(_net_7417), .c(n7224), .d(_net_7449), .o(n11645) );
ao22f01 g4915 ( .a(n7229), .b(_net_7513), .c(n7228), .d(_net_7481), .o(n11646) );
na02f01 g4916 ( .a(n11646), .b(n11645), .o(n8967) );
in01f01 g4917 ( .a(_net_7466), .o(n11648) );
na02f01 g4918 ( .a(n7883_1), .b(n6869), .o(n11649) );
oa12f01 g4919 ( .a(n11649), .b(n6869), .c(n11648), .o(n8976) );
in01f01 g4920 ( .a(_net_7581), .o(n11651) );
na02f01 g4921 ( .a(n7519), .b(n698), .o(n11652) );
oa12f01 g4922 ( .a(n11652), .b(n7519), .c(n11651), .o(n8986) );
na02f01 g4923 ( .a(n7440), .b(_net_7813), .o(n11654) );
oa12f01 g4924 ( .a(n11654), .b(n7440), .c(n10191), .o(n8995) );
na02f01 g4925 ( .a(n7440), .b(_net_7794), .o(n11656) );
oa12f01 g4926 ( .a(n11656), .b(n7440), .c(n9966_1), .o(n9000) );
na02f01 g4927 ( .a(n9915), .b(n9306), .o(n11658) );
na02f01 g4928 ( .a(n9914_1), .b(_net_7783), .o(n11659) );
na02f01 g4929 ( .a(n11659), .b(n11658), .o(n11660) );
oa22f01 g4930 ( .a(n11660), .b(n9913), .c(n9313), .d(n9306), .o(n9005) );
na02f01 g4931 ( .a(n7306), .b(_net_6018), .o(n11662) );
na02f01 g4932 ( .a(n7293), .b(net_218), .o(n11663) );
ao22f01 g4933 ( .a(n7297_1), .b(net_181), .c(n7296), .d(net_255), .o(n11664) );
ao22f01 g4934 ( .a(n7298), .b(_net_7745), .c(n7291), .d(_net_7716), .o(n11665) );
na04f01 g4935 ( .a(n11665), .b(n11664), .c(n11663), .d(n11662), .o(n9030) );
ao22f01 g4936 ( .a(n6738), .b(_net_7552), .c(n6736_1), .d(_net_7616), .o(n11667) );
ao22f01 g4937 ( .a(n6739), .b(_net_7648), .c(n6734), .d(_net_7584), .o(n11668) );
na02f01 g4938 ( .a(n11668), .b(n11667), .o(n9042) );
in01f01 g4939 ( .a(_net_7423), .o(n11670) );
na02f01 g4940 ( .a(n7550), .b(n634), .o(n11671) );
oa12f01 g4941 ( .a(n11671), .b(n7550), .c(n11670), .o(n9052) );
in01f01 g4942 ( .a(_net_115), .o(n11673) );
na02f01 g4943 ( .a(net_311), .b(_net_154), .o(n11674) );
oa12f01 g4944 ( .a(n11674), .b(n11673), .c(_net_154), .o(n9074) );
ao22f01 g4945 ( .a(n6736_1), .b(net_7642), .c(n6734), .d(net_7610), .o(n11676) );
ao22f01 g4946 ( .a(n6739), .b(net_7674), .c(n6738), .d(_net_7578), .o(n11677) );
na02f01 g4947 ( .a(n11677), .b(n11676), .o(n9096) );
na02f01 g4948 ( .a(n7440), .b(_net_7809), .o(n11679) );
oa12f01 g4949 ( .a(n11679), .b(n7440), .c(n8236), .o(n9101) );
in01f01 g4950 ( .a(_net_7716), .o(n11681) );
na02f01 g4951 ( .a(n7207_1), .b(_net_7818), .o(n11682) );
oa12f01 g4952 ( .a(n11682), .b(n7207_1), .c(n11681), .o(n9106) );
na02f01 g4953 ( .a(n7440), .b(_net_7812), .o(n11684) );
oa12f01 g4954 ( .a(n11684), .b(n7440), .c(n7143), .o(n9115) );
in01f01 g4955 ( .a(_net_7558), .o(n11686) );
na02f01 g4956 ( .a(n7644_1), .b(n7519), .o(n11687) );
oa12f01 g4957 ( .a(n11687), .b(n7519), .c(n11686), .o(n9124) );
in01f01 g4958 ( .a(_net_7660), .o(n11689) );
na02f01 g4959 ( .a(n8043), .b(n7446_1), .o(n11690) );
oa12f01 g4960 ( .a(n11690), .b(n7446_1), .c(n11689), .o(n9129) );
ao22f01 g4961 ( .a(n6877), .b(_net_7256), .c(n6876_1), .d(_net_7320), .o(n11692) );
ao22f01 g4962 ( .a(n6881_1), .b(_net_7288), .c(n6880), .d(_net_7352), .o(n11693) );
na02f01 g4963 ( .a(n11693), .b(n11692), .o(n9151) );
in01f01 g4964 ( .a(_net_7259), .o(n11695) );
na02f01 g4965 ( .a(n7033), .b(n6901), .o(n11696) );
oa12f01 g4966 ( .a(n11696), .b(n6901), .c(n11695), .o(n9156) );
in01f01 g4967 ( .a(_net_6187), .o(n11698) );
no02f01 g4968 ( .a(_net_392), .b(n11698), .o(n9173) );
in01f01 g4969 ( .a(_net_7260), .o(n11700) );
na02f01 g4970 ( .a(n10089_1), .b(n6901), .o(n11701) );
oa12f01 g4971 ( .a(n11701), .b(n6901), .c(n11700), .o(n9187) );
ao22f01 g4972 ( .a(n6877), .b(_net_7266), .c(n6876_1), .d(_net_7330), .o(n11703) );
ao22f01 g4973 ( .a(n6881_1), .b(_net_7298), .c(n6880), .d(_net_7362), .o(n11704) );
na02f01 g4974 ( .a(n11704), .b(n11703), .o(n9192) );
no02f01 g4975 ( .a(n6739), .b(n8349), .o(n11706) );
no03f01 g4976 ( .a(_net_7682), .b(n6733), .c(n6735), .o(n11707) );
no02f01 g4977 ( .a(n11707), .b(n11706), .o(n11708) );
oa22f01 g4978 ( .a(n11708), .b(n10455), .c(n10456), .d(n8349), .o(n9201) );
in01f01 g4979 ( .a(_net_5986), .o(n11710) );
na02f01 g4980 ( .a(n7348), .b(_net_7795), .o(n11711) );
oa12f01 g4981 ( .a(n11711), .b(n7348), .c(n11710), .o(n9206) );
in01f01 g4982 ( .a(n9347), .o(n11713) );
no02f01 g4983 ( .a(n11713), .b(x940), .o(n9211) );
no02f01 g4984 ( .a(n9283), .b(n6945), .o(n11715) );
no02f01 g4985 ( .a(n9292), .b(n6934_1), .o(n11716) );
in01f01 g4986 ( .a(_net_6094), .o(n11717) );
oa22f01 g4987 ( .a(n10132_1), .b(n6916), .c(n6932), .d(n11717), .o(n11718) );
no03f01 g4988 ( .a(n11718), .b(n11716), .c(n11715), .o(n11719) );
in01f01 g4989 ( .a(net_6613), .o(n11720) );
in01f01 g4990 ( .a(net_6581), .o(n11721) );
oa22f01 g4991 ( .a(n7058_1), .b(n11721), .c(n7057), .d(n11720), .o(n11722) );
in01f01 g4992 ( .a(net_6677), .o(n11723) );
in01f01 g4993 ( .a(net_6645), .o(n11724) );
oa22f01 g4994 ( .a(n7063), .b(n11723), .c(n7062_1), .d(n11724), .o(n11725) );
no02f01 g4995 ( .a(n11725), .b(n11722), .o(n11726) );
na02f01 g4996 ( .a(n11726), .b(n11719), .o(n9220) );
in01f01 g4997 ( .a(_net_7701), .o(n11728) );
na02f01 g4998 ( .a(n7207_1), .b(_net_7803), .o(n11729) );
oa12f01 g4999 ( .a(n11729), .b(n7207_1), .c(n11728), .o(n9233) );
na02f01 g5000 ( .a(_net_6405), .b(n8088_1), .o(n11731) );
na03f01 g5001 ( .a(n11731), .b(n8090), .c(n6910_1), .o(n9258) );
in01f01 g5002 ( .a(_net_7515), .o(n11733) );
na02f01 g5003 ( .a(n8193), .b(n7626_1), .o(n11734) );
oa12f01 g5004 ( .a(n11734), .b(n7626_1), .c(n11733), .o(n9263) );
no02f01 g5005 ( .a(n7228), .b(n7224), .o(n11736) );
oa22f01 g5006 ( .a(n11736), .b(n8872), .c(n8873_1), .d(n7227), .o(n9272) );
na02f01 g5007 ( .a(n8162), .b(n7124), .o(n11738) );
ao22f01 g5008 ( .a(n8159), .b(n7137), .c(n7119), .d(_net_6106), .o(n11739) );
na02f01 g5009 ( .a(n11739), .b(n11738), .o(n9277) );
no02f01 g5010 ( .a(n6843), .b(n6824), .o(n11741) );
no02f01 g5011 ( .a(n7612), .b(n6826_1), .o(n11742) );
in01f01 g5012 ( .a(_net_6137), .o(n11743) );
oa22f01 g5013 ( .a(n8397), .b(n6836_1), .c(n6844), .d(n11743), .o(n11744) );
no03f01 g5014 ( .a(n11744), .b(n11742), .c(n11741), .o(n11745) );
in01f01 g5015 ( .a(net_6886), .o(n11746) );
in01f01 g5016 ( .a(net_6854), .o(n11747) );
oa22f01 g5017 ( .a(n6850_1), .b(n11747), .c(n6849), .d(n11746), .o(n11748) );
in01f01 g5018 ( .a(net_6918), .o(n11749) );
in01f01 g5019 ( .a(net_6950), .o(n11750) );
oa22f01 g5020 ( .a(n6855_1), .b(n11750), .c(n6854), .d(n11749), .o(n11751) );
no02f01 g5021 ( .a(n11751), .b(n11748), .o(n11752) );
na02f01 g5022 ( .a(n11752), .b(n11745), .o(n9282) );
in01f01 g5023 ( .a(_net_7516), .o(n11754) );
na02f01 g5024 ( .a(n9872), .b(n7626_1), .o(n11755) );
oa12f01 g5025 ( .a(n11755), .b(n7626_1), .c(n11754), .o(n9307) );
in01f01 g5026 ( .a(_net_7726), .o(n11757) );
ao12f01 g5027 ( .a(n7343), .b(n11757), .c(n7190_1), .o(n9312) );
ao22f01 g5028 ( .a(n7225), .b(_net_7427), .c(n7224), .d(net_7459), .o(n11759) );
ao22f01 g5029 ( .a(n7229), .b(net_7523), .c(n7228), .d(net_7491), .o(n11760) );
na02f01 g5030 ( .a(n11760), .b(n11759), .o(n9321) );
no02f01 g5031 ( .a(n10938), .b(n9893), .o(n9330) );
in01f01 g5032 ( .a(net_6003), .o(n11763) );
in01f01 g5033 ( .a(_net_7725), .o(n11764) );
ao12f01 g5034 ( .a(n7343), .b(n11764), .c(n11763), .o(n9335) );
in01f01 g5035 ( .a(_net_7504), .o(n11766) );
na02f01 g5036 ( .a(n8141), .b(n7626_1), .o(n11767) );
oa12f01 g5037 ( .a(n11767), .b(n7626_1), .c(n11766), .o(n9352) );
in01f01 g5038 ( .a(_net_7569), .o(n11769) );
na02f01 g5039 ( .a(n9318), .b(n7519), .o(n11770) );
oa12f01 g5040 ( .a(n11770), .b(n7519), .c(n11769), .o(n9410) );
na02f01 g5041 ( .a(n6933), .b(_net_6085), .o(n11772) );
na02f01 g5042 ( .a(n8009), .b(n6917), .o(n11773) );
na02f01 g5043 ( .a(n11773), .b(n11772), .o(n9415) );
in01f01 g5044 ( .a(_net_7317), .o(n11775) );
na02f01 g5045 ( .a(n7183), .b(n7150), .o(n11776) );
oa12f01 g5046 ( .a(n11776), .b(n7150), .c(n11775), .o(n9420) );
in01f01 g5047 ( .a(_net_7745), .o(n11778) );
in01f01 g5048 ( .a(_net_288), .o(n11779) );
ao12f01 g5049 ( .a(n7343), .b(n11779), .c(n11778), .o(n9436) );
ao22f01 g5050 ( .a(n7288_1), .b(net_6035), .c(n7286), .d(net_274), .o(n11781) );
ao22f01 g5051 ( .a(n7298), .b(_net_7727), .c(n7291), .d(_net_7698), .o(n11782) );
na02f01 g5052 ( .a(n7302_1), .b(_net_121), .o(n11783) );
na03f01 g5053 ( .a(n7308), .b(net_200), .c(x1322), .o(n11784) );
na02f01 g5054 ( .a(n7296), .b(net_237), .o(n11785) );
na03f01 g5055 ( .a(n7308), .b(net_163), .c(n6800), .o(n11786) );
na03f01 g5056 ( .a(n11786), .b(n11785), .c(n11784), .o(n11787) );
ao12f01 g5057 ( .a(n11787), .b(n7306), .c(_net_5991), .o(n11788) );
na04f01 g5058 ( .a(n11788), .b(n11783), .c(n11782), .d(n11781), .o(n9441) );
in01f01 g5059 ( .a(_net_6319), .o(n11790) );
no02f01 g5060 ( .a(_net_392), .b(n11790), .o(n9449) );
ao12f01 g5061 ( .a(n7067_1), .b(_net_6693), .c(_net_6690), .o(n11792) );
oa12f01 g5062 ( .a(n11792), .b(_net_6693), .c(_net_6690), .o(n11793) );
na02f01 g5063 ( .a(n7665), .b(n548), .o(n11794) );
oa12f01 g5064 ( .a(n9971_1), .b(n11794), .c(n11793), .o(n9454) );
in01f01 g5065 ( .a(_net_7415), .o(n11796) );
na02f01 g5066 ( .a(n7550), .b(n7504), .o(n11797) );
oa12f01 g5067 ( .a(n11797), .b(n7550), .c(n11796), .o(n9487) );
in01f01 g5068 ( .a(_net_7282), .o(n11799) );
na02f01 g5069 ( .a(n8731), .b(n7180), .o(n11800) );
oa12f01 g5070 ( .a(n11800), .b(n7180), .c(n11799), .o(n9492) );
in01f01 g5071 ( .a(_net_7597), .o(n11802) );
na02f01 g5072 ( .a(n7428), .b(n6968), .o(n11803) );
oa12f01 g5073 ( .a(n11803), .b(n6968), .c(n11802), .o(n9497) );
in01f01 g5074 ( .a(_net_7617), .o(n11805) );
na02f01 g5075 ( .a(n8246), .b(n7400_1), .o(n11806) );
oa12f01 g5076 ( .a(n11806), .b(n7400_1), .c(n11805), .o(n9507) );
in01f01 g5077 ( .a(_net_7616), .o(n11808) );
na02f01 g5078 ( .a(n8842), .b(n7400_1), .o(n11809) );
oa12f01 g5079 ( .a(n11809), .b(n7400_1), .c(n11808), .o(n9512) );
ao22f01 g5080 ( .a(n7225), .b(_net_7425), .c(n7224), .d(net_7457), .o(n11811) );
ao22f01 g5081 ( .a(n7229), .b(net_7521), .c(n7228), .d(net_7489), .o(n11812) );
na02f01 g5082 ( .a(n11812), .b(n11811), .o(n9533) );
ao22f01 g5083 ( .a(net_7739), .b(net_7710), .c(net_7737), .d(net_7708), .o(n11814) );
ao22f01 g5084 ( .a(net_7740), .b(net_7711), .c(net_7742), .d(net_7713), .o(n11815) );
ao22f01 g5085 ( .a(_net_7705), .b(_net_7734), .c(_net_7736), .d(_net_7707), .o(n11816) );
ao22f01 g5086 ( .a(net_7709), .b(net_7738), .c(_net_7733), .d(_net_7704), .o(n11817) );
na04f01 g5087 ( .a(n11817), .b(n11816), .c(n11815), .d(n11814), .o(n11818) );
na02f01 g5088 ( .a(_net_7745), .b(_net_7716), .o(n11819) );
ao22f01 g5089 ( .a(_net_7717), .b(_net_7746), .c(_net_7719), .d(_net_7748), .o(n11820) );
ao22f01 g5090 ( .a(net_7715), .b(net_7744), .c(net_7714), .d(net_7743), .o(n11821) );
ao22f01 g5091 ( .a(net_7712), .b(net_7741), .c(_net_7718), .d(_net_7747), .o(n11822) );
na04f01 g5092 ( .a(n11822), .b(n11821), .c(n11820), .d(n11819), .o(n11823) );
no02f01 g5093 ( .a(n11823), .b(n11818), .o(n11824) );
ao22f01 g5094 ( .a(_net_7723), .b(_net_7694), .c(net_7691), .d(_net_7720), .o(n11825) );
ao22f01 g5095 ( .a(_net_7693), .b(_net_7722), .c(_net_7721), .d(_net_7692), .o(n11826) );
ao22f01 g5096 ( .a(_net_7695), .b(_net_7724), .c(_net_7727), .d(_net_7698), .o(n11827) );
na03f01 g5097 ( .a(n11827), .b(n11826), .c(n11825), .o(n11828) );
ao22f01 g5098 ( .a(_net_7702), .b(_net_7731), .c(_net_7700), .d(_net_7729), .o(n11829) );
ao22f01 g5099 ( .a(_net_7735), .b(_net_7706), .c(_net_7703), .d(_net_7732), .o(n11830) );
ao22f01 g5100 ( .a(_net_7726), .b(_net_7697), .c(_net_7699), .d(_net_7728), .o(n11831) );
ao22f01 g5101 ( .a(_net_7725), .b(_net_7696), .c(_net_7701), .d(_net_7730), .o(n11832) );
na04f01 g5102 ( .a(n11832), .b(n11831), .c(n11830), .d(n11829), .o(n11833) );
no02f01 g5103 ( .a(n11833), .b(n11828), .o(n11834) );
na02f01 g5104 ( .a(n11834), .b(n11824), .o(n9546) );
in01f01 g5105 ( .a(net_7756), .o(n11836) );
na04f01 g5106 ( .a(_net_6017), .b(_net_7791), .c(net_303), .d(n11836), .o(n11837) );
ao12f01 g5107 ( .a(n11837), .b(net_306), .c(_net_6018), .o(n9554) );
no04f01 g5108 ( .a(n10024), .b(n7292_1), .c(x1215), .d(x1322), .o(n9559) );
na02f01 g5109 ( .a(n7348), .b(_net_7821), .o(n11840) );
oa12f01 g5110 ( .a(n11840), .b(n7348), .c(n7692), .o(n9564) );
in01f01 g5111 ( .a(_net_7509), .o(n11842) );
na02f01 g5112 ( .a(n8633), .b(n7626_1), .o(n11843) );
oa12f01 g5113 ( .a(n11843), .b(n7626_1), .c(n11842), .o(n9569) );
no03f01 g5114 ( .a(n8236), .b(_net_293), .c(n9540), .o(n11845) );
no02f01 g5115 ( .a(n8236), .b(n7653), .o(n11846) );
ao22f01 g5116 ( .a(n11846), .b(n10197), .c(n11845), .d(n10201), .o(n11847) );
ao12f01 g5117 ( .a(n8236), .b(_net_266), .c(n7653), .o(n11848) );
no03f01 g5118 ( .a(n8236), .b(_net_293), .c(_net_294), .o(n11849) );
ao22f01 g5119 ( .a(n11849), .b(n10199), .c(n11848), .d(n10192), .o(n11850) );
na02f01 g5120 ( .a(n11850), .b(n11847), .o(n9574) );
in01f01 g5121 ( .a(_net_7506), .o(n11852) );
na02f01 g5122 ( .a(n7626_1), .b(n6891), .o(n11853) );
oa12f01 g5123 ( .a(n11853), .b(n7626_1), .c(n11852), .o(n9583) );
no03f01 g5124 ( .a(n9339_1), .b(n6976), .c(_net_6032), .o(n11855) );
no02f01 g5125 ( .a(n6976), .b(n7316_1), .o(n11856) );
ao22f01 g5126 ( .a(n11856), .b(n9345), .c(n11855), .d(n9343_1), .o(n11857) );
ao12f01 g5127 ( .a(n6976), .b(n7316_1), .c(_net_5978), .o(n11858) );
no03f01 g5128 ( .a(_net_6033), .b(n6976), .c(_net_6032), .o(n11859) );
ao22f01 g5129 ( .a(n11859), .b(n9341), .c(n11858), .d(n9335_1), .o(n11860) );
na02f01 g5130 ( .a(n11860), .b(n11857), .o(n9592) );
ao12f01 g5131 ( .a(n7012), .b(n10472), .c(n10471), .o(n11862) );
no02f01 g5132 ( .a(n8052), .b(n6997), .o(n11863) );
in01f01 g5133 ( .a(_net_6153), .o(n11864) );
oa22f01 g5134 ( .a(n8060), .b(n6980), .c(n6995_1), .d(n11864), .o(n11865) );
no03f01 g5135 ( .a(n11865), .b(n11863), .c(n11862), .o(n11866) );
in01f01 g5136 ( .a(net_6985), .o(n11867) );
in01f01 g5137 ( .a(net_7017), .o(n11868) );
oa22f01 g5138 ( .a(n8075_1), .b(n11867), .c(n8074), .d(n11868), .o(n11869) );
in01f01 g5139 ( .a(net_7081), .o(n11870) );
in01f01 g5140 ( .a(net_7049), .o(n11871) );
oa22f01 g5141 ( .a(n8080_1), .b(n11870), .c(n8079), .d(n11871), .o(n11872) );
no02f01 g5142 ( .a(n11872), .b(n11869), .o(n11873) );
na02f01 g5143 ( .a(n11873), .b(n11866), .o(n9597) );
in01f01 g5144 ( .a(_net_7324), .o(n11875) );
na02f01 g5145 ( .a(n10089_1), .b(n7150), .o(n11876) );
oa12f01 g5146 ( .a(n11876), .b(n7150), .c(n11875), .o(n9602) );
in01f01 g5147 ( .a(n8177), .o(n11878) );
no03f01 g5148 ( .a(n9819_1), .b(n8178), .c(n11878), .o(n9616) );
in01f01 g5149 ( .a(_net_7436), .o(n11880) );
na02f01 g5150 ( .a(n7952), .b(n7197), .o(n11881) );
oa12f01 g5151 ( .a(n11881), .b(n7197), .c(n11880), .o(n9633) );
in01f01 g5152 ( .a(_net_7414), .o(n11883) );
na02f01 g5153 ( .a(n8994), .b(n7550), .o(n11884) );
oa12f01 g5154 ( .a(n11884), .b(n7550), .c(n11883), .o(n9638) );
in01f01 g5155 ( .a(_net_7327), .o(n11886) );
na02f01 g5156 ( .a(n7994_1), .b(n7150), .o(n11887) );
oa12f01 g5157 ( .a(n11887), .b(n7150), .c(n11886), .o(n9655) );
in01f01 g5158 ( .a(_net_7656), .o(n11889) );
na02f01 g5159 ( .a(n9881), .b(n7446_1), .o(n11890) );
oa12f01 g5160 ( .a(n11890), .b(n7446_1), .c(n11889), .o(n9664) );
in01f01 g5161 ( .a(_net_7588), .o(n11892) );
na02f01 g5162 ( .a(n8426_1), .b(n6968), .o(n11893) );
oa12f01 g5163 ( .a(n11893), .b(n6968), .c(n11892), .o(n9673) );
no04f01 g5164 ( .a(n8925), .b(n8915), .c(n6867_1), .d(_net_7532), .o(n9678) );
in01f01 g5165 ( .a(_net_7560), .o(n11896) );
na02f01 g5166 ( .a(n9881), .b(n7519), .o(n11897) );
oa12f01 g5167 ( .a(n11897), .b(n7519), .c(n11896), .o(n9683) );
na02f01 g5168 ( .a(n8124), .b(_net_6693), .o(n11899) );
na03f01 g5169 ( .a(n8123), .b(n8121_1), .c(n9973), .o(n11900) );
na02f01 g5170 ( .a(n8936), .b(net_6691), .o(n11901) );
na03f01 g5171 ( .a(n8935), .b(n8934_1), .c(n7153), .o(n11902) );
ao22f01 g5172 ( .a(n11902), .b(n11901), .c(n6944), .d(_net_6687), .o(n11903) );
na02f01 g5173 ( .a(n10364), .b(n7663), .o(n11904) );
na03f01 g5174 ( .a(n10363), .b(n10362), .c(_net_6692), .o(n11905) );
na03f01 g5175 ( .a(n11905), .b(n11904), .c(n11903), .o(n11906) );
ao12f01 g5176 ( .a(n11906), .b(n11900), .c(n11899), .o(n9700) );
na02f01 g5177 ( .a(n10421), .b(_net_6406), .o(n11908) );
no04f01 g5178 ( .a(n11908), .b(n10424), .c(n11878), .d(n8090), .o(n9709) );
no02f01 g5179 ( .a(n8406), .b(n6824), .o(n11910) );
no02f01 g5180 ( .a(n11539), .b(n6826_1), .o(n11911) );
ao22f01 g5181 ( .a(n6811), .b(net_6848), .c(n6808), .d(net_6912), .o(n11912) );
ao22f01 g5182 ( .a(n6816), .b(net_6880), .c(n6814), .d(net_6944), .o(n11913) );
ao12f01 g5183 ( .a(n6836_1), .b(n11913), .c(n11912), .o(n11914) );
in01f01 g5184 ( .a(_net_6143), .o(n11915) );
no02f01 g5185 ( .a(n6844), .b(n11915), .o(n11916) );
no04f01 g5186 ( .a(n11916), .b(n11914), .c(n11911), .d(n11910), .o(n11917) );
in01f01 g5187 ( .a(net_6860), .o(n11918) );
in01f01 g5188 ( .a(net_6892), .o(n11919) );
oa22f01 g5189 ( .a(n6850_1), .b(n11918), .c(n6849), .d(n11919), .o(n11920) );
in01f01 g5190 ( .a(net_6924), .o(n11921) );
in01f01 g5191 ( .a(net_6956), .o(n11922) );
oa22f01 g5192 ( .a(n6855_1), .b(n11922), .c(n6854), .d(n11921), .o(n11923) );
no02f01 g5193 ( .a(n11923), .b(n11920), .o(n11924) );
na02f01 g5194 ( .a(n11924), .b(n11917), .o(n9714) );
no02f01 g5195 ( .a(n9757), .b(n7721), .o(n11926) );
no02f01 g5196 ( .a(n9766), .b(n7592), .o(n11927) );
in01f01 g5197 ( .a(_net_6174), .o(n11928) );
oa22f01 g5198 ( .a(n11480), .b(n7574), .c(n7590), .d(n11928), .o(n11929) );
no03f01 g5199 ( .a(n11929), .b(n11927), .c(n11926), .o(n11930) );
in01f01 g5200 ( .a(net_7153), .o(n11931) );
in01f01 g5201 ( .a(net_7121), .o(n11932) );
oa22f01 g5202 ( .a(n7740), .b(n11932), .c(n7739), .d(n11931), .o(n11933) );
in01f01 g5203 ( .a(net_7217), .o(n11934) );
in01f01 g5204 ( .a(net_7185), .o(n11935) );
oa22f01 g5205 ( .a(n7745), .b(n11934), .c(n7744), .d(n11935), .o(n11936) );
no02f01 g5206 ( .a(n11936), .b(n11933), .o(n11937) );
na02f01 g5207 ( .a(n11937), .b(n11930), .o(n9719) );
no02f01 g5208 ( .a(n7026), .b(net_7378), .o(n11939) );
in01f01 g5209 ( .a(n11939), .o(n11940) );
no02f01 g5210 ( .a(n11940), .b(n9437), .o(n11941) );
no02f01 g5211 ( .a(n11939), .b(n9438), .o(n11942) );
oa12f01 g5212 ( .a(n9197), .b(n11942), .c(n11941), .o(n11943) );
no02f01 g5213 ( .a(n11942), .b(n11941), .o(n11944) );
na02f01 g5214 ( .a(n11944), .b(n3464), .o(n11945) );
na02f01 g5215 ( .a(n11945), .b(n11943), .o(n9733) );
ao22f01 g5216 ( .a(n6877), .b(_net_7264), .c(n6876_1), .d(_net_7328), .o(n11947) );
ao22f01 g5217 ( .a(n6881_1), .b(_net_7296), .c(n6880), .d(_net_7360), .o(n11948) );
na02f01 g5218 ( .a(n11948), .b(n11947), .o(n9742) );
in01f01 g5219 ( .a(_net_7576), .o(n11950) );
na02f01 g5220 ( .a(n2404), .b(n7519), .o(n11951) );
oa12f01 g5221 ( .a(n11951), .b(n7519), .c(n11950), .o(n9763) );
in01f01 g5222 ( .a(_net_7283), .o(n11953) );
na02f01 g5223 ( .a(n7659), .b(n7180), .o(n11954) );
oa12f01 g5224 ( .a(n11954), .b(n7180), .c(n11953), .o(n9768) );
in01f01 g5225 ( .a(_net_6002), .o(n11956) );
na02f01 g5226 ( .a(n7348), .b(_net_7808), .o(n11957) );
oa12f01 g5227 ( .a(n11957), .b(n7348), .c(n11956), .o(n9773) );
in01f01 g5228 ( .a(_net_7566), .o(n11959) );
na02f01 g5229 ( .a(n9373_1), .b(n7519), .o(n11960) );
oa12f01 g5230 ( .a(n11960), .b(n7519), .c(n11959), .o(n9787) );
na02f01 g5231 ( .a(n7348), .b(_net_7798), .o(n11962) );
oa12f01 g5232 ( .a(n11962), .b(n7348), .c(n7535_1), .o(n9792) );
na02f01 g5233 ( .a(n7028), .b(_net_7384), .o(n11964) );
na02f01 g5234 ( .a(n7029), .b(n9441_1), .o(n11965) );
na03f01 g5235 ( .a(n11965), .b(n11964), .c(n9852), .o(n11966) );
na03f01 g5236 ( .a(_net_7383), .b(_net_7381), .c(_net_7382), .o(n11967) );
na02f01 g5237 ( .a(n11967), .b(n9441_1), .o(n11968) );
in01f01 g5238 ( .a(n11967), .o(n11969) );
na02f01 g5239 ( .a(n11969), .b(_net_7384), .o(n11970) );
na03f01 g5240 ( .a(n11970), .b(n11968), .c(n9858_1), .o(n11971) );
na02f01 g5241 ( .a(n9860), .b(_net_7384), .o(n11972) );
na03f01 g5242 ( .a(n11972), .b(n11971), .c(n11966), .o(n9801) );
in01f01 g5243 ( .a(_net_5859), .o(n11974) );
in01f01 g5244 ( .a(x1062), .o(n11975) );
na03f01 g5245 ( .a(n11385), .b(net_7772), .c(n11975), .o(n11976) );
oa12f01 g5246 ( .a(n11976), .b(n11974), .c(x1062), .o(n9814) );
na02f01 g5247 ( .a(n7852), .b(n7194_1), .o(n11978) );
no02f01 g5248 ( .a(_net_7533), .b(n7846), .o(n11979) );
no02f01 g5249 ( .a(n7194_1), .b(_net_7532), .o(n11980) );
oa12f01 g5250 ( .a(n7845_1), .b(n11980), .c(n11979), .o(n11981) );
na02f01 g5251 ( .a(n7854), .b(_net_7533), .o(n11982) );
na03f01 g5252 ( .a(n11982), .b(n11981), .c(n11978), .o(n9819) );
oa12f01 g5253 ( .a(n7027_1), .b(n9854), .c(n7026), .o(n11984) );
na03f01 g5254 ( .a(n11984), .b(n11967), .c(n9858_1), .o(n11985) );
na02f01 g5255 ( .a(n7179), .b(n7149), .o(n11986) );
ao22f01 g5256 ( .a(n11986), .b(n9852), .c(n9860), .d(_net_7383), .o(n11987) );
na02f01 g5257 ( .a(n11987), .b(n11985), .o(n9824) );
in01f01 g5258 ( .a(_net_7421), .o(n11989) );
na02f01 g5259 ( .a(n1277), .b(n7550), .o(n11990) );
oa12f01 g5260 ( .a(n11990), .b(n7550), .c(n11989), .o(n9849) );
na02f01 g5261 ( .a(n9260), .b(n10421), .o(n11992) );
oa12f01 g5262 ( .a(_net_6407), .b(n9259), .c(n9258_1), .o(n11993) );
na03f01 g5263 ( .a(n11993), .b(n11992), .c(n6910_1), .o(n9858) );
no02f01 g5264 ( .a(_net_7097), .b(n8385), .o(n11995) );
no02f01 g5265 ( .a(n8760), .b(net_7096), .o(n11996) );
no02f01 g5266 ( .a(n11996), .b(n11995), .o(n11997) );
oa22f01 g5267 ( .a(n11997), .b(n10574), .c(n10578), .d(n8760), .o(n9863) );
in01f01 g5268 ( .a(n9665), .o(n11999) );
na02f01 g5269 ( .a(n9664_1), .b(n9663), .o(n12000) );
na02f01 g5270 ( .a(n12000), .b(n11999), .o(n12001) );
oa22f01 g5271 ( .a(n12001), .b(n9411), .c(n9409), .d(n9663), .o(n9880) );
oa12f01 g5272 ( .a(n7124), .b(n10744), .c(n10741), .o(n12003) );
ao22f01 g5273 ( .a(n11582), .b(n8159), .c(n7119), .d(_net_6111), .o(n12004) );
na02f01 g5274 ( .a(n11415), .b(n11414), .o(n12005) );
ao22f01 g5275 ( .a(n12005), .b(n8167), .c(n8183_1), .d(n8164), .o(n12006) );
na03f01 g5276 ( .a(n12006), .b(n12004), .c(n12003), .o(n9889) );
in01f01 g5277 ( .a(_net_287), .o(n12008) );
na02f01 g5278 ( .a(_net_225), .b(_net_227), .o(n12009) );
na02f01 g5279 ( .a(n12009), .b(n12008), .o(n9894) );
na02f01 g5280 ( .a(n7298), .b(net_7740), .o(n12011) );
ao22f01 g5281 ( .a(n7306), .b(_net_6010), .c(n7291), .d(net_7711), .o(n12012) );
na02f01 g5282 ( .a(n7302_1), .b(net_150), .o(n12013) );
na02f01 g5283 ( .a(n7296), .b(net_250), .o(n12014) );
na03f01 g5284 ( .a(n7308), .b(_net_176), .c(n6800), .o(n12015) );
na03f01 g5285 ( .a(n7308), .b(_net_213), .c(x1322), .o(n12016) );
na03f01 g5286 ( .a(n12016), .b(n12015), .c(n12014), .o(n12017) );
ao12f01 g5287 ( .a(n12017), .b(n7286), .c(_net_293), .o(n12018) );
na04f01 g5288 ( .a(n12018), .b(n12013), .c(n12012), .d(n12011), .o(n9907) );
oa12f01 g5289 ( .a(n11779), .b(n7851), .c(n7410), .o(n9939) );
in01f01 g5290 ( .a(_net_7348), .o(n12021) );
na02f01 g5291 ( .a(n7030), .b(n6904), .o(n12022) );
oa12f01 g5292 ( .a(n12022), .b(n7030), .c(n12021), .o(n9949) );
in01f01 g5293 ( .a(_net_7402), .o(n12024) );
na02f01 g5294 ( .a(n7883_1), .b(n7550), .o(n12025) );
oa12f01 g5295 ( .a(n12025), .b(n7550), .c(n12024), .o(n9966) );
no02f01 g5296 ( .a(n10554), .b(n6764), .o(n12027) );
no02f01 g5297 ( .a(n9225_1), .b(n6766), .o(n12028) );
in01f01 g5298 ( .a(_net_6076), .o(n12029) );
oa22f01 g5299 ( .a(n9233_1), .b(n6775), .c(n6784), .d(n12029), .o(n12030) );
no03f01 g5300 ( .a(n12030), .b(n12028), .c(n12027), .o(n12031) );
in01f01 g5301 ( .a(net_6448), .o(n12032) );
in01f01 g5302 ( .a(net_6480), .o(n12033) );
oa22f01 g5303 ( .a(n6790), .b(n12032), .c(n6789), .d(n12033), .o(n12034) );
in01f01 g5304 ( .a(net_6512), .o(n12035) );
in01f01 g5305 ( .a(net_6544), .o(n12036) );
oa22f01 g5306 ( .a(n6795), .b(n12036), .c(n6794), .d(n12035), .o(n12037) );
no02f01 g5307 ( .a(n12037), .b(n12034), .o(n12038) );
na02f01 g5308 ( .a(n12038), .b(n12031), .o(n9971) );
no02f01 g5309 ( .a(n11636), .b(_net_7788), .o(n12040) );
no03f01 g5310 ( .a(n12040), .b(n10533), .c(n7358), .o(n9981) );
in01f01 g5311 ( .a(_net_7717), .o(n12042) );
na02f01 g5312 ( .a(n7207_1), .b(_net_7819), .o(n12043) );
oa12f01 g5313 ( .a(n12043), .b(n7207_1), .c(n12042), .o(n9997) );
na02f01 g5314 ( .a(n7440), .b(_net_7793), .o(n12045) );
oa12f01 g5315 ( .a(n12045), .b(n7440), .c(n8094), .o(n10019) );
in01f01 g5316 ( .a(_net_7582), .o(n12047) );
na02f01 g5317 ( .a(n3604), .b(n7519), .o(n12048) );
oa12f01 g5318 ( .a(n12048), .b(n7519), .c(n12047), .o(n10032) );
na02f01 g5319 ( .a(n7348), .b(_net_7817), .o(n12050) );
oa12f01 g5320 ( .a(n12050), .b(n7348), .c(n6819), .o(n10037) );
in01f01 g5321 ( .a(_net_6202), .o(n12052) );
no02f01 g5322 ( .a(_net_392), .b(n12052), .o(n10042) );
in01f01 g5323 ( .a(_net_7287), .o(n12054) );
na02f01 g5324 ( .a(n8022), .b(n7180), .o(n12055) );
oa12f01 g5325 ( .a(n12055), .b(n7180), .c(n12054), .o(n10052) );
in01f01 g5326 ( .a(n10633), .o(n12057) );
no02f01 g5327 ( .a(n12057), .b(x1034), .o(n10061) );
ao22f01 g5328 ( .a(n7306), .b(_net_5995), .c(n7291), .d(_net_7699), .o(n12059) );
ao22f01 g5329 ( .a(n7288_1), .b(_net_6039), .c(n7286), .d(_net_278), .o(n12060) );
na02f01 g5330 ( .a(n7302_1), .b(_net_122), .o(n12061) );
na03f01 g5331 ( .a(n7308), .b(_net_201), .c(x1322), .o(n12062) );
na02f01 g5332 ( .a(n7296), .b(net_238), .o(n12063) );
na03f01 g5333 ( .a(n7308), .b(net_164), .c(n6800), .o(n12064) );
na03f01 g5334 ( .a(n12064), .b(n12063), .c(n12062), .o(n12065) );
ao12f01 g5335 ( .a(n12065), .b(n7298), .c(_net_7728), .o(n12066) );
na04f01 g5336 ( .a(n12066), .b(n12061), .c(n12060), .d(n12059), .o(n10066) );
in01f01 g5337 ( .a(_net_7251), .o(n12068) );
na02f01 g5338 ( .a(n7659), .b(n6901), .o(n12069) );
oa12f01 g5339 ( .a(n12069), .b(n6901), .c(n12068), .o(n10074) );
na02f01 g5340 ( .a(n8861), .b(n7754), .o(n12071) );
no02f01 g5341 ( .a(n6754), .b(n7749), .o(n12072) );
no02f01 g5342 ( .a(n6779_1), .b(_net_6555), .o(n12073) );
no02f01 g5343 ( .a(n12073), .b(n12072), .o(n12074) );
ao22f01 g5344 ( .a(n12074), .b(n8859), .c(n8862), .d(_net_6555), .o(n12075) );
na02f01 g5345 ( .a(n12075), .b(n12071), .o(n10079) );
oa12f01 g5346 ( .a(n8213), .b(n6832), .c(n6829), .o(n12077) );
ao22f01 g5347 ( .a(n8211_1), .b(_net_6131), .c(n9200), .d(n10704), .o(n12078) );
na02f01 g5348 ( .a(n11913), .b(n11912), .o(n12079) );
ao22f01 g5349 ( .a(n12079), .b(n9207), .c(n10708), .d(n9205), .o(n12080) );
na03f01 g5350 ( .a(n12080), .b(n12078), .c(n12077), .o(n10084) );
no02f01 g5351 ( .a(n10436), .b(n7721), .o(n12082) );
no02f01 g5352 ( .a(n10439), .b(n7592), .o(n12083) );
in01f01 g5353 ( .a(_net_6183), .o(n12084) );
no02f01 g5354 ( .a(n9074_1), .b(n9071), .o(n12085) );
oa22f01 g5355 ( .a(n12085), .b(n7574), .c(n7590), .d(n12084), .o(n12086) );
no03f01 g5356 ( .a(n12086), .b(n12083), .c(n12082), .o(n12087) );
in01f01 g5357 ( .a(net_7162), .o(n12088) );
in01f01 g5358 ( .a(net_7130), .o(n12089) );
oa22f01 g5359 ( .a(n7740), .b(n12089), .c(n7739), .d(n12088), .o(n12090) );
in01f01 g5360 ( .a(net_7194), .o(n12091) );
in01f01 g5361 ( .a(net_7226), .o(n12092) );
oa22f01 g5362 ( .a(n7745), .b(n12092), .c(n7744), .d(n12091), .o(n12093) );
no02f01 g5363 ( .a(n12093), .b(n12090), .o(n12094) );
na02f01 g5364 ( .a(n12094), .b(n12087), .o(n10089) );
in01f01 g5365 ( .a(_net_7264), .o(n12096) );
na02f01 g5366 ( .a(n7437_1), .b(n6901), .o(n12097) );
oa12f01 g5367 ( .a(n12097), .b(n6901), .c(n12096), .o(n10094) );
in01f01 g5368 ( .a(_net_7479), .o(n12099) );
na02f01 g5369 ( .a(n7504), .b(n6869), .o(n12100) );
oa12f01 g5370 ( .a(n12100), .b(n6869), .c(n12099), .o(n10099) );
ao22f01 g5371 ( .a(n6736_1), .b(_net_7634), .c(n6734), .d(_net_7602), .o(n12102) );
ao22f01 g5372 ( .a(n6739), .b(_net_7666), .c(n6738), .d(_net_7570), .o(n12103) );
na02f01 g5373 ( .a(n12103), .b(n12102), .o(n10116) );
in01f01 g5374 ( .a(_net_7356), .o(n12105) );
na02f01 g5375 ( .a(n10089_1), .b(n7030), .o(n12106) );
oa12f01 g5376 ( .a(n12106), .b(n7030), .c(n12105), .o(n10128) );
no02f01 g5377 ( .a(n9766), .b(n7721), .o(n12108) );
no02f01 g5378 ( .a(n11480), .b(n7592), .o(n12109) );
in01f01 g5379 ( .a(_net_6176), .o(n12110) );
oa22f01 g5380 ( .a(n7935), .b(n7574), .c(n7590), .d(n12110), .o(n12111) );
no03f01 g5381 ( .a(n12111), .b(n12109), .c(n12108), .o(n12112) );
in01f01 g5382 ( .a(net_7123), .o(n12113) );
in01f01 g5383 ( .a(net_7155), .o(n12114) );
oa22f01 g5384 ( .a(n7740), .b(n12113), .c(n7739), .d(n12114), .o(n12115) );
in01f01 g5385 ( .a(net_7219), .o(n12116) );
in01f01 g5386 ( .a(net_7187), .o(n12117) );
oa22f01 g5387 ( .a(n7745), .b(n12116), .c(n7744), .d(n12117), .o(n12118) );
no02f01 g5388 ( .a(n12118), .b(n12115), .o(n12119) );
na02f01 g5389 ( .a(n12119), .b(n12112), .o(n10137) );
na02f01 g5390 ( .a(n7917), .b(n7575), .o(n12121) );
oa12f01 g5391 ( .a(n12121), .b(n7590), .c(n11532), .o(n10150) );
bf01f01 g5392 ( .a(_net_5857), .o(x124) );
bf01f01 g5393 ( .a(_net_5852), .o(x84) );
bf01f01 g5394 ( .a(_net_5859), .o(x131) );
bf01f01 g5395 ( .a(x130657), .o(x145) );
bf01f01 g5396 ( .a(_net_5850), .o(x63) );
bf01f01 g5397 ( .a(_net_5853), .o(x96) );
bf01f01 g5398 ( .a(_net_5855), .o(x106) );
bf01f01 g5399 ( .a(_net_5854), .o(x101) );
bf01f01 g5400 ( .a(_net_5856), .o(x114) );
bf01f01 g5401 ( .a(_net_5851), .o(x77) );
bf01f01 g5402 ( .a(net_7807), .o(n276) );
bf01f01 g5403 ( .a(_net_6104), .o(n286) );
bf01f01 g5404 ( .a(net_6453), .o(n291) );
bf01f01 g5405 ( .a(_net_7820), .o(n305) );
bf01f01 g5406 ( .a(net_6704), .o(n310) );
bf01f01 g5407 ( .a(net_7802), .o(n324) );
bf01f01 g5408 ( .a(net_133), .o(n334) );
bf01f01 g5409 ( .a(_net_6168), .o(n339) );
bf01f01 g5410 ( .a(_net_6080), .o(n344) );
bf01f01 g5411 ( .a(net_6474), .o(n349) );
bf01f01 g5412 ( .a(x1542), .o(n352) );
bf01f01 g5413 ( .a(net_7114), .o(n357) );
bf01f01 g5414 ( .a(_net_7819), .o(n361) );
bf01f01 g5415 ( .a(net_6996), .o(n366) );
bf01f01 g5416 ( .a(_net_7820), .o(n395) );
bf01f01 g5417 ( .a(net_6395), .o(n405) );
bf01f01 g5418 ( .a(_net_6117), .o(n410) );
bf01f01 g5419 ( .a(_net_7795), .o(n415) );
bf01f01 g5420 ( .a(_net_7819), .o(n424) );
bf01f01 g5421 ( .a(_net_7806), .o(n429) );
bf01f01 g5422 ( .a(net_7713), .o(n434) );
bf01f01 g5423 ( .a(_net_7815), .o(n438) );
bf01f01 g5424 ( .a(net_7000), .o(n443) );
bf01f01 g5425 ( .a(x1527), .o(n451) );
bf01f01 g5426 ( .a(_net_7798), .o(n455) );
bf01f01 g5427 ( .a(net_7388), .o(n470) );
bf01f01 g5428 ( .a(net_6397), .o(n474) );
bf01f01 g5429 ( .a(_net_7818), .o(n479) );
bf01f01 g5430 ( .a(net_6870), .o(n484) );
bf01f01 g5431 ( .a(_net_7794), .o(n488) );
bf01f01 g5432 ( .a(_net_7822), .o(n493) );
bf01f01 g5433 ( .a(net_6059), .o(n498) );
bf01f01 g5434 ( .a(_net_6091), .o(n503) );
bf01f01 g5435 ( .a(_net_6112), .o(n508) );
bf01f01 g5436 ( .a(_net_7794), .o(n556) );
bf01f01 g5437 ( .a(_net_7808), .o(n566) );
bf01f01 g5438 ( .a(net_152), .o(n571) );
bf01f01 g5439 ( .a(x1587), .o(n580) );
bf01f01 g5440 ( .a(_net_6177), .o(n585) );
bf01f01 g5441 ( .a(net_6400), .o(n590) );
bf01f01 g5442 ( .a(_net_7800), .o(n610) );
bf01f01 g5443 ( .a(net_7246), .o(n625) );
bf01f01 g5444 ( .a(net_6383), .o(n664) );
bf01f01 g5445 ( .a(net_6440), .o(n669) );
bf01f01 g5446 ( .a(_net_7823), .o(n678) );
bf01f01 g5447 ( .a(_net_7796), .o(n683) );
bf01f01 g5448 ( .a(_net_6127), .o(n703) );
bf01f01 g5449 ( .a(net_6396), .o(n722) );
bf01f01 g5450 ( .a(net_147), .o(n741) );
bf01f01 g5451 ( .a(_net_5976), .o(n751) );
bf01f01 g5452 ( .a(net_6468), .o(n761) );
bf01f01 g5453 ( .a(x806), .o(n774) );
bf01f01 g5454 ( .a(net_6385), .o(n779) );
bf01f01 g5455 ( .a(net_7802), .o(n783) );
bf01f01 g5456 ( .a(net_7134), .o(n798) );
bf01f01 g5457 ( .a(net_7133), .o(n802) );
bf01f01 g5458 ( .a(net_6399), .o(n811) );
bf01f01 g5459 ( .a(_net_6084), .o(n815) );
bf01f01 g5460 ( .a(net_7396), .o(n830) );
bf01f01 g5461 ( .a(_net_7818), .o(n839) );
bf01f01 g5462 ( .a(net_6381), .o(n844) );
bf01f01 g5463 ( .a(net_7390), .o(n854) );
bf01f01 g5464 ( .a(_net_7794), .o(n857) );
bf01f01 g5465 ( .a(net_6711), .o(n867) );
bf01f01 g5466 ( .a(_net_7818), .o(n870) );
bf01f01 g5467 ( .a(_net_7816), .o(n880) );
bf01f01 g5468 ( .a(net_6616), .o(n890) );
bf01f01 g5469 ( .a(net_6382), .o(n894) );
bf01f01 g5470 ( .a(net_6739), .o(n899) );
bf01f01 g5471 ( .a(_net_7800), .o(n907) );
bf01f01 g5472 ( .a(_net_7806), .o(n911) );
bf01f01 g5473 ( .a(net_6746), .o(n916) );
bf01f01 g5474 ( .a(_net_6160), .o(n920) );
bf01f01 g5475 ( .a(net_7799), .o(n935) );
bf01f01 g5476 ( .a(net_6979), .o(n940) );
bf01f01 g5477 ( .a(x1467), .o(n948) );
bf01f01 g5478 ( .a(net_6989), .o(n953) );
bf01f01 g5479 ( .a(_net_7823), .o(n956) );
bf01f01 g5480 ( .a(_net_7813), .o(n976) );
bf01f01 g5481 ( .a(net_6999), .o(n981) );
bf01f01 g5482 ( .a(net_388), .o(n1000) );
bf01f01 g5483 ( .a(net_6391), .o(n1005) );
bf01f01 g5484 ( .a(net_6998), .o(n1020) );
bf01f01 g5485 ( .a(net_6386), .o(n1053) );
bf01f01 g5486 ( .a(_net_7812), .o(n1062) );
bf01f01 g5487 ( .a(net_7004), .o(n1077) );
bf01f01 g5488 ( .a(net_7010), .o(n1081) );
bf01f01 g5489 ( .a(net_6461), .o(n1085) );
bf01f01 g5490 ( .a(net_6832), .o(n1089) );
bf01f01 g5491 ( .a(net_6977), .o(n1093) );
bf01f01 g5492 ( .a(_net_7801), .o(n1097) );
bf01f01 g5493 ( .a(net_6856), .o(n1102) );
bf01f01 g5494 ( .a(_net_6183), .o(n1111) );
bf01f01 g5495 ( .a(net_6847), .o(n1121) );
bf01f01 g5496 ( .a(_net_7809), .o(n1130) );
bf01f01 g5497 ( .a(net_6986), .o(n1140) );
bf01f01 g5498 ( .a(_net_6099), .o(n1144) );
bf01f01 g5499 ( .a(_net_7815), .o(n1148) );
bf01f01 g5500 ( .a(_net_6066), .o(n1158) );
bf01f01 g5501 ( .a(net_6398), .o(n1168) );
bf01f01 g5502 ( .a(net_144), .o(n1183) );
bf01f01 g5503 ( .a(net_6400), .o(n1187) );
bf01f01 g5504 ( .a(_net_7823), .o(n1191) );
bf01f01 g5505 ( .a(_net_7822), .o(n1195) );
bf01f01 g5506 ( .a(_net_6064), .o(n1200) );
bf01f01 g5507 ( .a(_net_7814), .o(n1205) );
bf01f01 g5508 ( .a(net_6845), .o(n1210) );
bf01f01 g5509 ( .a(net_6608), .o(n1224) );
bf01f01 g5510 ( .a(_net_7795), .o(n1232) );
no02f01 g5511 ( .a(n6966), .b(n7599_1), .o(n1236) );
bf01f01 g5512 ( .a(_net_7820), .o(n1240) );
bf01f01 g5513 ( .a(net_6395), .o(n1244) );
bf01f01 g5514 ( .a(_net_7794), .o(n1248) );
bf01f01 g5515 ( .a(net_7019), .o(n1258) );
bf01f01 g5516 ( .a(_net_6158), .o(n1262) );
bf01f01 g5517 ( .a(net_7119), .o(n1287) );
bf01f01 g5518 ( .a(net_6574), .o(n1291) );
bf01f01 g5519 ( .a(_net_7803), .o(n1300) );
bf01f01 g5520 ( .a(net_7395), .o(n1305) );
bf01f01 g5521 ( .a(_net_7812), .o(n1318) );
bf01f01 g5522 ( .a(_net_7798), .o(n1322) );
bf01f01 g5523 ( .a(_net_7820), .o(n1326) );
bf01f01 g5524 ( .a(net_6859), .o(n1331) );
bf01f01 g5525 ( .a(net_6877), .o(n1355) );
bf01f01 g5526 ( .a(net_7234), .o(n1359) );
bf01f01 g5527 ( .a(_net_5960), .o(n1378) );
bf01f01 g5528 ( .a(net_6694), .o(n1383) );
bf01f01 g5529 ( .a(net_6400), .o(n1386) );
bf01f01 g5530 ( .a(_net_7794), .o(n1400) );
bf01f01 g5531 ( .a(_net_7815), .o(n1414) );
bf01f01 g5532 ( .a(_net_7809), .o(n1423) );
bf01f01 g5533 ( .a(net_6745), .o(n1438) );
bf01f01 g5534 ( .a(_net_7813), .o(n1446) );
bf01f01 g5535 ( .a(_net_7803), .o(n1455) );
bf01f01 g5536 ( .a(_net_6132), .o(n1460) );
bf01f01 g5537 ( .a(_net_7821), .o(n1465) );
bf01f01 g5538 ( .a(net_6392), .o(n1469) );
bf01f01 g5539 ( .a(net_6612), .o(n1474) );
bf01f01 g5540 ( .a(_net_6106), .o(n1478) );
bf01f01 g5541 ( .a(x1417), .o(n1482) );
bf01f01 g5542 ( .a(_net_7803), .o(n1491) );
bf01f01 g5543 ( .a(net_7550), .o(n1506) );
bf01f01 g5544 ( .a(_net_7824), .o(n1510) );
bf01f01 g5545 ( .a(net_6619), .o(n1515) );
bf01f01 g5546 ( .a(net_7106), .o(n1524) );
bf01f01 g5547 ( .a(_net_6179), .o(n1528) );
bf01f01 g5548 ( .a(net_7247), .o(n1538) );
bf01f01 g5549 ( .a(net_7146), .o(n1551) );
bf01f01 g5550 ( .a(net_7126), .o(n1560) );
bf01f01 g5551 ( .a(net_6482), .o(n1564) );
bf01f01 g5552 ( .a(net_6888), .o(n1568) );
bf01f01 g5553 ( .a(net_6388), .o(n1577) );
bf01f01 g5554 ( .a(net_6584), .o(n1587) );
bf01f01 g5555 ( .a(net_6387), .o(n1591) );
bf01f01 g5556 ( .a(net_6732), .o(n1596) );
bf01f01 g5557 ( .a(_net_7814), .o(n1615) );
bf01f01 g5558 ( .a(_net_7796), .o(n1619) );
bf01f01 g5559 ( .a(_net_7810), .o(n1629) );
bf01f01 g5560 ( .a(net_7124), .o(n1649) );
bf01f01 g5561 ( .a(net_135), .o(n1653) );
bf01f01 g5562 ( .a(net_6061), .o(n1663) );
bf01f01 g5563 ( .a(_net_5980), .o(n1668) );
bf01f01 g5564 ( .a(net_6723), .o(n1673) );
bf01f01 g5565 ( .a(_net_7824), .o(n1681) );
bf01f01 g5566 ( .a(_net_7817), .o(n1686) );
bf01f01 g5567 ( .a(_net_7805), .o(n1691) );
bf01f01 g5568 ( .a(net_6432), .o(n1701) );
bf01f01 g5569 ( .a(_net_7805), .o(n1704) );
bf01f01 g5570 ( .a(_net_7800), .o(n1709) );
bf01f01 g5571 ( .a(_net_7803), .o(n1718) );
bf01f01 g5572 ( .a(_net_7818), .o(n1722) );
bf01f01 g5573 ( .a(_net_7809), .o(n1732) );
bf01f01 g5574 ( .a(_net_7796), .o(n1756) );
bf01f01 g5575 ( .a(net_6570), .o(n1761) );
bf01f01 g5576 ( .a(_net_7821), .o(n1765) );
bf01f01 g5577 ( .a(net_6602), .o(n1775) );
bf01f01 g5578 ( .a(net_7551), .o(n1779) );
bf01f01 g5579 ( .a(_net_7800), .o(n1782) );
bf01f01 g5580 ( .a(_net_6120), .o(n1797) );
bf01f01 g5581 ( .a(_net_6175), .o(n1817) );
bf01f01 g5582 ( .a(_net_6093), .o(n1822) );
bf01f01 g5583 ( .a(_net_6072), .o(n1827) );
bf01f01 g5584 ( .a(x1432), .o(n1836) );
bf01f01 g5585 ( .a(x1382), .o(n1855) );
bf01f01 g5586 ( .a(net_6699), .o(n1865) );
bf01f01 g5587 ( .a(net_6599), .o(n1874) );
bf01f01 g5588 ( .a(_net_6082), .o(n1903) );
bf01f01 g5589 ( .a(_net_7816), .o(n1913) );
bf01f01 g5590 ( .a(net_7116), .o(n1918) );
bf01f01 g5591 ( .a(net_6995), .o(n1932) );
bf01f01 g5592 ( .a(net_6433), .o(n1941) );
bf01f01 g5593 ( .a(_net_7817), .o(n1954) );
bf01f01 g5594 ( .a(_net_6150), .o(n1964) );
bf01f01 g5595 ( .a(_net_7803), .o(n1973) );
bf01f01 g5596 ( .a(_net_7804), .o(n1978) );
bf01f01 g5597 ( .a(_net_6098), .o(n1983) );
bf01f01 g5598 ( .a(net_6737), .o(n1998) );
bf01f01 g5599 ( .a(_net_6107), .o(n2002) );
bf01f01 g5600 ( .a(_net_7815), .o(n2007) );
bf01f01 g5601 ( .a(_net_7818), .o(n2011) );
bf01f01 g5602 ( .a(_net_6122), .o(n2031) );
bf01f01 g5603 ( .a(net_6394), .o(n2036) );
bf01f01 g5604 ( .a(net_7391), .o(n2051) );
bf01f01 g5605 ( .a(net_7799), .o(n2074) );
bf01f01 g5606 ( .a(_net_5968), .o(n2079) );
bf01f01 g5607 ( .a(_net_7796), .o(n2088) );
bf01f01 g5608 ( .a(_net_7793), .o(n2093) );
bf01f01 g5609 ( .a(net_6709), .o(n2098) );
bf01f01 g5610 ( .a(net_6741), .o(n2102) );
bf01f01 g5611 ( .a(net_6056), .o(n2106) );
bf01f01 g5612 ( .a(net_7003), .o(n2111) );
bf01f01 g5613 ( .a(net_6452), .o(n2115) );
bf01f01 g5614 ( .a(net_6603), .o(n2119) );
bf01f01 g5615 ( .a(_net_7809), .o(n2122) );
bf01f01 g5616 ( .a(_net_6114), .o(n2127) );
bf01f01 g5617 ( .a(net_7147), .o(n2132) );
bf01f01 g5618 ( .a(net_6730), .o(n2136) );
bf01f01 g5619 ( .a(_net_7809), .o(n2144) );
bf01f01 g5620 ( .a(net_7144), .o(n2149) );
no02f01 g5621 ( .a(n6966), .b(n7250), .o(n2152) );
bf01f01 g5622 ( .a(_net_6140), .o(n2157) );
bf01f01 g5623 ( .a(net_6443), .o(n2186) );
bf01f01 g5624 ( .a(_net_7813), .o(n2189) );
bf01f01 g5625 ( .a(_net_7796), .o(n2203) );
bf01f01 g5626 ( .a(net_6456), .o(n2218) );
no02f01 g5627 ( .a(n6966), .b(n7351), .o(n2260) );
bf01f01 g5628 ( .a(net_6397), .o(n2284) );
bf01f01 g5629 ( .a(_net_7805), .o(n2288) );
bf01f01 g5630 ( .a(_net_6170), .o(n2293) );
bf01f01 g5631 ( .a(_net_7824), .o(n2307) );
bf01f01 g5632 ( .a(_net_7800), .o(n2316) );
bf01f01 g5633 ( .a(net_7159), .o(n2321) );
bf01f01 g5634 ( .a(net_6398), .o(n2324) );
bf01f01 g5635 ( .a(_net_7820), .o(n2338) );
bf01f01 g5636 ( .a(_net_7806), .o(n2342) );
bf01f01 g5637 ( .a(net_6849), .o(n2347) );
bf01f01 g5638 ( .a(net_142), .o(n2350) );
bf01f01 g5639 ( .a(_net_6101), .o(n2355) );
bf01f01 g5640 ( .a(_net_7812), .o(n2360) );
bf01f01 g5641 ( .a(net_6593), .o(n2370) );
bf01f01 g5642 ( .a(net_6397), .o(n2373) );
no02f01 g5643 ( .a(n6867_1), .b(n7978), .o(n2381) );
bf01f01 g5644 ( .a(net_6576), .o(n2391) );
bf01f01 g5645 ( .a(_net_7793), .o(n2399) );
bf01f01 g5646 ( .a(_net_7818), .o(n2417) );
bf01f01 g5647 ( .a(net_7016), .o(n2422) );
bf01f01 g5648 ( .a(net_6833), .o(n2426) );
bf01f01 g5649 ( .a(net_7240), .o(n2440) );
bf01f01 g5650 ( .a(net_6392), .o(n2448) );
bf01f01 g5651 ( .a(_net_7824), .o(n2452) );
bf01f01 g5652 ( .a(net_6426), .o(n2462) );
bf01f01 g5653 ( .a(_net_7818), .o(n2465) );
bf01f01 g5654 ( .a(_net_7810), .o(n2474) );
bf01f01 g5655 ( .a(net_7799), .o(n2488) );
bf01f01 g5656 ( .a(net_6435), .o(n2493) );
bf01f01 g5657 ( .a(_net_7805), .o(n2496) );
no02f01 g5658 ( .a(n6966), .b(n7351), .o(n2500) );
bf01f01 g5659 ( .a(_net_7795), .o(n2519) );
bf01f01 g5660 ( .a(_net_7797), .o(n2539) );
bf01f01 g5661 ( .a(net_7807), .o(n2543) );
no02f01 g5662 ( .a(n6899_1), .b(n7069), .o(n2547) );
bf01f01 g5663 ( .a(_net_7819), .o(n2556) );
bf01f01 g5664 ( .a(net_6390), .o(n2561) );
bf01f01 g5665 ( .a(_net_7798), .o(n2570) );
bf01f01 g5666 ( .a(net_6390), .o(n2594) );
bf01f01 g5667 ( .a(_net_7797), .o(n2597) );
bf01f01 g5668 ( .a(_net_7822), .o(n2601) );
bf01f01 g5669 ( .a(_net_7818), .o(n2605) );
bf01f01 g5670 ( .a(_net_6181), .o(n2610) );
bf01f01 g5671 ( .a(net_6967), .o(n2615) );
bf01f01 g5672 ( .a(_net_7793), .o(n2618) );
bf01f01 g5673 ( .a(_net_7822), .o(n2622) );
bf01f01 g5674 ( .a(_net_6126), .o(n2627) );
bf01f01 g5675 ( .a(_net_6145), .o(n2642) );
bf01f01 g5676 ( .a(net_6588), .o(n2647) );
bf01f01 g5677 ( .a(net_6606), .o(n2656) );
bf01f01 g5678 ( .a(net_149), .o(n2660) );
bf01f01 g5679 ( .a(_net_6134), .o(n2670) );
bf01f01 g5680 ( .a(net_6890), .o(n2675) );
bf01f01 g5681 ( .a(net_6964), .o(n2679) );
bf01f01 g5682 ( .a(_net_7822), .o(n2682) );
bf01f01 g5683 ( .a(net_7393), .o(n2692) );
bf01f01 g5684 ( .a(net_6981), .o(n2701) );
bf01f01 g5685 ( .a(net_6434), .o(n2705) );
bf01f01 g5686 ( .a(net_6969), .o(n2709) );
bf01f01 g5687 ( .a(net_6381), .o(n2727) );
bf01f01 g5688 ( .a(net_7708), .o(n2737) );
bf01f01 g5689 ( .a(net_6586), .o(n2741) );
bf01f01 g5690 ( .a(net_6725), .o(n2745) );
bf01f01 g5691 ( .a(_net_7823), .o(n2748) );
bf01f01 g5692 ( .a(_net_7823), .o(n2762) );
bf01f01 g5693 ( .a(net_7108), .o(n2767) );
bf01f01 g5694 ( .a(net_6880), .o(n2781) );
no02f01 g5695 ( .a(n6899_1), .b(n7509_1), .o(n2784) );
bf01f01 g5696 ( .a(_net_7801), .o(n2788) );
bf01f01 g5697 ( .a(net_7802), .o(n2792) );
bf01f01 g5698 ( .a(_net_7797), .o(n2801) );
bf01f01 g5699 ( .a(x1374), .o(n2805) );
bf01f01 g5700 ( .a(_net_7812), .o(n2814) );
bf01f01 g5701 ( .a(net_6579), .o(n2819) );
bf01f01 g5702 ( .a(net_7024), .o(n2823) );
bf01f01 g5703 ( .a(net_7153), .o(n2827) );
bf01f01 g5704 ( .a(_net_7801), .o(n2840) );
bf01f01 g5705 ( .a(net_7236), .o(n2860) );
bf01f01 g5706 ( .a(_net_6070), .o(n2864) );
bf01f01 g5707 ( .a(net_6478), .o(n2869) );
bf01f01 g5708 ( .a(net_6578), .o(n2873) );
bf01f01 g5709 ( .a(_net_6068), .o(n2877) );
bf01f01 g5710 ( .a(net_7547), .o(n2882) );
bf01f01 g5711 ( .a(_net_7816), .o(n2885) );
bf01f01 g5712 ( .a(_net_5972), .o(n2895) );
no02f01 g5713 ( .a(n6867_1), .b(n6974_1), .o(n2904) );
bf01f01 g5714 ( .a(_net_7814), .o(n2908) );
bf01f01 g5715 ( .a(net_7022), .o(n2922) );
bf01f01 g5716 ( .a(net_6755), .o(n2926) );
bf01f01 g5717 ( .a(net_390), .o(n2935) );
bf01f01 g5718 ( .a(_net_7816), .o(n2939) );
bf01f01 g5719 ( .a(net_7158), .o(n2944) );
bf01f01 g5720 ( .a(_net_6142), .o(n2963) );
bf01f01 g5721 ( .a(net_6392), .o(n2967) );
bf01f01 g5722 ( .a(net_7007), .o(n2972) );
bf01f01 g5723 ( .a(net_6438), .o(n2996) );
bf01f01 g5724 ( .a(net_7105), .o(n3030) );
bf01f01 g5725 ( .a(_net_7806), .o(n3033) );
bf01f01 g5726 ( .a(_net_7809), .o(n3037) );
bf01f01 g5727 ( .a(net_7136), .o(n3052) );
bf01f01 g5728 ( .a(net_7121), .o(n3061) );
bf01f01 g5729 ( .a(_net_7806), .o(n3069) );
bf01f01 g5730 ( .a(net_6717), .o(n3074) );
bf01f01 g5731 ( .a(net_7799), .o(n3082) );
bf01f01 g5732 ( .a(net_6706), .o(n3102) );
bf01f01 g5733 ( .a(net_6396), .o(n3105) );
bf01f01 g5734 ( .a(net_6473), .o(n3110) );
bf01f01 g5735 ( .a(net_6743), .o(n3114) );
bf01f01 g5736 ( .a(_net_7824), .o(n3117) );
no02f01 g5737 ( .a(n6966), .b(n7599_1), .o(n3121) );
bf01f01 g5738 ( .a(net_7387), .o(n3126) );
bf01f01 g5739 ( .a(_net_7809), .o(n3134) );
bf01f01 g5740 ( .a(_net_7819), .o(n3143) );
bf01f01 g5741 ( .a(_net_7805), .o(n3152) );
bf01f01 g5742 ( .a(net_6751), .o(n3162) );
in01f01 g5743 ( .a(n7343), .o(n3165) );
bf01f01 g5744 ( .a(_net_7815), .o(n3174) );
bf01f01 g5745 ( .a(net_6450), .o(n3178) );
bf01f01 g5746 ( .a(_net_7798), .o(n3186) );
bf01f01 g5747 ( .a(net_6861), .o(n3190) );
bf01f01 g5748 ( .a(net_7536), .o(n3199) );
bf01f01 g5749 ( .a(_net_7793), .o(n3207) );
bf01f01 g5750 ( .a(net_139), .o(n3226) );
bf01f01 g5751 ( .a(x1443), .o(n3235) );
bf01f01 g5752 ( .a(_net_7822), .o(n3244) );
bf01f01 g5753 ( .a(_net_6083), .o(n3249) );
bf01f01 g5754 ( .a(x1366), .o(n3258) );
bf01f01 g5755 ( .a(net_7799), .o(n3272) );
no02f01 g5756 ( .a(n6867_1), .b(n8170_1), .o(n3276) );
bf01f01 g5757 ( .a(_net_7795), .o(n3280) );
bf01f01 g5758 ( .a(net_7710), .o(n3290) );
bf01f01 g5759 ( .a(_net_7793), .o(n3299) );
bf01f01 g5760 ( .a(_net_7809), .o(n3303) );
bf01f01 g5761 ( .a(net_6883), .o(n3318) );
no02f01 g5762 ( .a(n6899_1), .b(n7173), .o(n3325) );
bf01f01 g5763 ( .a(net_6868), .o(n3330) );
no02f01 g5764 ( .a(n6899_1), .b(n7254), .o(n3333) );
bf01f01 g5765 ( .a(_net_6063), .o(n3343) );
bf01f01 g5766 ( .a(net_7140), .o(n3348) );
bf01f01 g5767 ( .a(_net_6071), .o(n3361) );
bf01f01 g5768 ( .a(_net_7821), .o(n3365) );
no02f01 g5769 ( .a(n6867_1), .b(n7650), .o(n3374) );
bf01f01 g5770 ( .a(net_6698), .o(n3379) );
bf01f01 g5771 ( .a(net_6485), .o(n3383) );
bf01f01 g5772 ( .a(net_7807), .o(n3386) );
bf01f01 g5773 ( .a(x1424), .o(n3390) );
bf01f01 g5774 ( .a(net_6386), .o(n3404) );
bf01f01 g5775 ( .a(_net_7820), .o(n3408) );
bf01f01 g5776 ( .a(net_148), .o(n3413) );
bf01f01 g5777 ( .a(net_7248), .o(n3418) );
in01f01 g5778 ( .a(n7343), .o(n3431) );
bf01f01 g5779 ( .a(net_7120), .o(n3436) );
bf01f01 g5780 ( .a(net_6389), .o(n3445) );
bf01f01 g5781 ( .a(_net_6173), .o(n3450) );
bf01f01 g5782 ( .a(_net_7811), .o(n3469) );
bf01f01 g5783 ( .a(_net_6136), .o(n3479) );
bf01f01 g5784 ( .a(net_7241), .o(n3494) );
bf01f01 g5785 ( .a(_net_7803), .o(n3497) );
bf01f01 g5786 ( .a(_net_263), .o(n3502) );
bf01f01 g5787 ( .a(_net_7793), .o(n3511) );
bf01f01 g5788 ( .a(_net_7800), .o(n3520) );
bf01f01 g5789 ( .a(net_150), .o(n3524) );
bf01f01 g5790 ( .a(_net_7815), .o(n3528) );
bf01f01 g5791 ( .a(net_6384), .o(n3532) );
bf01f01 g5792 ( .a(_net_6078), .o(n3537) );
bf01f01 g5793 ( .a(net_6885), .o(n3542) );
bf01f01 g5794 ( .a(net_6385), .o(n3555) );
bf01f01 g5795 ( .a(_net_7810), .o(n3559) );
bf01f01 g5796 ( .a(net_6873), .o(n3564) );
no02f01 g5797 ( .a(n6966), .b(n8514), .o(n3567) );
bf01f01 g5798 ( .a(net_6476), .o(n3587) );
bf01f01 g5799 ( .a(_net_7803), .o(n3590) );
bf01f01 g5800 ( .a(net_6583), .o(n3600) );
bf01f01 g5801 ( .a(_net_7812), .o(n3618) );
bf01f01 g5802 ( .a(_net_6124), .o(n3623) );
in01f01 g5803 ( .a(n7343), .o(n3642) );
bf01f01 g5804 ( .a(net_7157), .o(n3651) );
bf01f01 g5805 ( .a(net_6591), .o(n3655) );
bf01f01 g5806 ( .a(net_6394), .o(n3658) );
no02f01 g5807 ( .a(n6867_1), .b(n8173), .o(n3661) );
bf01f01 g5808 ( .a(_net_7794), .o(n3670) );
bf01f01 g5809 ( .a(_net_7801), .o(n3679) );
bf01f01 g5810 ( .a(net_6605), .o(n3689) );
bf01f01 g5811 ( .a(net_6976), .o(n3703) );
bf01f01 g5812 ( .a(net_6721), .o(n3707) );
bf01f01 g5813 ( .a(net_6486), .o(n3716) );
bf01f01 g5814 ( .a(_net_6092), .o(n3720) );
bf01f01 g5815 ( .a(net_6881), .o(n3725) );
bf01f01 g5816 ( .a(_net_7813), .o(n3729) );
bf01f01 g5817 ( .a(x1550), .o(n3733) );
bf01f01 g5818 ( .a(_net_6129), .o(n3747) );
bf01f01 g5819 ( .a(_net_6069), .o(n3752) );
bf01f01 g5820 ( .a(net_6391), .o(n3756) );
bf01f01 g5821 ( .a(net_6442), .o(n3761) );
bf01f01 g5822 ( .a(net_6991), .o(n3770) );
bf01f01 g5823 ( .a(_net_7796), .o(n3773) );
bf01f01 g5824 ( .a(_net_7798), .o(n3777) );
bf01f01 g5825 ( .a(_net_7804), .o(n3791) );
bf01f01 g5826 ( .a(net_7149), .o(n3801) );
bf01f01 g5827 ( .a(net_7714), .o(n3805) );
bf01f01 g5828 ( .a(net_6429), .o(n3809) );
bf01f01 g5829 ( .a(net_6394), .o(n3817) );
bf01f01 g5830 ( .a(_net_6076), .o(n3822) );
bf01f01 g5831 ( .a(net_7802), .o(n3831) );
bf01f01 g5832 ( .a(net_6829), .o(n3851) );
bf01f01 g5833 ( .a(net_6595), .o(n3855) );
bf01f01 g5834 ( .a(net_6850), .o(n3864) );
bf01f01 g5835 ( .a(_net_7806), .o(n3867) );
bf01f01 g5836 ( .a(net_7799), .o(n3881) );
bf01f01 g5837 ( .a(net_6855), .o(n3896) );
bf01f01 g5838 ( .a(net_7799), .o(n3899) );
bf01f01 g5839 ( .a(net_7239), .o(n3904) );
bf01f01 g5840 ( .a(_net_7814), .o(n3917) );
bf01f01 g5841 ( .a(_net_7823), .o(n3936) );
bf01f01 g5842 ( .a(net_6384), .o(n3945) );
bf01f01 g5843 ( .a(_net_7822), .o(n3949) );
bf01f01 g5844 ( .a(_net_7815), .o(n3953) );
bf01f01 g5845 ( .a(net_6387), .o(n3957) );
bf01f01 g5846 ( .a(_net_6176), .o(n3962) );
bf01f01 g5847 ( .a(net_7537), .o(n3972) );
bf01f01 g5848 ( .a(_net_7815), .o(n3985) );
bf01f01 g5849 ( .a(net_6392), .o(n3989) );
bf01f01 g5850 ( .a(_net_7795), .o(n3993) );
bf01f01 g5851 ( .a(_net_7817), .o(n4002) );
bf01f01 g5852 ( .a(net_6852), .o(n4007) );
bf01f01 g5853 ( .a(_net_6103), .o(n4011) );
bf01f01 g5854 ( .a(_net_7813), .o(n4020) );
bf01f01 g5855 ( .a(_net_7804), .o(n4024) );
bf01f01 g5856 ( .a(_net_7821), .o(n4033) );
bf01f01 g5857 ( .a(_net_7793), .o(n4037) );
bf01f01 g5858 ( .a(net_6390), .o(n4046) );
bf01f01 g5859 ( .a(net_6613), .o(n4051) );
bf01f01 g5860 ( .a(net_7711), .o(n4055) );
bf01f01 g5861 ( .a(net_7013), .o(n4059) );
bf01f01 g5862 ( .a(net_6444), .o(n4068) );
bf01f01 g5863 ( .a(_net_7814), .o(n4071) );
bf01f01 g5864 ( .a(net_6399), .o(n4075) );
no02f01 g5865 ( .a(n6966), .b(n7188), .o(n4079) );
bf01f01 g5866 ( .a(_net_7798), .o(n4098) );
bf01f01 g5867 ( .a(_net_7813), .o(n4102) );
bf01f01 g5868 ( .a(net_6867), .o(n4112) );
bf01f01 g5869 ( .a(net_7400), .o(n4131) );
bf01f01 g5870 ( .a(net_6592), .o(n4145) );
bf01f01 g5871 ( .a(_net_7793), .o(n4148) );
bf01f01 g5872 ( .a(net_145), .o(n4153) );
bf01f01 g5873 ( .a(net_6714), .o(n4158) );
bf01f01 g5874 ( .a(net_6382), .o(n4161) );
bf01f01 g5875 ( .a(_net_6087), .o(n4176) );
bf01f01 g5876 ( .a(net_7123), .o(n4191) );
bf01f01 g5877 ( .a(_net_7822), .o(n4194) );
bf01f01 g5878 ( .a(net_6447), .o(n4199) );
bf01f01 g5879 ( .a(_net_7808), .o(n4207) );
bf01f01 g5880 ( .a(_net_7814), .o(n4221) );
bf01f01 g5881 ( .a(net_5858), .o(n4231) );
bf01f01 g5882 ( .a(_net_7813), .o(n4235) );
bf01f01 g5883 ( .a(net_7398), .o(n4245) );
bf01f01 g5884 ( .a(net_6391), .o(n4253) );
bf01f01 g5885 ( .a(_net_7816), .o(n4258) );
bf01f01 g5886 ( .a(_net_7796), .o(n4267) );
bf01f01 g5887 ( .a(net_6387), .o(n4271) );
bf01f01 g5888 ( .a(_net_7794), .o(n4280) );
bf01f01 g5889 ( .a(x1459), .o(n4284) );
bf01f01 g5890 ( .a(net_6753), .o(n4309) );
bf01f01 g5891 ( .a(net_6471), .o(n4318) );
bf01f01 g5892 ( .a(net_6387), .o(n4326) );
bf01f01 g5893 ( .a(net_6978), .o(n4330) );
no02f01 g5894 ( .a(n6966), .b(n8899_1), .o(n4333) );
bf01f01 g5895 ( .a(_net_7808), .o(n4338) );
bf01f01 g5896 ( .a(_net_7791), .o(n4343) );
no02f01 g5897 ( .a(n6966), .b(n7891), .o(n4352) );
bf01f01 g5898 ( .a(net_6863), .o(n4362) );
bf01f01 g5899 ( .a(_net_7797), .o(n4365) );
bf01f01 g5900 ( .a(_net_7811), .o(n4370) );
bf01f01 g5901 ( .a(_net_7818), .o(n4374) );
bf01f01 g5902 ( .a(net_6974), .o(n4384) );
bf01f01 g5903 ( .a(net_6431), .o(n4388) );
bf01f01 g5904 ( .a(net_6564), .o(n4397) );
bf01f01 g5905 ( .a(net_7162), .o(n4401) );
bf01f01 g5906 ( .a(net_7111), .o(n4410) );
bf01f01 g5907 ( .a(_net_6151), .o(n4419) );
no02f01 g5908 ( .a(n6899_1), .b(n7507), .o(n4428) );
bf01f01 g5909 ( .a(net_6886), .o(n4448) );
no02f01 g5910 ( .a(n6899_1), .b(n7173), .o(n4451) );
in01f01 g5911 ( .a(n7343), .o(n4459) );
bf01f01 g5912 ( .a(_net_6147), .o(n4469) );
bf01f01 g5913 ( .a(_net_7797), .o(n4473) );
bf01f01 g5914 ( .a(net_6448), .o(n4478) );
bf01f01 g5915 ( .a(net_7129), .o(n4487) );
bf01f01 g5916 ( .a(net_386), .o(n4496) );
bf01f01 g5917 ( .a(_net_7808), .o(n4505) );
bf01f01 g5918 ( .a(_net_7801), .o(n4524) );
bf01f01 g5919 ( .a(_net_7794), .o(n4548) );
bf01f01 g5920 ( .a(_net_7809), .o(n4558) );
bf01f01 g5921 ( .a(_net_7796), .o(n4562) );
bf01f01 g5922 ( .a(net_131), .o(n4567) );
bf01f01 g5923 ( .a(_net_6109), .o(n4577) );
bf01f01 g5924 ( .a(_net_7812), .o(n4581) );
bf01f01 g5925 ( .a(_net_7801), .o(n4600) );
bf01f01 g5926 ( .a(_net_7805), .o(n4604) );
bf01f01 g5927 ( .a(_net_7811), .o(n4613) );
bf01f01 g5928 ( .a(net_7807), .o(n4617) );
bf01f01 g5929 ( .a(_net_6097), .o(n4622) );
bf01f01 g5930 ( .a(_net_7821), .o(n4631) );
bf01f01 g5931 ( .a(_net_6171), .o(n4651) );
bf01f01 g5932 ( .a(_net_7795), .o(n4660) );
bf01f01 g5933 ( .a(net_6736), .o(n4665) );
bf01f01 g5934 ( .a(net_6581), .o(n4669) );
bf01f01 g5935 ( .a(x1564), .o(n4681) );
bf01f01 g5936 ( .a(net_6393), .o(n4686) );
no02f01 g5937 ( .a(n6899_1), .b(n7560), .o(n4690) );
no02f01 g5938 ( .a(n6867_1), .b(n6974_1), .o(n4694) );
bf01f01 g5939 ( .a(net_6993), .o(n4699) );
bf01f01 g5940 ( .a(net_7142), .o(n4713) );
bf01f01 g5941 ( .a(_net_7817), .o(n4717) );
bf01f01 g5942 ( .a(_net_6095), .o(n4722) );
bf01f01 g5943 ( .a(net_6735), .o(n4742) );
bf01f01 g5944 ( .a(net_7807), .o(n4745) );
bf01f01 g5945 ( .a(_net_6138), .o(n4750) );
bf01f01 g5946 ( .a(_net_6153), .o(n4755) );
bf01f01 g5947 ( .a(net_137), .o(n4765) );
no02f01 g5948 ( .a(n6867_1), .b(n7203_1), .o(n4769) );
bf01f01 g5949 ( .a(net_7545), .o(n4774) );
bf01f01 g5950 ( .a(net_6449), .o(n4778) );
bf01f01 g5951 ( .a(_net_6156), .o(n4782) );
bf01f01 g5952 ( .a(net_7799), .o(n4791) );
bf01f01 g5953 ( .a(_net_7803), .o(n4795) );
bf01f01 g5954 ( .a(net_7014), .o(n4805) );
bf01f01 g5955 ( .a(net_7128), .o(n4814) );
no02f01 g5956 ( .a(n6899_1), .b(n8826_1), .o(n4822) );
bf01f01 g5957 ( .a(net_6567), .o(n4827) );
bf01f01 g5958 ( .a(_net_7820), .o(n4834) );
bf01f01 g5959 ( .a(_net_7814), .o(n4838) );
bf01f01 g5960 ( .a(_net_6074), .o(n4848) );
bf01f01 g5961 ( .a(net_6875), .o(n4853) );
bf01f01 g5962 ( .a(_net_6402), .o(n4862) );
bf01f01 g5963 ( .a(_net_7819), .o(n4867) );
bf01f01 g5964 ( .a(net_6384), .o(n4881) );
bf01f01 g5965 ( .a(_net_7801), .o(n4890) );
bf01f01 g5966 ( .a(net_7154), .o(n4895) );
bf01f01 g5967 ( .a(_net_6143), .o(n4899) );
bf01f01 g5968 ( .a(net_7001), .o(n4904) );
bf01f01 g5969 ( .a(net_6573), .o(n4913) );
bf01f01 g5970 ( .a(_net_7823), .o(n4931) );
bf01f01 g5971 ( .a(_net_7812), .o(n4940) );
bf01f01 g5972 ( .a(net_7807), .o(n4944) );
bf01f01 g5973 ( .a(_net_7818), .o(n4947) );
bf01f01 g5974 ( .a(net_6718), .o(n4957) );
bf01f01 g5975 ( .a(_net_7823), .o(n4965) );
bf01f01 g5976 ( .a(_net_7811), .o(n4969) );
bf01f01 g5977 ( .a(net_6484), .o(n4979) );
bf01f01 g5978 ( .a(net_6858), .o(n4983) );
bf01f01 g5979 ( .a(_net_6065), .o(n4996) );
bf01f01 g5980 ( .a(net_6617), .o(n5001) );
bf01f01 g5981 ( .a(net_6854), .o(n5005) );
bf01f01 g5982 ( .a(net_6386), .o(n5008) );
bf01f01 g5983 ( .a(net_7539), .o(n5023) );
bf01f01 g5984 ( .a(_net_7819), .o(n5031) );
bf01f01 g5985 ( .a(_net_7817), .o(n5035) );
bf01f01 g5986 ( .a(net_7399), .o(n5045) );
no02f01 g5987 ( .a(n6966), .b(n7891), .o(n5048) );
bf01f01 g5988 ( .a(net_6970), .o(n5053) );
no02f01 g5989 ( .a(n6899_1), .b(n7254), .o(n5056) );
bf01f01 g5990 ( .a(_net_6115), .o(n5066) );
bf01f01 g5991 ( .a(_net_7801), .o(n5070) );
bf01f01 g5992 ( .a(net_7011), .o(n5090) );
bf01f01 g5993 ( .a(net_6399), .o(n5098) );
bf01f01 g5994 ( .a(net_6391), .o(n5121) );
bf01f01 g5995 ( .a(net_6589), .o(n5126) );
bf01f01 g5996 ( .a(net_6985), .o(n5139) );
bf01f01 g5997 ( .a(net_6572), .o(n5148) );
bf01f01 g5998 ( .a(_net_7821), .o(n5151) );
bf01f01 g5999 ( .a(net_6428), .o(n5156) );
bf01f01 g6000 ( .a(_net_7793), .o(n5159) );
bf01f01 g6001 ( .a(_net_7808), .o(n5173) );
bf01f01 g6002 ( .a(net_6841), .o(n5178) );
bf01f01 g6003 ( .a(x1519), .o(n5181) );
bf01f01 g6004 ( .a(net_7691), .o(n5186) );
bf01f01 g6005 ( .a(_net_7794), .o(n5189) );
bf01f01 g6006 ( .a(net_7802), .o(n5193) );
bf01f01 g6007 ( .a(_net_7811), .o(n5202) );
bf01f01 g6008 ( .a(net_6569), .o(n5217) );
bf01f01 g6009 ( .a(net_6857), .o(n5221) );
bf01f01 g6010 ( .a(_net_7806), .o(n5234) );
bf01f01 g6011 ( .a(net_6487), .o(n5239) );
bf01f01 g6012 ( .a(_net_7814), .o(n5242) );
bf01f01 g6013 ( .a(_net_7797), .o(n5246) );
bf01f01 g6014 ( .a(net_6843), .o(n5261) );
bf01f01 g6015 ( .a(_net_7798), .o(n5269) );
bf01f01 g6016 ( .a(net_6395), .o(n5288) );
bf01f01 g6017 ( .a(net_6965), .o(n5298) );
bf01f01 g6018 ( .a(_net_6128), .o(n5302) );
bf01f01 g6019 ( .a(net_7006), .o(n5312) );
bf01f01 g6020 ( .a(net_6844), .o(n5326) );
bf01f01 g6021 ( .a(net_7002), .o(n5335) );
bf01f01 g6022 ( .a(_net_6161), .o(n5339) );
bf01f01 g6023 ( .a(net_6987), .o(n5349) );
bf01f01 g6024 ( .a(net_6454), .o(n5358) );
bf01f01 g6025 ( .a(net_6460), .o(n5362) );
bf01f01 g6026 ( .a(net_6860), .o(n5366) );
bf01f01 g6027 ( .a(net_143), .o(n5375) );
bf01f01 g6028 ( .a(net_6729), .o(n5380) );
bf01f01 g6029 ( .a(_net_7819), .o(n5383) );
bf01f01 g6030 ( .a(net_7021), .o(n5393) );
bf01f01 g6031 ( .a(net_7151), .o(n5402) );
bf01f01 g6032 ( .a(_net_7804), .o(n5415) );
bf01f01 g6033 ( .a(_net_7797), .o(n5424) );
bf01f01 g6034 ( .a(_net_7801), .o(n5433) );
bf01f01 g6035 ( .a(net_6395), .o(n5437) );
bf01f01 g6036 ( .a(_net_7824), .o(n5441) );
bf01f01 g6037 ( .a(net_6436), .o(n5451) );
bf01f01 g6038 ( .a(_net_6075), .o(n5460) );
no02f01 g6039 ( .a(n6899_1), .b(n7246), .o(n5464) );
bf01f01 g6040 ( .a(net_6610), .o(n5469) );
no02f01 g6041 ( .a(n6966), .b(n7520), .o(n5472) );
bf01f01 g6042 ( .a(_net_7815), .o(n5481) );
bf01f01 g6043 ( .a(net_387), .o(n5486) );
bf01f01 g6044 ( .a(net_6575), .o(n5500) );
bf01f01 g6045 ( .a(net_7100), .o(n5504) );
bf01f01 g6046 ( .a(net_6024), .o(n5513) );
bf01f01 g6047 ( .a(net_7018), .o(n5521) );
bf01f01 g6048 ( .a(net_6839), .o(n5539) );
bf01f01 g6049 ( .a(_net_7808), .o(n5547) );
bf01f01 g6050 ( .a(net_6398), .o(n5556) );
bf01f01 g6051 ( .a(_net_7824), .o(n5560) );
bf01f01 g6052 ( .a(net_6620), .o(n5575) );
bf01f01 g6053 ( .a(net_7546), .o(n5584) );
bf01f01 g6054 ( .a(net_7235), .o(n5588) );
no02f01 g6055 ( .a(n6966), .b(n8514), .o(n5591) );
bf01f01 g6056 ( .a(_net_6172), .o(n5606) );
bf01f01 g6057 ( .a(_net_7796), .o(n5610) );
bf01f01 g6058 ( .a(_net_7813), .o(n5613) );
bf01f01 g6059 ( .a(_net_6067), .o(n5618) );
bf01f01 g6060 ( .a(net_6983), .o(n5648) );
bf01f01 g6061 ( .a(_net_7800), .o(n5651) );
bf01f01 g6062 ( .a(_net_7795), .o(n5655) );
bf01f01 g6063 ( .a(_net_7813), .o(n5664) );
bf01f01 g6064 ( .a(net_6727), .o(n5679) );
bf01f01 g6065 ( .a(_net_7795), .o(n5682) );
bf01f01 g6066 ( .a(x1358), .o(n5686) );
bf01f01 g6067 ( .a(net_6609), .o(n5696) );
bf01f01 g6068 ( .a(_net_7810), .o(n5704) );
bf01f01 g6069 ( .a(_net_7806), .o(n5713) );
bf01f01 g6070 ( .a(_net_7796), .o(n5717) );
bf01f01 g6071 ( .a(net_6598), .o(n5727) );
bf01f01 g6072 ( .a(net_7107), .o(n5731) );
bf01f01 g6073 ( .a(net_7026), .o(n5735) );
bf01f01 g6074 ( .a(net_7244), .o(n5744) );
bf01f01 g6075 ( .a(_net_6131), .o(n5758) );
bf01f01 g6076 ( .a(net_6560), .o(n5763) );
bf01f01 g6077 ( .a(net_6590), .o(n5767) );
bf01f01 g6078 ( .a(net_6480), .o(n5771) );
bf01f01 g6079 ( .a(_net_7812), .o(n5779) );
bf01f01 g6080 ( .a(net_6388), .o(n5783) );
bf01f01 g6081 ( .a(_net_7814), .o(n5787) );
bf01f01 g6082 ( .a(net_7802), .o(n5796) );
bf01f01 g6083 ( .a(net_7012), .o(n5801) );
bf01f01 g6084 ( .a(net_6437), .o(n5805) );
bf01f01 g6085 ( .a(net_7113), .o(n5824) );
bf01f01 g6086 ( .a(net_6878), .o(n5833) );
bf01f01 g6087 ( .a(net_7802), .o(n5836) );
bf01f01 g6088 ( .a(_net_7793), .o(n5840) );
bf01f01 g6089 ( .a(net_6479), .o(n5860) );
bf01f01 g6090 ( .a(net_7102), .o(n5864) );
no02f01 g6091 ( .a(n6899_1), .b(n7560), .o(n5867) );
bf01f01 g6092 ( .a(_net_6144), .o(n5872) );
bf01f01 g6093 ( .a(_net_7822), .o(n5876) );
bf01f01 g6094 ( .a(net_6720), .o(n5881) );
bf01f01 g6095 ( .a(net_6391), .o(n5894) );
bf01f01 g6096 ( .a(net_7790), .o(n5903) );
bf01f01 g6097 ( .a(_net_6180), .o(n5908) );
bf01f01 g6098 ( .a(_net_7811), .o(n5912) );
bf01f01 g6099 ( .a(net_6971), .o(n5917) );
bf01f01 g6100 ( .a(_net_7795), .o(n5920) );
bf01f01 g6101 ( .a(net_6580), .o(n5930) );
bf01f01 g6102 ( .a(net_7127), .o(n5934) );
bf01f01 g6103 ( .a(net_6887), .o(n5943) );
bf01f01 g6104 ( .a(net_6562), .o(n5947) );
bf01f01 g6105 ( .a(net_6973), .o(n5951) );
bf01f01 g6106 ( .a(_net_6079), .o(n5955) );
bf01f01 g6107 ( .a(x1557), .o(n5964) );
bf01f01 g6108 ( .a(_net_7821), .o(n5968) );
bf01f01 g6109 ( .a(net_6618), .o(n5978) );
bf01f01 g6110 ( .a(net_7712), .o(n6002) );
bf01f01 g6111 ( .a(net_7115), .o(n6006) );
bf01f01 g6112 ( .a(net_7802), .o(n6009) );
bf01f01 g6113 ( .a(net_5861), .o(n6014) );
bf01f01 g6114 ( .a(_net_6118), .o(n6019) );
bf01f01 g6115 ( .a(net_7125), .o(n6034) );
bf01f01 g6116 ( .a(net_6733), .o(n6043) );
bf01f01 g6117 ( .a(_net_6166), .o(n6047) );
bf01f01 g6118 ( .a(_net_7805), .o(n6056) );
bf01f01 g6119 ( .a(net_6466), .o(n6066) );
bf01f01 g6120 ( .a(_net_7800), .o(n6069) );
bf01f01 g6121 ( .a(x1572), .o(n6078) );
bf01f01 g6122 ( .a(_net_6139), .o(n6098) );
bf01f01 g6123 ( .a(_net_7798), .o(n6102) );
bf01f01 g6124 ( .a(_net_7824), .o(n6106) );
no02f01 g6125 ( .a(n6899_1), .b(n7895), .o(n6110) );
bf01f01 g6126 ( .a(net_7807), .o(n6114) );
bf01f01 g6127 ( .a(_net_7803), .o(n6128) );
bf01f01 g6128 ( .a(x1479), .o(n6132) );
bf01f01 g6129 ( .a(net_6384), .o(n6136) );
bf01f01 g6130 ( .a(net_6594), .o(n6145) );
bf01f01 g6131 ( .a(_net_7800), .o(n6148) );
bf01f01 g6132 ( .a(net_6892), .o(n6158) );
bf01f01 g6133 ( .a(_net_7816), .o(n6161) );
bf01f01 g6134 ( .a(_net_6105), .o(n6176) );
bf01f01 g6135 ( .a(_net_6113), .o(n6181) );
bf01f01 g6136 ( .a(_net_7813), .o(n6195) );
bf01f01 g6137 ( .a(net_6397), .o(n6204) );
bf01f01 g6138 ( .a(net_7385), .o(n6214) );
no02f01 g6139 ( .a(n6966), .b(n7142_1), .o(n6222) );
in01f01 g6140 ( .a(n7343), .o(n6231) );
bf01f01 g6141 ( .a(net_7799), .o(n6235) );
bf01f01 g6142 ( .a(net_6400), .o(n6239) );
bf01f01 g6143 ( .a(net_6697), .o(n6254) );
bf01f01 g6144 ( .a(net_6750), .o(n6258) );
bf01f01 g6145 ( .a(x1534), .o(n6261) );
bf01f01 g6146 ( .a(_net_5964), .o(n6276) );
bf01f01 g6147 ( .a(net_146), .o(n6285) );
bf01f01 g6148 ( .a(net_7130), .o(n6299) );
no02f01 g6149 ( .a(n6867_1), .b(n9980), .o(n6302) );
bf01f01 g6150 ( .a(net_6393), .o(n6306) );
bf01f01 g6151 ( .a(net_7770), .o(n6316) );
bf01f01 g6152 ( .a(net_389), .o(n6319) );
bf01f01 g6153 ( .a(net_7161), .o(n6329) );
bf01f01 g6154 ( .a(net_6396), .o(n6332) );
bf01f01 g6155 ( .a(net_6469), .o(n6342) );
bf01f01 g6156 ( .a(_net_7794), .o(n6350) );
bf01f01 g6157 ( .a(net_6747), .o(n6354) );
bf01f01 g6158 ( .a(_net_7817), .o(n6357) );
bf01f01 g6159 ( .a(net_6439), .o(n6367) );
bf01f01 g6160 ( .a(net_7117), .o(n6386) );
bf01f01 g6161 ( .a(_net_6165), .o(n6390) );
bf01f01 g6162 ( .a(net_6398), .o(n6399) );
bf01f01 g6163 ( .a(net_6738), .o(n6403) );
bf01f01 g6164 ( .a(net_6481), .o(n6407) );
bf01f01 g6165 ( .a(_net_7806), .o(n6415) );
bf01f01 g6166 ( .a(_net_7795), .o(n6419) );
bf01f01 g6167 ( .a(net_6382), .o(n6423) );
bf01f01 g6168 ( .a(net_7802), .o(n6441) );
bf01f01 g6169 ( .a(net_6702), .o(n6446) );
bf01f01 g6170 ( .a(_net_6152), .o(n6460) );
bf01f01 g6171 ( .a(_net_7817), .o(n6464) );
bf01f01 g6172 ( .a(net_6980), .o(n6469) );
bf01f01 g6173 ( .a(_net_7812), .o(n6472) );
bf01f01 g6174 ( .a(net_7148), .o(n6477) );
bf01f01 g6175 ( .a(_net_7796), .o(n6480) );
bf01f01 g6176 ( .a(net_6462), .o(n6485) );
bf01f01 g6177 ( .a(net_7242), .o(n6489) );
bf01f01 g6178 ( .a(_net_6159), .o(n6498) );
bf01f01 g6179 ( .a(net_7807), .o(n6502) );
bf01f01 g6180 ( .a(net_6563), .o(n6507) );
bf01f01 g6181 ( .a(net_6604), .o(n6511) );
bf01f01 g6182 ( .a(net_6836), .o(n6515) );
bf01f01 g6183 ( .a(net_6866), .o(n6519) );
bf01f01 g6184 ( .a(x1501), .o(n6522) );
bf01f01 g6185 ( .a(net_6385), .o(n6531) );
no02f01 g6186 ( .a(n6966), .b(n8812), .o(n6535) );
bf01f01 g6187 ( .a(net_7397), .o(n6550) );
bf01f01 g6188 ( .a(net_6713), .o(n6554) );
bf01f01 g6189 ( .a(net_6846), .o(n6563) );
bf01f01 g6190 ( .a(net_6381), .o(n6566) );
no02f01 g6191 ( .a(n6867_1), .b(n7650), .o(n6574) );
bf01f01 g6192 ( .a(net_132), .o(n6578) );
bf01f01 g6193 ( .a(_net_7817), .o(n6586) );
bf01f01 g6194 ( .a(_net_6096), .o(n6611) );
bf01f01 g6195 ( .a(_net_7817), .o(n6615) );
bf01f01 g6196 ( .a(_net_7793), .o(n6619) );
bf01f01 g6197 ( .a(_net_6085), .o(n6629) );
bf01f01 g6198 ( .a(_net_7817), .o(n6638) );
bf01f01 g6199 ( .a(net_7145), .o(n6648) );
no02f01 g6200 ( .a(n6966), .b(n8812), .o(n6656) );
bf01f01 g6201 ( .a(net_6424), .o(n6661) );
bf01f01 g6202 ( .a(net_6390), .o(n6669) );
bf01f01 g6203 ( .a(net_6834), .o(n6674) );
bf01f01 g6204 ( .a(net_6708), .o(n6678) );
bf01f01 g6205 ( .a(net_6997), .o(n6687) );
bf01f01 g6206 ( .a(_net_6157), .o(n6700) );
bf01f01 g6207 ( .a(_net_7794), .o(n6704) );
bf01f01 g6208 ( .a(_net_7793), .o(n6713) );
bf01f01 g6209 ( .a(_net_7796), .o(n6717) );
bf01f01 g6210 ( .a(_net_7810), .o(n6732) );
bf01f01 g6211 ( .a(net_7799), .o(n6736) );
bf01f01 g6212 ( .a(net_7549), .o(n6746) );
bf01f01 g6213 ( .a(_net_7810), .o(n6749) );
bf01f01 g6214 ( .a(_net_7794), .o(n6752) );
bf01f01 g6215 ( .a(net_6389), .o(n6756) );
bf01f01 g6216 ( .a(net_6728), .o(n6761) );
bf01f01 g6217 ( .a(net_6830), .o(n6770) );
bf01f01 g6218 ( .a(_net_7824), .o(n6783) );
bf01f01 g6219 ( .a(net_7394), .o(n6793) );
bf01f01 g6220 ( .a(_net_7801), .o(n6796) );
bf01f01 g6221 ( .a(net_6990), .o(n6806) );
bf01f01 g6222 ( .a(net_7799), .o(n6809) );
bf01f01 g6223 ( .a(_net_7798), .o(n6813) );
bf01f01 g6224 ( .a(net_6392), .o(n6822) );
bf01f01 g6225 ( .a(_net_7809), .o(n6826) );
bf01f01 g6226 ( .a(net_7025), .o(n6836) );
bf01f01 g6227 ( .a(net_6470), .o(n6860) );
bf01f01 g6228 ( .a(_net_7796), .o(n6863) );
bf01f01 g6229 ( .a(_net_7823), .o(n6867) );
bf01f01 g6230 ( .a(net_7807), .o(n6876) );
bf01f01 g6231 ( .a(net_6712), .o(n6886) );
bf01f01 g6232 ( .a(net_7009), .o(n6895) );
bf01f01 g6233 ( .a(net_6607), .o(n6899) );
bf01f01 g6234 ( .a(net_6395), .o(n6902) );
bf01f01 g6235 ( .a(_net_7804), .o(n6906) );
bf01f01 g6236 ( .a(_net_7818), .o(n6910) );
no02f01 g6237 ( .a(n6899_1), .b(n8964), .o(n6919) );
bf01f01 g6238 ( .a(net_7150), .o(n6934) );
bf01f01 g6239 ( .a(net_6390), .o(n6947) );
bf01f01 g6240 ( .a(net_6587), .o(n6957) );
bf01f01 g6241 ( .a(_net_7812), .o(n6960) );
bf01f01 g6242 ( .a(net_7245), .o(n6974) );
bf01f01 g6243 ( .a(_net_7816), .o(n6977) );
bf01f01 g6244 ( .a(_net_6146), .o(n6982) );
bf01f01 g6245 ( .a(net_7802), .o(n6986) );
bf01f01 g6246 ( .a(_net_7800), .o(n6990) );
bf01f01 g6247 ( .a(net_6621), .o(n7005) );
bf01f01 g6248 ( .a(net_6597), .o(n7009) );
bf01f01 g6249 ( .a(net_7802), .o(n7027) );
bf01f01 g6250 ( .a(net_6388), .o(n7036) );
bf01f01 g6251 ( .a(net_6889), .o(n7041) );
bf01f01 g6252 ( .a(_net_6182), .o(n7045) );
bf01f01 g6253 ( .a(net_6393), .o(n7049) );
bf01f01 g6254 ( .a(_net_7804), .o(n7062) );
bf01f01 g6255 ( .a(net_6872), .o(n7082) );
no02f01 g6256 ( .a(n6867_1), .b(n7175), .o(n7085) );
bf01f01 g6257 ( .a(_net_7811), .o(n7089) );
bf01f01 g6258 ( .a(net_6398), .o(n7093) );
bf01f01 g6259 ( .a(net_7152), .o(n7098) );
bf01f01 g6260 ( .a(_net_7821), .o(n7111) );
bf01f01 g6261 ( .a(_net_6133), .o(n7116) );
bf01f01 g6262 ( .a(_net_7803), .o(n7120) );
bf01f01 g6263 ( .a(net_6561), .o(n7125) );
bf01f01 g6264 ( .a(_net_7798), .o(n7128) );
no02f01 g6265 ( .a(n6867_1), .b(n9870), .o(n7142) );
bf01f01 g6266 ( .a(_net_6073), .o(n7147) );
bf01f01 g6267 ( .a(_net_7816), .o(n7151) );
bf01f01 g6268 ( .a(_net_7824), .o(n7155) );
bf01f01 g6269 ( .a(net_6862), .o(n7160) );
bf01f01 g6270 ( .a(net_141), .o(n7167) );
bf01f01 g6271 ( .a(net_7543), .o(n7182) );
no02f01 g6272 ( .a(n6899_1), .b(n8229), .o(n7185) );
bf01f01 g6273 ( .a(net_6430), .o(n7190) );
bf01f01 g6274 ( .a(net_7238), .o(n7199) );
bf01f01 g6275 ( .a(net_6477), .o(n7203) );
bf01f01 g6276 ( .a(net_6559), .o(n7212) );
bf01f01 g6277 ( .a(_net_7823), .o(n7230) );
bf01f01 g6278 ( .a(x1486), .o(n7249) );
bf01f01 g6279 ( .a(_net_7804), .o(n7252) );
bf01f01 g6280 ( .a(net_7792), .o(n7256) );
bf01f01 g6281 ( .a(_net_7797), .o(n7260) );
bf01f01 g6282 ( .a(_net_7816), .o(n7284) );
bf01f01 g6283 ( .a(net_6397), .o(n7288) );
bf01f01 g6284 ( .a(x1406), .o(n7292) );
bf01f01 g6285 ( .a(net_6869), .o(n7312) );
bf01f01 g6286 ( .a(_net_6178), .o(n7316) );
bf01f01 g6287 ( .a(net_6715), .o(n7326) );
bf01f01 g6288 ( .a(_net_6088), .o(n7330) );
bf01f01 g6289 ( .a(net_5860), .o(n7335) );
bf01f01 g6290 ( .a(_net_7803), .o(n7344) );
bf01f01 g6291 ( .a(net_6058), .o(n7349) );
bf01f01 g6292 ( .a(net_7008), .o(n7359) );
bf01f01 g6293 ( .a(_net_6121), .o(n7368) );
bf01f01 g6294 ( .a(_net_7798), .o(n7372) );
bf01f01 g6295 ( .a(net_134), .o(n7376) );
bf01f01 g6296 ( .a(net_7118), .o(n7391) );
bf01f01 g6297 ( .a(_net_7808), .o(n7404) );
bf01f01 g6298 ( .a(_net_7819), .o(n7408) );
bf01f01 g6299 ( .a(net_6994), .o(n7413) );
bf01f01 g6300 ( .a(_net_6081), .o(n7417) );
bf01f01 g6301 ( .a(_net_6149), .o(n7427) );
bf01f01 g6302 ( .a(net_6700), .o(n7442) );
bf01f01 g6303 ( .a(net_6696), .o(n7446) );
bf01f01 g6304 ( .a(net_6740), .o(n7450) );
bf01f01 g6305 ( .a(_net_7814), .o(n7463) );
bf01f01 g6306 ( .a(_net_6141), .o(n7468) );
bf01f01 g6307 ( .a(_net_7810), .o(n7482) );
bf01f01 g6308 ( .a(net_6726), .o(n7492) );
bf01f01 g6309 ( .a(net_6383), .o(n7505) );
bf01f01 g6310 ( .a(_net_7809), .o(n7509) );
bf01f01 g6311 ( .a(_net_7823), .o(n7513) );
bf01f01 g6312 ( .a(_net_7809), .o(n7522) );
bf01f01 g6313 ( .a(net_6451), .o(n7527) );
bf01f01 g6314 ( .a(_net_7808), .o(n7530) );
bf01f01 g6315 ( .a(net_6757), .o(n7535) );
bf01f01 g6316 ( .a(_net_6090), .o(n7553) );
bf01f01 g6317 ( .a(x1345), .o(n7567) );
bf01f01 g6318 ( .a(_net_6123), .o(n7577) );
bf01f01 g6319 ( .a(_net_7814), .o(n7581) );
no02f01 g6320 ( .a(n6867_1), .b(n10215), .o(n7599) );
bf01f01 g6321 ( .a(net_6716), .o(n7604) );
bf01f01 g6322 ( .a(net_7392), .o(n7618) );
no02f01 g6323 ( .a(n6867_1), .b(n8845_1), .o(n7626) );
no02f01 g6324 ( .a(n6966), .b(n7188), .o(n7635) );
bf01f01 g6325 ( .a(net_6396), .o(n7644) );
bf01f01 g6326 ( .a(net_7139), .o(n7654) );
bf01f01 g6327 ( .a(net_6467), .o(n7658) );
no02f01 g6328 ( .a(n6867_1), .b(n9980), .o(n7661) );
bf01f01 g6329 ( .a(net_6748), .o(n7700) );
bf01f01 g6330 ( .a(_net_6108), .o(n7704) );
bf01f01 g6331 ( .a(_net_226), .o(n7714) );
bf01f01 g6332 ( .a(net_6837), .o(n7719) );
no02f01 g6333 ( .a(n6867_1), .b(n10215), .o(n7732) );
bf01f01 g6334 ( .a(net_6441), .o(n7756) );
bf01f01 g6335 ( .a(net_7143), .o(n7760) );
bf01f01 g6336 ( .a(net_7160), .o(n7764) );
bf01f01 g6337 ( .a(net_6396), .o(n7776) );
bf01f01 g6338 ( .a(_net_7824), .o(n7779) );
bf01f01 g6339 ( .a(net_6710), .o(n7784) );
bf01f01 g6340 ( .a(_net_7800), .o(n7802) );
bf01f01 g6341 ( .a(_net_7815), .o(n7806) );
bf01f01 g6342 ( .a(_net_7797), .o(n7810) );
bf01f01 g6343 ( .a(net_6734), .o(n7815) );
bf01f01 g6344 ( .a(net_6386), .o(n7818) );
bf01f01 g6345 ( .a(_net_7801), .o(n7826) );
bf01f01 g6346 ( .a(net_6566), .o(n7831) );
bf01f01 g6347 ( .a(_net_6135), .o(n7840) );
bf01f01 g6348 ( .a(net_6382), .o(n7848) );
bf01f01 g6349 ( .a(net_6393), .o(n7867) );
bf01f01 g6350 ( .a(_net_7800), .o(n7871) );
bf01f01 g6351 ( .a(net_6874), .o(n7875) );
no02f01 g6352 ( .a(n6966), .b(n8899_1), .o(n7878) );
bf01f01 g6353 ( .a(_net_6148), .o(n7883) );
bf01f01 g6354 ( .a(net_7249), .o(n7893) );
bf01f01 g6355 ( .a(_net_7822), .o(n7906) );
bf01f01 g6356 ( .a(_net_6167), .o(n7916) );
bf01f01 g6357 ( .a(net_6386), .o(n7920) );
no02f01 g6358 ( .a(n6867_1), .b(n8170_1), .o(n7924) );
bf01f01 g6359 ( .a(net_6568), .o(n7929) );
bf01f01 g6360 ( .a(_net_7798), .o(n7937) );
bf01f01 g6361 ( .a(net_7540), .o(n7942) );
bf01f01 g6362 ( .a(net_6390), .o(n7945) );
bf01f01 g6363 ( .a(net_6724), .o(n7955) );
bf01f01 g6364 ( .a(net_138), .o(n7958) );
bf01f01 g6365 ( .a(_net_7811), .o(n7962) );
bf01f01 g6366 ( .a(net_6992), .o(n7967) );
no02f01 g6367 ( .a(n6867_1), .b(n7601), .o(n7970) );
bf01f01 g6368 ( .a(_net_7821), .o(n7989) );
bf01f01 g6369 ( .a(net_6585), .o(n7994) );
bf01f01 g6370 ( .a(_net_7820), .o(n7997) );
bf01f01 g6371 ( .a(net_6975), .o(n8002) );
bf01f01 g6372 ( .a(net_6394), .o(n8005) );
bf01f01 g6373 ( .a(net_7131), .o(n8015) );
bf01f01 g6374 ( .a(_net_7815), .o(n8028) );
in01f01 g6375 ( .a(n7343), .o(n8042) );
bf01f01 g6376 ( .a(_net_6169), .o(n8047) );
bf01f01 g6377 ( .a(net_6399), .o(n8051) );
bf01f01 g6378 ( .a(net_6988), .o(n8056) );
bf01f01 g6379 ( .a(_net_7819), .o(n8059) );
bf01f01 g6380 ( .a(net_6968), .o(n8064) );
bf01f01 g6381 ( .a(_net_7813), .o(n8067) );
bf01f01 g6382 ( .a(net_6614), .o(n8072) );
bf01f01 g6383 ( .a(_net_7824), .o(n8075) );
bf01f01 g6384 ( .a(net_6596), .o(n8085) );
bf01f01 g6385 ( .a(_net_7808), .o(n8088) );
bf01f01 g6386 ( .a(_net_7801), .o(n8092) );
bf01f01 g6387 ( .a(_net_7801), .o(n8116) );
bf01f01 g6388 ( .a(_net_7795), .o(n8125) );
bf01f01 g6389 ( .a(net_7141), .o(n8140) );
bf01f01 g6390 ( .a(net_6571), .o(n8144) );
bf01f01 g6391 ( .a(_net_7808), .o(n8147) );
no02f01 g6392 ( .a(n6899_1), .b(n8229), .o(n8156) );
bf01f01 g6393 ( .a(net_7715), .o(n8166) );
bf01f01 g6394 ( .a(_net_7820), .o(n8174) );
bf01f01 g6395 ( .a(net_7802), .o(n8183) );
bf01f01 g6396 ( .a(net_6835), .o(n8188) );
bf01f01 g6397 ( .a(_net_7816), .o(n8206) );
bf01f01 g6398 ( .a(net_6389), .o(n8220) );
bf01f01 g6399 ( .a(_net_7810), .o(n8228) );
bf01f01 g6400 ( .a(net_7807), .o(n8232) );
bf01f01 g6401 ( .a(net_6385), .o(n8241) );
bf01f01 g6402 ( .a(net_7799), .o(n8245) );
bf01f01 g6403 ( .a(net_6388), .o(n8249) );
no02f01 g6404 ( .a(n6966), .b(n7142_1), .o(n8262) );
bf01f01 g6405 ( .a(net_7799), .o(n8266) );
bf01f01 g6406 ( .a(_net_6116), .o(n8271) );
bf01f01 g6407 ( .a(net_6615), .o(n8276) );
bf01f01 g6408 ( .a(net_7538), .o(n8280) );
bf01f01 g6409 ( .a(_net_6125), .o(n8289) );
bf01f01 g6410 ( .a(_net_7810), .o(n8303) );
bf01f01 g6411 ( .a(_net_7811), .o(n8307) );
bf01f01 g6412 ( .a(_net_7816), .o(n8311) );
bf01f01 g6413 ( .a(net_6853), .o(n8316) );
bf01f01 g6414 ( .a(net_7138), .o(n8320) );
bf01f01 g6415 ( .a(_net_6100), .o(n8329) );
bf01f01 g6416 ( .a(net_6851), .o(n8334) );
bf01f01 g6417 ( .a(_net_7806), .o(n8337) );
bf01f01 g6418 ( .a(_net_7812), .o(n8340) );
bf01f01 g6419 ( .a(net_7023), .o(n8350) );
bf01f01 g6420 ( .a(net_6427), .o(n8359) );
no02f01 g6421 ( .a(n6966), .b(n7276), .o(n8362) );
bf01f01 g6422 ( .a(net_6425), .o(n8392) );
bf01f01 g6423 ( .a(net_7104), .o(n8401) );
bf01f01 g6424 ( .a(net_7137), .o(n8415) );
bf01f01 g6425 ( .a(net_6392), .o(n8418) );
bf01f01 g6426 ( .a(net_7237), .o(n8422) );
bf01f01 g6427 ( .a(net_6387), .o(n8430) );
bf01f01 g6428 ( .a(net_391), .o(n8438) );
no02f01 g6429 ( .a(n6899_1), .b(n7509_1), .o(n8447) );
no02f01 g6430 ( .a(n6867_1), .b(n7601), .o(n8451) );
bf01f01 g6431 ( .a(_net_7813), .o(n8455) );
bf01f01 g6432 ( .a(_net_7823), .o(n8459) );
bf01f01 g6433 ( .a(net_6742), .o(n8464) );
bf01f01 g6434 ( .a(_net_7804), .o(n8467) );
bf01f01 g6435 ( .a(net_6754), .o(n8477) );
bf01f01 g6436 ( .a(net_7020), .o(n8491) );
bf01f01 g6437 ( .a(_net_7810), .o(n8494) );
bf01f01 g6438 ( .a(net_6622), .o(n8504) );
bf01f01 g6439 ( .a(net_6744), .o(n8513) );
bf01f01 g6440 ( .a(net_6838), .o(n8522) );
bf01f01 g6441 ( .a(_net_7806), .o(n8535) );
bf01f01 g6442 ( .a(_net_7804), .o(n8544) );
bf01f01 g6443 ( .a(net_6707), .o(n8549) );
bf01f01 g6444 ( .a(_net_7795), .o(n8552) );
bf01f01 g6445 ( .a(_net_7824), .o(n8561) );
bf01f01 g6446 ( .a(_net_7797), .o(n8565) );
bf01f01 g6447 ( .a(net_6475), .o(n8575) );
bf01f01 g6448 ( .a(net_6385), .o(n8578) );
bf01f01 g6449 ( .a(net_6695), .o(n8598) );
bf01f01 g6450 ( .a(net_6463), .o(n8612) );
bf01f01 g6451 ( .a(net_6831), .o(n8621) );
bf01f01 g6452 ( .a(_net_7814), .o(n8628) );
bf01f01 g6453 ( .a(_net_7821), .o(n8632) );
bf01f01 g6454 ( .a(net_6013), .o(n8637) );
bf01f01 g6455 ( .a(net_6756), .o(n8641) );
bf01f01 g6456 ( .a(net_6865), .o(n8650) );
bf01f01 g6457 ( .a(net_6577), .o(n8654) );
bf01f01 g6458 ( .a(net_6600), .o(n8658) );
no02f01 g6459 ( .a(n6899_1), .b(n8964), .o(n8666) );
bf01f01 g6460 ( .a(net_6891), .o(n8681) );
bf01f01 g6461 ( .a(net_6722), .o(n8685) );
bf01f01 g6462 ( .a(x1451), .o(n8698) );
no02f01 g6463 ( .a(n6867_1), .b(n8845_1), .o(n8711) );
bf01f01 g6464 ( .a(net_6388), .o(n8715) );
no02f01 g6465 ( .a(n6899_1), .b(n7895), .o(n8734) );
bf01f01 g6466 ( .a(net_7389), .o(n8739) );
bf01f01 g6467 ( .a(net_140), .o(n8757) );
bf01f01 g6468 ( .a(net_7110), .o(n8767) );
bf01f01 g6469 ( .a(x1390), .o(n8784) );
bf01f01 g6470 ( .a(_net_7808), .o(n8788) );
bf01f01 g6471 ( .a(net_6882), .o(n8793) );
bf01f01 g6472 ( .a(net_6457), .o(n8797) );
bf01f01 g6473 ( .a(_net_7808), .o(n8800) );
bf01f01 g6474 ( .a(net_6982), .o(n8805) );
bf01f01 g6475 ( .a(_net_7797), .o(n8813) );
bf01f01 g6476 ( .a(net_7542), .o(n8823) );
bf01f01 g6477 ( .a(_net_7822), .o(n8826) );
bf01f01 g6478 ( .a(_net_7811), .o(n8835) );
bf01f01 g6479 ( .a(x1494), .o(n8864) );
bf01f01 g6480 ( .a(net_151), .o(n8873) );
bf01f01 g6481 ( .a(net_6389), .o(n8877) );
bf01f01 g6482 ( .a(net_6060), .o(n8882) );
bf01f01 g6483 ( .a(_net_7819), .o(n8886) );
bf01f01 g6484 ( .a(net_7132), .o(n8891) );
no02f01 g6485 ( .a(n6899_1), .b(n7507), .o(n8899) );
bf01f01 g6486 ( .a(_net_7822), .o(n8903) );
bf01f01 g6487 ( .a(_net_6119), .o(n8908) );
bf01f01 g6488 ( .a(_net_7804), .o(n8912) );
bf01f01 g6489 ( .a(_net_7809), .o(n8926) );
bf01f01 g6490 ( .a(net_7243), .o(n8931) );
no02f01 g6491 ( .a(n6899_1), .b(n8826_1), .o(n8934) );
bf01f01 g6492 ( .a(net_6458), .o(n8939) );
bf01f01 g6493 ( .a(_net_6086), .o(n8943) );
bf01f01 g6494 ( .a(_net_6130), .o(n8958) );
bf01f01 g6495 ( .a(net_7544), .o(n8963) );
bf01f01 g6496 ( .a(net_7807), .o(n8971) );
bf01f01 g6497 ( .a(_net_6154), .o(n8981) );
bf01f01 g6498 ( .a(net_6386), .o(n8990) );
bf01f01 g6499 ( .a(net_6582), .o(n9010) );
bf01f01 g6500 ( .a(net_7017), .o(n9014) );
bf01f01 g6501 ( .a(net_136), .o(n9017) );
bf01f01 g6502 ( .a(net_6445), .o(n9022) );
bf01f01 g6503 ( .a(_net_7800), .o(n9025) );
bf01f01 g6504 ( .a(net_6864), .o(n9034) );
bf01f01 g6505 ( .a(_net_7805), .o(n9037) );
bf01f01 g6506 ( .a(_net_189), .o(n9047) );
bf01f01 g6507 ( .a(net_6966), .o(n9057) );
no02f01 g6508 ( .a(n6899_1), .b(n7069), .o(n9060) );
bf01f01 g6509 ( .a(net_6984), .o(n9065) );
bf01f01 g6510 ( .a(_net_6110), .o(n9069) );
bf01f01 g6511 ( .a(net_7101), .o(n9079) );
bf01f01 g6512 ( .a(_net_7817), .o(n9082) );
bf01f01 g6513 ( .a(_net_7819), .o(n9086) );
bf01f01 g6514 ( .a(_net_6094), .o(n9091) );
bf01f01 g6515 ( .a(x1511), .o(n9110) );
bf01f01 g6516 ( .a(net_7155), .o(n9120) );
bf01f01 g6517 ( .a(_net_6137), .o(n9134) );
bf01f01 g6518 ( .a(_net_7793), .o(n9138) );
bf01f01 g6519 ( .a(net_6876), .o(n9143) );
bf01f01 g6520 ( .a(_net_7803), .o(n9146) );
bf01f01 g6521 ( .a(net_6393), .o(n9160) );
bf01f01 g6522 ( .a(_net_7811), .o(n9164) );
bf01f01 g6523 ( .a(net_6565), .o(n9169) );
bf01f01 g6524 ( .a(_net_6077), .o(n9178) );
bf01f01 g6525 ( .a(_net_7797), .o(n9182) );
bf01f01 g6526 ( .a(net_6383), .o(n9196) );
no02f01 g6527 ( .a(n6899_1), .b(n7246), .o(n9215) );
bf01f01 g6528 ( .a(net_7156), .o(n9225) );
no02f01 g6529 ( .a(n6867_1), .b(n7978), .o(n9228) );
bf01f01 g6530 ( .a(net_6705), .o(n9238) );
bf01f01 g6531 ( .a(net_6483), .o(n9242) );
bf01f01 g6532 ( .a(_net_7800), .o(n9245) );
bf01f01 g6533 ( .a(net_6701), .o(n9250) );
bf01f01 g6534 ( .a(net_7103), .o(n9254) );
bf01f01 g6535 ( .a(net_7807), .o(n9267) );
bf01f01 g6536 ( .a(net_6848), .o(n9287) );
bf01f01 g6537 ( .a(_net_7820), .o(n9290) );
bf01f01 g6538 ( .a(_net_7816), .o(n9294) );
no02f01 g6539 ( .a(n6966), .b(n10317), .o(n9298) );
no02f01 g6540 ( .a(n6867_1), .b(n7203_1), .o(n9302) );
no02f01 g6541 ( .a(n6899_1), .b(n7514), .o(n9316) );
bf01f01 g6542 ( .a(net_6749), .o(n9326) );
bf01f01 g6543 ( .a(_net_7800), .o(n9339) );
bf01f01 g6544 ( .a(_net_7808), .o(n9343) );
bf01f01 g6545 ( .a(net_7541), .o(n9348) );
bf01f01 g6546 ( .a(_net_7794), .o(n9356) );
bf01f01 g6547 ( .a(net_6464), .o(n9361) );
bf01f01 g6548 ( .a(_net_6089), .o(n9365) );
bf01f01 g6549 ( .a(net_7099), .o(n9370) );
bf01f01 g6550 ( .a(_net_7810), .o(n9373) );
bf01f01 g6551 ( .a(_net_7820), .o(n9377) );
bf01f01 g6552 ( .a(_net_7821), .o(n9381) );
bf01f01 g6553 ( .a(_net_7805), .o(n9385) );
bf01f01 g6554 ( .a(net_6601), .o(n9390) );
bf01f01 g6555 ( .a(_net_7804), .o(n9393) );
bf01f01 g6556 ( .a(_net_6102), .o(n9398) );
bf01f01 g6557 ( .a(x0), .o(n9402) );
bf01f01 g6558 ( .a(_net_7808), .o(n9405) );
bf01f01 g6559 ( .a(net_6459), .o(n9425) );
bf01f01 g6560 ( .a(_net_7808), .o(n9428) );
bf01f01 g6561 ( .a(_net_7810), .o(n9431) );
bf01f01 g6562 ( .a(net_6731), .o(n9445) );
bf01f01 g6563 ( .a(net_7709), .o(n9459) );
bf01f01 g6564 ( .a(_net_7816), .o(n9462) );
bf01f01 g6565 ( .a(net_6972), .o(n9467) );
bf01f01 g6566 ( .a(net_6394), .o(n9470) );
bf01f01 g6567 ( .a(net_6842), .o(n9475) );
no02f01 g6568 ( .a(n6867_1), .b(n9870), .o(n9478) );
bf01f01 g6569 ( .a(net_6611), .o(n9483) );
bf01f01 g6570 ( .a(_net_6163), .o(n9502) );
bf01f01 g6571 ( .a(net_6871), .o(n9517) );
bf01f01 g6572 ( .a(net_6391), .o(n9520) );
bf01f01 g6573 ( .a(net_7015), .o(n9525) );
bf01f01 g6574 ( .a(_net_7805), .o(n9528) );
bf01f01 g6575 ( .a(_net_7817), .o(n9537) );
bf01f01 g6576 ( .a(_net_7813), .o(n9541) );
no02f01 g6577 ( .a(n6867_1), .b(n7175), .o(n9549) );
bf01f01 g6578 ( .a(net_6840), .o(n9579) );
bf01f01 g6579 ( .a(net_6455), .o(n9588) );
bf01f01 g6580 ( .a(_net_7821), .o(n9606) );
bf01f01 g6581 ( .a(_net_6111), .o(n9611) );
bf01f01 g6582 ( .a(_net_7820), .o(n9620) );
bf01f01 g6583 ( .a(_net_7803), .o(n9624) );
bf01f01 g6584 ( .a(net_153), .o(n9628) );
bf01f01 g6585 ( .a(_net_7814), .o(n9642) );
bf01f01 g6586 ( .a(net_7386), .o(n9647) );
bf01f01 g6587 ( .a(net_7548), .o(n9651) );
bf01f01 g6588 ( .a(net_7005), .o(n9660) );
bf01f01 g6589 ( .a(net_6383), .o(n9668) );
bf01f01 g6590 ( .a(net_6392), .o(n9687) );
bf01f01 g6591 ( .a(net_6703), .o(n9692) );
bf01f01 g6592 ( .a(net_6381), .o(n9695) );
bf01f01 g6593 ( .a(_net_7804), .o(n9704) );
bf01f01 g6594 ( .a(_net_6162), .o(n9724) );
bf01f01 g6595 ( .a(net_6472), .o(n9729) );
bf01f01 g6596 ( .a(x1398), .o(n9737) );
bf01f01 g6597 ( .a(_net_7812), .o(n9746) );
bf01f01 g6598 ( .a(_net_7795), .o(n9750) );
no02f01 g6599 ( .a(n6867_1), .b(n8173), .o(n9754) );
no02f01 g6600 ( .a(n6966), .b(n7276), .o(n9758) );
bf01f01 g6601 ( .a(net_7027), .o(n9783) );
bf01f01 g6602 ( .a(_net_7810), .o(n9796) );
bf01f01 g6603 ( .a(net_6399), .o(n9805) );
bf01f01 g6604 ( .a(net_6388), .o(n9809) );
no02f01 g6605 ( .a(n6966), .b(n7520), .o(n9828) );
bf01f01 g6606 ( .a(net_7135), .o(n9833) );
bf01f01 g6607 ( .a(net_7122), .o(n9837) );
bf01f01 g6608 ( .a(net_6396), .o(n9840) );
bf01f01 g6609 ( .a(net_6387), .o(n9844) );
no02f01 g6610 ( .a(n6966), .b(n10317), .o(n9853) );
bf01f01 g6611 ( .a(_net_7811), .o(n9867) );
bf01f01 g6612 ( .a(_net_7797), .o(n9871) );
bf01f01 g6613 ( .a(_net_7806), .o(n9875) );
bf01f01 g6614 ( .a(net_7109), .o(n9885) );
bf01f01 g6615 ( .a(net_6752), .o(n9899) );
bf01f01 g6616 ( .a(_net_7798), .o(n9902) );
bf01f01 g6617 ( .a(net_6446), .o(n9911) );
bf01f01 g6618 ( .a(_net_7819), .o(n9914) );
bf01f01 g6619 ( .a(x1580), .o(n9918) );
bf01f01 g6620 ( .a(net_6719), .o(n9923) );
bf01f01 g6621 ( .a(net_6389), .o(n9926) );
bf01f01 g6622 ( .a(net_6393), .o(n9930) );
bf01f01 g6623 ( .a(net_6465), .o(n9935) );
bf01f01 g6624 ( .a(_net_6174), .o(n9944) );
in01f01 g6625 ( .a(n7343), .o(n9953) );
bf01f01 g6626 ( .a(net_6389), .o(n9957) );
bf01f01 g6627 ( .a(_net_7804), .o(n9961) );
bf01f01 g6628 ( .a(net_6057), .o(n9976) );
bf01f01 g6629 ( .a(net_6380), .o(n9985) );
bf01f01 g6630 ( .a(_net_7805), .o(n9988) );
bf01f01 g6631 ( .a(_net_7805), .o(n9992) );
bf01f01 g6632 ( .a(_net_7812), .o(n10001) );
bf01f01 g6633 ( .a(_net_6062), .o(n10006) );
bf01f01 g6634 ( .a(net_7802), .o(n10010) );
bf01f01 g6635 ( .a(x1351), .o(n10014) );
bf01f01 g6636 ( .a(net_130), .o(n10023) );
bf01f01 g6637 ( .a(net_6879), .o(n10028) );
bf01f01 g6638 ( .a(_net_6155), .o(n10047) );
no02f01 g6639 ( .a(n6966), .b(n7250), .o(n10056) );
bf01f01 g6640 ( .a(net_6884), .o(n10070) );
bf01f01 g6641 ( .a(_net_7815), .o(n10103) );
bf01f01 g6642 ( .a(_net_7818), .o(n10107) );
bf01f01 g6643 ( .a(net_7112), .o(n10112) );
bf01f01 g6644 ( .a(_net_7815), .o(n10120) );
bf01f01 g6645 ( .a(_net_7811), .o(n10124) );
bf01f01 g6646 ( .a(_net_7805), .o(n10132) );
bf01f01 g6647 ( .a(x1595), .o(n10141) );
no02f01 g6648 ( .a(n6899_1), .b(n7514), .o(n10145) );
bf01f01 g6649 ( .a(net_7807), .o(n10154) );
bf01f01 g6650 ( .a(_net_7806), .o(n10158) );
ms00f80 l0001 ( .d(n266), .o(net_249), .ck(clk) );
ms00f80 l0002 ( .d(n271), .o(net_254), .ck(clk) );
ms00f80 l0003 ( .d(n276), .o(net_6907), .ck(clk) );
ms00f80 l0004 ( .d(n281), .o(_net_6082), .ck(clk) );
ms00f80 l0005 ( .d(n286), .o(net_6300), .ck(clk) );
ms00f80 l0006 ( .d(n291), .o(net_6453), .ck(clk) );
ms00f80 l0007 ( .d(n295), .o(_net_6032), .ck(clk) );
ms00f80 l0008 ( .d(n300), .o(_net_6133), .ck(clk) );
ms00f80 l0009 ( .d(n305), .o(net_7222), .ck(clk) );
ms00f80 l0010 ( .d(n310), .o(net_6704), .ck(clk) );
ms00f80 l0011 ( .d(n314), .o(_net_7481), .ck(clk) );
ms00f80 l0012 ( .d(n319), .o(_net_175), .ck(clk) );
ms00f80 l0013 ( .d(n324), .o(net_7204), .ck(clk) );
ms00f80 l0014 ( .d(n329), .o(_net_6062), .ck(clk) );
ms00f80 l0015 ( .d(n334), .o(net_6227), .ck(clk) );
ms00f80 l0016 ( .d(n339), .o(net_6364), .ck(clk) );
ms00f80 l0017 ( .d(n344), .o(net_6256), .ck(clk) );
ms00f80 l0018 ( .d(n349), .o(net_6474), .ck(clk) );
ms00f80 l0019 ( .d(n352), .o(_net_7800), .ck(clk) );
ms00f80 l0020 ( .d(n357), .o(net_7114), .ck(clk) );
ms00f80 l0021 ( .d(n361), .o(net_6784), .ck(clk) );
ms00f80 l0022 ( .d(n366), .o(net_6996), .ck(clk) );
ms00f80 l0023 ( .d(n370), .o(_net_7474), .ck(clk) );
ms00f80 l0024 ( .d(n375), .o(_net_7252), .ck(clk) );
ms00f80 l0025 ( .d(n380), .o(_net_298), .ck(clk) );
ms00f80 l0026 ( .d(n385), .o(_net_6404), .ck(clk) );
ms00f80 l0027 ( .d(n390), .o(_net_6088), .ck(clk) );
ms00f80 l0028 ( .d(n395), .o(net_7055), .ck(clk) );
ms00f80 l0029 ( .d(n400), .o(_net_7595), .ck(clk) );
ms00f80 l0030 ( .d(n405), .o(net_6396), .ck(clk) );
ms00f80 l0031 ( .d(n410), .o(net_6313), .ck(clk) );
ms00f80 l0032 ( .d(n415), .o(net_7062), .ck(clk) );
ms00f80 l0033 ( .d(n420), .o(net_7525), .ck(clk) );
ms00f80 l0034 ( .d(n424), .o(net_6514), .ck(clk) );
ms00f80 l0035 ( .d(n429), .o(net_6803), .ck(clk) );
ms00f80 l0036 ( .d(n434), .o(net_7713), .ck(clk) );
ms00f80 l0037 ( .d(n438), .o(net_6510), .ck(clk) );
ms00f80 l0038 ( .d(n443), .o(net_7000), .ck(clk) );
ms00f80 l0039 ( .d(n447), .o(_net_6150), .ck(clk) );
ms00f80 l0040 ( .d(n451), .o(net_7802), .ck(clk) );
ms00f80 l0041 ( .d(n455), .o(net_6628), .ck(clk) );
ms00f80 l0042 ( .d(n460), .o(_net_7355), .ck(clk) );
ms00f80 l0043 ( .d(n465), .o(_net_6100), .ck(clk) );
ms00f80 l0044 ( .d(n470), .o(net_7388), .ck(clk) );
ms00f80 l0045 ( .d(n474), .o(net_362), .ck(clk) );
ms00f80 l0046 ( .d(n479), .o(net_6783), .ck(clk) );
ms00f80 l0047 ( .d(n484), .o(net_6870), .ck(clk) );
ms00f80 l0048 ( .d(n488), .o(net_7196), .ck(clk) );
ms00f80 l0049 ( .d(n493), .o(net_7224), .ck(clk) );
ms00f80 l0050 ( .d(n498), .o(_net_6194), .ck(clk) );
ms00f80 l0051 ( .d(n503), .o(net_6267), .ck(clk) );
ms00f80 l0052 ( .d(n508), .o(net_6308), .ck(clk) );
ms00f80 l0053 ( .d(n513), .o(net_6691), .ck(clk) );
ms00f80 l0054 ( .d(n518), .o(net_7369), .ck(clk) );
ms00f80 l0055 ( .d(n523), .o(_net_6079), .ck(clk) );
ms00f80 l0056 ( .d(n528), .o(_net_7689), .ck(clk) );
ms00f80 l0057 ( .d(n533), .o(_net_6104), .ck(clk) );
ms00f80 l0058 ( .d(n538), .o(_net_7603), .ck(clk) );
ms00f80 l0059 ( .d(n543), .o(_net_7316), .ck(clk) );
ms00f80 l0060 ( .d(n548), .o(_net_5965), .ck(clk) );
ms00f80 l0061 ( .d(n553), .o(x14), .ck(clk) );
ms00f80 l0062 ( .d(n556), .o(net_6791), .ck(clk) );
ms00f80 l0063 ( .d(n561), .o(_net_6294), .ck(clk) );
ms00f80 l0064 ( .d(n566), .o(net_6773), .ck(clk) );
ms00f80 l0065 ( .d(n571), .o(net_6218), .ck(clk) );
ms00f80 l0066 ( .d(n576), .o(net_7342), .ck(clk) );
ms00f80 l0067 ( .d(n580), .o(_net_7794), .ck(clk) );
ms00f80 l0068 ( .d(n585), .o(net_6373), .ck(clk) );
ms00f80 l0069 ( .d(n590), .o(net_365), .ck(clk) );
ms00f80 l0070 ( .d(n595), .o(net_7492), .ck(clk) );
ms00f80 l0071 ( .d(n600), .o(_net_7285), .ck(clk) );
ms00f80 l0072 ( .d(n605), .o(_net_6210), .ck(clk) );
ms00f80 l0073 ( .d(n610), .o(net_6900), .ck(clk) );
ms00f80 l0074 ( .d(n615), .o(net_7604), .ck(clk) );
ms00f80 l0075 ( .d(n620), .o(_net_6004), .ck(clk) );
ms00f80 l0076 ( .d(n625), .o(net_7246), .ck(clk) );
ms00f80 l0077 ( .d(n629), .o(_net_7441), .ck(clk) );
ms00f80 l0078 ( .d(n634), .o(net_7487), .ck(clk) );
ms00f80 l0079 ( .d(n639), .o(_net_7694), .ck(clk) );
ms00f80 l0080 ( .d(n644), .o(_net_7094), .ck(clk) );
ms00f80 l0081 ( .d(n649), .o(_net_212), .ck(clk) );
ms00f80 l0082 ( .d(n654), .o(_net_7753), .ck(clk) );
ms00f80 l0083 ( .d(n659), .o(net_160), .ck(clk) );
ms00f80 l0084 ( .d(n664), .o(net_6384), .ck(clk) );
ms00f80 l0085 ( .d(n669), .o(net_6440), .ck(clk) );
ms00f80 l0086 ( .d(n673), .o(_net_6208), .ck(clk) );
ms00f80 l0087 ( .d(n678), .o(net_6653), .ck(clk) );
ms00f80 l0088 ( .d(n683), .o(net_6491), .ck(clk) );
ms00f80 l0089 ( .d(n688), .o(_net_7330), .ck(clk) );
ms00f80 l0090 ( .d(n693), .o(_net_7271), .ck(clk) );
ms00f80 l0091 ( .d(n698), .o(net_7645), .ck(clk) );
ms00f80 l0092 ( .d(n703), .o(net_6323), .ck(clk) );
ms00f80 l0093 ( .d(n708), .o(_net_7300), .ck(clk) );
ms00f80 l0094 ( .d(n713), .o(net_7774), .ck(clk) );
ms00f80 l0095 ( .d(n718), .o(net_7637), .ck(clk) );
ms00f80 l0096 ( .d(n722), .o(net_361), .ck(clk) );
ms00f80 l0097 ( .d(n727), .o(net_236), .ck(clk) );
ms00f80 l0098 ( .d(n732), .o(x561), .ck(clk) );
ms00f80 l0099 ( .d(n736), .o(_net_6037), .ck(clk) );
ms00f80 l0100 ( .d(n741), .o(net_6213), .ck(clk) );
ms00f80 l0101 ( .d(n746), .o(net_235), .ck(clk) );
ms00f80 l0102 ( .d(n751), .o(net_7758), .ck(clk) );
ms00f80 l0103 ( .d(n756), .o(_net_6147), .ck(clk) );
ms00f80 l0104 ( .d(n761), .o(net_6468), .ck(clk) );
ms00f80 l0105 ( .d(n765), .o(_net_113), .ck(clk) );
ms00f80 l0106 ( .d(n770), .o(_net_7732), .ck(clk) );
ms00f80 l0107 ( .d(n774), .o(net_6380), .ck(clk) );
ms00f80 l0108 ( .d(n779), .o(net_6386), .ck(clk) );
ms00f80 l0109 ( .d(n783), .o(net_139), .ck(clk) );
ms00f80 l0110 ( .d(n788), .o(_net_6012), .ck(clk) );
ms00f80 l0111 ( .d(n793), .o(net_7607), .ck(clk) );
ms00f80 l0112 ( .d(n798), .o(net_7134), .ck(clk) );
ms00f80 l0113 ( .d(n802), .o(net_7133), .ck(clk) );
ms00f80 l0114 ( .d(n806), .o(_net_7786), .ck(clk) );
ms00f80 l0115 ( .d(n811), .o(net_6400), .ck(clk) );
ms00f80 l0116 ( .d(n815), .o(net_6260), .ck(clk) );
ms00f80 l0117 ( .d(n820), .o(_net_121), .ck(clk) );
ms00f80 l0118 ( .d(n825), .o(_net_120), .ck(clk) );
ms00f80 l0119 ( .d(n830), .o(net_7396), .ck(clk) );
ms00f80 l0120 ( .d(n834), .o(net_220), .ck(clk) );
ms00f80 l0121 ( .d(n839), .o(net_6545), .ck(clk) );
ms00f80 l0122 ( .d(n844), .o(net_326), .ck(clk) );
ms00f80 l0123 ( .d(n849), .o(net_171), .ck(clk) );
ms00f80 l0124 ( .d(n854), .o(net_7390), .ck(clk) );
ms00f80 l0125 ( .d(n857), .o(net_6521), .ck(clk) );
ms00f80 l0126 ( .d(n862), .o(_net_6086), .ck(clk) );
ms00f80 l0127 ( .d(n867), .o(net_6711), .ck(clk) );
ms00f80 l0128 ( .d(n870), .o(net_6815), .ck(clk) );
ms00f80 l0129 ( .d(n875), .o(net_7312), .ck(clk) );
ms00f80 l0130 ( .d(n880), .o(net_6646), .ck(clk) );
ms00f80 l0131 ( .d(n885), .o(_net_6008), .ck(clk) );
ms00f80 l0132 ( .d(n890), .o(net_6616), .ck(clk) );
ms00f80 l0133 ( .d(n894), .o(net_347), .ck(clk) );
ms00f80 l0134 ( .d(n899), .o(net_6739), .ck(clk) );
ms00f80 l0135 ( .d(n903), .o(_net_7439), .ck(clk) );
ms00f80 l0136 ( .d(n907), .o(net_7067), .ck(clk) );
ms00f80 l0137 ( .d(n911), .o(net_7073), .ck(clk) );
ms00f80 l0138 ( .d(n916), .o(net_6746), .ck(clk) );
ms00f80 l0139 ( .d(n920), .o(net_6356), .ck(clk) );
ms00f80 l0140 ( .d(n925), .o(_net_7354), .ck(clk) );
ms00f80 l0141 ( .d(n930), .o(_net_7632), .ck(clk) );
ms00f80 l0142 ( .d(n935), .o(net_7066), .ck(clk) );
ms00f80 l0143 ( .d(n940), .o(net_6979), .ck(clk) );
ms00f80 l0144 ( .d(n944), .o(_net_5851), .ck(clk) );
ms00f80 l0145 ( .d(n948), .o(_net_7809), .ck(clk) );
ms00f80 l0146 ( .d(n953), .o(net_6989), .ck(clk) );
ms00f80 l0147 ( .d(n956), .o(net_7058), .ck(clk) );
ms00f80 l0148 ( .d(n961), .o(_net_7629), .ck(clk) );
ms00f80 l0149 ( .d(n966), .o(net_204), .ck(clk) );
ms00f80 l0150 ( .d(n971), .o(_net_7296), .ck(clk) );
ms00f80 l0151 ( .d(n976), .o(net_150), .ck(clk) );
ms00f80 l0152 ( .d(n981), .o(net_6999), .ck(clk) );
ms00f80 l0153 ( .d(n985), .o(_net_282), .ck(clk) );
ms00f80 l0154 ( .d(n990), .o(_net_7653), .ck(clk) );
ms00f80 l0155 ( .d(n995), .o(_net_5856), .ck(clk) );
ms00f80 l0156 ( .d(n1000), .o(net_391), .ck(clk) );
ms00f80 l0157 ( .d(n1005), .o(net_6392), .ck(clk) );
ms00f80 l0158 ( .d(n1010), .o(_net_7621), .ck(clk) );
ms00f80 l0159 ( .d(n1015), .o(_net_6120), .ck(clk) );
ms00f80 l0160 ( .d(n1020), .o(net_6998), .ck(clk) );
ms00f80 l0161 ( .d(n1024), .o(_net_7447), .ck(clk) );
ms00f80 l0162 ( .d(n1029), .o(net_7334), .ck(clk) );
ms00f80 l0163 ( .d(n1034), .o(net_7311), .ck(clk) );
ms00f80 l0164 ( .d(n1039), .o(_net_6220), .ck(clk) );
ms00f80 l0165 ( .d(n1044), .o(_net_7281), .ck(clk) );
ms00f80 l0166 ( .d(n1049), .o(_net_7578), .ck(clk) );
ms00f80 l0167 ( .d(n1053), .o(net_351), .ck(clk) );
ms00f80 l0168 ( .d(n1058), .o(x657), .ck(clk) );
ms00f80 l0169 ( .d(n1062), .o(net_6944), .ck(clk) );
ms00f80 l0170 ( .d(n1067), .o(net_5992), .ck(clk) );
ms00f80 l0171 ( .d(n1072), .o(_net_6286), .ck(clk) );
ms00f80 l0172 ( .d(n1077), .o(net_7004), .ck(clk) );
ms00f80 l0173 ( .d(n1081), .o(net_7010), .ck(clk) );
ms00f80 l0174 ( .d(n1085), .o(net_6461), .ck(clk) );
ms00f80 l0175 ( .d(n1089), .o(net_6832), .ck(clk) );
ms00f80 l0176 ( .d(n1093), .o(net_6977), .ck(clk) );
ms00f80 l0177 ( .d(n1097), .o(net_6901), .ck(clk) );
ms00f80 l0178 ( .d(n1102), .o(net_6856), .ck(clk) );
ms00f80 l0179 ( .d(n1106), .o(_net_7412), .ck(clk) );
ms00f80 l0180 ( .d(n1111), .o(net_6379), .ck(clk) );
ms00f80 l0181 ( .d(n1116), .o(net_6060), .ck(clk) );
ms00f80 l0182 ( .d(n1121), .o(net_6847), .ck(clk) );
ms00f80 l0183 ( .d(n1125), .o(_net_7274), .ck(clk) );
ms00f80 l0184 ( .d(n1130), .o(net_6671), .ck(clk) );
ms00f80 l0185 ( .d(n1135), .o(_net_7299), .ck(clk) );
ms00f80 l0186 ( .d(n1140), .o(net_6986), .ck(clk) );
ms00f80 l0187 ( .d(n1144), .o(net_6275), .ck(clk) );
ms00f80 l0188 ( .d(n1148), .o(net_6677), .ck(clk) );
ms00f80 l0189 ( .d(n1153), .o(_net_6167), .ck(clk) );
ms00f80 l0190 ( .d(n1158), .o(net_6242), .ck(clk) );
ms00f80 l0191 ( .d(n1163), .o(net_7611), .ck(clk) );
ms00f80 l0192 ( .d(n1168), .o(net_363), .ck(clk) );
ms00f80 l0193 ( .d(n1173), .o(net_7523), .ck(clk) );
ms00f80 l0194 ( .d(n1178), .o(_net_6135), .ck(clk) );
ms00f80 l0195 ( .d(n1183), .o(net_6238), .ck(clk) );
ms00f80 l0196 ( .d(n1187), .o(net_345), .ck(clk) );
ms00f80 l0197 ( .d(n1191), .o(net_6788), .ck(clk) );
ms00f80 l0198 ( .d(n1195), .o(net_6922), .ck(clk) );
ms00f80 l0199 ( .d(n1200), .o(net_6240), .ck(clk) );
ms00f80 l0200 ( .d(n1205), .o(net_7081), .ck(clk) );
ms00f80 l0201 ( .d(n1210), .o(net_6845), .ck(clk) );
ms00f80 l0202 ( .d(n1214), .o(_net_7503), .ck(clk) );
ms00f80 l0203 ( .d(n1219), .o(_net_7428), .ck(clk) );
ms00f80 l0204 ( .d(n1224), .o(net_6608), .ck(clk) );
ms00f80 l0205 ( .d(n1228), .o(_net_7730), .ck(clk) );
ms00f80 l0206 ( .d(n1232), .o(net_132), .ck(clk) );
ms00f80 l0207 ( .d(n1236), .o(net_7675), .ck(clk) );
ms00f80 l0208 ( .d(n1240), .o(net_6952), .ck(clk) );
ms00f80 l0209 ( .d(n1244), .o(net_360), .ck(clk) );
ms00f80 l0210 ( .d(n1248), .o(net_6759), .ck(clk) );
ms00f80 l0211 ( .d(n1253), .o(_net_7512), .ck(clk) );
ms00f80 l0212 ( .d(n1258), .o(net_7019), .ck(clk) );
ms00f80 l0213 ( .d(n1262), .o(net_6354), .ck(clk) );
ms00f80 l0214 ( .d(n1267), .o(_net_7590), .ck(clk) );
ms00f80 l0215 ( .d(n1272), .o(_net_273), .ck(clk) );
ms00f80 l0216 ( .d(n1277), .o(net_7453), .ck(clk) );
ms00f80 l0217 ( .d(n1282), .o(_net_299), .ck(clk) );
ms00f80 l0218 ( .d(n1287), .o(net_7119), .ck(clk) );
ms00f80 l0219 ( .d(n1291), .o(net_6574), .ck(clk) );
ms00f80 l0220 ( .d(n1295), .o(_net_7315), .ck(clk) );
ms00f80 l0221 ( .d(n1300), .o(net_7070), .ck(clk) );
ms00f80 l0222 ( .d(n1305), .o(net_7395), .ck(clk) );
ms00f80 l0223 ( .d(n1309), .o(_net_5966), .ck(clk) );
ms00f80 l0224 ( .d(n1314), .o(_net_6000), .ck(clk) );
ms00f80 l0225 ( .d(n1318), .o(net_7182), .ck(clk) );
ms00f80 l0226 ( .d(n1322), .o(net_7200), .ck(clk) );
ms00f80 l0227 ( .d(n1326), .o(net_6515), .ck(clk) );
ms00f80 l0228 ( .d(n1331), .o(net_6859), .ck(clk) );
ms00f80 l0229 ( .d(n1335), .o(_net_5991), .ck(clk) );
ms00f80 l0230 ( .d(n1340), .o(_net_7707), .ck(clk) );
ms00f80 l0231 ( .d(n1345), .o(net_6961), .ck(clk) );
ms00f80 l0232 ( .d(n1350), .o(net_7303), .ck(clk) );
ms00f80 l0233 ( .d(n1355), .o(net_6877), .ck(clk) );
ms00f80 l0234 ( .d(n1359), .o(net_7234), .ck(clk) );
ms00f80 l0235 ( .d(n1363), .o(_net_213), .ck(clk) );
ms00f80 l0236 ( .d(n1368), .o(net_6025), .ck(clk) );
ms00f80 l0237 ( .d(n1373), .o(_net_5997), .ck(clk) );
ms00f80 l0238 ( .d(n1378), .o(net_7750), .ck(clk) );
ms00f80 l0239 ( .d(n1383), .o(net_6694), .ck(clk) );
ms00f80 l0240 ( .d(n1386), .o(net_325), .ck(clk) );
ms00f80 l0241 ( .d(n1391), .o(_net_7658), .ck(clk) );
ms00f80 l0242 ( .d(n1396), .o(net_6190), .ck(clk) );
ms00f80 l0243 ( .d(n1400), .o(net_6624), .ck(clk) );
ms00f80 l0244 ( .d(n1405), .o(_net_6182), .ck(clk) );
ms00f80 l0245 ( .d(n1410), .o(_net_5960), .ck(clk) );
ms00f80 l0246 ( .d(n1414), .o(net_7217), .ck(clk) );
ms00f80 l0247 ( .d(n1419), .o(_net_7253), .ck(clk) );
ms00f80 l0248 ( .d(n1423), .o(net_6941), .ck(clk) );
ms00f80 l0249 ( .d(n1428), .o(_net_7497), .ck(clk) );
ms00f80 l0250 ( .d(n1433), .o(_net_7768), .ck(clk) );
ms00f80 l0251 ( .d(n1438), .o(net_6745), .ck(clk) );
ms00f80 l0252 ( .d(n1442), .o(_net_7565), .ck(clk) );
ms00f80 l0253 ( .d(n1446), .o(net_6913), .ck(clk) );
ms00f80 l0254 ( .d(n1451), .o(_net_6044), .ck(clk) );
ms00f80 l0255 ( .d(n1455), .o(net_6633), .ck(clk) );
ms00f80 l0256 ( .d(n1460), .o(net_6328), .ck(clk) );
ms00f80 l0257 ( .d(n1465), .o(net_6953), .ck(clk) );
ms00f80 l0258 ( .d(n1469), .o(net_357), .ck(clk) );
ms00f80 l0259 ( .d(n1474), .o(net_6612), .ck(clk) );
ms00f80 l0260 ( .d(n1478), .o(net_6302), .ck(clk) );
ms00f80 l0261 ( .d(n1482), .o(_net_7815), .ck(clk) );
ms00f80 l0262 ( .d(n1487), .o(_net_7746), .ck(clk) );
ms00f80 l0263 ( .d(n1491), .o(net_6768), .ck(clk) );
ms00f80 l0264 ( .d(n1496), .o(net_6059), .ck(clk) );
ms00f80 l0265 ( .d(n1501), .o(_net_7698), .ck(clk) );
ms00f80 l0266 ( .d(n1506), .o(net_7550), .ck(clk) );
ms00f80 l0267 ( .d(n1510), .o(net_7091), .ck(clk) );
ms00f80 l0268 ( .d(n1515), .o(net_6619), .ck(clk) );
ms00f80 l0269 ( .d(n1519), .o(_net_6095), .ck(clk) );
ms00f80 l0270 ( .d(n1524), .o(net_7106), .ck(clk) );
ms00f80 l0271 ( .d(n1528), .o(net_6375), .ck(clk) );
ms00f80 l0272 ( .d(n1533), .o(net_203), .ck(clk) );
ms00f80 l0273 ( .d(n1538), .o(net_7247), .ck(clk) );
ms00f80 l0274 ( .d(n1542), .o(x287), .ck(clk) );
ms00f80 l0275 ( .d(n1546), .o(_net_7534), .ck(clk) );
ms00f80 l0276 ( .d(n1551), .o(net_7146), .ck(clk) );
ms00f80 l0277 ( .d(n1555), .o(_net_7406), .ck(clk) );
ms00f80 l0278 ( .d(n1560), .o(net_7126), .ck(clk) );
ms00f80 l0279 ( .d(n1564), .o(net_6482), .ck(clk) );
ms00f80 l0280 ( .d(n1568), .o(net_6888), .ck(clk) );
ms00f80 l0281 ( .d(n1572), .o(net_258), .ck(clk) );
ms00f80 l0282 ( .d(n1577), .o(net_353), .ck(clk) );
ms00f80 l0283 ( .d(n1582), .o(_net_7535), .ck(clk) );
ms00f80 l0284 ( .d(n1587), .o(net_6584), .ck(clk) );
ms00f80 l0285 ( .d(n1591), .o(net_352), .ck(clk) );
ms00f80 l0286 ( .d(n1596), .o(net_6732), .ck(clk) );
ms00f80 l0287 ( .d(n1600), .o(_net_7759), .ck(clk) );
ms00f80 l0288 ( .d(n1605), .o(net_165), .ck(clk) );
ms00f80 l0289 ( .d(n1610), .o(_net_7498), .ck(clk) );
ms00f80 l0290 ( .d(n1615), .o(net_6914), .ck(clk) );
ms00f80 l0291 ( .d(n1619), .o(net_7198), .ck(clk) );
ms00f80 l0292 ( .d(n1624), .o(_net_7696), .ck(clk) );
ms00f80 l0293 ( .d(n1629), .o(net_6537), .ck(clk) );
ms00f80 l0294 ( .d(n1634), .o(_net_7570), .ck(clk) );
ms00f80 l0295 ( .d(n1639), .o(net_7308), .ck(clk) );
ms00f80 l0296 ( .d(n1644), .o(net_260), .ck(clk) );
ms00f80 l0297 ( .d(n1649), .o(net_7124), .ck(clk) );
ms00f80 l0298 ( .d(n1653), .o(net_6229), .ck(clk) );
ms00f80 l0299 ( .d(n1658), .o(net_245), .ck(clk) );
ms00f80 l0300 ( .d(n1663), .o(net_6197), .ck(clk) );
ms00f80 l0301 ( .d(n1668), .o(net_7760), .ck(clk) );
ms00f80 l0302 ( .d(n1673), .o(net_6723), .ck(clk) );
ms00f80 l0303 ( .d(n1677), .o(_net_6042), .ck(clk) );
ms00f80 l0304 ( .d(n1681), .o(net_6654), .ck(clk) );
ms00f80 l0305 ( .d(n1686), .o(net_6512), .ck(clk) );
ms00f80 l0306 ( .d(n1691), .o(net_6770), .ck(clk) );
ms00f80 l0307 ( .d(n1696), .o(_net_6168), .ck(clk) );
ms00f80 l0308 ( .d(n1701), .o(net_6432), .ck(clk) );
ms00f80 l0309 ( .d(n1704), .o(net_6500), .ck(clk) );
ms00f80 l0310 ( .d(n1709), .o(net_7170), .ck(clk) );
ms00f80 l0311 ( .d(n1714), .o(_net_7358), .ck(clk) );
ms00f80 l0312 ( .d(n1718), .o(net_6903), .ck(clk) );
ms00f80 l0313 ( .d(n1722), .o(net_7220), .ck(clk) );
ms00f80 l0314 ( .d(n1727), .o(_net_6180), .ck(clk) );
ms00f80 l0315 ( .d(n1732), .o(net_6806), .ck(clk) );
ms00f80 l0316 ( .d(n1737), .o(_net_7468), .ck(clk) );
ms00f80 l0317 ( .d(n1742), .o(_net_5996), .ck(clk) );
ms00f80 l0318 ( .d(n1747), .o(_net_6077), .ck(clk) );
ms00f80 l0319 ( .d(n1752), .o(net_7495), .ck(clk) );
ms00f80 l0320 ( .d(n1756), .o(net_6896), .ck(clk) );
ms00f80 l0321 ( .d(n1761), .o(net_6570), .ck(clk) );
ms00f80 l0322 ( .d(n1765), .o(net_7223), .ck(clk) );
ms00f80 l0323 ( .d(n1770), .o(_net_5985), .ck(clk) );
ms00f80 l0324 ( .d(n1775), .o(net_6602), .ck(clk) );
ms00f80 l0325 ( .d(n1779), .o(net_7551), .ck(clk) );
ms00f80 l0326 ( .d(n1782), .o(net_7035), .ck(clk) );
ms00f80 l0327 ( .d(n1787), .o(_net_6296), .ck(clk) );
ms00f80 l0328 ( .d(n1792), .o(net_7742), .ck(clk) );
ms00f80 l0329 ( .d(n1797), .o(net_6316), .ck(clk) );
ms00f80 l0330 ( .d(n1802), .o(_net_6185), .ck(clk) );
ms00f80 l0331 ( .d(n1807), .o(_net_7328), .ck(clk) );
ms00f80 l0332 ( .d(n1812), .o(_net_7359), .ck(clk) );
ms00f80 l0333 ( .d(n1817), .o(net_6371), .ck(clk) );
ms00f80 l0334 ( .d(n1822), .o(net_6269), .ck(clk) );
ms00f80 l0335 ( .d(n1827), .o(net_6248), .ck(clk) );
ms00f80 l0336 ( .d(n1832), .o(_net_7650), .ck(clk) );
ms00f80 l0337 ( .d(n1836), .o(_net_7813), .ck(clk) );
ms00f80 l0338 ( .d(n1841), .o(_net_6087), .ck(clk) );
ms00f80 l0339 ( .d(n1846), .o(_net_6292), .ck(clk) );
ms00f80 l0340 ( .d(n1851), .o(net_6223), .ck(clk) );
ms00f80 l0341 ( .d(n1855), .o(_net_7819), .ck(clk) );
ms00f80 l0342 ( .d(n1860), .o(net_7767), .ck(clk) );
ms00f80 l0343 ( .d(n1865), .o(net_6699), .ck(clk) );
ms00f80 l0344 ( .d(n1869), .o(_net_7255), .ck(clk) );
ms00f80 l0345 ( .d(n1874), .o(net_6599), .ck(clk) );
ms00f80 l0346 ( .d(n1878), .o(_net_7600), .ck(clk) );
ms00f80 l0347 ( .d(n1883), .o(_net_6067), .ck(clk) );
ms00f80 l0348 ( .d(n1888), .o(_net_7628), .ck(clk) );
ms00f80 l0349 ( .d(n1893), .o(_net_6155), .ck(clk) );
ms00f80 l0350 ( .d(n1898), .o(net_6053), .ck(clk) );
ms00f80 l0351 ( .d(n1903), .o(net_6258), .ck(clk) );
ms00f80 l0352 ( .d(n1908), .o(_net_7379), .ck(clk) );
ms00f80 l0353 ( .d(n1913), .o(net_6543), .ck(clk) );
ms00f80 l0354 ( .d(n1918), .o(net_7116), .ck(clk) );
ms00f80 l0355 ( .d(n1922), .o(_net_6070), .ck(clk) );
ms00f80 l0356 ( .d(n1927), .o(_net_6690), .ck(clk) );
ms00f80 l0357 ( .d(n1932), .o(net_6995), .ck(clk) );
ms00f80 l0358 ( .d(n1936), .o(net_241), .ck(clk) );
ms00f80 l0359 ( .d(n1941), .o(net_6433), .ck(clk) );
ms00f80 l0360 ( .d(n1945), .o(_net_7472), .ck(clk) );
ms00f80 l0361 ( .d(n1950), .o(_net_7532), .ck(clk) );
ms00f80 l0362 ( .d(n1954), .o(net_7052), .ck(clk) );
ms00f80 l0363 ( .d(n1959), .o(_net_129), .ck(clk) );
ms00f80 l0364 ( .d(n1964), .o(net_6346), .ck(clk) );
ms00f80 l0365 ( .d(n1969), .o(_net_7594), .ck(clk) );
ms00f80 l0366 ( .d(n1973), .o(net_6800), .ck(clk) );
ms00f80 l0367 ( .d(n1978), .o(net_7174), .ck(clk) );
ms00f80 l0368 ( .d(n1983), .o(net_6274), .ck(clk) );
ms00f80 l0369 ( .d(n1988), .o(_net_6108), .ck(clk) );
ms00f80 l0370 ( .d(n1993), .o(net_7520), .ck(clk) );
ms00f80 l0371 ( .d(n1998), .o(net_6737), .ck(clk) );
ms00f80 l0372 ( .d(n2002), .o(net_6303), .ck(clk) );
ms00f80 l0373 ( .d(n2007), .o(net_6812), .ck(clk) );
ms00f80 l0374 ( .d(n2011), .o(net_7188), .ck(clk) );
ms00f80 l0375 ( .d(n2016), .o(_net_7426), .ck(clk) );
ms00f80 l0376 ( .d(n2021), .o(net_7790), .ck(clk) );
ms00f80 l0377 ( .d(n2026), .o(_net_6107), .ck(clk) );
ms00f80 l0378 ( .d(n2031), .o(net_6318), .ck(clk) );
ms00f80 l0379 ( .d(n2036), .o(net_319), .ck(clk) );
ms00f80 l0380 ( .d(n2041), .o(_net_7483), .ck(clk) );
ms00f80 l0381 ( .d(n2046), .o(_net_7093), .ck(clk) );
ms00f80 l0382 ( .d(n2051), .o(net_7391), .ck(clk) );
ms00f80 l0383 ( .d(n2055), .o(_net_7465), .ck(clk) );
ms00f80 l0384 ( .d(n2060), .o(_net_7352), .ck(clk) );
ms00f80 l0385 ( .d(n2065), .o(_net_6125), .ck(clk) );
ms00f80 l0386 ( .d(n2070), .o(_net_6827), .ck(clk) );
ms00f80 l0387 ( .d(n2074), .o(net_7201), .ck(clk) );
ms00f80 l0388 ( .d(n2079), .o(net_7754), .ck(clk) );
ms00f80 l0389 ( .d(n2084), .o(net_7371), .ck(clk) );
ms00f80 l0390 ( .d(n2088), .o(net_7063), .ck(clk) );
ms00f80 l0391 ( .d(n2093), .o(net_6893), .ck(clk) );
ms00f80 l0392 ( .d(n2098), .o(net_6709), .ck(clk) );
ms00f80 l0393 ( .d(n2102), .o(net_6741), .ck(clk) );
ms00f80 l0394 ( .d(n2106), .o(net_6191), .ck(clk) );
ms00f80 l0395 ( .d(n2111), .o(net_7003), .ck(clk) );
ms00f80 l0396 ( .d(n2115), .o(net_6452), .ck(clk) );
ms00f80 l0397 ( .d(n2119), .o(net_6603), .ck(clk) );
ms00f80 l0398 ( .d(n2122), .o(net_7076), .ck(clk) );
ms00f80 l0399 ( .d(n2127), .o(net_6310), .ck(clk) );
ms00f80 l0400 ( .d(n2132), .o(net_7147), .ck(clk) );
ms00f80 l0401 ( .d(n2136), .o(net_6730), .ck(clk) );
ms00f80 l0402 ( .d(n2140), .o(_net_7683), .ck(clk) );
ms00f80 l0403 ( .d(n2144), .o(net_7179), .ck(clk) );
ms00f80 l0404 ( .d(n2149), .o(net_7144), .ck(clk) );
ms00f80 l0405 ( .d(n2152), .o(net_7613), .ck(clk) );
ms00f80 l0406 ( .d(n2157), .o(net_6336), .ck(clk) );
ms00f80 l0407 ( .d(n2162), .o(_net_7554), .ck(clk) );
ms00f80 l0408 ( .d(n2167), .o(_net_7649), .ck(clk) );
ms00f80 l0409 ( .d(n2172), .o(_net_6963), .ck(clk) );
ms00f80 l0410 ( .d(n2177), .o(x397), .ck(clk) );
ms00f80 l0411 ( .d(n2181), .o(_net_7763), .ck(clk) );
ms00f80 l0412 ( .d(n2186), .o(net_6443), .ck(clk) );
ms00f80 l0413 ( .d(n2189), .o(net_6540), .ck(clk) );
ms00f80 l0414 ( .d(n2194), .o(_net_6177), .ck(clk) );
ms00f80 l0415 ( .d(n2199), .o(_net_7229), .ck(clk) );
ms00f80 l0416 ( .d(n2203), .o(net_6658), .ck(clk) );
ms00f80 l0417 ( .d(n2208), .o(_net_5963), .ck(clk) );
ms00f80 l0418 ( .d(n2213), .o(_net_6016), .ck(clk) );
ms00f80 l0419 ( .d(n2218), .o(net_6456), .ck(clk) );
ms00f80 l0420 ( .d(n2222), .o(net_6556), .ck(clk) );
ms00f80 l0421 ( .d(n2227), .o(_net_6960), .ck(clk) );
ms00f80 l0422 ( .d(n2232), .o(_net_263), .ck(clk) );
ms00f80 l0423 ( .d(n2237), .o(_net_6184), .ck(clk) );
ms00f80 l0424 ( .d(n2242), .o(_net_7724), .ck(clk) );
ms00f80 l0425 ( .d(n2247), .o(x494), .ck(clk) );
ms00f80 l0426 ( .d(n2251), .o(_net_6401), .ck(clk) );
ms00f80 l0427 ( .d(n2256), .o(net_7458), .ck(clk) );
ms00f80 l0428 ( .d(n2260), .o(net_7671), .ck(clk) );
ms00f80 l0429 ( .d(n2265), .o(_net_7401), .ck(clk) );
ms00f80 l0430 ( .d(n2270), .o(_net_5977), .ck(clk) );
ms00f80 l0431 ( .d(n2275), .o(_net_6139), .ck(clk) );
ms00f80 l0432 ( .d(n2280), .o(_net_7748), .ck(clk) );
ms00f80 l0433 ( .d(n2284), .o(net_322), .ck(clk) );
ms00f80 l0434 ( .d(n2288), .o(net_142), .ck(clk) );
ms00f80 l0435 ( .d(n2293), .o(net_6366), .ck(clk) );
ms00f80 l0436 ( .d(n2298), .o(_net_6015), .ck(clk) );
ms00f80 l0437 ( .d(n2303), .o(_net_6187), .ck(clk) );
ms00f80 l0438 ( .d(n2307), .o(net_7194), .ck(clk) );
ms00f80 l0439 ( .d(n2312), .o(_net_7556), .ck(clk) );
ms00f80 l0440 ( .d(n2316), .o(net_6035), .ck(clk) );
ms00f80 l0441 ( .d(n2321), .o(net_7159), .ck(clk) );
ms00f80 l0442 ( .d(n2324), .o(net_323), .ck(clk) );
ms00f80 l0443 ( .d(n2329), .o(_net_6134), .ck(clk) );
ms00f80 l0444 ( .d(n2334), .o(_net_7747), .ck(clk) );
ms00f80 l0445 ( .d(n2338), .o(net_6920), .ck(clk) );
ms00f80 l0446 ( .d(n2342), .o(net_6501), .ck(clk) );
ms00f80 l0447 ( .d(n2347), .o(net_6849), .ck(clk) );
ms00f80 l0448 ( .d(n2350), .o(net_6236), .ck(clk) );
ms00f80 l0449 ( .d(n2355), .o(net_6277), .ck(clk) );
ms00f80 l0450 ( .d(n2360), .o(net_6912), .ck(clk) );
ms00f80 l0451 ( .d(n2365), .o(_net_6163), .ck(clk) );
ms00f80 l0452 ( .d(n2370), .o(net_6593), .ck(clk) );
ms00f80 l0453 ( .d(n2373), .o(net_6398), .ck(clk) );
ms00f80 l0454 ( .d(n2377), .o(_net_7720), .ck(clk) );
ms00f80 l0455 ( .d(n2381), .o(net_7527), .ck(clk) );
ms00f80 l0456 ( .d(n2386), .o(_net_6169), .ck(clk) );
ms00f80 l0457 ( .d(n2391), .o(net_6576), .ck(clk) );
ms00f80 l0458 ( .d(n2395), .o(net_183), .ck(clk) );
ms00f80 l0459 ( .d(n2399), .o(net_6758), .ck(clk) );
ms00f80 l0460 ( .d(n2404), .o(net_7608), .ck(clk) );
ms00f80 l0461 ( .d(n2409), .o(_net_7511), .ck(clk) );
ms00f80 l0462 ( .d(n2414), .o(x699), .ck(clk) );
ms00f80 l0463 ( .d(n2417), .o(net_6680), .ck(clk) );
ms00f80 l0464 ( .d(n2422), .o(net_7016), .ck(clk) );
ms00f80 l0465 ( .d(n2426), .o(net_6833), .ck(clk) );
ms00f80 l0466 ( .d(n2430), .o(_net_7431), .ck(clk) );
ms00f80 l0467 ( .d(n2435), .o(_net_279), .ck(clk) );
ms00f80 l0468 ( .d(n2440), .o(net_7240), .ck(clk) );
ms00f80 l0469 ( .d(n2444), .o(_net_5972), .ck(clk) );
ms00f80 l0470 ( .d(n2448), .o(net_377), .ck(clk) );
ms00f80 l0471 ( .d(n2452), .o(net_6821), .ck(clk) );
ms00f80 l0472 ( .d(n2457), .o(_net_5984), .ck(clk) );
ms00f80 l0473 ( .d(n2462), .o(net_6426), .ck(clk) );
ms00f80 l0474 ( .d(n2465), .o(net_6918), .ck(clk) );
ms00f80 l0475 ( .d(n2470), .o(_net_6118), .ck(clk) );
ms00f80 l0476 ( .d(n2474), .o(net_6672), .ck(clk) );
ms00f80 l0477 ( .d(n2479), .o(_net_7294), .ck(clk) );
ms00f80 l0478 ( .d(n2484), .o(net_224), .ck(clk) );
ms00f80 l0479 ( .d(n2488), .o(net_6764), .ck(clk) );
ms00f80 l0480 ( .d(n2493), .o(net_6435), .ck(clk) );
ms00f80 l0481 ( .d(n2496), .o(net_7207), .ck(clk) );
ms00f80 l0482 ( .d(n2500), .o(net_7639), .ck(clk) );
ms00f80 l0483 ( .d(n2505), .o(_net_7704), .ck(clk) );
ms00f80 l0484 ( .d(n2510), .o(net_252), .ck(clk) );
ms00f80 l0485 ( .d(n2515), .o(net_6014), .ck(clk) );
ms00f80 l0486 ( .d(n2519), .o(net_6522), .ck(clk) );
ms00f80 l0487 ( .d(n2524), .o(net_179), .ck(clk) );
ms00f80 l0488 ( .d(n2529), .o(_net_7419), .ck(clk) );
ms00f80 l0489 ( .d(n2534), .o(_net_6160), .ck(clk) );
ms00f80 l0490 ( .d(n2539), .o(net_134), .ck(clk) );
ms00f80 l0491 ( .d(n2543), .o(net_6939), .ck(clk) );
ms00f80 l0492 ( .d(n2547), .o(net_7337), .ck(clk) );
ms00f80 l0493 ( .d(n2552), .o(_net_7445), .ck(clk) );
ms00f80 l0494 ( .d(n2556), .o(net_6951), .ck(clk) );
ms00f80 l0495 ( .d(n2561), .o(net_300), .ck(clk) );
ms00f80 l0496 ( .d(n2566), .o(_net_7663), .ck(clk) );
ms00f80 l0497 ( .d(n2570), .o(net_6898), .ck(clk) );
ms00f80 l0498 ( .d(n2575), .o(_net_176), .ck(clk) );
ms00f80 l0499 ( .d(n2580), .o(net_207), .ck(clk) );
ms00f80 l0500 ( .d(n2585), .o(net_7779), .ck(clk) );
ms00f80 l0501 ( .d(n2590), .o(net_7096), .ck(clk) );
ms00f80 l0502 ( .d(n2594), .o(net_6391), .ck(clk) );
ms00f80 l0503 ( .d(n2597), .o(net_7032), .ck(clk) );
ms00f80 l0504 ( .d(n2601), .o(net_6517), .ck(clk) );
ms00f80 l0505 ( .d(n2605), .o(net_6513), .ck(clk) );
ms00f80 l0506 ( .d(n2610), .o(net_6377), .ck(clk) );
ms00f80 l0507 ( .d(n2615), .o(net_6967), .ck(clk) );
ms00f80 l0508 ( .d(n2618), .o(net_7060), .ck(clk) );
ms00f80 l0509 ( .d(n2622), .o(net_7089), .ck(clk) );
ms00f80 l0510 ( .d(n2627), .o(net_6322), .ck(clk) );
ms00f80 l0511 ( .d(n2632), .o(_net_7765), .ck(clk) );
ms00f80 l0512 ( .d(n2637), .o(net_257), .ck(clk) );
ms00f80 l0513 ( .d(n2642), .o(net_6341), .ck(clk) );
ms00f80 l0514 ( .d(n2647), .o(net_6588), .ck(clk) );
ms00f80 l0515 ( .d(n2651), .o(net_187), .ck(clk) );
ms00f80 l0516 ( .d(n2656), .o(net_6606), .ck(clk) );
ms00f80 l0517 ( .d(n2660), .o(net_6215), .ck(clk) );
ms00f80 l0518 ( .d(n2665), .o(_net_6121), .ck(clk) );
ms00f80 l0519 ( .d(n2670), .o(net_6330), .ck(clk) );
ms00f80 l0520 ( .d(n2675), .o(net_6890), .ck(clk) );
ms00f80 l0521 ( .d(n2679), .o(net_6964), .ck(clk) );
ms00f80 l0522 ( .d(n2682), .o(net_7057), .ck(clk) );
ms00f80 l0523 ( .d(n2687), .o(net_7777), .ck(clk) );
ms00f80 l0524 ( .d(n2692), .o(net_7393), .ck(clk) );
ms00f80 l0525 ( .d(n2696), .o(_net_6822), .ck(clk) );
ms00f80 l0526 ( .d(n2701), .o(net_6981), .ck(clk) );
ms00f80 l0527 ( .d(n2705), .o(net_6434), .ck(clk) );
ms00f80 l0528 ( .d(n2709), .o(net_6969), .ck(clk) );
ms00f80 l0529 ( .d(n2713), .o(_net_126), .ck(clk) );
ms00f80 l0530 ( .d(n2718), .o(net_238), .ck(clk) );
ms00f80 l0531 ( .d(n2723), .o(_net_280), .ck(clk) );
ms00f80 l0532 ( .d(n2727), .o(net_346), .ck(clk) );
ms00f80 l0533 ( .d(n2732), .o(_net_7314), .ck(clk) );
ms00f80 l0534 ( .d(n2737), .o(net_7708), .ck(clk) );
ms00f80 l0535 ( .d(n2741), .o(net_6586), .ck(clk) );
ms00f80 l0536 ( .d(n2745), .o(net_6725), .ck(clk) );
ms00f80 l0537 ( .d(n2748), .o(net_6955), .ck(clk) );
ms00f80 l0538 ( .d(n2753), .o(net_163), .ck(clk) );
ms00f80 l0539 ( .d(n2758), .o(_net_6097), .ck(clk) );
ms00f80 l0540 ( .d(n2762), .o(net_7225), .ck(clk) );
ms00f80 l0541 ( .d(n2767), .o(net_7108), .ck(clk) );
ms00f80 l0542 ( .d(n2771), .o(_net_6022), .ck(clk) );
ms00f80 l0543 ( .d(n2776), .o(_net_5978), .ck(clk) );
ms00f80 l0544 ( .d(n2781), .o(net_6880), .ck(clk) );
ms00f80 l0545 ( .d(n2784), .o(net_7343), .ck(clk) );
ms00f80 l0546 ( .d(n2788), .o(net_6496), .ck(clk) );
ms00f80 l0547 ( .d(n2792), .o(net_6664), .ck(clk) );
ms00f80 l0548 ( .d(n2797), .o(net_232), .ck(clk) );
ms00f80 l0549 ( .d(n2801), .o(net_6524), .ck(clk) );
ms00f80 l0550 ( .d(n2805), .o(_net_7820), .ck(clk) );
ms00f80 l0551 ( .d(n2810), .o(_net_214), .ck(clk) );
ms00f80 l0552 ( .d(n2814), .o(net_6539), .ck(clk) );
ms00f80 l0553 ( .d(n2819), .o(net_6579), .ck(clk) );
ms00f80 l0554 ( .d(n2823), .o(net_7024), .ck(clk) );
ms00f80 l0555 ( .d(n2827), .o(net_7153), .ck(clk) );
ms00f80 l0556 ( .d(n2831), .o(_net_6156), .ck(clk) );
ms00f80 l0557 ( .d(n2836), .o(_net_6029), .ck(clk) );
ms00f80 l0558 ( .d(n2840), .o(net_6631), .ck(clk) );
ms00f80 l0559 ( .d(n2845), .o(_net_7261), .ck(clk) );
ms00f80 l0560 ( .d(n2850), .o(net_7670), .ck(clk) );
ms00f80 l0561 ( .d(n2855), .o(_net_7501), .ck(clk) );
ms00f80 l0562 ( .d(n2860), .o(net_7236), .ck(clk) );
ms00f80 l0563 ( .d(n2864), .o(net_6246), .ck(clk) );
ms00f80 l0564 ( .d(n2869), .o(net_6478), .ck(clk) );
ms00f80 l0565 ( .d(n2873), .o(net_6578), .ck(clk) );
ms00f80 l0566 ( .d(n2877), .o(net_6244), .ck(clk) );
ms00f80 l0567 ( .d(n2882), .o(net_7547), .ck(clk) );
ms00f80 l0568 ( .d(n2885), .o(net_6813), .ck(clk) );
ms00f80 l0569 ( .d(n2890), .o(_net_7572), .ck(clk) );
ms00f80 l0570 ( .d(n2895), .o(net_7756), .ck(clk) );
ms00f80 l0571 ( .d(n2900), .o(_net_7722), .ck(clk) );
ms00f80 l0572 ( .d(n2904), .o(net_7461), .ck(clk) );
ms00f80 l0573 ( .d(n2908), .o(net_6946), .ck(clk) );
ms00f80 l0574 ( .d(n2913), .o(net_7336), .ck(clk) );
ms00f80 l0575 ( .d(n2918), .o(x315), .ck(clk) );
ms00f80 l0576 ( .d(n2922), .o(net_7022), .ck(clk) );
ms00f80 l0577 ( .d(n2926), .o(net_6755), .ck(clk) );
ms00f80 l0578 ( .d(n2930), .o(_net_6221), .ck(clk) );
ms00f80 l0579 ( .d(n2935), .o(_net_5920), .ck(clk) );
ms00f80 l0580 ( .d(n2939), .o(net_6781), .ck(clk) );
ms00f80 l0581 ( .d(n2944), .o(net_7158), .ck(clk) );
ms00f80 l0582 ( .d(n2948), .o(_net_5969), .ck(clk) );
ms00f80 l0583 ( .d(n2953), .o(_net_7552), .ck(clk) );
ms00f80 l0584 ( .d(n2958), .o(net_7457), .ck(clk) );
ms00f80 l0585 ( .d(n2963), .o(net_6338), .ck(clk) );
ms00f80 l0586 ( .d(n2967), .o(net_337), .ck(clk) );
ms00f80 l0587 ( .d(n2972), .o(net_7007), .ck(clk) );
ms00f80 l0588 ( .d(n2976), .o(_net_266), .ck(clk) );
ms00f80 l0589 ( .d(n2981), .o(_net_6553), .ck(clk) );
ms00f80 l0590 ( .d(n2986), .o(_net_6063), .ck(clk) );
ms00f80 l0591 ( .d(n2991), .o(_net_7531), .ck(clk) );
ms00f80 l0592 ( .d(n2996), .o(net_6438), .ck(clk) );
ms00f80 l0593 ( .d(n3000), .o(_net_6038), .ck(clk) );
ms00f80 l0594 ( .d(n3005), .o(_net_6090), .ck(clk) );
ms00f80 l0595 ( .d(n3010), .o(_net_7751), .ck(clk) );
ms00f80 l0596 ( .d(n3015), .o(net_7609), .ck(clk) );
ms00f80 l0597 ( .d(n3020), .o(_net_7320), .ck(clk) );
ms00f80 l0598 ( .d(n3025), .o(_net_173), .ck(clk) );
ms00f80 l0599 ( .d(n3030), .o(net_7105), .ck(clk) );
ms00f80 l0600 ( .d(n3033), .o(net_6906), .ck(clk) );
ms00f80 l0601 ( .d(n3037), .o(net_6909), .ck(clk) );
ms00f80 l0602 ( .d(n3042), .o(_net_6023), .ck(clk) );
ms00f80 l0603 ( .d(n3047), .o(_net_7667), .ck(clk) );
ms00f80 l0604 ( .d(n3052), .o(net_7136), .ck(clk) );
ms00f80 l0605 ( .d(n3056), .o(_net_226), .ck(clk) );
ms00f80 l0606 ( .d(n3061), .o(net_7121), .ck(clk) );
ms00f80 l0607 ( .d(n3065), .o(_net_184), .ck(clk) );
ms00f80 l0608 ( .d(n3069), .o(net_6938), .ck(clk) );
ms00f80 l0609 ( .d(n3074), .o(net_6717), .ck(clk) );
ms00f80 l0610 ( .d(n3078), .o(net_233), .ck(clk) );
ms00f80 l0611 ( .d(n3082), .o(net_6796), .ck(clk) );
ms00f80 l0612 ( .d(n3087), .o(_net_6688), .ck(clk) );
ms00f80 l0613 ( .d(n3092), .o(_net_6281), .ck(clk) );
ms00f80 l0614 ( .d(n3097), .o(_net_128), .ck(clk) );
ms00f80 l0615 ( .d(n3102), .o(net_6706), .ck(clk) );
ms00f80 l0616 ( .d(n3105), .o(net_303), .ck(clk) );
ms00f80 l0617 ( .d(n3110), .o(net_6473), .ck(clk) );
ms00f80 l0618 ( .d(n3114), .o(net_6743), .ck(clk) );
ms00f80 l0619 ( .d(n3117), .o(net_153), .ck(clk) );
ms00f80 l0620 ( .d(n3121), .o(net_7643), .ck(clk) );
ms00f80 l0621 ( .d(n3126), .o(net_7387), .ck(clk) );
ms00f80 l0622 ( .d(n3130), .o(_net_7410), .ck(clk) );
ms00f80 l0623 ( .d(n3134), .o(net_6639), .ck(clk) );
ms00f80 l0624 ( .d(n3139), .o(_net_7557), .ck(clk) );
ms00f80 l0625 ( .d(n3143), .o(net_6681), .ck(clk) );
ms00f80 l0626 ( .d(n3148), .o(_net_7449), .ck(clk) );
ms00f80 l0627 ( .d(n3152), .o(net_7040), .ck(clk) );
ms00f80 l0628 ( .d(n3157), .o(_net_7690), .ck(clk) );
ms00f80 l0629 ( .d(n3162), .o(net_6751), .ck(clk) );
ms00f80 l0630 ( .d(n3165), .o(net_7738), .ck(clk) );
ms00f80 l0631 ( .d(n3170), .o(_net_7470), .ck(clk) );
ms00f80 l0632 ( .d(n3174), .o(net_152), .ck(clk) );
ms00f80 l0633 ( .d(n3178), .o(net_6450), .ck(clk) );
ms00f80 l0634 ( .d(n3182), .o(_net_7350), .ck(clk) );
ms00f80 l0635 ( .d(n3186), .o(net_135), .ck(clk) );
ms00f80 l0636 ( .d(n3190), .o(net_6861), .ck(clk) );
ms00f80 l0637 ( .d(n3194), .o(_net_7277), .ck(clk) );
ms00f80 l0638 ( .d(n3199), .o(net_7536), .ck(clk) );
ms00f80 l0639 ( .d(n3203), .o(_net_178), .ck(clk) );
ms00f80 l0640 ( .d(n3207), .o(net_6488), .ck(clk) );
ms00f80 l0641 ( .d(n3212), .o(_net_7326), .ck(clk) );
ms00f80 l0642 ( .d(n3217), .o(_net_6110), .ck(clk) );
ms00f80 l0643 ( .d(n3222), .o(_net_7478), .ck(clk) );
ms00f80 l0644 ( .d(n3226), .o(net_6233), .ck(clk) );
ms00f80 l0645 ( .d(n3231), .o(_net_154), .ck(clk) );
ms00f80 l0646 ( .d(n3235), .o(_net_7812), .ck(clk) );
ms00f80 l0647 ( .d(n3240), .o(_net_6175), .ck(clk) );
ms00f80 l0648 ( .d(n3244), .o(net_6652), .ck(clk) );
ms00f80 l0649 ( .d(n3249), .o(_net_6259), .ck(clk) );
ms00f80 l0650 ( .d(n3254), .o(_net_272), .ck(clk) );
ms00f80 l0651 ( .d(n3258), .o(_net_7821), .ck(clk) );
ms00f80 l0652 ( .d(n3263), .o(_net_116), .ck(clk) );
ms00f80 l0653 ( .d(n3268), .o(_net_6102), .ck(clk) );
ms00f80 l0654 ( .d(n3272), .o(net_6661), .ck(clk) );
ms00f80 l0655 ( .d(n3276), .o(net_7488), .ck(clk) );
ms00f80 l0656 ( .d(n3280), .o(net_6760), .ck(clk) );
ms00f80 l0657 ( .d(n3285), .o(_net_6204), .ck(clk) );
ms00f80 l0658 ( .d(n3290), .o(net_7710), .ck(clk) );
ms00f80 l0659 ( .d(n3294), .o(_net_6083), .ck(clk) );
ms00f80 l0660 ( .d(n3299), .o(net_6623), .ck(clk) );
ms00f80 l0661 ( .d(n3303), .o(net_6536), .ck(clk) );
ms00f80 l0662 ( .d(n3308), .o(_net_7266), .ck(clk) );
ms00f80 l0663 ( .d(n3313), .o(_net_6171), .ck(clk) );
ms00f80 l0664 ( .d(n3318), .o(net_6883), .ck(clk) );
ms00f80 l0665 ( .d(n3322), .o(x447), .ck(clk) );
ms00f80 l0666 ( .d(n3325), .o(net_7310), .ck(clk) );
ms00f80 l0667 ( .d(n3330), .o(net_6868), .ck(clk) );
ms00f80 l0668 ( .d(n3333), .o(net_7344), .ck(clk) );
ms00f80 l0669 ( .d(n3338), .o(_net_6041), .ck(clk) );
ms00f80 l0670 ( .d(n3343), .o(_net_6199), .ck(clk) );
ms00f80 l0671 ( .d(n3348), .o(net_7140), .ck(clk) );
ms00f80 l0672 ( .d(n3352), .o(x589), .ck(clk) );
ms00f80 l0673 ( .d(n3356), .o(_net_7583), .ck(clk) );
ms00f80 l0674 ( .d(n3361), .o(net_6247), .ck(clk) );
ms00f80 l0675 ( .d(n3365), .o(net_6548), .ck(clk) );
ms00f80 l0676 ( .d(n3370), .o(_net_5980), .ck(clk) );
ms00f80 l0677 ( .d(n3374), .o(net_7517), .ck(clk) );
ms00f80 l0678 ( .d(n3379), .o(net_6698), .ck(clk) );
ms00f80 l0679 ( .d(n3383), .o(net_6485), .ck(clk) );
ms00f80 l0680 ( .d(n3386), .o(net_7042), .ck(clk) );
ms00f80 l0681 ( .d(n3390), .o(_net_7814), .ck(clk) );
ms00f80 l0682 ( .d(n3395), .o(_net_6142), .ck(clk) );
ms00f80 l0683 ( .d(n3400), .o(_net_7619), .ck(clk) );
ms00f80 l0684 ( .d(n3404), .o(net_371), .ck(clk) );
ms00f80 l0685 ( .d(n3408), .o(net_6547), .ck(clk) );
ms00f80 l0686 ( .d(n3413), .o(net_6214), .ck(clk) );
ms00f80 l0687 ( .d(n3418), .o(net_7248), .ck(clk) );
ms00f80 l0688 ( .d(n3422), .o(net_197), .ck(clk) );
ms00f80 l0689 ( .d(n3427), .o(_net_7618), .ck(clk) );
ms00f80 l0690 ( .d(n3431), .o(net_7743), .ck(clk) );
ms00f80 l0691 ( .d(n3436), .o(net_7120), .ck(clk) );
ms00f80 l0692 ( .d(n3440), .o(_net_211), .ck(clk) );
ms00f80 l0693 ( .d(n3445), .o(net_334), .ck(clk) );
ms00f80 l0694 ( .d(n3450), .o(net_6369), .ck(clk) );
ms00f80 l0695 ( .d(n3455), .o(x786), .ck(clk) );
ms00f80 l0696 ( .d(n3459), .o(_net_6075), .ck(clk) );
ms00f80 l0697 ( .d(n3464), .o(_net_191), .ck(clk) );
ms00f80 l0698 ( .d(n3469), .o(net_7213), .ck(clk) );
ms00f80 l0699 ( .d(n3474), .o(_net_6130), .ck(clk) );
ms00f80 l0700 ( .d(n3479), .o(net_6332), .ck(clk) );
ms00f80 l0701 ( .d(n3484), .o(_net_6290), .ck(clk) );
ms00f80 l0702 ( .d(n3489), .o(_net_7362), .ck(clk) );
ms00f80 l0703 ( .d(n3494), .o(net_7241), .ck(clk) );
ms00f80 l0704 ( .d(n3497), .o(net_140), .ck(clk) );
ms00f80 l0705 ( .d(n3502), .o(net_7766), .ck(clk) );
ms00f80 l0706 ( .d(n3507), .o(_net_6078), .ck(clk) );
ms00f80 l0707 ( .d(n3511), .o(net_7195), .ck(clk) );
ms00f80 l0708 ( .d(n3516), .o(_net_6687), .ck(clk) );
ms00f80 l0709 ( .d(n3520), .o(net_6765), .ck(clk) );
ms00f80 l0710 ( .d(n3524), .o(net_6216), .ck(clk) );
ms00f80 l0711 ( .d(n3528), .o(net_7082), .ck(clk) );
ms00f80 l0712 ( .d(n3532), .o(net_329), .ck(clk) );
ms00f80 l0713 ( .d(n3537), .o(net_6254), .ck(clk) );
ms00f80 l0714 ( .d(n3542), .o(net_6885), .ck(clk) );
ms00f80 l0715 ( .d(n3546), .o(net_7642), .ck(clk) );
ms00f80 l0716 ( .d(n3551), .o(net_7231), .ck(clk) );
ms00f80 l0717 ( .d(n3555), .o(net_310), .ck(clk) );
ms00f80 l0718 ( .d(n3559), .o(net_6505), .ck(clk) );
ms00f80 l0719 ( .d(n3564), .o(net_6873), .ck(clk) );
ms00f80 l0720 ( .d(n3567), .o(net_7672), .ck(clk) );
ms00f80 l0721 ( .d(n3572), .o(_net_7703), .ck(clk) );
ms00f80 l0722 ( .d(n3577), .o(_net_6408), .ck(clk) );
ms00f80 l0723 ( .d(n3582), .o(net_255), .ck(clk) );
ms00f80 l0724 ( .d(n3587), .o(net_6476), .ck(clk) );
ms00f80 l0725 ( .d(n3590), .o(net_6530), .ck(clk) );
ms00f80 l0726 ( .d(n3595), .o(_net_5962), .ck(clk) );
ms00f80 l0727 ( .d(n3600), .o(net_6583), .ck(clk) );
ms00f80 l0728 ( .d(n3604), .o(net_7678), .ck(clk) );
ms00f80 l0729 ( .d(n3609), .o(_net_6092), .ck(clk) );
ms00f80 l0730 ( .d(n3614), .o(_net_5988), .ck(clk) );
ms00f80 l0731 ( .d(n3618), .o(net_6674), .ck(clk) );
ms00f80 l0732 ( .d(n3623), .o(net_6320), .ck(clk) );
ms00f80 l0733 ( .d(n3628), .o(_net_7781), .ck(clk) );
ms00f80 l0734 ( .d(n3633), .o(_net_7665), .ck(clk) );
ms00f80 l0735 ( .d(n3638), .o(net_7378), .ck(clk) );
ms00f80 l0736 ( .d(n3642), .o(net_7737), .ck(clk) );
ms00f80 l0737 ( .d(n3647), .o(x217), .ck(clk) );
ms00f80 l0738 ( .d(n3651), .o(net_7157), .ck(clk) );
ms00f80 l0739 ( .d(n3655), .o(net_6591), .ck(clk) );
ms00f80 l0740 ( .d(n3658), .o(net_6395), .ck(clk) );
ms00f80 l0741 ( .d(n3661), .o(net_7490), .ck(clk) );
ms00f80 l0742 ( .d(n3666), .o(_net_7424), .ck(clk) );
ms00f80 l0743 ( .d(n3670), .o(net_7061), .ck(clk) );
ms00f80 l0744 ( .d(n3675), .o(_net_7728), .ck(clk) );
ms00f80 l0745 ( .d(n3679), .o(net_7171), .ck(clk) );
ms00f80 l0746 ( .d(n3684), .o(_net_5854), .ck(clk) );
ms00f80 l0747 ( .d(n3689), .o(net_6605), .ck(clk) );
ms00f80 l0748 ( .d(n3693), .o(_net_7250), .ck(clk) );
ms00f80 l0749 ( .d(n3698), .o(_net_5853), .ck(clk) );
ms00f80 l0750 ( .d(n3703), .o(net_6976), .ck(clk) );
ms00f80 l0751 ( .d(n3707), .o(net_6721), .ck(clk) );
ms00f80 l0752 ( .d(n3711), .o(net_7775), .ck(clk) );
ms00f80 l0753 ( .d(n3716), .o(net_6486), .ck(clk) );
ms00f80 l0754 ( .d(n3720), .o(net_6268), .ck(clk) );
ms00f80 l0755 ( .d(n3725), .o(net_6881), .ck(clk) );
ms00f80 l0756 ( .d(n3729), .o(net_7048), .ck(clk) );
ms00f80 l0757 ( .d(n3733), .o(net_7799), .ck(clk) );
ms00f80 l0758 ( .d(n3737), .o(_net_7444), .ck(clk) );
ms00f80 l0759 ( .d(n3742), .o(_net_7598), .ck(clk) );
ms00f80 l0760 ( .d(n3747), .o(net_6325), .ck(clk) );
ms00f80 l0761 ( .d(n3752), .o(net_6245), .ck(clk) );
ms00f80 l0762 ( .d(n3756), .o(net_336), .ck(clk) );
ms00f80 l0763 ( .d(n3761), .o(net_6442), .ck(clk) );
ms00f80 l0764 ( .d(n3765), .o(_net_290), .ck(clk) );
ms00f80 l0765 ( .d(n3770), .o(net_6991), .ck(clk) );
ms00f80 l0766 ( .d(n3773), .o(net_6928), .ck(clk) );
ms00f80 l0767 ( .d(n3777), .o(net_6525), .ck(clk) );
ms00f80 l0768 ( .d(n3782), .o(_net_7626), .ck(clk) );
ms00f80 l0769 ( .d(n3787), .o(_net_7092), .ck(clk) );
ms00f80 l0770 ( .d(n3791), .o(net_6666), .ck(clk) );
ms00f80 l0771 ( .d(n3796), .o(_net_7785), .ck(clk) );
ms00f80 l0772 ( .d(n3801), .o(net_7149), .ck(clk) );
ms00f80 l0773 ( .d(n3805), .o(net_7714), .ck(clk) );
ms00f80 l0774 ( .d(n3809), .o(net_6429), .ck(clk) );
ms00f80 l0775 ( .d(n3813), .o(net_182), .ck(clk) );
ms00f80 l0776 ( .d(n3817), .o(net_339), .ck(clk) );
ms00f80 l0777 ( .d(n3822), .o(net_6252), .ck(clk) );
ms00f80 l0778 ( .d(n3827), .o(net_286), .ck(clk) );
ms00f80 l0779 ( .d(n3831), .o(net_6799), .ck(clk) );
ms00f80 l0780 ( .d(n3836), .o(_net_6419), .ck(clk) );
ms00f80 l0781 ( .d(n3841), .o(_net_7652), .ck(clk) );
ms00f80 l0782 ( .d(n3846), .o(_net_6158), .ck(clk) );
ms00f80 l0783 ( .d(n3851), .o(net_6829), .ck(clk) );
ms00f80 l0784 ( .d(n3855), .o(net_6595), .ck(clk) );
ms00f80 l0785 ( .d(n3859), .o(_net_7290), .ck(clk) );
ms00f80 l0786 ( .d(n3864), .o(net_6850), .ck(clk) );
ms00f80 l0787 ( .d(n3867), .o(net_6636), .ck(clk) );
ms00f80 l0788 ( .d(n3872), .o(_net_188), .ck(clk) );
ms00f80 l0789 ( .d(n3877), .o(_net_6065), .ck(clk) );
ms00f80 l0790 ( .d(n3881), .o(net_6899), .ck(clk) );
ms00f80 l0791 ( .d(n3886), .o(_net_7574), .ck(clk) );
ms00f80 l0792 ( .d(n3891), .o(_net_123), .ck(clk) );
ms00f80 l0793 ( .d(n3896), .o(net_6855), .ck(clk) );
ms00f80 l0794 ( .d(n3899), .o(net_7034), .ck(clk) );
ms00f80 l0795 ( .d(n3904), .o(net_7239), .ck(clk) );
ms00f80 l0796 ( .d(n3908), .o(net_223), .ck(clk) );
ms00f80 l0797 ( .d(n3913), .o(_net_7270), .ck(clk) );
ms00f80 l0798 ( .d(n3917), .o(net_7184), .ck(clk) );
ms00f80 l0799 ( .d(n3922), .o(_net_6116), .ck(clk) );
ms00f80 l0800 ( .d(n3927), .o(_net_7563), .ck(clk) );
ms00f80 l0801 ( .d(n3932), .o(_net_7418), .ck(clk) );
ms00f80 l0802 ( .d(n3936), .o(net_6685), .ck(clk) );
ms00f80 l0803 ( .d(n3941), .o(_net_7591), .ck(clk) );
ms00f80 l0804 ( .d(n3945), .o(net_369), .ck(clk) );
ms00f80 l0805 ( .d(n3949), .o(net_6819), .ck(clk) );
ms00f80 l0806 ( .d(n3953), .o(net_7185), .ck(clk) );
ms00f80 l0807 ( .d(n3957), .o(net_372), .ck(clk) );
ms00f80 l0808 ( .d(n3962), .o(net_6372), .ck(clk) );
ms00f80 l0809 ( .d(n3967), .o(_net_7510), .ck(clk) );
ms00f80 l0810 ( .d(n3972), .o(net_7537), .ck(clk) );
ms00f80 l0811 ( .d(n3976), .o(_net_6202), .ck(clk) );
ms00f80 l0812 ( .d(n3981), .o(_net_6112), .ck(clk) );
ms00f80 l0813 ( .d(n3985), .o(net_7050), .ck(clk) );
ms00f80 l0814 ( .d(n3989), .o(net_309), .ck(clk) );
ms00f80 l0815 ( .d(n3993), .o(net_7165), .ck(clk) );
ms00f80 l0816 ( .d(n3998), .o(_net_7095), .ck(clk) );
ms00f80 l0817 ( .d(n4002), .o(net_6949), .ck(clk) );
ms00f80 l0818 ( .d(n4007), .o(net_6852), .ck(clk) );
ms00f80 l0819 ( .d(n4011), .o(net_6279), .ck(clk) );
ms00f80 l0820 ( .d(n4016), .o(_net_7733), .ck(clk) );
ms00f80 l0821 ( .d(n4020), .o(net_6810), .ck(clk) );
ms00f80 l0822 ( .d(n4024), .o(net_141), .ck(clk) );
ms00f80 l0823 ( .d(n4029), .o(_net_7601), .ck(clk) );
ms00f80 l0824 ( .d(n4033), .o(net_7191), .ck(clk) );
ms00f80 l0825 ( .d(n4037), .o(net_6790), .ck(clk) );
ms00f80 l0826 ( .d(n4042), .o(_net_7633), .ck(clk) );
ms00f80 l0827 ( .d(n4046), .o(net_355), .ck(clk) );
ms00f80 l0828 ( .d(n4051), .o(net_6613), .ck(clk) );
ms00f80 l0829 ( .d(n4055), .o(net_7711), .ck(clk) );
ms00f80 l0830 ( .d(n4059), .o(net_7013), .ck(clk) );
ms00f80 l0831 ( .d(n4063), .o(_net_7329), .ck(clk) );
ms00f80 l0832 ( .d(n4068), .o(net_6444), .ck(clk) );
ms00f80 l0833 ( .d(n4071), .o(net_6541), .ck(clk) );
ms00f80 l0834 ( .d(n4075), .o(net_364), .ck(clk) );
ms00f80 l0835 ( .d(n4079), .o(net_7636), .ck(clk) );
ms00f80 l0836 ( .d(n4084), .o(_net_294), .ck(clk) );
ms00f80 l0837 ( .d(n4089), .o(_net_6411), .ck(clk) );
ms00f80 l0838 ( .d(n4094), .o(_net_7404), .ck(clk) );
ms00f80 l0839 ( .d(n4098), .o(net_6493), .ck(clk) );
ms00f80 l0840 ( .d(n4102), .o(net_6778), .ck(clk) );
ms00f80 l0841 ( .d(n4107), .o(_net_7719), .ck(clk) );
ms00f80 l0842 ( .d(n4112), .o(net_6867), .ck(clk) );
ms00f80 l0843 ( .d(n4116), .o(_net_7364), .ck(clk) );
ms00f80 l0844 ( .d(n4121), .o(_net_276), .ck(clk) );
ms00f80 l0845 ( .d(n4126), .o(_net_7227), .ck(clk) );
ms00f80 l0846 ( .d(n4131), .o(net_7400), .ck(clk) );
ms00f80 l0847 ( .d(n4135), .o(_net_7232), .ck(clk) );
ms00f80 l0848 ( .d(n4140), .o(_net_7347), .ck(clk) );
ms00f80 l0849 ( .d(n4145), .o(net_6592), .ck(clk) );
ms00f80 l0850 ( .d(n4148), .o(net_7028), .ck(clk) );
ms00f80 l0851 ( .d(n4153), .o(_net_6239), .ck(clk) );
ms00f80 l0852 ( .d(n4158), .o(net_6714), .ck(clk) );
ms00f80 l0853 ( .d(n4161), .o(net_367), .ck(clk) );
ms00f80 l0854 ( .d(n4166), .o(_net_7437), .ck(clk) );
ms00f80 l0855 ( .d(n4171), .o(_net_7784), .ck(clk) );
ms00f80 l0856 ( .d(n4176), .o(net_6263), .ck(clk) );
ms00f80 l0857 ( .d(n4181), .o(net_234), .ck(clk) );
ms00f80 l0858 ( .d(n4186), .o(_net_7321), .ck(clk) );
ms00f80 l0859 ( .d(n4191), .o(net_7123), .ck(clk) );
ms00f80 l0860 ( .d(n4194), .o(net_6684), .ck(clk) );
ms00f80 l0861 ( .d(n4199), .o(net_6447), .ck(clk) );
ms00f80 l0862 ( .d(n4203), .o(_net_277), .ck(clk) );
ms00f80 l0863 ( .d(n4207), .o(net_7178), .ck(clk) );
ms00f80 l0864 ( .d(n4212), .o(net_206), .ck(clk) );
ms00f80 l0865 ( .d(n4217), .o(_net_7630), .ck(clk) );
ms00f80 l0866 ( .d(n4221), .o(net_7049), .ck(clk) );
ms00f80 l0867 ( .d(n4226), .o(_net_5968), .ck(clk) );
ms00f80 l0868 ( .d(n4231), .o(net_5858), .ck(clk) );
ms00f80 l0869 ( .d(n4235), .o(net_6643), .ck(clk) );
ms00f80 l0870 ( .d(n4240), .o(_net_7635), .ck(clk) );
ms00f80 l0871 ( .d(n4245), .o(net_7398), .ck(clk) );
ms00f80 l0872 ( .d(n4249), .o(_net_6152), .ck(clk) );
ms00f80 l0873 ( .d(n4253), .o(net_376), .ck(clk) );
ms00f80 l0874 ( .d(n4258), .o(net_296), .ck(clk) );
ms00f80 l0875 ( .d(n4263), .o(net_7338), .ck(clk) );
ms00f80 l0876 ( .d(n4267), .o(net_7031), .ck(clk) );
ms00f80 l0877 ( .d(n4271), .o(net_312), .ck(clk) );
ms00f80 l0878 ( .d(n4276), .o(_net_5981), .ck(clk) );
ms00f80 l0879 ( .d(n4280), .o(net_6926), .ck(clk) );
ms00f80 l0880 ( .d(n4284), .o(_net_7810), .ck(clk) );
ms00f80 l0881 ( .d(n4289), .o(_net_229), .ck(clk) );
ms00f80 l0882 ( .d(n4294), .o(_net_7318), .ck(clk) );
ms00f80 l0883 ( .d(n4299), .o(_net_6128), .ck(clk) );
ms00f80 l0884 ( .d(n4304), .o(_net_7688), .ck(clk) );
ms00f80 l0885 ( .d(n4309), .o(net_6753), .ck(clk) );
ms00f80 l0886 ( .d(n4313), .o(_net_6422), .ck(clk) );
ms00f80 l0887 ( .d(n4318), .o(net_6471), .ck(clk) );
ms00f80 l0888 ( .d(n4322), .o(_net_6050), .ck(clk) );
ms00f80 l0889 ( .d(n4326), .o(net_6388), .ck(clk) );
ms00f80 l0890 ( .d(n4330), .o(net_6978), .ck(clk) );
ms00f80 l0891 ( .d(n4333), .o(net_7641), .ck(clk) );
ms00f80 l0892 ( .d(n4338), .o(net_6805), .ck(clk) );
ms00f80 l0893 ( .d(n4343), .o(net_7771), .ck(clk) );
ms00f80 l0894 ( .d(n4348), .o(_net_7505), .ck(clk) );
ms00f80 l0895 ( .d(n4352), .o(net_7646), .ck(clk) );
ms00f80 l0896 ( .d(n4357), .o(_net_6009), .ck(clk) );
ms00f80 l0897 ( .d(n4362), .o(net_6863), .ck(clk) );
ms00f80 l0898 ( .d(n4365), .o(net_6762), .ck(clk) );
ms00f80 l0899 ( .d(n4370), .o(net_6641), .ck(clk) );
ms00f80 l0900 ( .d(n4374), .o(net_6950), .ck(clk) );
ms00f80 l0901 ( .d(n4379), .o(_net_7278), .ck(clk) );
ms00f80 l0902 ( .d(n4384), .o(net_6974), .ck(clk) );
ms00f80 l0903 ( .d(n4388), .o(net_6431), .ck(clk) );
ms00f80 l0904 ( .d(n4392), .o(_net_7301), .ck(clk) );
ms00f80 l0905 ( .d(n4397), .o(net_6564), .ck(clk) );
ms00f80 l0906 ( .d(n4401), .o(net_7162), .ck(clk) );
ms00f80 l0907 ( .d(n4405), .o(_net_265), .ck(clk) );
ms00f80 l0908 ( .d(n4410), .o(net_7111), .ck(clk) );
ms00f80 l0909 ( .d(n4414), .o(_net_7718), .ck(clk) );
ms00f80 l0910 ( .d(n4419), .o(net_6347), .ck(clk) );
ms00f80 l0911 ( .d(n4424), .o(_net_6045), .ck(clk) );
ms00f80 l0912 ( .d(n4428), .o(net_7366), .ck(clk) );
ms00f80 l0913 ( .d(n4433), .o(_net_7332), .ck(clk) );
ms00f80 l0914 ( .d(n4438), .o(_net_7403), .ck(clk) );
ms00f80 l0915 ( .d(n4443), .o(_net_6206), .ck(clk) );
ms00f80 l0916 ( .d(n4448), .o(net_6886), .ck(clk) );
ms00f80 l0917 ( .d(n4451), .o(net_7374), .ck(clk) );
ms00f80 l0918 ( .d(n4456), .o(x179), .ck(clk) );
ms00f80 l0919 ( .d(n4459), .o(net_7741), .ck(clk) );
ms00f80 l0920 ( .d(n4464), .o(_net_7323), .ck(clk) );
ms00f80 l0921 ( .d(n4469), .o(net_6343), .ck(clk) );
ms00f80 l0922 ( .d(n4473), .o(net_7199), .ck(clk) );
ms00f80 l0923 ( .d(n4478), .o(net_6448), .ck(clk) );
ms00f80 l0924 ( .d(n4482), .o(_net_6148), .ck(clk) );
ms00f80 l0925 ( .d(n4487), .o(net_7129), .ck(clk) );
ms00f80 l0926 ( .d(n4491), .o(_net_6018), .ck(clk) );
ms00f80 l0927 ( .d(n4496), .o(net_389), .ck(clk) );
ms00f80 l0928 ( .d(n4501), .o(net_155), .ck(clk) );
ms00f80 l0929 ( .d(n4505), .o(net_7075), .ck(clk) );
ms00f80 l0930 ( .d(n4510), .o(_net_7469), .ck(clk) );
ms00f80 l0931 ( .d(n4515), .o(_net_6173), .ck(clk) );
ms00f80 l0932 ( .d(n4520), .o(net_246), .ck(clk) );
ms00f80 l0933 ( .d(n4524), .o(net_138), .ck(clk) );
ms00f80 l0934 ( .d(n4529), .o(_net_6189), .ck(clk) );
ms00f80 l0935 ( .d(n4534), .o(net_6195), .ck(clk) );
ms00f80 l0936 ( .d(n4539), .o(_net_6172), .ck(clk) );
ms00f80 l0937 ( .d(n4544), .o(_net_7480), .ck(clk) );
ms00f80 l0938 ( .d(n4548), .o(net_6489), .ck(clk) );
ms00f80 l0939 ( .d(n4553), .o(_net_6165), .ck(clk) );
ms00f80 l0940 ( .d(n4558), .o(net_146), .ck(clk) );
ms00f80 l0941 ( .d(n4562), .o(net_6761), .ck(clk) );
ms00f80 l0942 ( .d(n4567), .o(net_6225), .ck(clk) );
ms00f80 l0943 ( .d(n4572), .o(_net_7475), .ck(clk) );
ms00f80 l0944 ( .d(n4577), .o(net_6305), .ck(clk) );
ms00f80 l0945 ( .d(n4581), .o(net_7079), .ck(clk) );
ms00f80 l0946 ( .d(n4586), .o(_net_6297), .ck(clk) );
ms00f80 l0947 ( .d(n4591), .o(_net_7233), .ck(clk) );
ms00f80 l0948 ( .d(n4596), .o(_net_7413), .ck(clk) );
ms00f80 l0949 ( .d(n4600), .o(net_7068), .ck(clk) );
ms00f80 l0950 ( .d(n4604), .o(net_6635), .ck(clk) );
ms00f80 l0951 ( .d(n4609), .o(_net_7586), .ck(clk) );
ms00f80 l0952 ( .d(n4613), .o(net_6776), .ck(clk) );
ms00f80 l0953 ( .d(n4617), .o(net_6637), .ck(clk) );
ms00f80 l0954 ( .d(n4622), .o(net_6273), .ck(clk) );
ms00f80 l0955 ( .d(n4627), .o(_net_7346), .ck(clk) );
ms00f80 l0956 ( .d(n4631), .o(net_6786), .ck(clk) );
ms00f80 l0957 ( .d(n4636), .o(net_253), .ck(clk) );
ms00f80 l0958 ( .d(n4641), .o(_net_6064), .ck(clk) );
ms00f80 l0959 ( .d(n4646), .o(_net_7269), .ck(clk) );
ms00f80 l0960 ( .d(n4651), .o(net_6367), .ck(clk) );
ms00f80 l0961 ( .d(n4656), .o(_net_7288), .ck(clk) );
ms00f80 l0962 ( .d(n4660), .o(net_7197), .ck(clk) );
ms00f80 l0963 ( .d(n4665), .o(net_6736), .ck(clk) );
ms00f80 l0964 ( .d(n4669), .o(net_6581), .ck(clk) );
ms00f80 l0965 ( .d(n4673), .o(net_6055), .ck(clk) );
ms00f80 l0966 ( .d(n4678), .o(x744), .ck(clk) );
ms00f80 l0967 ( .d(n4681), .o(_net_7797), .ck(clk) );
ms00f80 l0968 ( .d(n4686), .o(net_378), .ck(clk) );
ms00f80 l0969 ( .d(n4690), .o(net_7370), .ck(clk) );
ms00f80 l0970 ( .d(n4694), .o(net_7493), .ck(clk) );
ms00f80 l0971 ( .d(n4699), .o(net_6993), .ck(clk) );
ms00f80 l0972 ( .d(n4703), .o(_net_7749), .ck(clk) );
ms00f80 l0973 ( .d(n4708), .o(_net_6073), .ck(clk) );
ms00f80 l0974 ( .d(n4713), .o(net_7142), .ck(clk) );
ms00f80 l0975 ( .d(n4717), .o(net_6544), .ck(clk) );
ms00f80 l0976 ( .d(n4722), .o(net_6271), .ck(clk) );
ms00f80 l0977 ( .d(n4727), .o(_net_7692), .ck(clk) );
ms00f80 l0978 ( .d(n4732), .o(_net_7286), .ck(clk) );
ms00f80 l0979 ( .d(n4737), .o(_net_7382), .ck(clk) );
ms00f80 l0980 ( .d(n4742), .o(net_6735), .ck(clk) );
ms00f80 l0981 ( .d(n4745), .o(net_6502), .ck(clk) );
ms00f80 l0982 ( .d(n4750), .o(net_6334), .ck(clk) );
ms00f80 l0983 ( .d(n4755), .o(net_6349), .ck(clk) );
ms00f80 l0984 ( .d(n4760), .o(_net_7706), .ck(clk) );
ms00f80 l0985 ( .d(n4765), .o(net_6231), .ck(clk) );
ms00f80 l0986 ( .d(n4769), .o(net_7455), .ck(clk) );
ms00f80 l0987 ( .d(n4774), .o(net_7545), .ck(clk) );
ms00f80 l0988 ( .d(n4778), .o(net_6449), .ck(clk) );
ms00f80 l0989 ( .d(n4782), .o(net_6352), .ck(clk) );
ms00f80 l0990 ( .d(n4787), .o(_net_7559), .ck(clk) );
ms00f80 l0991 ( .d(n4791), .o(net_6931), .ck(clk) );
ms00f80 l0992 ( .d(n4795), .o(net_6935), .ck(clk) );
ms00f80 l0993 ( .d(n4800), .o(_net_7452), .ck(clk) );
ms00f80 l0994 ( .d(n4805), .o(net_7014), .ck(clk) );
ms00f80 l0995 ( .d(n4809), .o(_net_7655), .ck(clk) );
ms00f80 l0996 ( .d(n4814), .o(net_7128), .ck(clk) );
ms00f80 l0997 ( .d(n4818), .o(_net_7624), .ck(clk) );
ms00f80 l0998 ( .d(n4822), .o(net_7304), .ck(clk) );
ms00f80 l0999 ( .d(n4827), .o(net_6567), .ck(clk) );
ms00f80 l1000 ( .d(n4831), .o(x234), .ck(clk) );
ms00f80 l1001 ( .d(n4834), .o(net_6650), .ck(clk) );
ms00f80 l1002 ( .d(n4838), .o(net_6509), .ck(clk) );
ms00f80 l1003 ( .d(n4843), .o(_net_6019), .ck(clk) );
ms00f80 l1004 ( .d(n4848), .o(net_6250), .ck(clk) );
ms00f80 l1005 ( .d(n4853), .o(net_6875), .ck(clk) );
ms00f80 l1006 ( .d(n4857), .o(_net_5975), .ck(clk) );
ms00f80 l1007 ( .d(n4862), .o(net_6403), .ck(clk) );
ms00f80 l1008 ( .d(n4867), .o(net_7189), .ck(clk) );
ms00f80 l1009 ( .d(n4872), .o(_net_284), .ck(clk) );
ms00f80 l1010 ( .d(n4877), .o(_net_6406), .ck(clk) );
ms00f80 l1011 ( .d(n4881), .o(net_349), .ck(clk) );
ms00f80 l1012 ( .d(n4886), .o(net_202), .ck(clk) );
ms00f80 l1013 ( .d(n4890), .o(net_7203), .ck(clk) );
ms00f80 l1014 ( .d(n4895), .o(net_7154), .ck(clk) );
ms00f80 l1015 ( .d(n4899), .o(net_6339), .ck(clk) );
ms00f80 l1016 ( .d(n4904), .o(net_7001), .ck(clk) );
ms00f80 l1017 ( .d(n4908), .o(_net_5967), .ck(clk) );
ms00f80 l1018 ( .d(n4913), .o(net_6573), .ck(clk) );
ms00f80 l1019 ( .d(n4917), .o(_net_6011), .ck(clk) );
ms00f80 l1020 ( .d(n4922), .o(_net_5970), .ck(clk) );
ms00f80 l1021 ( .d(n4927), .o(_net_7782), .ck(clk) );
ms00f80 l1022 ( .d(n4931), .o(net_6820), .ck(clk) );
ms00f80 l1023 ( .d(n4936), .o(_net_7659), .ck(clk) );
ms00f80 l1024 ( .d(n4940), .o(net_7047), .ck(clk) );
ms00f80 l1025 ( .d(n4944), .o(net_144), .ck(clk) );
ms00f80 l1026 ( .d(n4947), .o(net_7085), .ck(clk) );
ms00f80 l1027 ( .d(n4952), .o(_net_295), .ck(clk) );
ms00f80 l1028 ( .d(n4957), .o(net_6718), .ck(clk) );
ms00f80 l1029 ( .d(n4961), .o(_net_7651), .ck(clk) );
ms00f80 l1030 ( .d(n4965), .o(net_6923), .ck(clk) );
ms00f80 l1031 ( .d(n4969), .o(net_6808), .ck(clk) );
ms00f80 l1032 ( .d(n4974), .o(_net_6157), .ck(clk) );
ms00f80 l1033 ( .d(n4979), .o(net_6484), .ck(clk) );
ms00f80 l1034 ( .d(n4983), .o(net_6858), .ck(clk) );
ms00f80 l1035 ( .d(n4987), .o(_net_7571), .ck(clk) );
ms00f80 l1036 ( .d(n4992), .o(x765), .ck(clk) );
ms00f80 l1037 ( .d(n4996), .o(net_6241), .ck(clk) );
ms00f80 l1038 ( .d(n5001), .o(net_6617), .ck(clk) );
ms00f80 l1039 ( .d(n5005), .o(net_6854), .ck(clk) );
ms00f80 l1040 ( .d(n5008), .o(net_331), .ck(clk) );
ms00f80 l1041 ( .d(n5013), .o(_net_7727), .ck(clk) );
ms00f80 l1042 ( .d(n5018), .o(_net_6693), .ck(clk) );
ms00f80 l1043 ( .d(n5023), .o(net_7539), .ck(clk) );
ms00f80 l1044 ( .d(n5027), .o(net_7518), .ck(clk) );
ms00f80 l1045 ( .d(n5031), .o(net_6546), .ck(clk) );
ms00f80 l1046 ( .d(n5035), .o(net_7219), .ck(clk) );
ms00f80 l1047 ( .d(n5040), .o(_net_6034), .ck(clk) );
ms00f80 l1048 ( .d(n5045), .o(net_7399), .ck(clk) );
ms00f80 l1049 ( .d(n5048), .o(net_7614), .ck(clk) );
ms00f80 l1050 ( .d(n5053), .o(net_6970), .ck(clk) );
ms00f80 l1051 ( .d(n5056), .o(net_7376), .ck(clk) );
ms00f80 l1052 ( .d(n5061), .o(_net_7507), .ck(clk) );
ms00f80 l1053 ( .d(n5066), .o(net_6311), .ck(clk) );
ms00f80 l1054 ( .d(n5070), .o(net_6663), .ck(clk) );
ms00f80 l1055 ( .d(n5075), .o(_net_7508), .ck(clk) );
ms00f80 l1056 ( .d(n5080), .o(_net_7514), .ck(clk) );
ms00f80 l1057 ( .d(n5085), .o(net_6057), .ck(clk) );
ms00f80 l1058 ( .d(n5090), .o(net_7011), .ck(clk) );
ms00f80 l1059 ( .d(n5094), .o(_net_7433), .ck(clk) );
ms00f80 l1060 ( .d(n5098), .o(net_324), .ck(clk) );
ms00f80 l1061 ( .d(n5103), .o(x379), .ck(clk) );
ms00f80 l1062 ( .d(n5107), .o(net_208), .ck(clk) );
ms00f80 l1063 ( .d(n5112), .o(_net_6415), .ck(clk) );
ms00f80 l1064 ( .d(n5117), .o(_net_227), .ck(clk) );
ms00f80 l1065 ( .d(n5121), .o(net_308), .ck(clk) );
ms00f80 l1066 ( .d(n5126), .o(net_6589), .ck(clk) );
ms00f80 l1067 ( .d(n5130), .o(x149), .ck(clk) );
ms00f80 l1068 ( .d(n5134), .o(net_218), .ck(clk) );
ms00f80 l1069 ( .d(n5139), .o(net_6985), .ck(clk) );
ms00f80 l1070 ( .d(n5143), .o(_net_7272), .ck(clk) );
ms00f80 l1071 ( .d(n5148), .o(net_6572), .ck(clk) );
ms00f80 l1072 ( .d(n5151), .o(net_6516), .ck(clk) );
ms00f80 l1073 ( .d(n5156), .o(net_6428), .ck(clk) );
ms00f80 l1074 ( .d(n5159), .o(net_130), .ck(clk) );
ms00f80 l1075 ( .d(n5164), .o(_net_271), .ck(clk) );
ms00f80 l1076 ( .d(n5169), .o(_net_7435), .ck(clk) );
ms00f80 l1077 ( .d(n5173), .o(net_6940), .ck(clk) );
ms00f80 l1078 ( .d(n5178), .o(net_6841), .ck(clk) );
ms00f80 l1079 ( .d(n5181), .o(_net_7803), .ck(clk) );
ms00f80 l1080 ( .d(n5186), .o(net_7691), .ck(clk) );
ms00f80 l1081 ( .d(n5189), .o(net_6656), .ck(clk) );
ms00f80 l1082 ( .d(n5193), .o(net_7037), .ck(clk) );
ms00f80 l1083 ( .d(n5198), .o(_net_6084), .ck(clk) );
ms00f80 l1084 ( .d(n5202), .o(net_6506), .ck(clk) );
ms00f80 l1085 ( .d(n5207), .o(_net_7686), .ck(clk) );
ms00f80 l1086 ( .d(n5212), .o(_net_6114), .ck(clk) );
ms00f80 l1087 ( .d(n5217), .o(net_6569), .ck(clk) );
ms00f80 l1088 ( .d(n5221), .o(net_6857), .ck(clk) );
ms00f80 l1089 ( .d(n5225), .o(_net_7593), .ck(clk) );
ms00f80 l1090 ( .d(n5230), .o(_net_7422), .ck(clk) );
ms00f80 l1091 ( .d(n5234), .o(net_7176), .ck(clk) );
ms00f80 l1092 ( .d(n5239), .o(net_6487), .ck(clk) );
ms00f80 l1093 ( .d(n5242), .o(net_6676), .ck(clk) );
ms00f80 l1094 ( .d(n5246), .o(net_6897), .ck(clk) );
ms00f80 l1095 ( .d(n5251), .o(_net_7297), .ck(clk) );
ms00f80 l1096 ( .d(n5256), .o(_net_7567), .ck(clk) );
ms00f80 l1097 ( .d(n5261), .o(net_6843), .ck(clk) );
ms00f80 l1098 ( .d(n5265), .o(_net_7416), .ck(clk) );
ms00f80 l1099 ( .d(n5269), .o(net_7168), .ck(clk) );
ms00f80 l1100 ( .d(n5274), .o(_net_7292), .ck(clk) );
ms00f80 l1101 ( .d(n5279), .o(_net_7731), .ck(clk) );
ms00f80 l1102 ( .d(n5284), .o(_net_6284), .ck(clk) );
ms00f80 l1103 ( .d(n5288), .o(net_320), .ck(clk) );
ms00f80 l1104 ( .d(n5293), .o(_net_7599), .ck(clk) );
ms00f80 l1105 ( .d(n5298), .o(net_6965), .ck(clk) );
ms00f80 l1106 ( .d(n5302), .o(net_6324), .ck(clk) );
ms00f80 l1107 ( .d(n5307), .o(_net_7411), .ck(clk) );
ms00f80 l1108 ( .d(n5312), .o(net_7006), .ck(clk) );
ms00f80 l1109 ( .d(n5316), .o(net_6061), .ck(clk) );
ms00f80 l1110 ( .d(n5321), .o(_net_7684), .ck(clk) );
ms00f80 l1111 ( .d(n5326), .o(net_6844), .ck(clk) );
ms00f80 l1112 ( .d(n5330), .o(_net_7662), .ck(clk) );
ms00f80 l1113 ( .d(n5335), .o(net_7002), .ck(clk) );
ms00f80 l1114 ( .d(n5339), .o(net_6357), .ck(clk) );
ms00f80 l1115 ( .d(n5344), .o(_net_6420), .ck(clk) );
ms00f80 l1116 ( .d(n5349), .o(net_6987), .ck(clk) );
ms00f80 l1117 ( .d(n5353), .o(_net_7280), .ck(clk) );
ms00f80 l1118 ( .d(n5358), .o(net_6454), .ck(clk) );
ms00f80 l1119 ( .d(n5362), .o(net_6460), .ck(clk) );
ms00f80 l1120 ( .d(n5366), .o(net_6860), .ck(clk) );
ms00f80 l1121 ( .d(n5370), .o(_net_7657), .ck(clk) );
ms00f80 l1122 ( .d(n5375), .o(net_6237), .ck(clk) );
ms00f80 l1123 ( .d(n5380), .o(net_6729), .ck(clk) );
ms00f80 l1124 ( .d(n5383), .o(net_6816), .ck(clk) );
ms00f80 l1125 ( .d(n5388), .o(_net_6096), .ck(clk) );
ms00f80 l1126 ( .d(n5393), .o(net_7021), .ck(clk) );
ms00f80 l1127 ( .d(n5397), .o(net_159), .ck(clk) );
ms00f80 l1128 ( .d(n5402), .o(net_7151), .ck(clk) );
ms00f80 l1129 ( .d(n5406), .o(_net_7429), .ck(clk) );
ms00f80 l1130 ( .d(n5411), .o(_net_7631), .ck(clk) );
ms00f80 l1131 ( .d(n5415), .o(net_7206), .ck(clk) );
ms00f80 l1132 ( .d(n5420), .o(_net_7295), .ck(clk) );
ms00f80 l1133 ( .d(n5424), .o(net_7167), .ck(clk) );
ms00f80 l1134 ( .d(n5429), .o(_net_6030), .ck(clk) );
ms00f80 l1135 ( .d(n5433), .o(net_6766), .ck(clk) );
ms00f80 l1136 ( .d(n5437), .o(net_380), .ck(clk) );
ms00f80 l1137 ( .d(n5441), .o(net_6551), .ck(clk) );
ms00f80 l1138 ( .d(n5446), .o(_net_119), .ck(clk) );
ms00f80 l1139 ( .d(n5451), .o(net_6436), .ck(clk) );
ms00f80 l1140 ( .d(n5455), .o(_net_5987), .ck(clk) );
ms00f80 l1141 ( .d(n5460), .o(net_6251), .ck(clk) );
ms00f80 l1142 ( .d(n5464), .o(net_7335), .ck(clk) );
ms00f80 l1143 ( .d(n5469), .o(net_6610), .ck(clk) );
ms00f80 l1144 ( .d(n5472), .o(net_7610), .ck(clk) );
ms00f80 l1145 ( .d(n5477), .o(_net_7587), .ck(clk) );
ms00f80 l1146 ( .d(n5481), .o(net_6915), .ck(clk) );
ms00f80 l1147 ( .d(n5486), .o(net_390), .ck(clk) );
ms00f80 l1148 ( .d(n5490), .o(_net_7513), .ck(clk) );
ms00f80 l1149 ( .d(n5495), .o(_net_270), .ck(clk) );
ms00f80 l1150 ( .d(n5500), .o(net_6575), .ck(clk) );
ms00f80 l1151 ( .d(n5504), .o(net_7100), .ck(clk) );
ms00f80 l1152 ( .d(n5508), .o(_net_7467), .ck(clk) );
ms00f80 l1153 ( .d(n5513), .o(net_6024), .ck(clk) );
ms00f80 l1154 ( .d(n5517), .o(x390), .ck(clk) );
ms00f80 l1155 ( .d(n5521), .o(net_7018), .ck(clk) );
ms00f80 l1156 ( .d(n5525), .o(x172), .ck(clk) );
ms00f80 l1157 ( .d(n5529), .o(net_7780), .ck(clk) );
ms00f80 l1158 ( .d(n5534), .o(_net_7721), .ck(clk) );
ms00f80 l1159 ( .d(n5539), .o(net_6839), .ck(clk) );
ms00f80 l1160 ( .d(n5543), .o(_net_7577), .ck(clk) );
ms00f80 l1161 ( .d(n5547), .o(net_6670), .ck(clk) );
ms00f80 l1162 ( .d(n5552), .o(net_7528), .ck(clk) );
ms00f80 l1163 ( .d(n5556), .o(net_343), .ck(clk) );
ms00f80 l1164 ( .d(n5560), .o(net_6789), .ck(clk) );
ms00f80 l1165 ( .d(n5565), .o(_net_7430), .ck(clk) );
ms00f80 l1166 ( .d(n5570), .o(_net_7502), .ck(clk) );
ms00f80 l1167 ( .d(n5575), .o(net_6620), .ck(clk) );
ms00f80 l1168 ( .d(n5579), .o(_net_7622), .ck(clk) );
ms00f80 l1169 ( .d(n5584), .o(net_7546), .ck(clk) );
ms00f80 l1170 ( .d(n5588), .o(net_7235), .ck(clk) );
ms00f80 l1171 ( .d(n5591), .o(net_7640), .ck(clk) );
ms00f80 l1172 ( .d(n5596), .o(_net_6162), .ck(clk) );
ms00f80 l1173 ( .d(n5601), .o(_net_7420), .ck(clk) );
ms00f80 l1174 ( .d(n5606), .o(net_6368), .ck(clk) );
ms00f80 l1175 ( .d(n5610), .o(net_133), .ck(clk) );
ms00f80 l1176 ( .d(n5613), .o(net_7080), .ck(clk) );
ms00f80 l1177 ( .d(n5618), .o(net_6243), .ck(clk) );
ms00f80 l1178 ( .d(n5623), .o(_net_6138), .ck(clk) );
ms00f80 l1179 ( .d(n5628), .o(net_7647), .ck(clk) );
ms00f80 l1180 ( .d(n5633), .o(_net_7736), .ck(clk) );
ms00f80 l1181 ( .d(n5638), .o(_net_6205), .ck(clk) );
ms00f80 l1182 ( .d(n5643), .o(_net_7634), .ck(clk) );
ms00f80 l1183 ( .d(n5648), .o(net_6983), .ck(clk) );
ms00f80 l1184 ( .d(n5651), .o(net_7202), .ck(clk) );
ms00f80 l1185 ( .d(n5655), .o(net_6490), .ck(clk) );
ms00f80 l1186 ( .d(n5660), .o(net_5849), .ck(clk) );
ms00f80 l1187 ( .d(n5664), .o(net_7215), .ck(clk) );
ms00f80 l1188 ( .d(n5669), .o(_net_7380), .ck(clk) );
ms00f80 l1189 ( .d(n5674), .o(_net_7564), .ck(clk) );
ms00f80 l1190 ( .d(n5679), .o(net_6727), .ck(clk) );
ms00f80 l1191 ( .d(n5682), .o(net_7030), .ck(clk) );
ms00f80 l1192 ( .d(n5686), .o(_net_7822), .ck(clk) );
ms00f80 l1193 ( .d(n5691), .o(_net_6283), .ck(clk) );
ms00f80 l1194 ( .d(n5696), .o(net_6609), .ck(clk) );
ms00f80 l1195 ( .d(n5700), .o(net_169), .ck(clk) );
ms00f80 l1196 ( .d(n5704), .o(net_6942), .ck(clk) );
ms00f80 l1197 ( .d(n5709), .o(net_6412), .ck(clk) );
ms00f80 l1198 ( .d(n5713), .o(net_6668), .ck(clk) );
ms00f80 l1199 ( .d(n5717), .o(net_6523), .ck(clk) );
ms00f80 l1200 ( .d(n5722), .o(_net_269), .ck(clk) );
ms00f80 l1201 ( .d(n5727), .o(net_6598), .ck(clk) );
ms00f80 l1202 ( .d(n5731), .o(net_7107), .ck(clk) );
ms00f80 l1203 ( .d(n5735), .o(net_7026), .ck(clk) );
ms00f80 l1204 ( .d(n5739), .o(_net_5998), .ck(clk) );
ms00f80 l1205 ( .d(n5744), .o(net_7244), .ck(clk) );
ms00f80 l1206 ( .d(n5748), .o(_net_6825), .ck(clk) );
ms00f80 l1207 ( .d(n5753), .o(_net_6414), .ck(clk) );
ms00f80 l1208 ( .d(n5758), .o(net_6327), .ck(clk) );
ms00f80 l1209 ( .d(n5763), .o(net_6560), .ck(clk) );
ms00f80 l1210 ( .d(n5767), .o(net_6590), .ck(clk) );
ms00f80 l1211 ( .d(n5771), .o(net_6480), .ck(clk) );
ms00f80 l1212 ( .d(n5775), .o(_net_6154), .ck(clk) );
ms00f80 l1213 ( .d(n5779), .o(net_6642), .ck(clk) );
ms00f80 l1214 ( .d(n5783), .o(net_373), .ck(clk) );
ms00f80 l1215 ( .d(n5787), .o(net_6779), .ck(clk) );
ms00f80 l1216 ( .d(n5792), .o(net_7529), .ck(clk) );
ms00f80 l1217 ( .d(n5796), .o(net_6632), .ck(clk) );
ms00f80 l1218 ( .d(n5801), .o(net_7012), .ck(clk) );
ms00f80 l1219 ( .d(n5805), .o(net_6437), .ck(clk) );
ms00f80 l1220 ( .d(n5809), .o(_net_7561), .ck(clk) );
ms00f80 l1221 ( .d(n5814), .o(net_7676), .ck(clk) );
ms00f80 l1222 ( .d(n5819), .o(net_247), .ck(clk) );
ms00f80 l1223 ( .d(n5824), .o(net_7113), .ck(clk) );
ms00f80 l1224 ( .d(n5828), .o(net_164), .ck(clk) );
ms00f80 l1225 ( .d(n5833), .o(net_6878), .ck(clk) );
ms00f80 l1226 ( .d(n5836), .o(net_6934), .ck(clk) );
ms00f80 l1227 ( .d(n5840), .o(net_6925), .ck(clk) );
ms00f80 l1228 ( .d(n5845), .o(net_259), .ck(clk) );
ms00f80 l1229 ( .d(n5850), .o(_net_7734), .ck(clk) );
ms00f80 l1230 ( .d(n5855), .o(net_6416), .ck(clk) );
ms00f80 l1231 ( .d(n5860), .o(net_6479), .ck(clk) );
ms00f80 l1232 ( .d(n5864), .o(net_7102), .ck(clk) );
ms00f80 l1233 ( .d(n5867), .o(net_7306), .ck(clk) );
ms00f80 l1234 ( .d(n5872), .o(net_6340), .ck(clk) );
ms00f80 l1235 ( .d(n5876), .o(net_6954), .ck(clk) );
ms00f80 l1236 ( .d(n5881), .o(net_6720), .ck(clk) );
ms00f80 l1237 ( .d(n5885), .o(_net_5982), .ck(clk) );
ms00f80 l1238 ( .d(n5890), .o(_net_283), .ck(clk) );
ms00f80 l1239 ( .d(n5894), .o(net_356), .ck(clk) );
ms00f80 l1240 ( .d(n5899), .o(_net_7407), .ck(clk) );
ms00f80 l1241 ( .d(n5903), .o(net_7792), .ck(clk) );
ms00f80 l1242 ( .d(n5908), .o(net_6376), .ck(clk) );
ms00f80 l1243 ( .d(n5912), .o(net_6538), .ck(clk) );
ms00f80 l1244 ( .d(n5917), .o(net_6971), .ck(clk) );
ms00f80 l1245 ( .d(n5920), .o(net_6927), .ck(clk) );
ms00f80 l1246 ( .d(n5925), .o(_net_6040), .ck(clk) );
ms00f80 l1247 ( .d(n5930), .o(net_6580), .ck(clk) );
ms00f80 l1248 ( .d(n5934), .o(net_7127), .ck(clk) );
ms00f80 l1249 ( .d(n5938), .o(_net_7553), .ck(clk) );
ms00f80 l1250 ( .d(n5943), .o(net_6887), .ck(clk) );
ms00f80 l1251 ( .d(n5947), .o(net_6562), .ck(clk) );
ms00f80 l1252 ( .d(n5951), .o(net_6973), .ck(clk) );
ms00f80 l1253 ( .d(n5955), .o(net_6255), .ck(clk) );
ms00f80 l1254 ( .d(n5960), .o(_net_6006), .ck(clk) );
ms00f80 l1255 ( .d(n5964), .o(_net_7798), .ck(clk) );
ms00f80 l1256 ( .d(n5968), .o(net_7056), .ck(clk) );
ms00f80 l1257 ( .d(n5973), .o(_net_7360), .ck(clk) );
ms00f80 l1258 ( .d(n5978), .o(net_6618), .ck(clk) );
ms00f80 l1259 ( .d(n5982), .o(_net_6689), .ck(clk) );
ms00f80 l1260 ( .d(n5987), .o(_net_6410), .ck(clk) );
ms00f80 l1261 ( .d(n5992), .o(_net_7357), .ck(clk) );
ms00f80 l1262 ( .d(n5997), .o(_net_6066), .ck(clk) );
ms00f80 l1263 ( .d(n6002), .o(net_7712), .ck(clk) );
ms00f80 l1264 ( .d(n6006), .o(net_7115), .ck(clk) );
ms00f80 l1265 ( .d(n6009), .o(net_6497), .ck(clk) );
ms00f80 l1266 ( .d(n6014), .o(net_5861), .ck(clk) );
ms00f80 l1267 ( .d(n6019), .o(net_6314), .ck(clk) );
ms00f80 l1268 ( .d(n6024), .o(_net_7596), .ck(clk) );
ms00f80 l1269 ( .d(n6029), .o(_net_6081), .ck(clk) );
ms00f80 l1270 ( .d(n6034), .o(net_7125), .ck(clk) );
ms00f80 l1271 ( .d(n6038), .o(net_251), .ck(clk) );
ms00f80 l1272 ( .d(n6043), .o(net_6733), .ck(clk) );
ms00f80 l1273 ( .d(n6047), .o(net_6362), .ck(clk) );
ms00f80 l1274 ( .d(n6052), .o(_net_6132), .ck(clk) );
ms00f80 l1275 ( .d(n6056), .o(net_6802), .ck(clk) );
ms00f80 l1276 ( .d(n6061), .o(_net_7482), .ck(clk) );
ms00f80 l1277 ( .d(n6066), .o(net_6466), .ck(clk) );
ms00f80 l1278 ( .d(n6069), .o(net_6630), .ck(clk) );
ms00f80 l1279 ( .d(n6074), .o(_net_6558), .ck(clk) );
ms00f80 l1280 ( .d(n6078), .o(_net_7796), .ck(clk) );
ms00f80 l1281 ( .d(n6083), .o(net_261), .ck(clk) );
ms00f80 l1282 ( .d(n6088), .o(net_6054), .ck(clk) );
ms00f80 l1283 ( .d(n6093), .o(_net_7405), .ck(clk) );
ms00f80 l1284 ( .d(n6098), .o(net_6335), .ck(clk) );
ms00f80 l1285 ( .d(n6102), .o(net_6763), .ck(clk) );
ms00f80 l1286 ( .d(n6106), .o(net_6686), .ck(clk) );
ms00f80 l1287 ( .d(n6110), .o(net_7372), .ck(clk) );
ms00f80 l1288 ( .d(n6114), .o(net_6804), .ck(clk) );
ms00f80 l1289 ( .d(n6119), .o(_net_6181), .ck(clk) );
ms00f80 l1290 ( .d(n6124), .o(_net_7729), .ck(clk) );
ms00f80 l1291 ( .d(n6128), .o(net_7038), .ck(clk) );
ms00f80 l1292 ( .d(n6132), .o(_net_7808), .ck(clk) );
ms00f80 l1293 ( .d(n6136), .o(net_6385), .ck(clk) );
ms00f80 l1294 ( .d(n6140), .o(_net_7681), .ck(clk) );
ms00f80 l1295 ( .d(n6145), .o(net_6594), .ck(clk) );
ms00f80 l1296 ( .d(n6148), .o(net_274), .ck(clk) );
ms00f80 l1297 ( .d(n6153), .o(_net_6293), .ck(clk) );
ms00f80 l1298 ( .d(n6158), .o(net_6892), .ck(clk) );
ms00f80 l1299 ( .d(n6161), .o(net_7083), .ck(clk) );
ms00f80 l1300 ( .d(n6166), .o(_net_6209), .ck(clk) );
ms00f80 l1301 ( .d(n6171), .o(_net_6071), .ck(clk) );
ms00f80 l1302 ( .d(n6176), .o(net_6301), .ck(clk) );
ms00f80 l1303 ( .d(n6181), .o(net_6309), .ck(clk) );
ms00f80 l1304 ( .d(n6186), .o(_net_6124), .ck(clk) );
ms00f80 l1305 ( .d(n6191), .o(_net_6149), .ck(clk) );
ms00f80 l1306 ( .d(n6195), .o(net_6508), .ck(clk) );
ms00f80 l1307 ( .d(n6200), .o(_net_7693), .ck(clk) );
ms00f80 l1308 ( .d(n6204), .o(net_382), .ck(clk) );
ms00f80 l1309 ( .d(n6209), .o(_net_7254), .ck(clk) );
ms00f80 l1310 ( .d(n6214), .o(net_7385), .ck(clk) );
ms00f80 l1311 ( .d(n6218), .o(_net_6099), .ck(clk) );
ms00f80 l1312 ( .d(n6222), .o(net_7679), .ck(clk) );
ms00f80 l1313 ( .d(n6227), .o(net_186), .ck(clk) );
ms00f80 l1314 ( .d(n6231), .o(net_7739), .ck(clk) );
ms00f80 l1315 ( .d(n6235), .o(net_6629), .ck(clk) );
ms00f80 l1316 ( .d(n6239), .o(net_385), .ck(clk) );
ms00f80 l1317 ( .d(n6244), .o(_net_210), .ck(clk) );
ms00f80 l1318 ( .d(n6249), .o(_net_201), .ck(clk) );
ms00f80 l1319 ( .d(n6254), .o(net_6697), .ck(clk) );
ms00f80 l1320 ( .d(n6258), .o(net_6750), .ck(clk) );
ms00f80 l1321 ( .d(n6261), .o(_net_7801), .ck(clk) );
ms00f80 l1322 ( .d(n6266), .o(_net_7434), .ck(clk) );
ms00f80 l1323 ( .d(n6271), .o(net_167), .ck(clk) );
ms00f80 l1324 ( .d(n6276), .o(net_7752), .ck(clk) );
ms00f80 l1325 ( .d(n6281), .o(_net_174), .ck(clk) );
ms00f80 l1326 ( .d(n6285), .o(net_6212), .ck(clk) );
ms00f80 l1327 ( .d(n6290), .o(x718), .ck(clk) );
ms00f80 l1328 ( .d(n6294), .o(_net_7789), .ck(clk) );
ms00f80 l1329 ( .d(n6299), .o(net_7130), .ck(clk) );
ms00f80 l1330 ( .d(n6302), .o(net_7454), .ck(clk) );
ms00f80 l1331 ( .d(n6306), .o(net_302), .ck(clk) );
ms00f80 l1332 ( .d(n6311), .o(_net_5994), .ck(clk) );
ms00f80 l1333 ( .d(n6316), .o(net_7770), .ck(clk) );
ms00f80 l1334 ( .d(n6319), .o(_net_5922), .ck(clk) );
ms00f80 l1335 ( .d(n6324), .o(_net_6001), .ck(clk) );
ms00f80 l1336 ( .d(n6329), .o(net_7161), .ck(clk) );
ms00f80 l1337 ( .d(n6332), .o(net_381), .ck(clk) );
ms00f80 l1338 ( .d(n6337), .o(_net_6074), .ck(clk) );
ms00f80 l1339 ( .d(n6342), .o(net_6469), .ck(clk) );
ms00f80 l1340 ( .d(n6346), .o(_net_7353), .ck(clk) );
ms00f80 l1341 ( .d(n6350), .o(net_131), .ck(clk) );
ms00f80 l1342 ( .d(n6354), .o(net_6747), .ck(clk) );
ms00f80 l1343 ( .d(n6357), .o(net_6679), .ck(clk) );
ms00f80 l1344 ( .d(n6362), .o(_net_7440), .ck(clk) );
ms00f80 l1345 ( .d(n6367), .o(net_6439), .ck(clk) );
ms00f80 l1346 ( .d(n6371), .o(_net_7098), .ck(clk) );
ms00f80 l1347 ( .d(n6376), .o(net_7341), .ck(clk) );
ms00f80 l1348 ( .d(n6381), .o(_net_7661), .ck(clk) );
ms00f80 l1349 ( .d(n6386), .o(net_7117), .ck(clk) );
ms00f80 l1350 ( .d(n6390), .o(net_6361), .ck(clk) );
ms00f80 l1351 ( .d(n6395), .o(_net_6101), .ck(clk) );
ms00f80 l1352 ( .d(n6399), .o(net_6399), .ck(clk) );
ms00f80 l1353 ( .d(n6403), .o(net_6738), .ck(clk) );
ms00f80 l1354 ( .d(n6407), .o(net_6481), .ck(clk) );
ms00f80 l1355 ( .d(n6411), .o(_net_7438), .ck(clk) );
ms00f80 l1356 ( .d(n6415), .o(net_7208), .ck(clk) );
ms00f80 l1357 ( .d(n6419), .o(net_6625), .ck(clk) );
ms00f80 l1358 ( .d(n6423), .o(net_6383), .ck(clk) );
ms00f80 l1359 ( .d(n6427), .o(net_6826), .ck(clk) );
ms00f80 l1360 ( .d(n6432), .o(net_156), .ck(clk) );
ms00f80 l1361 ( .d(n6437), .o(net_7462), .ck(clk) );
ms00f80 l1362 ( .d(n6441), .o(net_7069), .ck(clk) );
ms00f80 l1363 ( .d(n6446), .o(net_6702), .ck(clk) );
ms00f80 l1364 ( .d(n6450), .o(_net_6692), .ck(clk) );
ms00f80 l1365 ( .d(n6455), .o(_net_7257), .ck(clk) );
ms00f80 l1366 ( .d(n6460), .o(net_6348), .ck(clk) );
ms00f80 l1367 ( .d(n6464), .o(net_6647), .ck(clk) );
ms00f80 l1368 ( .d(n6469), .o(net_6980), .ck(clk) );
ms00f80 l1369 ( .d(n6472), .o(net_6777), .ck(clk) );
ms00f80 l1370 ( .d(n6477), .o(net_7148), .ck(clk) );
ms00f80 l1371 ( .d(n6480), .o(net_6626), .ck(clk) );
ms00f80 l1372 ( .d(n6485), .o(net_6462), .ck(clk) );
ms00f80 l1373 ( .d(n6489), .o(net_7242), .ck(clk) );
ms00f80 l1374 ( .d(n6493), .o(net_205), .ck(clk) );
ms00f80 l1375 ( .d(n6498), .o(net_6355), .ck(clk) );
ms00f80 l1376 ( .d(n6502), .o(net_7074), .ck(clk) );
ms00f80 l1377 ( .d(n6507), .o(net_6563), .ck(clk) );
ms00f80 l1378 ( .d(n6511), .o(net_6604), .ck(clk) );
ms00f80 l1379 ( .d(n6515), .o(net_6836), .ck(clk) );
ms00f80 l1380 ( .d(n6519), .o(net_6866), .ck(clk) );
ms00f80 l1381 ( .d(n6522), .o(_net_7805), .ck(clk) );
ms00f80 l1382 ( .d(n6527), .o(_net_5857), .ck(clk) );
ms00f80 l1383 ( .d(n6531), .o(net_330), .ck(clk) );
ms00f80 l1384 ( .d(n6535), .o(net_7606), .ck(clk) );
ms00f80 l1385 ( .d(n6540), .o(_net_6126), .ck(clk) );
ms00f80 l1386 ( .d(n6545), .o(_net_118), .ck(clk) );
ms00f80 l1387 ( .d(n6550), .o(net_7397), .ck(clk) );
ms00f80 l1388 ( .d(n6554), .o(net_6713), .ck(clk) );
ms00f80 l1389 ( .d(n6558), .o(_net_7654), .ck(clk) );
ms00f80 l1390 ( .d(n6563), .o(net_6846), .ck(clk) );
ms00f80 l1391 ( .d(n6566), .o(net_6382), .ck(clk) );
ms00f80 l1392 ( .d(n6570), .o(_net_6146), .ck(clk) );
ms00f80 l1393 ( .d(n6574), .o(net_7485), .ck(clk) );
ms00f80 l1394 ( .d(n6578), .o(net_6226), .ck(clk) );
ms00f80 l1395 ( .d(n6583), .o(net_386), .ck(clk) );
ms00f80 l1396 ( .d(n6586), .o(net_6814), .ck(clk) );
ms00f80 l1397 ( .d(n6591), .o(net_157), .ck(clk) );
ms00f80 l1398 ( .d(n6596), .o(_net_6119), .ck(clk) );
ms00f80 l1399 ( .d(n6601), .o(_net_7448), .ck(clk) );
ms00f80 l1400 ( .d(n6606), .o(_net_5976), .ck(clk) );
ms00f80 l1401 ( .d(n6611), .o(net_6272), .ck(clk) );
ms00f80 l1402 ( .d(n6615), .o(net_6917), .ck(clk) );
ms00f80 l1403 ( .d(n6619), .o(net_7163), .ck(clk) );
ms00f80 l1404 ( .d(n6624), .o(net_168), .ck(clk) );
ms00f80 l1405 ( .d(n6629), .o(net_6261), .ck(clk) );
ms00f80 l1406 ( .d(n6634), .o(_net_6170), .ck(clk) );
ms00f80 l1407 ( .d(n6638), .o(net_7187), .ck(clk) );
ms00f80 l1408 ( .d(n6643), .o(net_6003), .ck(clk) );
ms00f80 l1409 ( .d(n6648), .o(net_7145), .ck(clk) );
ms00f80 l1410 ( .d(n6652), .o(_net_124), .ck(clk) );
ms00f80 l1411 ( .d(n6656), .o(net_7638), .ck(clk) );
ms00f80 l1412 ( .d(n6661), .o(net_6424), .ck(clk) );
ms00f80 l1413 ( .d(n6665), .o(_net_6129), .ck(clk) );
ms00f80 l1414 ( .d(n6669), .o(net_315), .ck(clk) );
ms00f80 l1415 ( .d(n6674), .o(net_6834), .ck(clk) );
ms00f80 l1416 ( .d(n6678), .o(net_6708), .ck(clk) );
ms00f80 l1417 ( .d(n6682), .o(_net_278), .ck(clk) );
ms00f80 l1418 ( .d(n6687), .o(net_6997), .ck(clk) );
ms00f80 l1419 ( .d(n6691), .o(x681), .ck(clk) );
ms00f80 l1420 ( .d(n6695), .o(_net_7623), .ck(clk) );
ms00f80 l1421 ( .d(n6700), .o(net_6353), .ck(clk) );
ms00f80 l1422 ( .d(n6704), .o(net_7029), .ck(clk) );
ms00f80 l1423 ( .d(n6709), .o(_net_7279), .ck(clk) );
ms00f80 l1424 ( .d(n6713), .o(net_6655), .ck(clk) );
ms00f80 l1425 ( .d(n6717), .o(net_6793), .ck(clk) );
ms00f80 l1426 ( .d(n6722), .o(net_7345), .ck(clk) );
ms00f80 l1427 ( .d(n6727), .o(_net_6113), .ck(clk) );
ms00f80 l1428 ( .d(n6732), .o(net_7180), .ck(clk) );
ms00f80 l1429 ( .d(n6736), .o(net_136), .ck(clk) );
ms00f80 l1430 ( .d(n6741), .o(_net_7620), .ck(clk) );
ms00f80 l1431 ( .d(n6746), .o(net_7549), .ck(clk) );
ms00f80 l1432 ( .d(n6749), .o(net_147), .ck(clk) );
ms00f80 l1433 ( .d(n6752), .o(net_6894), .ck(clk) );
ms00f80 l1434 ( .d(n6756), .o(net_314), .ck(clk) );
ms00f80 l1435 ( .d(n6761), .o(net_6728), .ck(clk) );
ms00f80 l1436 ( .d(n6765), .o(_net_6136), .ck(clk) );
ms00f80 l1437 ( .d(n6770), .o(net_6830), .ck(clk) );
ms00f80 l1438 ( .d(n6774), .o(_net_6117), .ck(clk) );
ms00f80 l1439 ( .d(n6779), .o(_net_7723), .ck(clk) );
ms00f80 l1440 ( .d(n6783), .o(net_6519), .ck(clk) );
ms00f80 l1441 ( .d(n6788), .o(_net_7446), .ck(clk) );
ms00f80 l1442 ( .d(n6793), .o(net_7394), .ck(clk) );
ms00f80 l1443 ( .d(n6796), .o(net_6933), .ck(clk) );
ms00f80 l1444 ( .d(n6801), .o(_net_7258), .ck(clk) );
ms00f80 l1445 ( .d(n6806), .o(net_6990), .ck(clk) );
ms00f80 l1446 ( .d(n6809), .o(net_6526), .ck(clk) );
ms00f80 l1447 ( .d(n6813), .o(net_7033), .ck(clk) );
ms00f80 l1448 ( .d(n6818), .o(_net_7700), .ck(clk) );
ms00f80 l1449 ( .d(n6822), .o(net_301), .ck(clk) );
ms00f80 l1450 ( .d(n6826), .o(net_7044), .ck(clk) );
ms00f80 l1451 ( .d(n6831), .o(_net_7584), .ck(clk) );
ms00f80 l1452 ( .d(n6836), .o(net_7025), .ck(clk) );
ms00f80 l1453 ( .d(n6840), .o(_net_5993), .ck(clk) );
ms00f80 l1454 ( .d(n6845), .o(_net_7325), .ck(clk) );
ms00f80 l1455 ( .d(n6850), .o(net_240), .ck(clk) );
ms00f80 l1456 ( .d(n6855), .o(_net_5990), .ck(clk) );
ms00f80 l1457 ( .d(n6860), .o(net_6470), .ck(clk) );
ms00f80 l1458 ( .d(n6863), .o(net_7166), .ck(clk) );
ms00f80 l1459 ( .d(n6867), .o(net_7193), .ck(clk) );
ms00f80 l1460 ( .d(n6872), .o(net_216), .ck(clk) );
ms00f80 l1461 ( .d(n6876), .o(net_7209), .ck(clk) );
ms00f80 l1462 ( .d(n6881), .o(_net_6161), .ck(clk) );
ms00f80 l1463 ( .d(n6886), .o(net_6712), .ck(clk) );
ms00f80 l1464 ( .d(n6890), .o(_net_7427), .ck(clk) );
ms00f80 l1465 ( .d(n6895), .o(net_7009), .ck(clk) );
ms00f80 l1466 ( .d(n6899), .o(net_6607), .ck(clk) );
ms00f80 l1467 ( .d(n6902), .o(net_340), .ck(clk) );
ms00f80 l1468 ( .d(n6906), .o(net_6904), .ck(clk) );
ms00f80 l1469 ( .d(n6910), .o(net_7053), .ck(clk) );
ms00f80 l1470 ( .d(n6915), .o(_net_215), .ck(clk) );
ms00f80 l1471 ( .d(n6919), .o(net_7309), .ck(clk) );
ms00f80 l1472 ( .d(n6924), .o(_net_7443), .ck(clk) );
ms00f80 l1473 ( .d(n6929), .o(net_244), .ck(clk) );
ms00f80 l1474 ( .d(n6934), .o(net_7150), .ck(clk) );
ms00f80 l1475 ( .d(n6938), .o(_net_114), .ck(clk) );
ms00f80 l1476 ( .d(n6943), .o(_net_7589), .ck(clk) );
ms00f80 l1477 ( .d(n6947), .o(net_375), .ck(clk) );
ms00f80 l1478 ( .d(n6952), .o(_net_7500), .ck(clk) );
ms00f80 l1479 ( .d(n6957), .o(net_6587), .ck(clk) );
ms00f80 l1480 ( .d(n6960), .o(net_149), .ck(clk) );
ms00f80 l1481 ( .d(n6964), .o(_net_6098), .ck(clk) );
ms00f80 l1482 ( .d(n6969), .o(net_194), .ck(clk) );
ms00f80 l1483 ( .d(n6974), .o(net_7245), .ck(clk) );
ms00f80 l1484 ( .d(n6977), .o(net_7051), .ck(clk) );
ms00f80 l1485 ( .d(n6982), .o(net_6342), .ck(clk) );
ms00f80 l1486 ( .d(n6986), .o(net_7172), .ck(clk) );
ms00f80 l1487 ( .d(n6990), .o(net_6495), .ck(clk) );
ms00f80 l1488 ( .d(n6995), .o(_net_7256), .ck(clk) );
ms00f80 l1489 ( .d(n7000), .o(_net_281), .ck(clk) );
ms00f80 l1490 ( .d(n7005), .o(net_6621), .ck(clk) );
ms00f80 l1491 ( .d(n7009), .o(net_6597), .ck(clk) );
ms00f80 l1492 ( .d(n7013), .o(_net_7408), .ck(clk) );
ms00f80 l1493 ( .d(n7018), .o(_net_6140), .ck(clk) );
ms00f80 l1494 ( .d(n7023), .o(net_222), .ck(clk) );
ms00f80 l1495 ( .d(n7027), .o(net_6902), .ck(clk) );
ms00f80 l1496 ( .d(n7032), .o(_net_7298), .ck(clk) );
ms00f80 l1497 ( .d(n7036), .o(net_306), .ck(clk) );
ms00f80 l1498 ( .d(n7041), .o(net_6889), .ck(clk) );
ms00f80 l1499 ( .d(n7045), .o(net_6378), .ck(clk) );
ms00f80 l1500 ( .d(n7049), .o(net_6394), .ck(clk) );
ms00f80 l1501 ( .d(n7053), .o(_net_7579), .ck(clk) );
ms00f80 l1502 ( .d(n7058), .o(_net_7268), .ck(clk) );
ms00f80 l1503 ( .d(n7062), .o(net_6769), .ck(clk) );
ms00f80 l1504 ( .d(n7067), .o(_net_6122), .ck(clk) );
ms00f80 l1505 ( .d(n7072), .o(_net_7761), .ck(clk) );
ms00f80 l1506 ( .d(n7077), .o(_net_6285), .ck(clk) );
ms00f80 l1507 ( .d(n7082), .o(net_6872), .ck(clk) );
ms00f80 l1508 ( .d(n7085), .o(net_7460), .ck(clk) );
ms00f80 l1509 ( .d(n7089), .o(net_6673), .ck(clk) );
ms00f80 l1510 ( .d(n7093), .o(net_383), .ck(clk) );
ms00f80 l1511 ( .d(n7098), .o(net_7152), .ck(clk) );
ms00f80 l1512 ( .d(n7102), .o(_net_193), .ck(clk) );
ms00f80 l1513 ( .d(n7107), .o(net_7769), .ck(clk) );
ms00f80 l1514 ( .d(n7111), .o(net_7088), .ck(clk) );
ms00f80 l1515 ( .d(n7116), .o(net_6329), .ck(clk) );
ms00f80 l1516 ( .d(n7120), .o(net_6498), .ck(clk) );
ms00f80 l1517 ( .d(n7125), .o(net_6561), .ck(clk) );
ms00f80 l1518 ( .d(n7128), .o(net_6660), .ck(clk) );
ms00f80 l1519 ( .d(n7133), .o(_net_7705), .ck(clk) );
ms00f80 l1520 ( .d(n7138), .o(_net_5848), .ck(clk) );
ms00f80 l1521 ( .d(n7142), .o(net_7496), .ck(clk) );
ms00f80 l1522 ( .d(n7147), .o(net_6249), .ck(clk) );
ms00f80 l1523 ( .d(n7151), .o(net_6948), .ck(clk) );
ms00f80 l1524 ( .d(n7155), .o(net_7226), .ck(clk) );
ms00f80 l1525 ( .d(n7160), .o(net_6862), .ck(clk) );
ms00f80 l1526 ( .d(n7164), .o(x195), .ck(clk) );
ms00f80 l1527 ( .d(n7167), .o(net_6235), .ck(clk) );
ms00f80 l1528 ( .d(n7172), .o(_net_5979), .ck(clk) );
ms00f80 l1529 ( .d(n7177), .o(net_161), .ck(clk) );
ms00f80 l1530 ( .d(n7182), .o(net_7543), .ck(clk) );
ms00f80 l1531 ( .d(n7185), .o(net_7307), .ck(clk) );
ms00f80 l1532 ( .d(n7190), .o(net_6430), .ck(clk) );
ms00f80 l1533 ( .d(n7194), .o(_net_6554), .ck(clk) );
ms00f80 l1534 ( .d(n7199), .o(net_7238), .ck(clk) );
ms00f80 l1535 ( .d(n7203), .o(net_6477), .ck(clk) );
ms00f80 l1536 ( .d(n7207), .o(_net_6080), .ck(clk) );
ms00f80 l1537 ( .d(n7212), .o(net_6559), .ck(clk) );
ms00f80 l1538 ( .d(n7216), .o(_net_7361), .ck(clk) );
ms00f80 l1539 ( .d(n7221), .o(net_6211), .ck(clk) );
ms00f80 l1540 ( .d(n7226), .o(_net_6200), .ck(clk) );
ms00f80 l1541 ( .d(n7230), .o(net_7090), .ck(clk) );
ms00f80 l1542 ( .d(n7235), .o(_net_6295), .ck(clk) );
ms00f80 l1543 ( .d(n7240), .o(_net_6145), .ck(clk) );
ms00f80 l1544 ( .d(n7245), .o(_net_6423), .ck(clk) );
ms00f80 l1545 ( .d(n7249), .o(net_7807), .ck(clk) );
ms00f80 l1546 ( .d(n7252), .o(net_6801), .ck(clk) );
ms00f80 l1547 ( .d(n7256), .o(_net_7791), .ck(clk) );
ms00f80 l1548 ( .d(n7260), .o(net_6627), .ck(clk) );
ms00f80 l1549 ( .d(n7265), .o(_net_6402), .ck(clk) );
ms00f80 l1550 ( .d(n7270), .o(_net_6151), .ck(clk) );
ms00f80 l1551 ( .d(n7275), .o(_net_6291), .ck(clk) );
ms00f80 l1552 ( .d(n7280), .o(_net_6026), .ck(clk) );
ms00f80 l1553 ( .d(n7284), .o(net_6511), .ck(clk) );
ms00f80 l1554 ( .d(n7288), .o(net_342), .ck(clk) );
ms00f80 l1555 ( .d(n7292), .o(_net_7816), .ck(clk) );
ms00f80 l1556 ( .d(n7297), .o(_net_6028), .ck(clk) );
ms00f80 l1557 ( .d(n7302), .o(_net_6288), .ck(clk) );
ms00f80 l1558 ( .d(n7307), .o(_net_7697), .ck(clk) );
ms00f80 l1559 ( .d(n7312), .o(net_6869), .ck(clk) );
ms00f80 l1560 ( .d(n7316), .o(net_6374), .ck(clk) );
ms00f80 l1561 ( .d(n7321), .o(_net_7365), .ck(clk) );
ms00f80 l1562 ( .d(n7326), .o(net_6715), .ck(clk) );
ms00f80 l1563 ( .d(n7330), .o(net_6264), .ck(clk) );
ms00f80 l1564 ( .d(n7335), .o(net_5860), .ck(clk) );
ms00f80 l1565 ( .d(n7340), .o(_net_6179), .ck(clk) );
ms00f80 l1566 ( .d(n7344), .o(net_7173), .ck(clk) );
ms00f80 l1567 ( .d(n7349), .o(net_6193), .ck(clk) );
ms00f80 l1568 ( .d(n7354), .o(net_250), .ck(clk) );
ms00f80 l1569 ( .d(n7359), .o(net_7008), .ck(clk) );
ms00f80 l1570 ( .d(n7363), .o(net_185), .ck(clk) );
ms00f80 l1571 ( .d(n7368), .o(net_6317), .ck(clk) );
ms00f80 l1572 ( .d(n7372), .o(net_7065), .ck(clk) );
ms00f80 l1573 ( .d(n7376), .o(net_6228), .ck(clk) );
ms00f80 l1574 ( .d(n7381), .o(_net_7666), .ck(clk) );
ms00f80 l1575 ( .d(n7386), .o(_net_6105), .ck(clk) );
ms00f80 l1576 ( .d(n7391), .o(net_7118), .ck(clk) );
ms00f80 l1577 ( .d(n7395), .o(_net_117), .ck(clk) );
ms00f80 l1578 ( .d(n7400), .o(_net_7473), .ck(clk) );
ms00f80 l1579 ( .d(n7404), .o(net_6503), .ck(clk) );
ms00f80 l1580 ( .d(n7408), .o(net_7054), .ck(clk) );
ms00f80 l1581 ( .d(n7413), .o(net_6994), .ck(clk) );
ms00f80 l1582 ( .d(n7417), .o(net_6257), .ck(clk) );
ms00f80 l1583 ( .d(n7422), .o(_net_6957), .ck(clk) );
ms00f80 l1584 ( .d(n7427), .o(net_6345), .ck(clk) );
ms00f80 l1585 ( .d(n7432), .o(_net_7757), .ck(clk) );
ms00f80 l1586 ( .d(n7437), .o(_net_6069), .ck(clk) );
ms00f80 l1587 ( .d(n7442), .o(net_6700), .ck(clk) );
ms00f80 l1588 ( .d(n7446), .o(net_6696), .ck(clk) );
ms00f80 l1589 ( .d(n7450), .o(net_6740), .ck(clk) );
ms00f80 l1590 ( .d(n7454), .o(_net_6007), .ck(clk) );
ms00f80 l1591 ( .d(n7459), .o(_net_7263), .ck(clk) );
ms00f80 l1592 ( .d(n7463), .o(net_7216), .ck(clk) );
ms00f80 l1593 ( .d(n7468), .o(net_6337), .ck(clk) );
ms00f80 l1594 ( .d(n7473), .o(_net_6222), .ck(clk) );
ms00f80 l1595 ( .d(n7478), .o(_net_7351), .ck(clk) );
ms00f80 l1596 ( .d(n7482), .o(net_7077), .ck(clk) );
ms00f80 l1597 ( .d(n7487), .o(_net_6962), .ck(clk) );
ms00f80 l1598 ( .d(n7492), .o(net_6726), .ck(clk) );
ms00f80 l1599 ( .d(n7496), .o(_net_6068), .ck(clk) );
ms00f80 l1600 ( .d(n7501), .o(_net_264), .ck(clk) );
ms00f80 l1601 ( .d(n7505), .o(net_348), .ck(clk) );
ms00f80 l1602 ( .d(n7509), .o(net_6774), .ck(clk) );
ms00f80 l1603 ( .d(n7513), .o(net_6550), .ck(clk) );
ms00f80 l1604 ( .d(n7518), .o(_net_7471), .ck(clk) );
ms00f80 l1605 ( .d(n7522), .o(net_7211), .ck(clk) );
ms00f80 l1606 ( .d(n7527), .o(net_6451), .ck(clk) );
ms00f80 l1607 ( .d(n7530), .o(net_7210), .ck(clk) );
ms00f80 l1608 ( .d(n7535), .o(net_6757), .ck(clk) );
ms00f80 l1609 ( .d(n7539), .o(x476), .ck(clk) );
ms00f80 l1610 ( .d(n7543), .o(_net_177), .ck(clk) );
ms00f80 l1611 ( .d(n7548), .o(net_243), .ck(clk) );
ms00f80 l1612 ( .d(n7553), .o(net_6266), .ck(clk) );
ms00f80 l1613 ( .d(n7558), .o(_net_7381), .ck(clk) );
ms00f80 l1614 ( .d(n7563), .o(_net_7293), .ck(clk) );
ms00f80 l1615 ( .d(n7567), .o(_net_7824), .ck(clk) );
ms00f80 l1616 ( .d(n7572), .o(_net_6127), .ck(clk) );
ms00f80 l1617 ( .d(n7577), .o(_net_6319), .ck(clk) );
ms00f80 l1618 ( .d(n7581), .o(net_6811), .ck(clk) );
ms00f80 l1619 ( .d(n7586), .o(_net_6033), .ck(clk) );
ms00f80 l1620 ( .d(n7591), .o(_net_127), .ck(clk) );
ms00f80 l1621 ( .d(n7596), .o(x187), .ck(clk) );
ms00f80 l1622 ( .d(n7599), .o(net_7494), .ck(clk) );
ms00f80 l1623 ( .d(n7604), .o(net_6716), .ck(clk) );
ms00f80 l1624 ( .d(n7608), .o(_net_6959), .ck(clk) );
ms00f80 l1625 ( .d(n7613), .o(net_199), .ck(clk) );
ms00f80 l1626 ( .d(n7618), .o(net_7392), .ck(clk) );
ms00f80 l1627 ( .d(n7622), .o(_net_6207), .ck(clk) );
ms00f80 l1628 ( .d(n7626), .o(net_7489), .ck(clk) );
ms00f80 l1629 ( .d(n7631), .o(_net_7331), .ck(clk) );
ms00f80 l1630 ( .d(n7635), .o(net_7668), .ck(clk) );
ms00f80 l1631 ( .d(n7640), .o(_net_5999), .ck(clk) );
ms00f80 l1632 ( .d(n7644), .o(net_341), .ck(clk) );
ms00f80 l1633 ( .d(n7649), .o(net_6299), .ck(clk) );
ms00f80 l1634 ( .d(n7654), .o(net_7139), .ck(clk) );
ms00f80 l1635 ( .d(n7658), .o(net_6467), .ck(clk) );
ms00f80 l1636 ( .d(n7661), .o(net_7486), .ck(clk) );
ms00f80 l1637 ( .d(n7666), .o(_net_7228), .ck(clk) );
ms00f80 l1638 ( .d(n7671), .o(_net_6091), .ck(clk) );
ms00f80 l1639 ( .d(n7676), .o(_net_6103), .ck(clk) );
ms00f80 l1640 ( .d(n7681), .o(_net_125), .ck(clk) );
ms00f80 l1641 ( .d(n7686), .o(net_231), .ck(clk) );
ms00f80 l1642 ( .d(n7691), .o(x38), .ck(clk) );
ms00f80 l1643 ( .d(n7695), .o(_net_5995), .ck(clk) );
ms00f80 l1644 ( .d(n7700), .o(net_6748), .ck(clk) );
ms00f80 l1645 ( .d(n7704), .o(net_6304), .ck(clk) );
ms00f80 l1646 ( .d(n7709), .o(net_6047), .ck(clk) );
ms00f80 l1647 ( .d(n7714), .o(net_7764), .ck(clk) );
ms00f80 l1648 ( .d(n7719), .o(net_6837), .ck(clk) );
ms00f80 l1649 ( .d(n7723), .o(_net_7273), .ck(clk) );
ms00f80 l1650 ( .d(n7728), .o(_net_7289), .ck(clk) );
ms00f80 l1651 ( .d(n7732), .o(net_7526), .ck(clk) );
ms00f80 l1652 ( .d(n7737), .o(x522), .ck(clk) );
ms00f80 l1653 ( .d(n7741), .o(_net_392), .ck(clk) );
ms00f80 l1654 ( .d(n7746), .o(_net_6828), .ck(clk) );
ms00f80 l1655 ( .d(n7751), .o(_net_7555), .ck(clk) );
ms00f80 l1656 ( .d(n7756), .o(net_6441), .ck(clk) );
ms00f80 l1657 ( .d(n7760), .o(net_7143), .ck(clk) );
ms00f80 l1658 ( .d(n7764), .o(net_7160), .ck(clk) );
ms00f80 l1659 ( .d(n7768), .o(_net_7699), .ck(clk) );
ms00f80 l1660 ( .d(n7773), .o(x420), .ck(clk) );
ms00f80 l1661 ( .d(n7776), .o(net_6397), .ck(clk) );
ms00f80 l1662 ( .d(n7779), .o(net_7059), .ck(clk) );
ms00f80 l1663 ( .d(n7784), .o(net_6710), .ck(clk) );
ms00f80 l1664 ( .d(n7788), .o(_net_6093), .ck(clk) );
ms00f80 l1665 ( .d(n7793), .o(_net_6049), .ck(clk) );
ms00f80 l1666 ( .d(n7798), .o(_net_7442), .ck(clk) );
ms00f80 l1667 ( .d(n7802), .o(net_6797), .ck(clk) );
ms00f80 l1668 ( .d(n7806), .o(net_6947), .ck(clk) );
ms00f80 l1669 ( .d(n7810), .o(net_6659), .ck(clk) );
ms00f80 l1670 ( .d(n7815), .o(net_6734), .ck(clk) );
ms00f80 l1671 ( .d(n7818), .o(net_6387), .ck(clk) );
ms00f80 l1672 ( .d(n7822), .o(_net_5974), .ck(clk) );
ms00f80 l1673 ( .d(n7826), .o(net_6528), .ck(clk) );
ms00f80 l1674 ( .d(n7831), .o(net_6566), .ck(clk) );
ms00f80 l1675 ( .d(n7835), .o(_net_7276), .ck(clk) );
ms00f80 l1676 ( .d(n7840), .o(net_6331), .ck(clk) );
ms00f80 l1677 ( .d(n7845), .o(x264), .ck(clk) );
ms00f80 l1678 ( .d(n7848), .o(net_327), .ck(clk) );
ms00f80 l1679 ( .d(n7853), .o(net_200), .ck(clk) );
ms00f80 l1680 ( .d(n7858), .o(_net_5971), .ck(clk) );
ms00f80 l1681 ( .d(n7863), .o(_net_6409), .ck(clk) );
ms00f80 l1682 ( .d(n7867), .o(net_358), .ck(clk) );
ms00f80 l1683 ( .d(n7871), .o(net_137), .ck(clk) );
ms00f80 l1684 ( .d(n7875), .o(net_6874), .ck(clk) );
ms00f80 l1685 ( .d(n7878), .o(net_7673), .ck(clk) );
ms00f80 l1686 ( .d(n7883), .o(net_6344), .ck(clk) );
ms00f80 l1687 ( .d(n7888), .o(_net_7484), .ck(clk) );
ms00f80 l1688 ( .d(n7893), .o(net_7249), .ck(clk) );
ms00f80 l1689 ( .d(n7897), .o(_net_5850), .ck(clk) );
ms00f80 l1690 ( .d(n7902), .o(_net_6031), .ck(clk) );
ms00f80 l1691 ( .d(n7906), .o(net_7192), .ck(clk) );
ms00f80 l1692 ( .d(n7911), .o(_net_6552), .ck(clk) );
ms00f80 l1693 ( .d(n7916), .o(net_6363), .ck(clk) );
ms00f80 l1694 ( .d(n7920), .o(net_311), .ck(clk) );
ms00f80 l1695 ( .d(n7924), .o(net_7456), .ck(clk) );
ms00f80 l1696 ( .d(n7929), .o(net_6568), .ck(clk) );
ms00f80 l1697 ( .d(n7933), .o(net_237), .ck(clk) );
ms00f80 l1698 ( .d(n7937), .o(net_6930), .ck(clk) );
ms00f80 l1699 ( .d(n7942), .o(net_7540), .ck(clk) );
ms00f80 l1700 ( .d(n7945), .o(net_335), .ck(clk) );
ms00f80 l1701 ( .d(n7950), .o(net_6056), .ck(clk) );
ms00f80 l1702 ( .d(n7955), .o(net_6724), .ck(clk) );
ms00f80 l1703 ( .d(n7958), .o(net_6232), .ck(clk) );
ms00f80 l1704 ( .d(n7962), .o(net_7078), .ck(clk) );
ms00f80 l1705 ( .d(n7967), .o(net_6992), .ck(clk) );
ms00f80 l1706 ( .d(n7970), .o(net_7491), .ck(clk) );
ms00f80 l1707 ( .d(n7975), .o(_net_5855), .ck(clk) );
ms00f80 l1708 ( .d(n7980), .o(net_158), .ck(clk) );
ms00f80 l1709 ( .d(n7985), .o(_net_7425), .ck(clk) );
ms00f80 l1710 ( .d(n7989), .o(net_6651), .ck(clk) );
ms00f80 l1711 ( .d(n7994), .o(net_6585), .ck(clk) );
ms00f80 l1712 ( .d(n7997), .o(net_7087), .ck(clk) );
ms00f80 l1713 ( .d(n8002), .o(net_6975), .ck(clk) );
ms00f80 l1714 ( .d(n8005), .o(net_379), .ck(clk) );
ms00f80 l1715 ( .d(n8010), .o(_net_5852), .ck(clk) );
ms00f80 l1716 ( .d(n8015), .o(net_7131), .ck(clk) );
ms00f80 l1717 ( .d(n8019), .o(_net_291), .ck(clk) );
ms00f80 l1718 ( .d(n8024), .o(_net_6287), .ck(clk) );
ms00f80 l1719 ( .d(n8028), .o(net_6542), .ck(clk) );
ms00f80 l1720 ( .d(n8033), .o(_net_6072), .ck(clk) );
ms00f80 l1721 ( .d(n8038), .o(net_7680), .ck(clk) );
ms00f80 l1722 ( .d(n8042), .o(net_7744), .ck(clk) );
ms00f80 l1723 ( .d(n8047), .o(net_6365), .ck(clk) );
ms00f80 l1724 ( .d(n8051), .o(net_344), .ck(clk) );
ms00f80 l1725 ( .d(n8056), .o(net_6988), .ck(clk) );
ms00f80 l1726 ( .d(n8059), .o(net_6919), .ck(clk) );
ms00f80 l1727 ( .d(n8064), .o(net_6968), .ck(clk) );
ms00f80 l1728 ( .d(n8067), .o(net_6675), .ck(clk) );
ms00f80 l1729 ( .d(n8072), .o(net_6614), .ck(clk) );
ms00f80 l1730 ( .d(n8075), .o(net_6924), .ck(clk) );
ms00f80 l1731 ( .d(n8080), .o(_net_7262), .ck(clk) );
ms00f80 l1732 ( .d(n8085), .o(net_6596), .ck(clk) );
ms00f80 l1733 ( .d(n8088), .o(net_285), .ck(clk) );
ms00f80 l1734 ( .d(n8092), .o(net_7036), .ck(clk) );
ms00f80 l1735 ( .d(n8097), .o(_net_7573), .ck(clk) );
ms00f80 l1736 ( .d(n8102), .o(_net_7499), .ck(clk) );
ms00f80 l1737 ( .d(n8107), .o(_net_7417), .ck(clk) );
ms00f80 l1738 ( .d(n8112), .o(_net_6115), .ck(clk) );
ms00f80 l1739 ( .d(n8116), .o(net_6798), .ck(clk) );
ms00f80 l1740 ( .d(n8121), .o(_net_7562), .ck(clk) );
ms00f80 l1741 ( .d(n8125), .o(net_6895), .ck(clk) );
ms00f80 l1742 ( .d(n8130), .o(_net_7291), .ck(clk) );
ms00f80 l1743 ( .d(n8135), .o(_net_7592), .ck(clk) );
ms00f80 l1744 ( .d(n8140), .o(net_7141), .ck(clk) );
ms00f80 l1745 ( .d(n8144), .o(net_6571), .ck(clk) );
ms00f80 l1746 ( .d(n8147), .o(net_6638), .ck(clk) );
ms00f80 l1747 ( .d(n8152), .o(_net_262), .ck(clk) );
ms00f80 l1748 ( .d(n8156), .o(net_7339), .ck(clk) );
ms00f80 l1749 ( .d(n8161), .o(net_242), .ck(clk) );
ms00f80 l1750 ( .d(n8166), .o(net_7715), .ck(clk) );
ms00f80 l1751 ( .d(n8170), .o(_net_221), .ck(clk) );
ms00f80 l1752 ( .d(n8174), .o(net_6682), .ck(clk) );
ms00f80 l1753 ( .d(n8179), .o(_net_180), .ck(clk) );
ms00f80 l1754 ( .d(n8183), .o(net_6767), .ck(clk) );
ms00f80 l1755 ( .d(n8188), .o(net_6835), .ck(clk) );
ms00f80 l1756 ( .d(n8192), .o(_net_7275), .ck(clk) );
ms00f80 l1757 ( .d(n8197), .o(net_275), .ck(clk) );
ms00f80 l1758 ( .d(n8202), .o(_net_6159), .ck(clk) );
ms00f80 l1759 ( .d(n8206), .o(net_6678), .ck(clk) );
ms00f80 l1760 ( .d(n8211), .o(net_7772), .ck(clk) );
ms00f80 l1761 ( .d(n8216), .o(_net_7702), .ck(clk) );
ms00f80 l1762 ( .d(n8220), .o(net_6390), .ck(clk) );
ms00f80 l1763 ( .d(n8224), .o(_net_7755), .ck(clk) );
ms00f80 l1764 ( .d(n8228), .o(net_6910), .ck(clk) );
ms00f80 l1765 ( .d(n8232), .o(net_7177), .ck(clk) );
ms00f80 l1766 ( .d(n8237), .o(_net_7580), .ck(clk) );
ms00f80 l1767 ( .d(n8241), .o(net_370), .ck(clk) );
ms00f80 l1768 ( .d(n8245), .o(net_6494), .ck(clk) );
ms00f80 l1769 ( .d(n8249), .o(net_6389), .ck(clk) );
ms00f80 l1770 ( .d(n8253), .o(_net_7432), .ck(clk) );
ms00f80 l1771 ( .d(n8258), .o(net_196), .ck(clk) );
ms00f80 l1772 ( .d(n8262), .o(net_7615), .ck(clk) );
ms00f80 l1773 ( .d(n8266), .o(net_7169), .ck(clk) );
ms00f80 l1774 ( .d(n8271), .o(net_6312), .ck(clk) );
ms00f80 l1775 ( .d(n8276), .o(net_6615), .ck(clk) );
ms00f80 l1776 ( .d(n8280), .o(net_7538), .ck(clk) );
ms00f80 l1777 ( .d(n8284), .o(_net_6413), .ck(clk) );
ms00f80 l1778 ( .d(n8289), .o(net_6321), .ck(clk) );
ms00f80 l1779 ( .d(n8294), .o(_net_7648), .ck(clk) );
ms00f80 l1780 ( .d(n8299), .o(_net_6020), .ck(clk) );
ms00f80 l1781 ( .d(n8303), .o(net_7045), .ck(clk) );
ms00f80 l1782 ( .d(n8307), .o(net_7181), .ck(clk) );
ms00f80 l1783 ( .d(n8311), .o(net_7186), .ck(clk) );
ms00f80 l1784 ( .d(n8316), .o(net_6853), .ck(clk) );
ms00f80 l1785 ( .d(n8320), .o(net_7138), .ck(clk) );
ms00f80 l1786 ( .d(n8324), .o(_net_6201), .ck(clk) );
ms00f80 l1787 ( .d(n8329), .o(net_6276), .ck(clk) );
ms00f80 l1788 ( .d(n8334), .o(net_6851), .ck(clk) );
ms00f80 l1789 ( .d(n8337), .o(net_143), .ck(clk) );
ms00f80 l1790 ( .d(n8340), .o(net_6809), .ck(clk) );
ms00f80 l1791 ( .d(n8345), .o(_net_6123), .ck(clk) );
ms00f80 l1792 ( .d(n8350), .o(net_7023), .ck(clk) );
ms00f80 l1793 ( .d(n8354), .o(_net_6823), .ck(clk) );
ms00f80 l1794 ( .d(n8359), .o(net_6427), .ck(clk) );
ms00f80 l1795 ( .d(n8362), .o(net_7605), .ck(clk) );
ms00f80 l1796 ( .d(n8367), .o(_net_189), .ck(clk) );
ms00f80 l1797 ( .d(n8372), .o(_net_7685), .ck(clk) );
ms00f80 l1798 ( .d(n8377), .o(_net_7735), .ck(clk) );
ms00f80 l1799 ( .d(n8382), .o(_net_7602), .ck(clk) );
ms00f80 l1800 ( .d(n8387), .o(_net_6027), .ck(clk) );
ms00f80 l1801 ( .d(n8392), .o(net_6425), .ck(clk) );
ms00f80 l1802 ( .d(n8396), .o(_net_7568), .ck(clk) );
ms00f80 l1803 ( .d(n8401), .o(net_7104), .ck(clk) );
ms00f80 l1804 ( .d(n8405), .o(_net_6958), .ck(clk) );
ms00f80 l1805 ( .d(n8410), .o(_net_7333), .ck(clk) );
ms00f80 l1806 ( .d(n8415), .o(net_7137), .ck(clk) );
ms00f80 l1807 ( .d(n8418), .o(net_6393), .ck(clk) );
ms00f80 l1808 ( .d(n8422), .o(net_7237), .ck(clk) );
ms00f80 l1809 ( .d(n8426), .o(_net_6089), .ck(clk) );
ms00f80 l1810 ( .d(n8430), .o(net_332), .ck(clk) );
ms00f80 l1811 ( .d(n8435), .o(x342), .ck(clk) );
ms00f80 l1812 ( .d(n8438), .o(_net_5924), .ck(clk) );
ms00f80 l1813 ( .d(n8443), .o(_net_7687), .ck(clk) );
ms00f80 l1814 ( .d(n8447), .o(net_7375), .ck(clk) );
ms00f80 l1815 ( .d(n8451), .o(net_7459), .ck(clk) );
ms00f80 l1816 ( .d(n8455), .o(net_6945), .ck(clk) );
ms00f80 l1817 ( .d(n8459), .o(net_6518), .ck(clk) );
ms00f80 l1818 ( .d(n8464), .o(net_6742), .ck(clk) );
ms00f80 l1819 ( .d(n8467), .o(net_7039), .ck(clk) );
ms00f80 l1820 ( .d(n8472), .o(_net_5961), .ck(clk) );
ms00f80 l1821 ( .d(n8477), .o(net_6754), .ck(clk) );
ms00f80 l1822 ( .d(n8481), .o(_net_7450), .ck(clk) );
ms00f80 l1823 ( .d(n8486), .o(_net_6178), .ck(clk) );
ms00f80 l1824 ( .d(n8491), .o(net_7020), .ck(clk) );
ms00f80 l1825 ( .d(n8494), .o(net_7212), .ck(clk) );
ms00f80 l1826 ( .d(n8499), .o(_net_6039), .ck(clk) );
ms00f80 l1827 ( .d(n8504), .o(net_6622), .ck(clk) );
ms00f80 l1828 ( .d(n8508), .o(_net_6557), .ck(clk) );
ms00f80 l1829 ( .d(n8513), .o(net_6744), .ck(clk) );
ms00f80 l1830 ( .d(n8517), .o(_net_7575), .ck(clk) );
ms00f80 l1831 ( .d(n8522), .o(net_6838), .ck(clk) );
ms00f80 l1832 ( .d(n8526), .o(_net_7349), .ck(clk) );
ms00f80 l1833 ( .d(n8531), .o(_net_7284), .ck(clk) );
ms00f80 l1834 ( .d(n8535), .o(net_6771), .ck(clk) );
ms00f80 l1835 ( .d(n8540), .o(net_239), .ck(clk) );
ms00f80 l1836 ( .d(n8544), .o(net_6499), .ck(clk) );
ms00f80 l1837 ( .d(n8549), .o(net_6707), .ck(clk) );
ms00f80 l1838 ( .d(n8552), .o(net_6792), .ck(clk) );
ms00f80 l1839 ( .d(n8557), .o(net_166), .ck(clk) );
ms00f80 l1840 ( .d(n8561), .o(net_6956), .ck(clk) );
ms00f80 l1841 ( .d(n8565), .o(net_6794), .ck(clk) );
ms00f80 l1842 ( .d(n8570), .o(_net_122), .ck(clk) );
ms00f80 l1843 ( .d(n8575), .o(net_6475), .ck(clk) );
ms00f80 l1844 ( .d(n8578), .o(net_350), .ck(clk) );
ms00f80 l1845 ( .d(n8583), .o(_net_6282), .ck(clk) );
ms00f80 l1846 ( .d(n8588), .o(net_7778), .ck(clk) );
ms00f80 l1847 ( .d(n8593), .o(_net_7695), .ck(clk) );
ms00f80 l1848 ( .d(n8598), .o(net_6695), .ck(clk) );
ms00f80 l1849 ( .d(n8602), .o(_net_7319), .ck(clk) );
ms00f80 l1850 ( .d(n8607), .o(net_181), .ck(clk) );
ms00f80 l1851 ( .d(n8612), .o(net_6463), .ck(clk) );
ms00f80 l1852 ( .d(n8616), .o(net_6360), .ck(clk) );
ms00f80 l1853 ( .d(n8621), .o(net_6831), .ck(clk) );
ms00f80 l1854 ( .d(n8625), .o(net_388), .ck(clk) );
ms00f80 l1855 ( .d(n8628), .o(net_151), .ck(clk) );
ms00f80 l1856 ( .d(n8632), .o(net_6683), .ck(clk) );
ms00f80 l1857 ( .d(n8637), .o(net_6013), .ck(clk) );
ms00f80 l1858 ( .d(n8641), .o(net_6756), .ck(clk) );
ms00f80 l1859 ( .d(n8645), .o(_net_6141), .ck(clk) );
ms00f80 l1860 ( .d(n8650), .o(net_6865), .ck(clk) );
ms00f80 l1861 ( .d(n8654), .o(net_6577), .ck(clk) );
ms00f80 l1862 ( .d(n8658), .o(net_6600), .ck(clk) );
ms00f80 l1863 ( .d(n8662), .o(net_198), .ck(clk) );
ms00f80 l1864 ( .d(n8666), .o(net_7373), .ck(clk) );
ms00f80 l1865 ( .d(n8671), .o(_net_7267), .ck(clk) );
ms00f80 l1866 ( .d(n8676), .o(_net_6418), .ck(clk) );
ms00f80 l1867 ( .d(n8681), .o(net_6891), .ck(clk) );
ms00f80 l1868 ( .d(n8685), .o(net_6722), .ck(clk) );
ms00f80 l1869 ( .d(n8689), .o(_net_7627), .ck(clk) );
ms00f80 l1870 ( .d(n8694), .o(_net_6144), .ck(clk) );
ms00f80 l1871 ( .d(n8698), .o(_net_7811), .ck(clk) );
ms00f80 l1872 ( .d(n8703), .o(_net_6010), .ck(clk) );
ms00f80 l1873 ( .d(n8708), .o(x538), .ck(clk) );
ms00f80 l1874 ( .d(n8711), .o(net_7521), .ck(clk) );
ms00f80 l1875 ( .d(n8715), .o(net_333), .ck(clk) );
ms00f80 l1876 ( .d(n8720), .o(_net_7477), .ck(clk) );
ms00f80 l1877 ( .d(n8725), .o(_net_6824), .ck(clk) );
ms00f80 l1878 ( .d(n8730), .o(_net_6109), .ck(clk) );
ms00f80 l1879 ( .d(n8734), .o(net_7340), .ck(clk) );
ms00f80 l1880 ( .d(n8739), .o(net_7389), .ck(clk) );
ms00f80 l1881 ( .d(n8743), .o(_net_6043), .ck(clk) );
ms00f80 l1882 ( .d(n8748), .o(_net_7476), .ck(clk) );
ms00f80 l1883 ( .d(n8753), .o(_net_7585), .ck(clk) );
ms00f80 l1884 ( .d(n8757), .o(net_6234), .ck(clk) );
ms00f80 l1885 ( .d(n8762), .o(_net_6289), .ck(clk) );
ms00f80 l1886 ( .d(n8767), .o(net_7110), .ck(clk) );
ms00f80 l1887 ( .d(n8771), .o(net_387), .ck(clk) );
ms00f80 l1888 ( .d(n8775), .o(_net_7230), .ck(clk) );
ms00f80 l1889 ( .d(n8780), .o(_net_7265), .ck(clk) );
ms00f80 l1890 ( .d(n8784), .o(_net_7818), .ck(clk) );
ms00f80 l1891 ( .d(n8788), .o(net_6046), .ck(clk) );
ms00f80 l1892 ( .d(n8793), .o(net_6882), .ck(clk) );
ms00f80 l1893 ( .d(n8797), .o(net_6457), .ck(clk) );
ms00f80 l1894 ( .d(n8800), .o(net_7043), .ck(clk) );
ms00f80 l1895 ( .d(n8805), .o(net_6982), .ck(clk) );
ms00f80 l1896 ( .d(n8809), .o(net_6417), .ck(clk) );
ms00f80 l1897 ( .d(n8813), .o(net_7064), .ck(clk) );
ms00f80 l1898 ( .d(n8818), .o(_net_7409), .ck(clk) );
ms00f80 l1899 ( .d(n8823), .o(net_7542), .ck(clk) );
ms00f80 l1900 ( .d(n8826), .o(net_6787), .ck(clk) );
ms00f80 l1901 ( .d(n8831), .o(net_195), .ck(clk) );
ms00f80 l1902 ( .d(n8835), .o(net_7046), .ck(clk) );
ms00f80 l1903 ( .d(n8840), .o(_net_7664), .ck(clk) );
ms00f80 l1904 ( .d(n8845), .o(_net_6048), .ck(clk) );
ms00f80 l1905 ( .d(n8850), .o(_net_228), .ck(clk) );
ms00f80 l1906 ( .d(n8855), .o(_net_7363), .ck(clk) );
ms00f80 l1907 ( .d(n8860), .o(_net_7625), .ck(clk) );
ms00f80 l1908 ( .d(n8864), .o(_net_7806), .ck(clk) );
ms00f80 l1909 ( .d(n8869), .o(_net_6186), .ck(clk) );
ms00f80 l1910 ( .d(n8873), .o(net_6217), .ck(clk) );
ms00f80 l1911 ( .d(n8877), .o(net_307), .ck(clk) );
ms00f80 l1912 ( .d(n8882), .o(net_6196), .ck(clk) );
ms00f80 l1913 ( .d(n8886), .o(net_7086), .ck(clk) );
ms00f80 l1914 ( .d(n8891), .o(net_7132), .ck(clk) );
ms00f80 l1915 ( .d(n8895), .o(_net_6298), .ck(clk) );
ms00f80 l1916 ( .d(n8899), .o(net_7302), .ck(clk) );
ms00f80 l1917 ( .d(n8903), .o(net_6549), .ck(clk) );
ms00f80 l1918 ( .d(n8908), .o(net_6315), .ck(clk) );
ms00f80 l1919 ( .d(n8912), .o(net_6531), .ck(clk) );
ms00f80 l1920 ( .d(n8917), .o(_net_6166), .ck(clk) );
ms00f80 l1921 ( .d(n8922), .o(_net_7787), .ck(clk) );
ms00f80 l1922 ( .d(n8926), .o(net_6504), .ck(clk) );
ms00f80 l1923 ( .d(n8931), .o(net_7243), .ck(clk) );
ms00f80 l1924 ( .d(n8934), .o(net_7368), .ck(clk) );
ms00f80 l1925 ( .d(n8939), .o(net_6458), .ck(clk) );
ms00f80 l1926 ( .d(n8943), .o(net_6262), .ck(clk) );
ms00f80 l1927 ( .d(n8948), .o(_net_7322), .ck(clk) );
ms00f80 l1928 ( .d(n8953), .o(_net_7451), .ck(clk) );
ms00f80 l1929 ( .d(n8958), .o(net_6326), .ck(clk) );
ms00f80 l1930 ( .d(n8963), .o(net_7544), .ck(clk) );
ms00f80 l1931 ( .d(n8967), .o(_net_209), .ck(clk) );
ms00f80 l1932 ( .d(n8971), .o(net_6534), .ck(clk) );
ms00f80 l1933 ( .d(n8976), .o(_net_7466), .ck(clk) );
ms00f80 l1934 ( .d(n8981), .o(net_6350), .ck(clk) );
ms00f80 l1935 ( .d(n8986), .o(_net_7581), .ck(clk) );
ms00f80 l1936 ( .d(n8990), .o(net_304), .ck(clk) );
ms00f80 l1937 ( .d(n8995), .o(_net_293), .ck(clk) );
ms00f80 l1938 ( .d(n9000), .o(_net_268), .ck(clk) );
ms00f80 l1939 ( .d(n9005), .o(_net_7783), .ck(clk) );
ms00f80 l1940 ( .d(n9010), .o(net_6582), .ck(clk) );
ms00f80 l1941 ( .d(n9014), .o(net_7017), .ck(clk) );
ms00f80 l1942 ( .d(n9017), .o(net_6230), .ck(clk) );
ms00f80 l1943 ( .d(n9022), .o(net_6445), .ck(clk) );
ms00f80 l1944 ( .d(n9025), .o(net_6932), .ck(clk) );
ms00f80 l1945 ( .d(n9030), .o(x249), .ck(clk) );
ms00f80 l1946 ( .d(n9034), .o(net_6864), .ck(clk) );
ms00f80 l1947 ( .d(n9037), .o(net_6937), .ck(clk) );
ms00f80 l1948 ( .d(n9042), .o(net_230), .ck(clk) );
ms00f80 l1949 ( .d(n9047), .o(net_7762), .ck(clk) );
ms00f80 l1950 ( .d(n9052), .o(_net_7423), .ck(clk) );
ms00f80 l1951 ( .d(n9057), .o(net_6966), .ck(clk) );
ms00f80 l1952 ( .d(n9060), .o(net_7305), .ck(clk) );
ms00f80 l1953 ( .d(n9065), .o(net_6984), .ck(clk) );
ms00f80 l1954 ( .d(n9069), .o(net_6306), .ck(clk) );
ms00f80 l1955 ( .d(n9074), .o(_net_115), .ck(clk) );
ms00f80 l1956 ( .d(n9079), .o(net_7101), .ck(clk) );
ms00f80 l1957 ( .d(n9082), .o(net_7084), .ck(clk) );
ms00f80 l1958 ( .d(n9086), .o(net_6649), .ck(clk) );
ms00f80 l1959 ( .d(n9091), .o(net_6270), .ck(clk) );
ms00f80 l1960 ( .d(n9096), .o(net_256), .ck(clk) );
ms00f80 l1961 ( .d(n9101), .o(_net_289), .ck(clk) );
ms00f80 l1962 ( .d(n9106), .o(_net_7716), .ck(clk) );
ms00f80 l1963 ( .d(n9110), .o(_net_7804), .ck(clk) );
ms00f80 l1964 ( .d(n9115), .o(_net_292), .ck(clk) );
ms00f80 l1965 ( .d(n9120), .o(net_7155), .ck(clk) );
ms00f80 l1966 ( .d(n9124), .o(_net_7558), .ck(clk) );
ms00f80 l1967 ( .d(n9129), .o(_net_7660), .ck(clk) );
ms00f80 l1968 ( .d(n9134), .o(net_6333), .ck(clk) );
ms00f80 l1969 ( .d(n9138), .o(net_6520), .ck(clk) );
ms00f80 l1970 ( .d(n9143), .o(net_6876), .ck(clk) );
ms00f80 l1971 ( .d(n9146), .o(net_6665), .ck(clk) );
ms00f80 l1972 ( .d(n9151), .o(net_162), .ck(clk) );
ms00f80 l1973 ( .d(n9156), .o(_net_7259), .ck(clk) );
ms00f80 l1974 ( .d(n9160), .o(net_318), .ck(clk) );
ms00f80 l1975 ( .d(n9164), .o(net_6911), .ck(clk) );
ms00f80 l1976 ( .d(n9169), .o(net_6565), .ck(clk) );
ms00f80 l1977 ( .d(n9173), .o(_net_6188), .ck(clk) );
ms00f80 l1978 ( .d(n9178), .o(net_6253), .ck(clk) );
ms00f80 l1979 ( .d(n9182), .o(net_6492), .ck(clk) );
ms00f80 l1980 ( .d(n9187), .o(_net_7260), .ck(clk) );
ms00f80 l1981 ( .d(n9192), .o(_net_172), .ck(clk) );
ms00f80 l1982 ( .d(n9196), .o(net_328), .ck(clk) );
ms00f80 l1983 ( .d(n9201), .o(_net_7682), .ck(clk) );
ms00f80 l1984 ( .d(n9206), .o(_net_5986), .ck(clk) );
ms00f80 l1985 ( .d(n9211), .o(net_7776), .ck(clk) );
ms00f80 l1986 ( .d(n9215), .o(net_7367), .ck(clk) );
ms00f80 l1987 ( .d(n9220), .o(_net_6094), .ck(clk) );
ms00f80 l1988 ( .d(n9225), .o(net_7156), .ck(clk) );
ms00f80 l1989 ( .d(n9228), .o(net_7463), .ck(clk) );
ms00f80 l1990 ( .d(n9233), .o(_net_7701), .ck(clk) );
ms00f80 l1991 ( .d(n9238), .o(net_6705), .ck(clk) );
ms00f80 l1992 ( .d(n9242), .o(net_6483), .ck(clk) );
ms00f80 l1993 ( .d(n9245), .o(net_6527), .ck(clk) );
ms00f80 l1994 ( .d(n9250), .o(net_6701), .ck(clk) );
ms00f80 l1995 ( .d(n9254), .o(net_7103), .ck(clk) );
ms00f80 l1996 ( .d(n9258), .o(_net_6405), .ck(clk) );
ms00f80 l1997 ( .d(n9263), .o(_net_7515), .ck(clk) );
ms00f80 l1998 ( .d(n9267), .o(net_6669), .ck(clk) );
ms00f80 l1999 ( .d(n9272), .o(_net_7530), .ck(clk) );
ms00f80 l2000 ( .d(n9277), .o(_net_6106), .ck(clk) );
ms00f80 l2001 ( .d(n9282), .o(_net_6137), .ck(clk) );
ms00f80 l2002 ( .d(n9287), .o(net_6848), .ck(clk) );
ms00f80 l2003 ( .d(n9290), .o(net_7190), .ck(clk) );
ms00f80 l2004 ( .d(n9294), .o(net_7218), .ck(clk) );
ms00f80 l2005 ( .d(n9298), .o(net_7612), .ck(clk) );
ms00f80 l2006 ( .d(n9302), .o(net_7519), .ck(clk) );
ms00f80 l2007 ( .d(n9307), .o(_net_7516), .ck(clk) );
ms00f80 l2008 ( .d(n9312), .o(_net_7726), .ck(clk) );
ms00f80 l2009 ( .d(n9316), .o(net_7377), .ck(clk) );
ms00f80 l2010 ( .d(n9321), .o(net_219), .ck(clk) );
ms00f80 l2011 ( .d(n9326), .o(net_6749), .ck(clk) );
ms00f80 l2012 ( .d(n9330), .o(_net_5983), .ck(clk) );
ms00f80 l2013 ( .d(n9335), .o(_net_7725), .ck(clk) );
ms00f80 l2014 ( .d(n9339), .o(net_6662), .ck(clk) );
ms00f80 l2015 ( .d(n9343), .o(net_6535), .ck(clk) );
ms00f80 l2016 ( .d(n9348), .o(net_7541), .ck(clk) );
ms00f80 l2017 ( .d(n9352), .o(_net_7504), .ck(clk) );
ms00f80 l2018 ( .d(n9356), .o(net_7164), .ck(clk) );
ms00f80 l2019 ( .d(n9361), .o(net_6464), .ck(clk) );
ms00f80 l2020 ( .d(n9365), .o(net_6265), .ck(clk) );
ms00f80 l2021 ( .d(n9370), .o(net_7099), .ck(clk) );
ms00f80 l2022 ( .d(n9373), .o(net_6640), .ck(clk) );
ms00f80 l2023 ( .d(n9377), .o(net_6817), .ck(clk) );
ms00f80 l2024 ( .d(n9381), .o(net_6921), .ck(clk) );
ms00f80 l2025 ( .d(n9385), .o(net_7072), .ck(clk) );
ms00f80 l2026 ( .d(n9390), .o(net_6601), .ck(clk) );
ms00f80 l2027 ( .d(n9393), .o(net_6936), .ck(clk) );
ms00f80 l2028 ( .d(n9398), .o(net_6278), .ck(clk) );
ms00f80 l2029 ( .d(n9402), .o(x0), .ck(clk) );
ms00f80 l2030 ( .d(n9405), .o(net_6908), .ck(clk) );
ms00f80 l2031 ( .d(n9410), .o(_net_7569), .ck(clk) );
ms00f80 l2032 ( .d(n9415), .o(_net_6085), .ck(clk) );
ms00f80 l2033 ( .d(n9420), .o(_net_7317), .ck(clk) );
ms00f80 l2034 ( .d(n9425), .o(net_6459), .ck(clk) );
ms00f80 l2035 ( .d(n9428), .o(net_145), .ck(clk) );
ms00f80 l2036 ( .d(n9431), .o(net_6775), .ck(clk) );
ms00f80 l2037 ( .d(n9436), .o(_net_7745), .ck(clk) );
ms00f80 l2038 ( .d(n9441), .o(x638), .ck(clk) );
ms00f80 l2039 ( .d(n9445), .o(net_6731), .ck(clk) );
ms00f80 l2040 ( .d(n9449), .o(_net_6280), .ck(clk) );
ms00f80 l2041 ( .d(n9454), .o(_net_6005), .ck(clk) );
ms00f80 l2042 ( .d(n9459), .o(net_7709), .ck(clk) );
ms00f80 l2043 ( .d(n9462), .o(net_6916), .ck(clk) );
ms00f80 l2044 ( .d(n9467), .o(net_6972), .ck(clk) );
ms00f80 l2045 ( .d(n9470), .o(net_359), .ck(clk) );
ms00f80 l2046 ( .d(n9475), .o(net_6842), .ck(clk) );
ms00f80 l2047 ( .d(n9478), .o(net_7464), .ck(clk) );
ms00f80 l2048 ( .d(n9483), .o(net_6611), .ck(clk) );
ms00f80 l2049 ( .d(n9487), .o(_net_7415), .ck(clk) );
ms00f80 l2050 ( .d(n9492), .o(_net_7282), .ck(clk) );
ms00f80 l2051 ( .d(n9497), .o(_net_7597), .ck(clk) );
ms00f80 l2052 ( .d(n9502), .o(net_6359), .ck(clk) );
ms00f80 l2053 ( .d(n9507), .o(_net_7617), .ck(clk) );
ms00f80 l2054 ( .d(n9512), .o(_net_7616), .ck(clk) );
ms00f80 l2055 ( .d(n9517), .o(net_6871), .ck(clk) );
ms00f80 l2056 ( .d(n9520), .o(net_316), .ck(clk) );
ms00f80 l2057 ( .d(n9525), .o(net_7015), .ck(clk) );
ms00f80 l2058 ( .d(n9528), .o(net_6667), .ck(clk) );
ms00f80 l2059 ( .d(n9533), .o(_net_217), .ck(clk) );
ms00f80 l2060 ( .d(n9537), .o(net_6782), .ck(clk) );
ms00f80 l2061 ( .d(n9541), .o(net_7183), .ck(clk) );
ms00f80 l2062 ( .d(n9546), .o(x138), .ck(clk) );
ms00f80 l2063 ( .d(n9549), .o(net_7524), .ck(clk) );
ms00f80 l2064 ( .d(n9554), .o(net_6058), .ck(clk) );
ms00f80 l2065 ( .d(n9559), .o(_net_190), .ck(clk) );
ms00f80 l2066 ( .d(n9564), .o(_net_6021), .ck(clk) );
ms00f80 l2067 ( .d(n9569), .o(_net_7509), .ck(clk) );
ms00f80 l2068 ( .d(n9574), .o(net_297), .ck(clk) );
ms00f80 l2069 ( .d(n9579), .o(net_6840), .ck(clk) );
ms00f80 l2070 ( .d(n9583), .o(_net_7506), .ck(clk) );
ms00f80 l2071 ( .d(n9588), .o(net_6455), .ck(clk) );
ms00f80 l2072 ( .d(n9592), .o(net_6036), .ck(clk) );
ms00f80 l2073 ( .d(n9597), .o(_net_6153), .ck(clk) );
ms00f80 l2074 ( .d(n9602), .o(_net_7324), .ck(clk) );
ms00f80 l2075 ( .d(n9606), .o(net_6818), .ck(clk) );
ms00f80 l2076 ( .d(n9611), .o(net_6307), .ck(clk) );
ms00f80 l2077 ( .d(n9616), .o(_net_6052), .ck(clk) );
ms00f80 l2078 ( .d(n9620), .o(net_6785), .ck(clk) );
ms00f80 l2079 ( .d(n9624), .o(net_7205), .ck(clk) );
ms00f80 l2080 ( .d(n9628), .o(_net_6219), .ck(clk) );
ms00f80 l2081 ( .d(n9633), .o(_net_7436), .ck(clk) );
ms00f80 l2082 ( .d(n9638), .o(_net_7414), .ck(clk) );
ms00f80 l2083 ( .d(n9642), .o(net_6644), .ck(clk) );
ms00f80 l2084 ( .d(n9647), .o(net_7386), .ck(clk) );
ms00f80 l2085 ( .d(n9651), .o(net_7548), .ck(clk) );
ms00f80 l2086 ( .d(n9655), .o(_net_7327), .ck(clk) );
ms00f80 l2087 ( .d(n9660), .o(net_7005), .ck(clk) );
ms00f80 l2088 ( .d(n9664), .o(_net_7656), .ck(clk) );
ms00f80 l2089 ( .d(n9668), .o(net_368), .ck(clk) );
ms00f80 l2090 ( .d(n9673), .o(_net_7588), .ck(clk) );
ms00f80 l2091 ( .d(n9678), .o(_net_225), .ck(clk) );
ms00f80 l2092 ( .d(n9683), .o(_net_7560), .ck(clk) );
ms00f80 l2093 ( .d(n9687), .o(net_317), .ck(clk) );
ms00f80 l2094 ( .d(n9692), .o(net_6703), .ck(clk) );
ms00f80 l2095 ( .d(n9695), .o(net_366), .ck(clk) );
ms00f80 l2096 ( .d(n9700), .o(_net_5964), .ck(clk) );
ms00f80 l2097 ( .d(n9704), .o(net_6634), .ck(clk) );
ms00f80 l2098 ( .d(n9709), .o(_net_6051), .ck(clk) );
ms00f80 l2099 ( .d(n9714), .o(_net_6143), .ck(clk) );
ms00f80 l2100 ( .d(n9719), .o(_net_6174), .ck(clk) );
ms00f80 l2101 ( .d(n9724), .o(net_6358), .ck(clk) );
ms00f80 l2102 ( .d(n9729), .o(net_6472), .ck(clk) );
ms00f80 l2103 ( .d(n9733), .o(_net_192), .ck(clk) );
ms00f80 l2104 ( .d(n9737), .o(_net_7817), .ck(clk) );
ms00f80 l2105 ( .d(n9742), .o(net_170), .ck(clk) );
ms00f80 l2106 ( .d(n9746), .o(net_7214), .ck(clk) );
ms00f80 l2107 ( .d(n9750), .o(net_6657), .ck(clk) );
ms00f80 l2108 ( .d(n9754), .o(net_7522), .ck(clk) );
ms00f80 l2109 ( .d(n9758), .o(net_7669), .ck(clk) );
ms00f80 l2110 ( .d(n9763), .o(_net_7576), .ck(clk) );
ms00f80 l2111 ( .d(n9768), .o(_net_7283), .ck(clk) );
ms00f80 l2112 ( .d(n9773), .o(_net_6002), .ck(clk) );
ms00f80 l2113 ( .d(n9778), .o(_net_5973), .ck(clk) );
ms00f80 l2114 ( .d(n9783), .o(net_7027), .ck(clk) );
ms00f80 l2115 ( .d(n9787), .o(_net_7566), .ck(clk) );
ms00f80 l2116 ( .d(n9792), .o(_net_5989), .ck(clk) );
ms00f80 l2117 ( .d(n9796), .o(net_6807), .ck(clk) );
ms00f80 l2118 ( .d(n9801), .o(_net_7384), .ck(clk) );
ms00f80 l2119 ( .d(n9805), .o(net_384), .ck(clk) );
ms00f80 l2120 ( .d(n9809), .o(net_313), .ck(clk) );
ms00f80 l2121 ( .d(n9814), .o(_net_5859), .ck(clk) );
ms00f80 l2122 ( .d(n9819), .o(_net_7533), .ck(clk) );
ms00f80 l2123 ( .d(n9824), .o(_net_7383), .ck(clk) );
ms00f80 l2124 ( .d(n9828), .o(net_7674), .ck(clk) );
ms00f80 l2125 ( .d(n9833), .o(net_7135), .ck(clk) );
ms00f80 l2126 ( .d(n9837), .o(net_7122), .ck(clk) );
ms00f80 l2127 ( .d(n9840), .o(net_321), .ck(clk) );
ms00f80 l2128 ( .d(n9844), .o(net_305), .ck(clk) );
ms00f80 l2129 ( .d(n9849), .o(_net_7421), .ck(clk) );
ms00f80 l2130 ( .d(n9853), .o(net_7644), .ck(clk) );
ms00f80 l2131 ( .d(n9858), .o(_net_6407), .ck(clk) );
ms00f80 l2132 ( .d(n9863), .o(_net_7097), .ck(clk) );
ms00f80 l2133 ( .d(n9867), .o(net_6943), .ck(clk) );
ms00f80 l2134 ( .d(n9871), .o(net_6929), .ck(clk) );
ms00f80 l2135 ( .d(n9875), .o(net_6533), .ck(clk) );
ms00f80 l2136 ( .d(n9880), .o(_net_6421), .ck(clk) );
ms00f80 l2137 ( .d(n9885), .o(net_7109), .ck(clk) );
ms00f80 l2138 ( .d(n9889), .o(_net_6111), .ck(clk) );
ms00f80 l2139 ( .d(n9894), .o(_net_287), .ck(clk) );
ms00f80 l2140 ( .d(n9899), .o(net_6752), .ck(clk) );
ms00f80 l2141 ( .d(n9902), .o(net_6795), .ck(clk) );
ms00f80 l2142 ( .d(n9907), .o(x361), .ck(clk) );
ms00f80 l2143 ( .d(n9911), .o(net_6446), .ck(clk) );
ms00f80 l2144 ( .d(n9914), .o(net_7221), .ck(clk) );
ms00f80 l2145 ( .d(n9918), .o(_net_7795), .ck(clk) );
ms00f80 l2146 ( .d(n9923), .o(net_6719), .ck(clk) );
ms00f80 l2147 ( .d(n9926), .o(net_374), .ck(clk) );
ms00f80 l2148 ( .d(n9930), .o(net_338), .ck(clk) );
ms00f80 l2149 ( .d(n9935), .o(net_6465), .ck(clk) );
ms00f80 l2150 ( .d(n9939), .o(_net_288), .ck(clk) );
ms00f80 l2151 ( .d(n9944), .o(net_6370), .ck(clk) );
ms00f80 l2152 ( .d(n9949), .o(_net_7348), .ck(clk) );
ms00f80 l2153 ( .d(n9953), .o(net_7740), .ck(clk) );
ms00f80 l2154 ( .d(n9957), .o(net_354), .ck(clk) );
ms00f80 l2155 ( .d(n9961), .o(net_7071), .ck(clk) );
ms00f80 l2156 ( .d(n9966), .o(_net_7402), .ck(clk) );
ms00f80 l2157 ( .d(n9971), .o(_net_6076), .ck(clk) );
ms00f80 l2158 ( .d(n9976), .o(net_6192), .ck(clk) );
ms00f80 l2159 ( .d(n9981), .o(_net_7788), .ck(clk) );
ms00f80 l2160 ( .d(n9985), .o(net_6381), .ck(clk) );
ms00f80 l2161 ( .d(n9988), .o(net_6905), .ck(clk) );
ms00f80 l2162 ( .d(n9992), .o(net_7175), .ck(clk) );
ms00f80 l2163 ( .d(n9997), .o(_net_7717), .ck(clk) );
ms00f80 l2164 ( .d(n10001), .o(net_6507), .ck(clk) );
ms00f80 l2165 ( .d(n10006), .o(net_6198), .ck(clk) );
ms00f80 l2166 ( .d(n10010), .o(net_6529), .ck(clk) );
ms00f80 l2167 ( .d(n10014), .o(_net_7823), .ck(clk) );
ms00f80 l2168 ( .d(n10019), .o(_net_267), .ck(clk) );
ms00f80 l2169 ( .d(n10023), .o(net_6224), .ck(clk) );
ms00f80 l2170 ( .d(n10028), .o(net_6879), .ck(clk) );
ms00f80 l2171 ( .d(n10032), .o(_net_7582), .ck(clk) );
ms00f80 l2172 ( .d(n10037), .o(_net_6017), .ck(clk) );
ms00f80 l2173 ( .d(n10042), .o(_net_6203), .ck(clk) );
ms00f80 l2174 ( .d(n10047), .o(net_6351), .ck(clk) );
ms00f80 l2175 ( .d(n10052), .o(_net_7287), .ck(clk) );
ms00f80 l2176 ( .d(n10056), .o(net_7677), .ck(clk) );
ms00f80 l2177 ( .d(n10061), .o(net_7773), .ck(clk) );
ms00f80 l2178 ( .d(n10066), .o(x620), .ck(clk) );
ms00f80 l2179 ( .d(n10070), .o(net_6884), .ck(clk) );
ms00f80 l2180 ( .d(n10074), .o(_net_7251), .ck(clk) );
ms00f80 l2181 ( .d(n10079), .o(_net_6555), .ck(clk) );
ms00f80 l2182 ( .d(n10084), .o(_net_6131), .ck(clk) );
ms00f80 l2183 ( .d(n10089), .o(_net_6183), .ck(clk) );
ms00f80 l2184 ( .d(n10094), .o(_net_7264), .ck(clk) );
ms00f80 l2185 ( .d(n10099), .o(_net_7479), .ck(clk) );
ms00f80 l2186 ( .d(n10103), .o(net_6645), .ck(clk) );
ms00f80 l2187 ( .d(n10107), .o(net_6648), .ck(clk) );
ms00f80 l2188 ( .d(n10112), .o(net_7112), .ck(clk) );
ms00f80 l2189 ( .d(n10116), .o(net_248), .ck(clk) );
ms00f80 l2190 ( .d(n10120), .o(net_6780), .ck(clk) );
ms00f80 l2191 ( .d(n10124), .o(net_148), .ck(clk) );
ms00f80 l2192 ( .d(n10128), .o(_net_7356), .ck(clk) );
ms00f80 l2193 ( .d(n10132), .o(net_6532), .ck(clk) );
ms00f80 l2194 ( .d(n10137), .o(_net_6176), .ck(clk) );
ms00f80 l2195 ( .d(n10141), .o(_net_7793), .ck(clk) );
ms00f80 l2196 ( .d(n10145), .o(net_7313), .ck(clk) );
ms00f80 l2197 ( .d(n10150), .o(_net_6164), .ck(clk) );
ms00f80 l2198 ( .d(n10154), .o(net_6772), .ck(clk) );
ms00f80 l2199 ( .d(n10158), .o(net_7041), .ck(clk) );
vcc     t0 ( .o(n7265) );

endmodule
