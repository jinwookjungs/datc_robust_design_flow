// Written by verilog_parser.py of OpenDesign Flow Database.
// Date: 2019-06-04 13:24:09
// Format: ICCAD2015 placement contest

module ac97_ctrl (
clk,
x1006,
x1034,
x1062,
x1101,
x1126,
x1155,
x1193,
x1203,
x1209,
x1215,
x1231,
x1261,
x1286,
x130657,
x1322,
x1345,
x1351,
x1358,
x1366,
x1374,
x1382,
x1390,
x1398,
x1406,
x1417,
x1424,
x1432,
x1443,
x1451,
x1459,
x1467,
x1479,
x1486,
x1494,
x1501,
x1511,
x1519,
x1527,
x1534,
x1542,
x1550,
x1557,
x1564,
x1572,
x1580,
x1587,
x1595,
x806,
x837,
x868,
x889,
x906,
x940,
x977,
_net_6050,
_net_6051,
_net_6052,
net_275,
net_286,
net_300,
net_301,
net_302,
net_5849,
net_6047,
net_6053,
net_6054,
net_6055,
net_6190,
net_6191,
net_6192,
net_6193,
net_6195,
net_6196,
net_6197,
net_6198,
net_6211,
net_6212,
net_6213,
net_6214,
net_6215,
net_6216,
net_6217,
net_6218,
net_6223,
net_6224,
net_6225,
net_6226,
net_6227,
net_6228,
net_6229,
net_6230,
net_6231,
net_6232,
net_6233,
net_6234,
net_6235,
net_6236,
net_6237,
net_6238,
net_6240,
net_6241,
net_6242,
net_6243,
net_6244,
net_6245,
net_6246,
net_6247,
net_6248,
net_6249,
net_6250,
net_6251,
net_6252,
net_6253,
net_6254,
net_6255,
net_6256,
net_6257,
net_6258,
net_6260,
net_6261,
net_6262,
net_6263,
net_6264,
net_6265,
net_6266,
net_6267,
net_6268,
net_6269,
net_6270,
net_6271,
net_6272,
net_6273,
net_6274,
net_6275,
net_6276,
net_6277,
net_6278,
net_6279,
net_6299,
net_6300,
net_6301,
net_6302,
net_6303,
net_6304,
net_6305,
net_6306,
net_6307,
net_6308,
net_6309,
net_6310,
net_6311,
net_6312,
net_6313,
net_6314,
net_6315,
net_6316,
net_6317,
net_6318,
net_6320,
net_6321,
net_6322,
net_6323,
net_6324,
net_6325,
net_6326,
net_6327,
net_6328,
net_6329,
net_6330,
net_6331,
net_6332,
net_6333,
net_6334,
net_6335,
net_6336,
net_6337,
net_6338,
net_6339,
net_6340,
net_6341,
net_6342,
net_6343,
net_6344,
net_6345,
net_6346,
net_6347,
net_6348,
net_6349,
net_6350,
net_6351,
net_6352,
net_6353,
net_6354,
net_6355,
net_6356,
net_6357,
net_6358,
net_6359,
net_6360,
net_6361,
net_6362,
net_6363,
net_6364,
net_6365,
net_6366,
net_6367,
net_6368,
net_6369,
net_6370,
net_6371,
net_6372,
net_6373,
net_6374,
net_6375,
net_6376,
net_6377,
net_6378,
net_6379,
net_7762,
net_7764,
net_7766,
x0,
x101,
x106,
x114,
x124,
x131,
x138,
x14,
x145,
x149,
x172,
x179,
x187,
x195,
x217,
x234,
x249,
x264,
x287,
x30,
x315,
x342,
x361,
x379,
x38,
x390,
x397,
x420,
x447,
x476,
x494,
x522,
x538,
x561,
x589,
x620,
x63,
x638,
x657,
x681,
x699,
x718,
x744,
x765,
x77,
x786,
x84,
x96
);

// Start PIs
input clk;
input x1006;
input x1034;
input x1062;
input x1101;
input x1126;
input x1155;
input x1193;
input x1203;
input x1209;
input x1215;
input x1231;
input x1261;
input x1286;
input x130657;
input x1322;
input x1345;
input x1351;
input x1358;
input x1366;
input x1374;
input x1382;
input x1390;
input x1398;
input x1406;
input x1417;
input x1424;
input x1432;
input x1443;
input x1451;
input x1459;
input x1467;
input x1479;
input x1486;
input x1494;
input x1501;
input x1511;
input x1519;
input x1527;
input x1534;
input x1542;
input x1550;
input x1557;
input x1564;
input x1572;
input x1580;
input x1587;
input x1595;
input x806;
input x837;
input x868;
input x889;
input x906;
input x940;
input x977;

// Start POs
output _net_6050;
output _net_6051;
output _net_6052;
output net_275;
output net_286;
output net_300;
output net_301;
output net_302;
output net_5849;
output net_6047;
output net_6053;
output net_6054;
output net_6055;
output net_6190;
output net_6191;
output net_6192;
output net_6193;
output net_6195;
output net_6196;
output net_6197;
output net_6198;
output net_6211;
output net_6212;
output net_6213;
output net_6214;
output net_6215;
output net_6216;
output net_6217;
output net_6218;
output net_6223;
output net_6224;
output net_6225;
output net_6226;
output net_6227;
output net_6228;
output net_6229;
output net_6230;
output net_6231;
output net_6232;
output net_6233;
output net_6234;
output net_6235;
output net_6236;
output net_6237;
output net_6238;
output net_6240;
output net_6241;
output net_6242;
output net_6243;
output net_6244;
output net_6245;
output net_6246;
output net_6247;
output net_6248;
output net_6249;
output net_6250;
output net_6251;
output net_6252;
output net_6253;
output net_6254;
output net_6255;
output net_6256;
output net_6257;
output net_6258;
output net_6260;
output net_6261;
output net_6262;
output net_6263;
output net_6264;
output net_6265;
output net_6266;
output net_6267;
output net_6268;
output net_6269;
output net_6270;
output net_6271;
output net_6272;
output net_6273;
output net_6274;
output net_6275;
output net_6276;
output net_6277;
output net_6278;
output net_6279;
output net_6299;
output net_6300;
output net_6301;
output net_6302;
output net_6303;
output net_6304;
output net_6305;
output net_6306;
output net_6307;
output net_6308;
output net_6309;
output net_6310;
output net_6311;
output net_6312;
output net_6313;
output net_6314;
output net_6315;
output net_6316;
output net_6317;
output net_6318;
output net_6320;
output net_6321;
output net_6322;
output net_6323;
output net_6324;
output net_6325;
output net_6326;
output net_6327;
output net_6328;
output net_6329;
output net_6330;
output net_6331;
output net_6332;
output net_6333;
output net_6334;
output net_6335;
output net_6336;
output net_6337;
output net_6338;
output net_6339;
output net_6340;
output net_6341;
output net_6342;
output net_6343;
output net_6344;
output net_6345;
output net_6346;
output net_6347;
output net_6348;
output net_6349;
output net_6350;
output net_6351;
output net_6352;
output net_6353;
output net_6354;
output net_6355;
output net_6356;
output net_6357;
output net_6358;
output net_6359;
output net_6360;
output net_6361;
output net_6362;
output net_6363;
output net_6364;
output net_6365;
output net_6366;
output net_6367;
output net_6368;
output net_6369;
output net_6370;
output net_6371;
output net_6372;
output net_6373;
output net_6374;
output net_6375;
output net_6376;
output net_6377;
output net_6378;
output net_6379;
output net_7762;
output net_7764;
output net_7766;
output x0;
output x101;
output x106;
output x114;
output x124;
output x131;
output x138;
output x14;
output x145;
output x149;
output x172;
output x179;
output x187;
output x195;
output x217;
output x234;
output x249;
output x264;
output x287;
output x30;
output x315;
output x342;
output x361;
output x379;
output x38;
output x390;
output x397;
output x420;
output x447;
output x476;
output x494;
output x522;
output x538;
output x561;
output x589;
output x620;
output x63;
output x638;
output x657;
output x681;
output x699;
output x718;
output x744;
output x765;
output x77;
output x786;
output x84;
output x96;

// Start wires
wire clk;
wire x1006;
wire x1034;
wire x1062;
wire x1101;
wire x1126;
wire x1155;
wire x1193;
wire x1203;
wire x1209;
wire x1215;
wire x1231;
wire x1261;
wire x1286;
wire x130657;
wire x1322;
wire x1345;
wire x1351;
wire x1358;
wire x1366;
wire x1374;
wire x1382;
wire x1390;
wire x1398;
wire x1406;
wire x1417;
wire x1424;
wire x1432;
wire x1443;
wire x1451;
wire x1459;
wire x1467;
wire x1479;
wire x1486;
wire x1494;
wire x1501;
wire x1511;
wire x1519;
wire x1527;
wire x1534;
wire x1542;
wire x1550;
wire x1557;
wire x1564;
wire x1572;
wire x1580;
wire x1587;
wire x1595;
wire x806;
wire x837;
wire x868;
wire x889;
wire x906;
wire x940;
wire x977;
wire _net_6050;
wire _net_6051;
wire _net_6052;
wire net_275;
wire net_286;
wire net_300;
wire net_301;
wire net_302;
wire net_5849;
wire net_6047;
wire net_6053;
wire net_6054;
wire net_6055;
wire net_6190;
wire net_6191;
wire net_6192;
wire net_6193;
wire net_6195;
wire net_6196;
wire net_6197;
wire net_6198;
wire net_6211;
wire net_6212;
wire net_6213;
wire net_6214;
wire net_6215;
wire net_6216;
wire net_6217;
wire net_6218;
wire net_6223;
wire net_6224;
wire net_6225;
wire net_6226;
wire net_6227;
wire net_6228;
wire net_6229;
wire net_6230;
wire net_6231;
wire net_6232;
wire net_6233;
wire net_6234;
wire net_6235;
wire net_6236;
wire net_6237;
wire net_6238;
wire net_6240;
wire net_6241;
wire net_6242;
wire net_6243;
wire net_6244;
wire net_6245;
wire net_6246;
wire net_6247;
wire net_6248;
wire net_6249;
wire net_6250;
wire net_6251;
wire net_6252;
wire net_6253;
wire net_6254;
wire net_6255;
wire net_6256;
wire net_6257;
wire net_6258;
wire net_6260;
wire net_6261;
wire net_6262;
wire net_6263;
wire net_6264;
wire net_6265;
wire net_6266;
wire net_6267;
wire net_6268;
wire net_6269;
wire net_6270;
wire net_6271;
wire net_6272;
wire net_6273;
wire net_6274;
wire net_6275;
wire net_6276;
wire net_6277;
wire net_6278;
wire net_6279;
wire net_6299;
wire net_6300;
wire net_6301;
wire net_6302;
wire net_6303;
wire net_6304;
wire net_6305;
wire net_6306;
wire net_6307;
wire net_6308;
wire net_6309;
wire net_6310;
wire net_6311;
wire net_6312;
wire net_6313;
wire net_6314;
wire net_6315;
wire net_6316;
wire net_6317;
wire net_6318;
wire net_6320;
wire net_6321;
wire net_6322;
wire net_6323;
wire net_6324;
wire net_6325;
wire net_6326;
wire net_6327;
wire net_6328;
wire net_6329;
wire net_6330;
wire net_6331;
wire net_6332;
wire net_6333;
wire net_6334;
wire net_6335;
wire net_6336;
wire net_6337;
wire net_6338;
wire net_6339;
wire net_6340;
wire net_6341;
wire net_6342;
wire net_6343;
wire net_6344;
wire net_6345;
wire net_6346;
wire net_6347;
wire net_6348;
wire net_6349;
wire net_6350;
wire net_6351;
wire net_6352;
wire net_6353;
wire net_6354;
wire net_6355;
wire net_6356;
wire net_6357;
wire net_6358;
wire net_6359;
wire net_6360;
wire net_6361;
wire net_6362;
wire net_6363;
wire net_6364;
wire net_6365;
wire net_6366;
wire net_6367;
wire net_6368;
wire net_6369;
wire net_6370;
wire net_6371;
wire net_6372;
wire net_6373;
wire net_6374;
wire net_6375;
wire net_6376;
wire net_6377;
wire net_6378;
wire net_6379;
wire net_7762;
wire net_7764;
wire net_7766;
wire x0;
wire x101;
wire x106;
wire x114;
wire x124;
wire x131;
wire x138;
wire x14;
wire x145;
wire x149;
wire x172;
wire x179;
wire x187;
wire x195;
wire x217;
wire x234;
wire x249;
wire x264;
wire x287;
wire x30;
wire x315;
wire x342;
wire x361;
wire x379;
wire x38;
wire x390;
wire x397;
wire x420;
wire x447;
wire x476;
wire x494;
wire x522;
wire x538;
wire x561;
wire x589;
wire x620;
wire x63;
wire x638;
wire x657;
wire x681;
wire x699;
wire x718;
wire x744;
wire x765;
wire x77;
wire x786;
wire x84;
wire x96;
wire _net_113;
wire _net_114;
wire _net_115;
wire _net_116;
wire _net_117;
wire _net_118;
wire _net_119;
wire _net_120;
wire _net_121;
wire _net_122;
wire _net_123;
wire _net_124;
wire _net_125;
wire _net_126;
wire _net_127;
wire _net_128;
wire _net_129;
wire _net_154;
wire _net_172;
wire _net_173;
wire _net_174;
wire _net_175;
wire _net_176;
wire _net_177;
wire _net_178;
wire _net_180;
wire _net_184;
wire _net_188;
wire _net_189;
wire _net_190;
wire _net_191;
wire _net_192;
wire _net_193;
wire _net_201;
wire _net_209;
wire _net_210;
wire _net_211;
wire _net_212;
wire _net_213;
wire _net_214;
wire _net_215;
wire _net_217;
wire _net_221;
wire _net_225;
wire _net_226;
wire _net_227;
wire _net_228;
wire _net_229;
wire _net_262;
wire _net_263;
wire _net_264;
wire _net_265;
wire _net_266;
wire _net_267;
wire _net_268;
wire _net_269;
wire _net_270;
wire _net_271;
wire _net_272;
wire _net_273;
wire _net_276;
wire _net_277;
wire _net_278;
wire _net_279;
wire _net_280;
wire _net_281;
wire _net_282;
wire _net_283;
wire _net_284;
wire _net_287;
wire _net_288;
wire _net_289;
wire _net_290;
wire _net_291;
wire _net_292;
wire _net_293;
wire _net_294;
wire _net_295;
wire _net_298;
wire _net_299;
wire _net_392;
wire _net_5848;
wire _net_5850;
wire _net_5851;
wire _net_5852;
wire _net_5853;
wire _net_5854;
wire _net_5855;
wire _net_5856;
wire _net_5857;
wire _net_5859;
wire _net_5920;
wire _net_5922;
wire _net_5924;
wire _net_5960;
wire _net_5961;
wire _net_5962;
wire _net_5963;
wire _net_5964;
wire _net_5965;
wire _net_5966;
wire _net_5967;
wire _net_5968;
wire _net_5969;
wire _net_5970;
wire _net_5971;
wire _net_5972;
wire _net_5973;
wire _net_5974;
wire _net_5975;
wire _net_5976;
wire _net_5977;
wire _net_5978;
wire _net_5979;
wire _net_5980;
wire _net_5981;
wire _net_5982;
wire _net_5983;
wire _net_5984;
wire _net_5985;
wire _net_5986;
wire _net_5987;
wire _net_5988;
wire _net_5989;
wire _net_5990;
wire _net_5991;
wire _net_5993;
wire _net_5994;
wire _net_5995;
wire _net_5996;
wire _net_5997;
wire _net_5998;
wire _net_5999;
wire _net_6000;
wire _net_6001;
wire _net_6002;
wire _net_6004;
wire _net_6005;
wire _net_6006;
wire _net_6007;
wire _net_6008;
wire _net_6009;
wire _net_6010;
wire _net_6011;
wire _net_6012;
wire _net_6015;
wire _net_6016;
wire _net_6017;
wire _net_6018;
wire _net_6019;
wire _net_6020;
wire _net_6021;
wire _net_6022;
wire _net_6023;
wire _net_6026;
wire _net_6027;
wire _net_6028;
wire _net_6029;
wire _net_6030;
wire _net_6031;
wire _net_6032;
wire _net_6033;
wire _net_6034;
wire _net_6037;
wire _net_6038;
wire _net_6039;
wire _net_6040;
wire _net_6041;
wire _net_6042;
wire _net_6043;
wire _net_6044;
wire _net_6045;
wire _net_6048;
wire _net_6049;
wire _net_6062;
wire _net_6063;
wire _net_6064;
wire _net_6065;
wire _net_6066;
wire _net_6067;
wire _net_6068;
wire _net_6069;
wire _net_6070;
wire _net_6071;
wire _net_6072;
wire _net_6073;
wire _net_6074;
wire _net_6075;
wire _net_6076;
wire _net_6077;
wire _net_6078;
wire _net_6079;
wire _net_6080;
wire _net_6081;
wire _net_6082;
wire _net_6083;
wire _net_6084;
wire _net_6085;
wire _net_6086;
wire _net_6087;
wire _net_6088;
wire _net_6089;
wire _net_6090;
wire _net_6091;
wire _net_6092;
wire _net_6093;
wire _net_6094;
wire _net_6095;
wire _net_6096;
wire _net_6097;
wire _net_6098;
wire _net_6099;
wire _net_6100;
wire _net_6101;
wire _net_6102;
wire _net_6103;
wire _net_6104;
wire _net_6105;
wire _net_6106;
wire _net_6107;
wire _net_6108;
wire _net_6109;
wire _net_6110;
wire _net_6111;
wire _net_6112;
wire _net_6113;
wire _net_6114;
wire _net_6115;
wire _net_6116;
wire _net_6117;
wire _net_6118;
wire _net_6119;
wire _net_6120;
wire _net_6121;
wire _net_6122;
wire _net_6123;
wire _net_6124;
wire _net_6125;
wire _net_6126;
wire _net_6127;
wire _net_6128;
wire _net_6129;
wire _net_6130;
wire _net_6131;
wire _net_6132;
wire _net_6133;
wire _net_6134;
wire _net_6135;
wire _net_6136;
wire _net_6137;
wire _net_6138;
wire _net_6139;
wire _net_6140;
wire _net_6141;
wire _net_6142;
wire _net_6143;
wire _net_6144;
wire _net_6145;
wire _net_6146;
wire _net_6147;
wire _net_6148;
wire _net_6149;
wire _net_6150;
wire _net_6151;
wire _net_6152;
wire _net_6153;
wire _net_6154;
wire _net_6155;
wire _net_6156;
wire _net_6157;
wire _net_6158;
wire _net_6159;
wire _net_6160;
wire _net_6161;
wire _net_6162;
wire _net_6163;
wire _net_6164;
wire _net_6165;
wire _net_6166;
wire _net_6167;
wire _net_6168;
wire _net_6169;
wire _net_6170;
wire _net_6171;
wire _net_6172;
wire _net_6173;
wire _net_6174;
wire _net_6175;
wire _net_6176;
wire _net_6177;
wire _net_6178;
wire _net_6179;
wire _net_6180;
wire _net_6181;
wire _net_6182;
wire _net_6183;
wire _net_6184;
wire _net_6185;
wire _net_6186;
wire _net_6187;
wire _net_6188;
wire _net_6189;
wire _net_6194;
wire _net_6199;
wire _net_6200;
wire _net_6201;
wire _net_6202;
wire _net_6203;
wire _net_6204;
wire _net_6205;
wire _net_6206;
wire _net_6207;
wire _net_6208;
wire _net_6209;
wire _net_6210;
wire _net_6219;
wire _net_6220;
wire _net_6221;
wire _net_6222;
wire _net_6239;
wire _net_6259;
wire _net_6280;
wire _net_6281;
wire _net_6282;
wire _net_6283;
wire _net_6284;
wire _net_6285;
wire _net_6286;
wire _net_6287;
wire _net_6288;
wire _net_6289;
wire _net_6290;
wire _net_6291;
wire _net_6292;
wire _net_6293;
wire _net_6294;
wire _net_6295;
wire _net_6296;
wire _net_6297;
wire _net_6298;
wire _net_6319;
wire _net_6401;
wire _net_6402;
wire _net_6404;
wire _net_6405;
wire _net_6406;
wire _net_6407;
wire _net_6408;
wire _net_6409;
wire _net_6410;
wire _net_6411;
wire _net_6413;
wire _net_6414;
wire _net_6415;
wire _net_6418;
wire _net_6419;
wire _net_6420;
wire _net_6421;
wire _net_6422;
wire _net_6423;
wire _net_6552;
wire _net_6553;
wire _net_6554;
wire _net_6555;
wire _net_6557;
wire _net_6558;
wire _net_6687;
wire _net_6688;
wire _net_6689;
wire _net_6690;
wire _net_6692;
wire _net_6693;
wire _net_6822;
wire _net_6823;
wire _net_6824;
wire _net_6825;
wire _net_6827;
wire _net_6828;
wire _net_6957;
wire _net_6958;
wire _net_6959;
wire _net_6960;
wire _net_6962;
wire _net_6963;
wire _net_7092;
wire _net_7093;
wire _net_7094;
wire _net_7095;
wire _net_7097;
wire _net_7098;
wire _net_7227;
wire _net_7228;
wire _net_7229;
wire _net_7230;
wire _net_7232;
wire _net_7233;
wire _net_7250;
wire _net_7251;
wire _net_7252;
wire _net_7253;
wire _net_7254;
wire _net_7255;
wire _net_7256;
wire _net_7257;
wire _net_7258;
wire _net_7259;
wire _net_7260;
wire _net_7261;
wire _net_7262;
wire _net_7263;
wire _net_7264;
wire _net_7265;
wire _net_7266;
wire _net_7267;
wire _net_7268;
wire _net_7269;
wire _net_7270;
wire _net_7271;
wire _net_7272;
wire _net_7273;
wire _net_7274;
wire _net_7275;
wire _net_7276;
wire _net_7277;
wire _net_7278;
wire _net_7279;
wire _net_7280;
wire _net_7281;
wire _net_7282;
wire _net_7283;
wire _net_7284;
wire _net_7285;
wire _net_7286;
wire _net_7287;
wire _net_7288;
wire _net_7289;
wire _net_7290;
wire _net_7291;
wire _net_7292;
wire _net_7293;
wire _net_7294;
wire _net_7295;
wire _net_7296;
wire _net_7297;
wire _net_7298;
wire _net_7299;
wire _net_7300;
wire _net_7301;
wire _net_7314;
wire _net_7315;
wire _net_7316;
wire _net_7317;
wire _net_7318;
wire _net_7319;
wire _net_7320;
wire _net_7321;
wire _net_7322;
wire _net_7323;
wire _net_7324;
wire _net_7325;
wire _net_7326;
wire _net_7327;
wire _net_7328;
wire _net_7329;
wire _net_7330;
wire _net_7331;
wire _net_7332;
wire _net_7333;
wire _net_7346;
wire _net_7347;
wire _net_7348;
wire _net_7349;
wire _net_7350;
wire _net_7351;
wire _net_7352;
wire _net_7353;
wire _net_7354;
wire _net_7355;
wire _net_7356;
wire _net_7357;
wire _net_7358;
wire _net_7359;
wire _net_7360;
wire _net_7361;
wire _net_7362;
wire _net_7363;
wire _net_7364;
wire _net_7365;
wire _net_7379;
wire _net_7380;
wire _net_7381;
wire _net_7382;
wire _net_7383;
wire _net_7384;
wire _net_7401;
wire _net_7402;
wire _net_7403;
wire _net_7404;
wire _net_7405;
wire _net_7406;
wire _net_7407;
wire _net_7408;
wire _net_7409;
wire _net_7410;
wire _net_7411;
wire _net_7412;
wire _net_7413;
wire _net_7414;
wire _net_7415;
wire _net_7416;
wire _net_7417;
wire _net_7418;
wire _net_7419;
wire _net_7420;
wire _net_7421;
wire _net_7422;
wire _net_7423;
wire _net_7424;
wire _net_7425;
wire _net_7426;
wire _net_7427;
wire _net_7428;
wire _net_7429;
wire _net_7430;
wire _net_7431;
wire _net_7432;
wire _net_7433;
wire _net_7434;
wire _net_7435;
wire _net_7436;
wire _net_7437;
wire _net_7438;
wire _net_7439;
wire _net_7440;
wire _net_7441;
wire _net_7442;
wire _net_7443;
wire _net_7444;
wire _net_7445;
wire _net_7446;
wire _net_7447;
wire _net_7448;
wire _net_7449;
wire _net_7450;
wire _net_7451;
wire _net_7452;
wire _net_7465;
wire _net_7466;
wire _net_7467;
wire _net_7468;
wire _net_7469;
wire _net_7470;
wire _net_7471;
wire _net_7472;
wire _net_7473;
wire _net_7474;
wire _net_7475;
wire _net_7476;
wire _net_7477;
wire _net_7478;
wire _net_7479;
wire _net_7480;
wire _net_7481;
wire _net_7482;
wire _net_7483;
wire _net_7484;
wire _net_7497;
wire _net_7498;
wire _net_7499;
wire _net_7500;
wire _net_7501;
wire _net_7502;
wire _net_7503;
wire _net_7504;
wire _net_7505;
wire _net_7506;
wire _net_7507;
wire _net_7508;
wire _net_7509;
wire _net_7510;
wire _net_7511;
wire _net_7512;
wire _net_7513;
wire _net_7514;
wire _net_7515;
wire _net_7516;
wire _net_7530;
wire _net_7531;
wire _net_7532;
wire _net_7533;
wire _net_7534;
wire _net_7535;
wire _net_7552;
wire _net_7553;
wire _net_7554;
wire _net_7555;
wire _net_7556;
wire _net_7557;
wire _net_7558;
wire _net_7559;
wire _net_7560;
wire _net_7561;
wire _net_7562;
wire _net_7563;
wire _net_7564;
wire _net_7565;
wire _net_7566;
wire _net_7567;
wire _net_7568;
wire _net_7569;
wire _net_7570;
wire _net_7571;
wire _net_7572;
wire _net_7573;
wire _net_7574;
wire _net_7575;
wire _net_7576;
wire _net_7577;
wire _net_7578;
wire _net_7579;
wire _net_7580;
wire _net_7581;
wire _net_7582;
wire _net_7583;
wire _net_7584;
wire _net_7585;
wire _net_7586;
wire _net_7587;
wire _net_7588;
wire _net_7589;
wire _net_7590;
wire _net_7591;
wire _net_7592;
wire _net_7593;
wire _net_7594;
wire _net_7595;
wire _net_7596;
wire _net_7597;
wire _net_7598;
wire _net_7599;
wire _net_7600;
wire _net_7601;
wire _net_7602;
wire _net_7603;
wire _net_7616;
wire _net_7617;
wire _net_7618;
wire _net_7619;
wire _net_7620;
wire _net_7621;
wire _net_7622;
wire _net_7623;
wire _net_7624;
wire _net_7625;
wire _net_7626;
wire _net_7627;
wire _net_7628;
wire _net_7629;
wire _net_7630;
wire _net_7631;
wire _net_7632;
wire _net_7633;
wire _net_7634;
wire _net_7635;
wire _net_7648;
wire _net_7649;
wire _net_7650;
wire _net_7651;
wire _net_7652;
wire _net_7653;
wire _net_7654;
wire _net_7655;
wire _net_7656;
wire _net_7657;
wire _net_7658;
wire _net_7659;
wire _net_7660;
wire _net_7661;
wire _net_7662;
wire _net_7663;
wire _net_7664;
wire _net_7665;
wire _net_7666;
wire _net_7667;
wire _net_7681;
wire _net_7682;
wire _net_7683;
wire _net_7684;
wire _net_7685;
wire _net_7686;
wire _net_7687;
wire _net_7688;
wire _net_7689;
wire _net_7690;
wire _net_7692;
wire _net_7693;
wire _net_7694;
wire _net_7695;
wire _net_7696;
wire _net_7697;
wire _net_7698;
wire _net_7699;
wire _net_7700;
wire _net_7701;
wire _net_7702;
wire _net_7703;
wire _net_7704;
wire _net_7705;
wire _net_7706;
wire _net_7707;
wire _net_7716;
wire _net_7717;
wire _net_7718;
wire _net_7719;
wire _net_7720;
wire _net_7721;
wire _net_7722;
wire _net_7723;
wire _net_7724;
wire _net_7725;
wire _net_7726;
wire _net_7727;
wire _net_7728;
wire _net_7729;
wire _net_7730;
wire _net_7731;
wire _net_7732;
wire _net_7733;
wire _net_7734;
wire _net_7735;
wire _net_7736;
wire _net_7745;
wire _net_7746;
wire _net_7747;
wire _net_7748;
wire _net_7749;
wire _net_7751;
wire _net_7753;
wire _net_7755;
wire _net_7757;
wire _net_7759;
wire _net_7761;
wire _net_7763;
wire _net_7765;
wire _net_7768;
wire _net_7781;
wire _net_7782;
wire _net_7783;
wire _net_7784;
wire _net_7785;
wire _net_7786;
wire _net_7787;
wire _net_7788;
wire _net_7789;
wire _net_7791;
wire _net_7793;
wire _net_7794;
wire _net_7795;
wire _net_7796;
wire _net_7797;
wire _net_7798;
wire _net_7800;
wire _net_7801;
wire _net_7803;
wire _net_7804;
wire _net_7805;
wire _net_7806;
wire _net_7808;
wire _net_7809;
wire _net_7810;
wire _net_7811;
wire _net_7812;
wire _net_7813;
wire _net_7814;
wire _net_7815;
wire _net_7816;
wire _net_7817;
wire _net_7818;
wire _net_7819;
wire _net_7820;
wire _net_7821;
wire _net_7822;
wire _net_7823;
wire _net_7824;
wire n1000;
wire n10000;
wire n10001;
wire n10001_1;
wire n10002;
wire n10003;
wire n10004;
wire n10005;
wire n10006;
wire n10006_1;
wire n10007;
wire n10009;
wire n10010;
wire n10010_1;
wire n10012;
wire n10013;
wire n10014;
wire n10014_1;
wire n10015;
wire n10016;
wire n10017;
wire n10018;
wire n10019;
wire n10019_1;
wire n10020;
wire n10021;
wire n10022;
wire n10023;
wire n10024;
wire n10026;
wire n10028;
wire n10028_1;
wire n10029;
wire n10031;
wire n10032;
wire n10032_1;
wire n10034;
wire n10035;
wire n10037;
wire n10037_1;
wire n10038;
wire n10040;
wire n10041;
wire n10042;
wire n10043;
wire n10044;
wire n10045;
wire n10046;
wire n10047;
wire n10047_1;
wire n10048;
wire n10049;
wire n1005;
wire n10050;
wire n10051;
wire n10052;
wire n10052_1;
wire n10053;
wire n10055;
wire n10056;
wire n10056_1;
wire n10057;
wire n10058;
wire n10059;
wire n10060;
wire n10061;
wire n10061_1;
wire n10062;
wire n10063;
wire n10064;
wire n10065;
wire n10066;
wire n10066_1;
wire n10068;
wire n10069;
wire n10070;
wire n10070_1;
wire n10071;
wire n10072;
wire n10074;
wire n10074_1;
wire n10075;
wire n10077;
wire n10078;
wire n10079;
wire n10080;
wire n10081;
wire n10083;
wire n10084;
wire n10084_1;
wire n10086;
wire n10087;
wire n10088;
wire n10089;
wire n10089_1;
wire n10090;
wire n10092;
wire n10093;
wire n10094;
wire n10095;
wire n10097;
wire n10098;
wire n10099;
wire n1010;
wire n10100;
wire n10101;
wire n10103;
wire n10103_1;
wire n10104;
wire n10106;
wire n10107;
wire n10107_1;
wire n10108;
wire n10109;
wire n10110;
wire n10112;
wire n10112_1;
wire n10113;
wire n10115;
wire n10116;
wire n10116_1;
wire n10117;
wire n10119;
wire n10120;
wire n10120_1;
wire n10122;
wire n10123;
wire n10124;
wire n10125;
wire n10126;
wire n10127;
wire n10128;
wire n10128_1;
wire n10129;
wire n10130;
wire n10131;
wire n10132;
wire n10132_1;
wire n10133;
wire n10134;
wire n10135;
wire n10136;
wire n10137;
wire n10137_1;
wire n10138;
wire n10139;
wire n10140;
wire n10141;
wire n10141_1;
wire n10142;
wire n10143;
wire n10145;
wire n10145_1;
wire n10146;
wire n10148;
wire n10149;
wire n1015;
wire n10150;
wire n10151;
wire n10152;
wire n10154;
wire n10154_1;
wire n10155;
wire n10157;
wire n10158;
wire n10158_1;
wire n10160;
wire n10161;
wire n10163;
wire n10164;
wire n10166;
wire n10167;
wire n10169;
wire n10170;
wire n10172;
wire n10174;
wire n10175;
wire n10177;
wire n10178;
wire n10179;
wire n10180;
wire n10181;
wire n10182;
wire n10183;
wire n10184;
wire n10186;
wire n10187;
wire n10188;
wire n10189;
wire n10191;
wire n10192;
wire n10193;
wire n10194;
wire n10195;
wire n10196;
wire n10197;
wire n10198;
wire n10199;
wire n1020;
wire n10200;
wire n10201;
wire n10202;
wire n10203;
wire n10204;
wire n10206;
wire n10207;
wire n10208;
wire n10210;
wire n10211;
wire n10214;
wire n10215;
wire n10217;
wire n10219;
wire n10220;
wire n10222;
wire n10223;
wire n10225;
wire n10226;
wire n10227;
wire n10228;
wire n10229;
wire n10230;
wire n10231;
wire n10232;
wire n10233;
wire n10234;
wire n10235;
wire n10236;
wire n10237;
wire n10239;
wire n1024;
wire n10240;
wire n10242;
wire n10243;
wire n10244;
wire n10245;
wire n10246;
wire n10247;
wire n10248;
wire n10249;
wire n10250;
wire n10251;
wire n10252;
wire n10253;
wire n10254;
wire n10255;
wire n10256;
wire n10257;
wire n10258;
wire n10259;
wire n10260;
wire n10262;
wire n10264;
wire n10266;
wire n10267;
wire n10270;
wire n10271;
wire n10272;
wire n10274;
wire n10275;
wire n10277;
wire n10279;
wire n10280;
wire n10283;
wire n10284;
wire n10286;
wire n10287;
wire n10289;
wire n1029;
wire n10290;
wire n10291;
wire n10292;
wire n10293;
wire n10294;
wire n10295;
wire n10297;
wire n10298;
wire n10299;
wire n10301;
wire n10302;
wire n10303;
wire n10304;
wire n10305;
wire n10306;
wire n10307;
wire n10308;
wire n10309;
wire n10310;
wire n10311;
wire n10312;
wire n10314;
wire n10315;
wire n10317;
wire n10319;
wire n10320;
wire n10322;
wire n10323;
wire n10325;
wire n10326;
wire n10328;
wire n10329;
wire n10331;
wire n10332;
wire n10333;
wire n10334;
wire n10336;
wire n10337;
wire n10338;
wire n10339;
wire n1034;
wire n10340;
wire n10341;
wire n10342;
wire n10343;
wire n10344;
wire n10346;
wire n10348;
wire n10349;
wire n10351;
wire n10352;
wire n10354;
wire n10355;
wire n10357;
wire n10359;
wire n10360;
wire n10362;
wire n10363;
wire n10364;
wire n10365;
wire n10366;
wire n10367;
wire n10369;
wire n10371;
wire n10372;
wire n10374;
wire n10375;
wire n10377;
wire n10378;
wire n10380;
wire n10381;
wire n10382;
wire n10383;
wire n10384;
wire n10385;
wire n10386;
wire n10387;
wire n10388;
wire n10389;
wire n1039;
wire n10390;
wire n10391;
wire n10393;
wire n10394;
wire n10396;
wire n10397;
wire n10398;
wire n10399;
wire n10400;
wire n10401;
wire n10402;
wire n10403;
wire n10404;
wire n10405;
wire n10406;
wire n10407;
wire n10409;
wire n10410;
wire n10412;
wire n10413;
wire n10414;
wire n10415;
wire n10416;
wire n10418;
wire n10419;
wire n10421;
wire n10422;
wire n10423;
wire n10424;
wire n10426;
wire n10427;
wire n10429;
wire n10430;
wire n10431;
wire n10432;
wire n10433;
wire n10434;
wire n10435;
wire n10436;
wire n10437;
wire n10438;
wire n10439;
wire n1044;
wire n10440;
wire n10441;
wire n10442;
wire n10443;
wire n10444;
wire n10445;
wire n10446;
wire n10447;
wire n10448;
wire n10450;
wire n10452;
wire n10453;
wire n10455;
wire n10456;
wire n10458;
wire n10460;
wire n10462;
wire n10463;
wire n10464;
wire n10465;
wire n10466;
wire n10468;
wire n10469;
wire n10471;
wire n10472;
wire n10473;
wire n10474;
wire n10475;
wire n10476;
wire n10477;
wire n10479;
wire n10480;
wire n10482;
wire n10483;
wire n10485;
wire n10486;
wire n10487;
wire n10488;
wire n10489;
wire n1049;
wire n10490;
wire n10491;
wire n10492;
wire n10493;
wire n10494;
wire n10495;
wire n10496;
wire n10497;
wire n10498;
wire n10499;
wire n10500;
wire n10501;
wire n10502;
wire n10503;
wire n10505;
wire n10506;
wire n10508;
wire n10509;
wire n10511;
wire n10512;
wire n10514;
wire n10515;
wire n10517;
wire n10518;
wire n10520;
wire n10521;
wire n10523;
wire n10524;
wire n10525;
wire n10526;
wire n10527;
wire n10528;
wire n10529;
wire n1053;
wire n10530;
wire n10532;
wire n10533;
wire n10534;
wire n10535;
wire n10536;
wire n10537;
wire n10539;
wire n10540;
wire n10541;
wire n10543;
wire n10544;
wire n10546;
wire n10547;
wire n10548;
wire n10549;
wire n10550;
wire n10551;
wire n10552;
wire n10553;
wire n10554;
wire n10555;
wire n10556;
wire n10557;
wire n10558;
wire n10559;
wire n10560;
wire n10561;
wire n10562;
wire n10563;
wire n10564;
wire n10565;
wire n10567;
wire n10568;
wire n10570;
wire n10571;
wire n10573;
wire n10574;
wire n10575;
wire n10576;
wire n10577;
wire n10578;
wire n1058;
wire n10580;
wire n10581;
wire n10583;
wire n10584;
wire n10585;
wire n10586;
wire n10587;
wire n10588;
wire n10589;
wire n10590;
wire n10591;
wire n10592;
wire n10593;
wire n10594;
wire n10595;
wire n10596;
wire n10597;
wire n10598;
wire n10599;
wire n10600;
wire n10601;
wire n10603;
wire n10604;
wire n10606;
wire n10607;
wire n10609;
wire n10610;
wire n10611;
wire n10613;
wire n10614;
wire n10616;
wire n10617;
wire n10619;
wire n1062;
wire n10620;
wire n10621;
wire n10622;
wire n10623;
wire n10624;
wire n10625;
wire n10626;
wire n10627;
wire n10628;
wire n10629;
wire n10630;
wire n10631;
wire n10632;
wire n10633;
wire n10634;
wire n10636;
wire n10637;
wire n10639;
wire n10640;
wire n10642;
wire n10643;
wire n10645;
wire n10646;
wire n10648;
wire n10649;
wire n10651;
wire n10652;
wire n10654;
wire n10655;
wire n10656;
wire n10657;
wire n10658;
wire n10659;
wire n10660;
wire n10661;
wire n10662;
wire n10663;
wire n10664;
wire n10665;
wire n10666;
wire n10667;
wire n10668;
wire n10669;
wire n1067;
wire n10670;
wire n10671;
wire n10672;
wire n10674;
wire n10675;
wire n10677;
wire n10678;
wire n10679;
wire n10680;
wire n10681;
wire n10682;
wire n10683;
wire n10684;
wire n10686;
wire n10687;
wire n10689;
wire n10690;
wire n10691;
wire n10692;
wire n10694;
wire n10695;
wire n10696;
wire n10697;
wire n10698;
wire n10699;
wire n10701;
wire n10702;
wire n10704;
wire n10705;
wire n10706;
wire n10707;
wire n10708;
wire n10709;
wire n10710;
wire n10711;
wire n10712;
wire n10713;
wire n10714;
wire n10715;
wire n10716;
wire n10717;
wire n10719;
wire n1072;
wire n10721;
wire n10722;
wire n10723;
wire n10724;
wire n10725;
wire n10726;
wire n10727;
wire n10728;
wire n10730;
wire n10731;
wire n10733;
wire n10734;
wire n10736;
wire n10737;
wire n10738;
wire n10739;
wire n10740;
wire n10741;
wire n10742;
wire n10743;
wire n10744;
wire n10745;
wire n10746;
wire n10747;
wire n10748;
wire n10749;
wire n10750;
wire n10751;
wire n10752;
wire n10753;
wire n10754;
wire n10755;
wire n10756;
wire n10757;
wire n10758;
wire n10759;
wire n10760;
wire n10761;
wire n10762;
wire n10763;
wire n10765;
wire n10766;
wire n10768;
wire n10769;
wire n1077;
wire n10770;
wire n10771;
wire n10772;
wire n10773;
wire n10774;
wire n10775;
wire n10776;
wire n10777;
wire n10778;
wire n10779;
wire n10781;
wire n10782;
wire n10783;
wire n10784;
wire n10785;
wire n10786;
wire n10787;
wire n10788;
wire n10789;
wire n10790;
wire n10791;
wire n10792;
wire n10794;
wire n10795;
wire n10797;
wire n10798;
wire n10800;
wire n10801;
wire n10803;
wire n10804;
wire n10806;
wire n10807;
wire n1081;
wire n10810;
wire n10811;
wire n10813;
wire n10814;
wire n10816;
wire n10817;
wire n10819;
wire n10820;
wire n10822;
wire n10823;
wire n10824;
wire n10825;
wire n10826;
wire n10827;
wire n10828;
wire n10829;
wire n10830;
wire n10831;
wire n10832;
wire n10833;
wire n10835;
wire n10836;
wire n10838;
wire n10839;
wire n10841;
wire n10842;
wire n10844;
wire n10845;
wire n10847;
wire n10848;
wire n1085;
wire n10850;
wire n10851;
wire n10853;
wire n10854;
wire n10856;
wire n10857;
wire n10858;
wire n10859;
wire n10860;
wire n10861;
wire n10862;
wire n10863;
wire n10864;
wire n10865;
wire n10866;
wire n10867;
wire n10869;
wire n10870;
wire n10872;
wire n10873;
wire n10875;
wire n10877;
wire n10878;
wire n10880;
wire n10881;
wire n10882;
wire n10883;
wire n10884;
wire n10885;
wire n10886;
wire n10887;
wire n10888;
wire n10889;
wire n1089;
wire n10890;
wire n10891;
wire n10893;
wire n10894;
wire n10896;
wire n10897;
wire n10899;
wire n10900;
wire n10902;
wire n10903;
wire n10905;
wire n10906;
wire n10907;
wire n10908;
wire n10909;
wire n10910;
wire n10911;
wire n10912;
wire n10913;
wire n10914;
wire n10915;
wire n10916;
wire n10917;
wire n10920;
wire n10922;
wire n10923;
wire n10925;
wire n10926;
wire n10928;
wire n10929;
wire n1093;
wire n10931;
wire n10933;
wire n10934;
wire n10935;
wire n10936;
wire n10938;
wire n10940;
wire n10941;
wire n10943;
wire n10944;
wire n10945;
wire n10947;
wire n10948;
wire n10949;
wire n10950;
wire n10951;
wire n10952;
wire n10953;
wire n10954;
wire n10955;
wire n10956;
wire n10957;
wire n10958;
wire n10960;
wire n10961;
wire n10963;
wire n10965;
wire n10967;
wire n10969;
wire n1097;
wire n10970;
wire n10972;
wire n10973;
wire n10974;
wire n10977;
wire n10978;
wire n10979;
wire n10980;
wire n10982;
wire n10985;
wire n10987;
wire n10989;
wire n10990;
wire n10992;
wire n10993;
wire n10995;
wire n10996;
wire n10997;
wire n10998;
wire n10999;
wire n11000;
wire n11001;
wire n11002;
wire n11003;
wire n11004;
wire n11005;
wire n11006;
wire n11008;
wire n11009;
wire n11011;
wire n11012;
wire n11014;
wire n11015;
wire n11017;
wire n11018;
wire n1102;
wire n11020;
wire n11021;
wire n11023;
wire n11024;
wire n11026;
wire n11027;
wire n11028;
wire n11029;
wire n11030;
wire n11031;
wire n11034;
wire n11035;
wire n11036;
wire n11037;
wire n11039;
wire n11040;
wire n11042;
wire n11043;
wire n11045;
wire n11047;
wire n11048;
wire n11050;
wire n11051;
wire n11052;
wire n11054;
wire n11055;
wire n11056;
wire n11057;
wire n1106;
wire n11060;
wire n11061;
wire n11063;
wire n11064;
wire n11065;
wire n11066;
wire n11067;
wire n11068;
wire n11069;
wire n11070;
wire n11072;
wire n11073;
wire n11075;
wire n11076;
wire n11078;
wire n11079;
wire n11080;
wire n11081;
wire n11083;
wire n11084;
wire n11086;
wire n11087;
wire n11089;
wire n11090;
wire n11092;
wire n11093;
wire n11095;
wire n11096;
wire n11097;
wire n11099;
wire n11100;
wire n11101;
wire n11103;
wire n11104;
wire n11106;
wire n11108;
wire n11109;
wire n1111;
wire n11111;
wire n11113;
wire n11115;
wire n11116;
wire n11118;
wire n11119;
wire n11120;
wire n11121;
wire n11122;
wire n11123;
wire n11124;
wire n11125;
wire n11126;
wire n11127;
wire n11128;
wire n11129;
wire n11130;
wire n11131;
wire n11133;
wire n11134;
wire n11135;
wire n11136;
wire n11137;
wire n11138;
wire n11139;
wire n11140;
wire n11141;
wire n11142;
wire n11143;
wire n11144;
wire n11146;
wire n11147;
wire n11149;
wire n11150;
wire n11152;
wire n11154;
wire n11155;
wire n11156;
wire n11157;
wire n11158;
wire n11159;
wire n1116;
wire n11161;
wire n11162;
wire n11164;
wire n11165;
wire n11167;
wire n11168;
wire n11169;
wire n11170;
wire n11171;
wire n11172;
wire n11173;
wire n11174;
wire n11177;
wire n11178;
wire n11179;
wire n11181;
wire n11182;
wire n11184;
wire n11185;
wire n11187;
wire n11188;
wire n11189;
wire n11190;
wire n11191;
wire n11192;
wire n11193;
wire n11194;
wire n11196;
wire n11197;
wire n11198;
wire n11199;
wire n11200;
wire n11201;
wire n11202;
wire n11203;
wire n11204;
wire n11205;
wire n11206;
wire n11207;
wire n11209;
wire n1121;
wire n11210;
wire n11211;
wire n11212;
wire n11214;
wire n11215;
wire n11217;
wire n11218;
wire n11219;
wire n11220;
wire n11221;
wire n11222;
wire n11223;
wire n11224;
wire n11225;
wire n11226;
wire n11227;
wire n11229;
wire n11231;
wire n11232;
wire n11234;
wire n11235;
wire n11236;
wire n11237;
wire n11239;
wire n11240;
wire n11243;
wire n11244;
wire n11246;
wire n11247;
wire n11249;
wire n1125;
wire n11250;
wire n11251;
wire n11253;
wire n11254;
wire n11256;
wire n11257;
wire n11258;
wire n11259;
wire n11261;
wire n11262;
wire n11264;
wire n11265;
wire n11267;
wire n11268;
wire n11269;
wire n11271;
wire n11272;
wire n11274;
wire n11275;
wire n11277;
wire n11278;
wire n11279;
wire n11280;
wire n11281;
wire n11282;
wire n11283;
wire n11284;
wire n11285;
wire n11286;
wire n11287;
wire n11288;
wire n11289;
wire n11290;
wire n11291;
wire n11293;
wire n11294;
wire n11296;
wire n11298;
wire n11299;
wire n1130;
wire n11300;
wire n11301;
wire n11302;
wire n11303;
wire n11304;
wire n11305;
wire n11306;
wire n11307;
wire n11308;
wire n11309;
wire n11311;
wire n11312;
wire n11314;
wire n11315;
wire n11317;
wire n11318;
wire n11320;
wire n11321;
wire n11323;
wire n11324;
wire n11325;
wire n11326;
wire n11327;
wire n11328;
wire n11329;
wire n11330;
wire n11331;
wire n11332;
wire n11333;
wire n11334;
wire n11336;
wire n11337;
wire n11339;
wire n11340;
wire n11342;
wire n11343;
wire n11346;
wire n11347;
wire n11349;
wire n1135;
wire n11350;
wire n11352;
wire n11353;
wire n11355;
wire n11356;
wire n11358;
wire n11359;
wire n11360;
wire n11361;
wire n11362;
wire n11363;
wire n11365;
wire n11366;
wire n11367;
wire n11368;
wire n11369;
wire n11370;
wire n11371;
wire n11372;
wire n11373;
wire n11374;
wire n11375;
wire n11376;
wire n11378;
wire n11379;
wire n11380;
wire n11381;
wire n11382;
wire n11383;
wire n11384;
wire n11385;
wire n11386;
wire n11388;
wire n11389;
wire n11392;
wire n11393;
wire n11395;
wire n11396;
wire n11398;
wire n11399;
wire n1140;
wire n11401;
wire n11402;
wire n11404;
wire n11405;
wire n11407;
wire n11408;
wire n11410;
wire n11412;
wire n11413;
wire n11414;
wire n11415;
wire n11416;
wire n11417;
wire n11418;
wire n11419;
wire n11420;
wire n11421;
wire n11422;
wire n11423;
wire n11424;
wire n11425;
wire n11426;
wire n11428;
wire n11429;
wire n11431;
wire n11433;
wire n11434;
wire n11435;
wire n11436;
wire n11438;
wire n1144;
wire n11440;
wire n11441;
wire n11443;
wire n11444;
wire n11445;
wire n11447;
wire n11448;
wire n11450;
wire n11451;
wire n11453;
wire n11454;
wire n11456;
wire n11457;
wire n11458;
wire n11459;
wire n11461;
wire n11462;
wire n11463;
wire n11464;
wire n11465;
wire n11466;
wire n11467;
wire n11468;
wire n11471;
wire n11472;
wire n11474;
wire n11475;
wire n11476;
wire n11477;
wire n11478;
wire n11479;
wire n1148;
wire n11480;
wire n11481;
wire n11482;
wire n11483;
wire n11484;
wire n11485;
wire n11486;
wire n11487;
wire n11488;
wire n11489;
wire n11490;
wire n11491;
wire n11492;
wire n11494;
wire n11495;
wire n11497;
wire n11498;
wire n11499;
wire n11501;
wire n11502;
wire n11504;
wire n11505;
wire n11507;
wire n11508;
wire n11510;
wire n11511;
wire n11513;
wire n11514;
wire n11516;
wire n11517;
wire n11519;
wire n11521;
wire n11523;
wire n11524;
wire n11526;
wire n11527;
wire n11529;
wire n1153;
wire n11530;
wire n11532;
wire n11534;
wire n11536;
wire n11537;
wire n11538;
wire n11539;
wire n11540;
wire n11541;
wire n11542;
wire n11543;
wire n11544;
wire n11545;
wire n11546;
wire n11547;
wire n11548;
wire n11550;
wire n11551;
wire n11553;
wire n11554;
wire n11556;
wire n11558;
wire n11559;
wire n11561;
wire n11562;
wire n11564;
wire n11566;
wire n11567;
wire n11568;
wire n11569;
wire n11570;
wire n11571;
wire n11572;
wire n11573;
wire n11575;
wire n11576;
wire n11578;
wire n11579;
wire n1158;
wire n11580;
wire n11582;
wire n11583;
wire n11584;
wire n11585;
wire n11586;
wire n11588;
wire n11589;
wire n11591;
wire n11592;
wire n11594;
wire n11595;
wire n11597;
wire n11599;
wire n11600;
wire n11602;
wire n11603;
wire n11604;
wire n11605;
wire n11606;
wire n11608;
wire n11609;
wire n11612;
wire n11613;
wire n11615;
wire n11616;
wire n11618;
wire n11619;
wire n11621;
wire n11623;
wire n11624;
wire n11626;
wire n11627;
wire n11629;
wire n1163;
wire n11631;
wire n11633;
wire n11634;
wire n11636;
wire n11637;
wire n11639;
wire n11640;
wire n11642;
wire n11643;
wire n11645;
wire n11646;
wire n11648;
wire n11649;
wire n11651;
wire n11652;
wire n11654;
wire n11656;
wire n11658;
wire n11659;
wire n11660;
wire n11662;
wire n11663;
wire n11664;
wire n11665;
wire n11667;
wire n11668;
wire n11670;
wire n11671;
wire n11673;
wire n11674;
wire n11676;
wire n11677;
wire n11679;
wire n1168;
wire n11681;
wire n11682;
wire n11684;
wire n11686;
wire n11687;
wire n11689;
wire n11690;
wire n11692;
wire n11693;
wire n11695;
wire n11696;
wire n11698;
wire n11700;
wire n11701;
wire n11703;
wire n11704;
wire n11706;
wire n11707;
wire n11708;
wire n11710;
wire n11711;
wire n11713;
wire n11715;
wire n11716;
wire n11717;
wire n11718;
wire n11719;
wire n11720;
wire n11721;
wire n11722;
wire n11723;
wire n11724;
wire n11725;
wire n11726;
wire n11728;
wire n11729;
wire n1173;
wire n11731;
wire n11733;
wire n11734;
wire n11736;
wire n11738;
wire n11739;
wire n11741;
wire n11742;
wire n11743;
wire n11744;
wire n11745;
wire n11746;
wire n11747;
wire n11748;
wire n11749;
wire n11750;
wire n11751;
wire n11752;
wire n11754;
wire n11755;
wire n11757;
wire n11759;
wire n11760;
wire n11763;
wire n11764;
wire n11766;
wire n11767;
wire n11769;
wire n11770;
wire n11772;
wire n11773;
wire n11775;
wire n11776;
wire n11778;
wire n11779;
wire n1178;
wire n11781;
wire n11782;
wire n11783;
wire n11784;
wire n11785;
wire n11786;
wire n11787;
wire n11788;
wire n11790;
wire n11792;
wire n11793;
wire n11794;
wire n11796;
wire n11797;
wire n11799;
wire n11800;
wire n11802;
wire n11803;
wire n11805;
wire n11806;
wire n11808;
wire n11809;
wire n11811;
wire n11812;
wire n11814;
wire n11815;
wire n11816;
wire n11817;
wire n11818;
wire n11819;
wire n11820;
wire n11821;
wire n11822;
wire n11823;
wire n11824;
wire n11825;
wire n11826;
wire n11827;
wire n11828;
wire n11829;
wire n1183;
wire n11830;
wire n11831;
wire n11832;
wire n11833;
wire n11834;
wire n11836;
wire n11837;
wire n11840;
wire n11842;
wire n11843;
wire n11845;
wire n11846;
wire n11847;
wire n11848;
wire n11849;
wire n11850;
wire n11852;
wire n11853;
wire n11855;
wire n11856;
wire n11857;
wire n11858;
wire n11859;
wire n11860;
wire n11862;
wire n11863;
wire n11864;
wire n11865;
wire n11866;
wire n11867;
wire n11868;
wire n11869;
wire n1187;
wire n11870;
wire n11871;
wire n11872;
wire n11873;
wire n11875;
wire n11876;
wire n11878;
wire n11880;
wire n11881;
wire n11883;
wire n11884;
wire n11886;
wire n11887;
wire n11889;
wire n11890;
wire n11892;
wire n11893;
wire n11896;
wire n11897;
wire n11899;
wire n11900;
wire n11901;
wire n11902;
wire n11903;
wire n11904;
wire n11905;
wire n11906;
wire n11908;
wire n1191;
wire n11910;
wire n11911;
wire n11912;
wire n11913;
wire n11914;
wire n11915;
wire n11916;
wire n11917;
wire n11918;
wire n11919;
wire n11920;
wire n11921;
wire n11922;
wire n11923;
wire n11924;
wire n11926;
wire n11927;
wire n11928;
wire n11929;
wire n11930;
wire n11931;
wire n11932;
wire n11933;
wire n11934;
wire n11935;
wire n11936;
wire n11937;
wire n11939;
wire n11940;
wire n11941;
wire n11942;
wire n11943;
wire n11944;
wire n11945;
wire n11947;
wire n11948;
wire n1195;
wire n11950;
wire n11951;
wire n11953;
wire n11954;
wire n11956;
wire n11957;
wire n11959;
wire n11960;
wire n11962;
wire n11964;
wire n11965;
wire n11966;
wire n11967;
wire n11968;
wire n11969;
wire n11970;
wire n11971;
wire n11972;
wire n11974;
wire n11975;
wire n11976;
wire n11978;
wire n11979;
wire n11980;
wire n11981;
wire n11982;
wire n11984;
wire n11985;
wire n11986;
wire n11987;
wire n11989;
wire n11990;
wire n11992;
wire n11993;
wire n11995;
wire n11996;
wire n11997;
wire n11999;
wire n1200;
wire n12000;
wire n12001;
wire n12003;
wire n12004;
wire n12005;
wire n12006;
wire n12008;
wire n12009;
wire n12011;
wire n12012;
wire n12013;
wire n12014;
wire n12015;
wire n12016;
wire n12017;
wire n12018;
wire n12021;
wire n12022;
wire n12024;
wire n12025;
wire n12027;
wire n12028;
wire n12029;
wire n12030;
wire n12031;
wire n12032;
wire n12033;
wire n12034;
wire n12035;
wire n12036;
wire n12037;
wire n12038;
wire n12040;
wire n12042;
wire n12043;
wire n12045;
wire n12047;
wire n12048;
wire n1205;
wire n12050;
wire n12052;
wire n12054;
wire n12055;
wire n12057;
wire n12059;
wire n12060;
wire n12061;
wire n12062;
wire n12063;
wire n12064;
wire n12065;
wire n12066;
wire n12068;
wire n12069;
wire n12071;
wire n12072;
wire n12073;
wire n12074;
wire n12075;
wire n12077;
wire n12078;
wire n12079;
wire n12080;
wire n12082;
wire n12083;
wire n12084;
wire n12085;
wire n12086;
wire n12087;
wire n12088;
wire n12089;
wire n12090;
wire n12091;
wire n12092;
wire n12093;
wire n12094;
wire n12096;
wire n12097;
wire n12099;
wire n1210;
wire n12100;
wire n12102;
wire n12103;
wire n12105;
wire n12106;
wire n12108;
wire n12109;
wire n12110;
wire n12111;
wire n12112;
wire n12113;
wire n12114;
wire n12115;
wire n12116;
wire n12117;
wire n12118;
wire n12119;
wire n12121;
wire n1214;
wire n1219;
wire n1224;
wire n1228;
wire n1232;
wire n1236;
wire n1240;
wire n1244;
wire n1248;
wire n1253;
wire n1258;
wire n1262;
wire n1267;
wire n1272;
wire n1277;
wire n1282;
wire n1287;
wire n1291;
wire n1295;
wire n1300;
wire n1305;
wire n1309;
wire n1314;
wire n1318;
wire n1322;
wire n1326;
wire n1331;
wire n1335;
wire n1340;
wire n1345;
wire n1350;
wire n1355;
wire n1359;
wire n1363;
wire n1368;
wire n1373;
wire n1378;
wire n1383;
wire n1386;
wire n1391;
wire n1396;
wire n1400;
wire n1405;
wire n1410;
wire n1414;
wire n1419;
wire n1423;
wire n1428;
wire n1433;
wire n1438;
wire n1442;
wire n1446;
wire n1451;
wire n1455;
wire n1460;
wire n1465;
wire n1469;
wire n1474;
wire n1478;
wire n1482;
wire n1487;
wire n1491;
wire n1496;
wire n1501;
wire n1506;
wire n1510;
wire n1515;
wire n1519;
wire n1524;
wire n1528;
wire n1533;
wire n1538;
wire n1542;
wire n1546;
wire n1551;
wire n1555;
wire n1560;
wire n1564;
wire n1568;
wire n1572;
wire n1577;
wire n1582;
wire n1587;
wire n1591;
wire n1596;
wire n1600;
wire n1605;
wire n1610;
wire n1615;
wire n1619;
wire n1624;
wire n1629;
wire n1634;
wire n1639;
wire n1644;
wire n1649;
wire n1653;
wire n1658;
wire n1663;
wire n1668;
wire n1673;
wire n1677;
wire n1681;
wire n1686;
wire n1691;
wire n1696;
wire n1701;
wire n1704;
wire n1709;
wire n1714;
wire n1718;
wire n1722;
wire n1727;
wire n1732;
wire n1737;
wire n1742;
wire n1747;
wire n1752;
wire n1756;
wire n1761;
wire n1765;
wire n1770;
wire n1775;
wire n1779;
wire n1782;
wire n1787;
wire n1792;
wire n1797;
wire n1802;
wire n1807;
wire n1812;
wire n1817;
wire n1822;
wire n1827;
wire n1832;
wire n1836;
wire n1841;
wire n1846;
wire n1851;
wire n1855;
wire n1860;
wire n1865;
wire n1869;
wire n1874;
wire n1878;
wire n1883;
wire n1888;
wire n1893;
wire n1898;
wire n1903;
wire n1908;
wire n1913;
wire n1918;
wire n1922;
wire n1927;
wire n1932;
wire n1936;
wire n1941;
wire n1945;
wire n1950;
wire n1954;
wire n1959;
wire n1964;
wire n1969;
wire n1973;
wire n1978;
wire n1983;
wire n1988;
wire n1993;
wire n1998;
wire n2002;
wire n2007;
wire n2011;
wire n2016;
wire n2021;
wire n2026;
wire n2031;
wire n2036;
wire n2041;
wire n2046;
wire n2051;
wire n2055;
wire n2060;
wire n2065;
wire n2070;
wire n2074;
wire n2079;
wire n2084;
wire n2088;
wire n2093;
wire n2098;
wire n2102;
wire n2106;
wire n2111;
wire n2115;
wire n2119;
wire n2122;
wire n2127;
wire n2132;
wire n2136;
wire n2140;
wire n2144;
wire n2149;
wire n2152;
wire n2157;
wire n2162;
wire n2167;
wire n2172;
wire n2177;
wire n2181;
wire n2186;
wire n2189;
wire n2194;
wire n2199;
wire n2203;
wire n2208;
wire n2213;
wire n2218;
wire n2222;
wire n2227;
wire n2232;
wire n2237;
wire n2242;
wire n2247;
wire n2251;
wire n2256;
wire n2260;
wire n2265;
wire n2270;
wire n2275;
wire n2280;
wire n2284;
wire n2288;
wire n2293;
wire n2298;
wire n2303;
wire n2307;
wire n2312;
wire n2316;
wire n2321;
wire n2324;
wire n2329;
wire n2334;
wire n2338;
wire n2342;
wire n2347;
wire n2350;
wire n2355;
wire n2360;
wire n2365;
wire n2370;
wire n2373;
wire n2377;
wire n2381;
wire n2386;
wire n2391;
wire n2395;
wire n2399;
wire n2404;
wire n2409;
wire n2414;
wire n2417;
wire n2422;
wire n2426;
wire n2430;
wire n2435;
wire n2440;
wire n2444;
wire n2448;
wire n2452;
wire n2457;
wire n2462;
wire n2465;
wire n2470;
wire n2474;
wire n2479;
wire n2484;
wire n2488;
wire n2493;
wire n2496;
wire n2500;
wire n2505;
wire n2510;
wire n2515;
wire n2519;
wire n2524;
wire n2529;
wire n2534;
wire n2539;
wire n2543;
wire n2547;
wire n2552;
wire n2556;
wire n2561;
wire n2566;
wire n2570;
wire n2575;
wire n2580;
wire n2585;
wire n2590;
wire n2594;
wire n2597;
wire n2601;
wire n2605;
wire n2610;
wire n2615;
wire n2618;
wire n2622;
wire n2627;
wire n2632;
wire n2637;
wire n2642;
wire n2647;
wire n2651;
wire n2656;
wire n266;
wire n2660;
wire n2665;
wire n2670;
wire n2675;
wire n2679;
wire n2682;
wire n2687;
wire n2692;
wire n2696;
wire n2701;
wire n2705;
wire n2709;
wire n271;
wire n2713;
wire n2718;
wire n2723;
wire n2727;
wire n2732;
wire n2737;
wire n2741;
wire n2745;
wire n2748;
wire n2753;
wire n2758;
wire n276;
wire n2762;
wire n2767;
wire n2771;
wire n2776;
wire n2781;
wire n2784;
wire n2788;
wire n2792;
wire n2797;
wire n2801;
wire n2805;
wire n281;
wire n2810;
wire n2814;
wire n2819;
wire n2823;
wire n2827;
wire n2831;
wire n2836;
wire n2840;
wire n2845;
wire n2850;
wire n2855;
wire n286;
wire n2860;
wire n2864;
wire n2869;
wire n2873;
wire n2877;
wire n2882;
wire n2885;
wire n2890;
wire n2895;
wire n2900;
wire n2904;
wire n2908;
wire n291;
wire n2913;
wire n2918;
wire n2922;
wire n2926;
wire n2930;
wire n2935;
wire n2939;
wire n2944;
wire n2948;
wire n295;
wire n2953;
wire n2958;
wire n2963;
wire n2967;
wire n2972;
wire n2976;
wire n2981;
wire n2986;
wire n2991;
wire n2996;
wire n300;
wire n3000;
wire n3005;
wire n3010;
wire n3015;
wire n3020;
wire n3025;
wire n3030;
wire n3033;
wire n3037;
wire n3042;
wire n3047;
wire n305;
wire n3052;
wire n3056;
wire n3061;
wire n3065;
wire n3069;
wire n3074;
wire n3078;
wire n3082;
wire n3087;
wire n3092;
wire n3097;
wire n310;
wire n3102;
wire n3105;
wire n3110;
wire n3114;
wire n3117;
wire n3121;
wire n3126;
wire n3130;
wire n3134;
wire n3139;
wire n314;
wire n3143;
wire n3148;
wire n3152;
wire n3157;
wire n3162;
wire n3165;
wire n3170;
wire n3174;
wire n3178;
wire n3182;
wire n3186;
wire n319;
wire n3190;
wire n3194;
wire n3199;
wire n3203;
wire n3207;
wire n3212;
wire n3217;
wire n3222;
wire n3226;
wire n3231;
wire n3235;
wire n324;
wire n3240;
wire n3244;
wire n3249;
wire n3254;
wire n3258;
wire n3263;
wire n3268;
wire n3272;
wire n3276;
wire n3280;
wire n3285;
wire n329;
wire n3290;
wire n3294;
wire n3299;
wire n3303;
wire n3308;
wire n3313;
wire n3318;
wire n3322;
wire n3325;
wire n3330;
wire n3333;
wire n3338;
wire n334;
wire n3343;
wire n3348;
wire n3352;
wire n3356;
wire n3361;
wire n3365;
wire n3370;
wire n3374;
wire n3379;
wire n3383;
wire n3386;
wire n339;
wire n3390;
wire n3395;
wire n3400;
wire n3404;
wire n3408;
wire n3413;
wire n3418;
wire n3422;
wire n3427;
wire n3431;
wire n3436;
wire n344;
wire n3440;
wire n3445;
wire n3450;
wire n3455;
wire n3459;
wire n3464;
wire n3469;
wire n3474;
wire n3479;
wire n3484;
wire n3489;
wire n349;
wire n3494;
wire n3497;
wire n3502;
wire n3507;
wire n3511;
wire n3516;
wire n352;
wire n3520;
wire n3524;
wire n3528;
wire n3532;
wire n3537;
wire n3542;
wire n3546;
wire n3551;
wire n3555;
wire n3559;
wire n3564;
wire n3567;
wire n357;
wire n3572;
wire n3577;
wire n3582;
wire n3587;
wire n3590;
wire n3595;
wire n3600;
wire n3604;
wire n3609;
wire n361;
wire n3614;
wire n3618;
wire n3623;
wire n3628;
wire n3633;
wire n3638;
wire n3642;
wire n3647;
wire n3651;
wire n3655;
wire n3658;
wire n366;
wire n3661;
wire n3666;
wire n3670;
wire n3675;
wire n3679;
wire n3684;
wire n3689;
wire n3693;
wire n3698;
wire n370;
wire n3703;
wire n3707;
wire n3711;
wire n3716;
wire n3720;
wire n3725;
wire n3729;
wire n3733;
wire n3737;
wire n3742;
wire n3747;
wire n375;
wire n3752;
wire n3756;
wire n3761;
wire n3765;
wire n3770;
wire n3773;
wire n3777;
wire n3782;
wire n3787;
wire n3791;
wire n3796;
wire n380;
wire n3801;
wire n3805;
wire n3809;
wire n3813;
wire n3817;
wire n3822;
wire n3827;
wire n3831;
wire n3836;
wire n3841;
wire n3846;
wire n385;
wire n3851;
wire n3855;
wire n3859;
wire n3864;
wire n3867;
wire n3872;
wire n3877;
wire n3881;
wire n3886;
wire n3891;
wire n3896;
wire n3899;
wire n390;
wire n3904;
wire n3908;
wire n3913;
wire n3917;
wire n3922;
wire n3927;
wire n3932;
wire n3936;
wire n3941;
wire n3945;
wire n3949;
wire n395;
wire n3953;
wire n3957;
wire n3962;
wire n3967;
wire n3972;
wire n3976;
wire n3981;
wire n3985;
wire n3989;
wire n3993;
wire n3998;
wire n400;
wire n4002;
wire n4007;
wire n4011;
wire n4016;
wire n4020;
wire n4024;
wire n4029;
wire n4033;
wire n4037;
wire n4042;
wire n4046;
wire n405;
wire n4051;
wire n4055;
wire n4059;
wire n4063;
wire n4068;
wire n4071;
wire n4075;
wire n4079;
wire n4084;
wire n4089;
wire n4094;
wire n4098;
wire n410;
wire n4102;
wire n4107;
wire n4112;
wire n4116;
wire n4121;
wire n4126;
wire n4131;
wire n4135;
wire n4140;
wire n4145;
wire n4148;
wire n415;
wire n4153;
wire n4158;
wire n4161;
wire n4166;
wire n4171;
wire n4176;
wire n4181;
wire n4186;
wire n4191;
wire n4194;
wire n4199;
wire n420;
wire n4203;
wire n4207;
wire n4212;
wire n4217;
wire n4221;
wire n4226;
wire n4231;
wire n4235;
wire n424;
wire n4240;
wire n4245;
wire n4249;
wire n4253;
wire n4258;
wire n4263;
wire n4267;
wire n4271;
wire n4276;
wire n4280;
wire n4284;
wire n4289;
wire n429;
wire n4294;
wire n4299;
wire n4304;
wire n4309;
wire n4313;
wire n4318;
wire n4322;
wire n4326;
wire n4330;
wire n4333;
wire n4338;
wire n434;
wire n4343;
wire n4348;
wire n4352;
wire n4357;
wire n4362;
wire n4365;
wire n4370;
wire n4374;
wire n4379;
wire n438;
wire n4384;
wire n4388;
wire n4392;
wire n4397;
wire n4401;
wire n4405;
wire n4410;
wire n4414;
wire n4419;
wire n4424;
wire n4428;
wire n443;
wire n4433;
wire n4438;
wire n4443;
wire n4448;
wire n4451;
wire n4456;
wire n4459;
wire n4464;
wire n4469;
wire n447;
wire n4473;
wire n4478;
wire n4482;
wire n4487;
wire n4491;
wire n4496;
wire n4501;
wire n4505;
wire n451;
wire n4510;
wire n4515;
wire n4520;
wire n4524;
wire n4529;
wire n4534;
wire n4539;
wire n4544;
wire n4548;
wire n455;
wire n4553;
wire n4558;
wire n4562;
wire n4567;
wire n4572;
wire n4577;
wire n4581;
wire n4586;
wire n4591;
wire n4596;
wire n460;
wire n4600;
wire n4604;
wire n4609;
wire n4613;
wire n4617;
wire n4622;
wire n4627;
wire n4631;
wire n4636;
wire n4641;
wire n4646;
wire n465;
wire n4651;
wire n4656;
wire n4660;
wire n4665;
wire n4669;
wire n4673;
wire n4678;
wire n4681;
wire n4686;
wire n4690;
wire n4694;
wire n4699;
wire n470;
wire n4703;
wire n4708;
wire n4713;
wire n4717;
wire n4722;
wire n4727;
wire n4732;
wire n4737;
wire n474;
wire n4742;
wire n4745;
wire n4750;
wire n4755;
wire n4760;
wire n4765;
wire n4769;
wire n4774;
wire n4778;
wire n4782;
wire n4787;
wire n479;
wire n4791;
wire n4795;
wire n4800;
wire n4805;
wire n4809;
wire n4814;
wire n4818;
wire n4822;
wire n4827;
wire n4831;
wire n4834;
wire n4838;
wire n484;
wire n4843;
wire n4848;
wire n4853;
wire n4857;
wire n4862;
wire n4867;
wire n4872;
wire n4877;
wire n488;
wire n4881;
wire n4886;
wire n4890;
wire n4895;
wire n4899;
wire n4904;
wire n4908;
wire n4913;
wire n4917;
wire n4922;
wire n4927;
wire n493;
wire n4931;
wire n4936;
wire n4940;
wire n4944;
wire n4947;
wire n4952;
wire n4957;
wire n4961;
wire n4965;
wire n4969;
wire n4974;
wire n4979;
wire n498;
wire n4983;
wire n4987;
wire n4992;
wire n4996;
wire n5001;
wire n5005;
wire n5008;
wire n5013;
wire n5018;
wire n5023;
wire n5027;
wire n503;
wire n5031;
wire n5035;
wire n5040;
wire n5045;
wire n5048;
wire n5053;
wire n5056;
wire n5061;
wire n5066;
wire n5070;
wire n5075;
wire n508;
wire n5080;
wire n5085;
wire n5090;
wire n5094;
wire n5098;
wire n5103;
wire n5107;
wire n5112;
wire n5117;
wire n5121;
wire n5126;
wire n513;
wire n5130;
wire n5134;
wire n5139;
wire n5143;
wire n5148;
wire n5151;
wire n5156;
wire n5159;
wire n5164;
wire n5169;
wire n5173;
wire n5178;
wire n518;
wire n5181;
wire n5186;
wire n5189;
wire n5193;
wire n5198;
wire n5202;
wire n5207;
wire n5212;
wire n5217;
wire n5221;
wire n5225;
wire n523;
wire n5230;
wire n5234;
wire n5239;
wire n5242;
wire n5246;
wire n5251;
wire n5256;
wire n5261;
wire n5265;
wire n5269;
wire n5274;
wire n5279;
wire n528;
wire n5284;
wire n5288;
wire n5293;
wire n5298;
wire n5302;
wire n5307;
wire n5312;
wire n5316;
wire n5321;
wire n5326;
wire n533;
wire n5330;
wire n5335;
wire n5339;
wire n5344;
wire n5349;
wire n5353;
wire n5358;
wire n5362;
wire n5366;
wire n5370;
wire n5375;
wire n538;
wire n5380;
wire n5383;
wire n5388;
wire n5393;
wire n5397;
wire n5402;
wire n5406;
wire n5411;
wire n5415;
wire n5420;
wire n5424;
wire n5429;
wire n543;
wire n5433;
wire n5437;
wire n5441;
wire n5446;
wire n5451;
wire n5455;
wire n5460;
wire n5464;
wire n5469;
wire n5472;
wire n5477;
wire n548;
wire n5481;
wire n5486;
wire n5490;
wire n5495;
wire n5500;
wire n5504;
wire n5508;
wire n5513;
wire n5517;
wire n5521;
wire n5525;
wire n5529;
wire n553;
wire n5534;
wire n5539;
wire n5543;
wire n5547;
wire n5552;
wire n5556;
wire n556;
wire n5560;
wire n5565;
wire n5570;
wire n5575;
wire n5579;
wire n5584;
wire n5588;
wire n5591;
wire n5596;
wire n5601;
wire n5606;
wire n561;
wire n5610;
wire n5613;
wire n5618;
wire n5623;
wire n5628;
wire n5633;
wire n5638;
wire n5643;
wire n5648;
wire n5651;
wire n5655;
wire n566;
wire n5660;
wire n5664;
wire n5669;
wire n5674;
wire n5679;
wire n5682;
wire n5686;
wire n5691;
wire n5696;
wire n5700;
wire n5704;
wire n5709;
wire n571;
wire n5713;
wire n5717;
wire n5722;
wire n5727;
wire n5731;
wire n5735;
wire n5739;
wire n5744;
wire n5748;
wire n5753;
wire n5758;
wire n576;
wire n5763;
wire n5767;
wire n5771;
wire n5775;
wire n5779;
wire n5783;
wire n5787;
wire n5792;
wire n5796;
wire n580;
wire n5801;
wire n5805;
wire n5809;
wire n5814;
wire n5819;
wire n5824;
wire n5828;
wire n5833;
wire n5836;
wire n5840;
wire n5845;
wire n585;
wire n5850;
wire n5855;
wire n5860;
wire n5864;
wire n5867;
wire n5872;
wire n5876;
wire n5881;
wire n5885;
wire n5890;
wire n5894;
wire n5899;
wire n590;
wire n5903;
wire n5908;
wire n5912;
wire n5917;
wire n5920;
wire n5925;
wire n5930;
wire n5934;
wire n5938;
wire n5943;
wire n5947;
wire n595;
wire n5951;
wire n5955;
wire n5960;
wire n5964;
wire n5968;
wire n5973;
wire n5978;
wire n5982;
wire n5987;
wire n5992;
wire n5997;
wire n600;
wire n6002;
wire n6006;
wire n6009;
wire n6014;
wire n6019;
wire n6024;
wire n6029;
wire n6034;
wire n6038;
wire n6043;
wire n6047;
wire n605;
wire n6052;
wire n6056;
wire n6061;
wire n6066;
wire n6069;
wire n6074;
wire n6078;
wire n6083;
wire n6088;
wire n6093;
wire n6098;
wire n610;
wire n6102;
wire n6106;
wire n6110;
wire n6114;
wire n6119;
wire n6124;
wire n6128;
wire n6132;
wire n6136;
wire n6140;
wire n6145;
wire n6148;
wire n615;
wire n6153;
wire n6158;
wire n6161;
wire n6166;
wire n6171;
wire n6176;
wire n6181;
wire n6186;
wire n6191;
wire n6195;
wire n620;
wire n6200;
wire n6204;
wire n6209;
wire n6214;
wire n6218;
wire n6222;
wire n6227;
wire n6231;
wire n6235;
wire n6239;
wire n6244;
wire n6249;
wire n625;
wire n6254;
wire n6258;
wire n6261;
wire n6266;
wire n6271;
wire n6276;
wire n6281;
wire n6285;
wire n629;
wire n6290;
wire n6294;
wire n6299;
wire n6302;
wire n6306;
wire n6311;
wire n6316;
wire n6319;
wire n6324;
wire n6329;
wire n6332;
wire n6337;
wire n634;
wire n6342;
wire n6346;
wire n6350;
wire n6354;
wire n6357;
wire n6362;
wire n6367;
wire n6371;
wire n6376;
wire n6381;
wire n6386;
wire n639;
wire n6390;
wire n6395;
wire n6399;
wire n6403;
wire n6407;
wire n6411;
wire n6415;
wire n6419;
wire n6423;
wire n6427;
wire n6432;
wire n6437;
wire n644;
wire n6441;
wire n6446;
wire n6450;
wire n6455;
wire n6460;
wire n6464;
wire n6469;
wire n6472;
wire n6477;
wire n6480;
wire n6485;
wire n6489;
wire n649;
wire n6493;
wire n6498;
wire n6502;
wire n6507;
wire n6511;
wire n6515;
wire n6519;
wire n6522;
wire n6527;
wire n6531;
wire n6535;
wire n654;
wire n6540;
wire n6545;
wire n6550;
wire n6554;
wire n6558;
wire n6563;
wire n6566;
wire n6570;
wire n6574;
wire n6578;
wire n6583;
wire n6586;
wire n659;
wire n6591;
wire n6596;
wire n6601;
wire n6606;
wire n6611;
wire n6615;
wire n6619;
wire n6624;
wire n6629;
wire n6634;
wire n6638;
wire n664;
wire n6643;
wire n6648;
wire n6652;
wire n6656;
wire n6661;
wire n6665;
wire n6669;
wire n6674;
wire n6678;
wire n6682;
wire n6687;
wire n669;
wire n6691;
wire n6695;
wire n6700;
wire n6704;
wire n6709;
wire n6713;
wire n6717;
wire n6722;
wire n6727;
wire n673;
wire n6730;
wire n6731;
wire n6732;
wire n6733;
wire n6734;
wire n6735;
wire n6736;
wire n6736_1;
wire n6737;
wire n6738;
wire n6739;
wire n6740;
wire n6741;
wire n6742;
wire n6743;
wire n6745;
wire n6746;
wire n6746_1;
wire n6747;
wire n6748;
wire n6749;
wire n6749_1;
wire n6750;
wire n6751;
wire n6752;
wire n6752_1;
wire n6753;
wire n6754;
wire n6755;
wire n6756;
wire n6756_1;
wire n6757;
wire n6758;
wire n6759;
wire n6760;
wire n6761;
wire n6761_1;
wire n6762;
wire n6763;
wire n6764;
wire n6765;
wire n6765_1;
wire n6766;
wire n6767;
wire n6768;
wire n6769;
wire n6770;
wire n6770_1;
wire n6771;
wire n6772;
wire n6773;
wire n6774;
wire n6774_1;
wire n6775;
wire n6776;
wire n6777;
wire n6778;
wire n6779;
wire n6779_1;
wire n678;
wire n6780;
wire n6781;
wire n6782;
wire n6783;
wire n6783_1;
wire n6784;
wire n6785;
wire n6786;
wire n6787;
wire n6788;
wire n6788_1;
wire n6789;
wire n6790;
wire n6791;
wire n6792;
wire n6793;
wire n6793_1;
wire n6794;
wire n6795;
wire n6796;
wire n6796_1;
wire n6797;
wire n6799;
wire n6800;
wire n6801;
wire n6801_1;
wire n6802;
wire n6803;
wire n6804;
wire n6806;
wire n6806_1;
wire n6807;
wire n6808;
wire n6809;
wire n6809_1;
wire n6810;
wire n6811;
wire n6812;
wire n6813;
wire n6813_1;
wire n6814;
wire n6815;
wire n6816;
wire n6817;
wire n6818;
wire n6818_1;
wire n6819;
wire n6820;
wire n6821;
wire n6822;
wire n6822_1;
wire n6823;
wire n6824;
wire n6825;
wire n6826;
wire n6826_1;
wire n6827;
wire n6828;
wire n6829;
wire n683;
wire n6830;
wire n6831;
wire n6831_1;
wire n6832;
wire n6833;
wire n6834;
wire n6835;
wire n6836;
wire n6836_1;
wire n6837;
wire n6838;
wire n6839;
wire n6840;
wire n6840_1;
wire n6841;
wire n6842;
wire n6843;
wire n6844;
wire n6845;
wire n6845_1;
wire n6846;
wire n6847;
wire n6848;
wire n6849;
wire n6850;
wire n6850_1;
wire n6851;
wire n6852;
wire n6853;
wire n6854;
wire n6855;
wire n6855_1;
wire n6856;
wire n6857;
wire n6859;
wire n6860;
wire n6860_1;
wire n6861;
wire n6862;
wire n6863;
wire n6863_1;
wire n6864;
wire n6865;
wire n6866;
wire n6867;
wire n6867_1;
wire n6868;
wire n6869;
wire n6870;
wire n6871;
wire n6872;
wire n6872_1;
wire n6873;
wire n6875;
wire n6876;
wire n6876_1;
wire n6877;
wire n6878;
wire n6879;
wire n688;
wire n6880;
wire n6881;
wire n6881_1;
wire n6882;
wire n6884;
wire n6885;
wire n6886;
wire n6886_1;
wire n6888;
wire n6889;
wire n6890;
wire n6890_1;
wire n6891;
wire n6892;
wire n6894;
wire n6895;
wire n6895_1;
wire n6896;
wire n6897;
wire n6898;
wire n6899;
wire n6899_1;
wire n6900;
wire n6901;
wire n6902;
wire n6902_1;
wire n6903;
wire n6904;
wire n6905;
wire n6906;
wire n6907;
wire n6908;
wire n6910;
wire n6910_1;
wire n6912;
wire n6913;
wire n6914;
wire n6915;
wire n6915_1;
wire n6916;
wire n6917;
wire n6918;
wire n6919;
wire n6919_1;
wire n6920;
wire n6921;
wire n6922;
wire n6923;
wire n6924;
wire n6924_1;
wire n6925;
wire n6926;
wire n6927;
wire n6928;
wire n6929;
wire n6929_1;
wire n693;
wire n6930;
wire n6931;
wire n6932;
wire n6933;
wire n6934;
wire n6934_1;
wire n6935;
wire n6936;
wire n6937;
wire n6938;
wire n6938_1;
wire n6939;
wire n6940;
wire n6941;
wire n6942;
wire n6943;
wire n6943_1;
wire n6944;
wire n6945;
wire n6946;
wire n6947;
wire n6947_1;
wire n6948;
wire n6949;
wire n6950;
wire n6951;
wire n6952;
wire n6952_1;
wire n6953;
wire n6954;
wire n6955;
wire n6956;
wire n6957;
wire n6958;
wire n6959;
wire n6960;
wire n6960_1;
wire n6961;
wire n6962;
wire n6963;
wire n6964;
wire n6964_1;
wire n6965;
wire n6966;
wire n6967;
wire n6968;
wire n6969;
wire n6969_1;
wire n6970;
wire n6971;
wire n6972;
wire n6974;
wire n6974_1;
wire n6976;
wire n6977;
wire n6977_1;
wire n6978;
wire n6979;
wire n698;
wire n6980;
wire n6981;
wire n6982;
wire n6982_1;
wire n6983;
wire n6984;
wire n6985;
wire n6986;
wire n6986_1;
wire n6987;
wire n6988;
wire n6989;
wire n6990;
wire n6990_1;
wire n6991;
wire n6992;
wire n6993;
wire n6994;
wire n6995;
wire n6995_1;
wire n6996;
wire n6997;
wire n6998;
wire n6999;
wire n7000;
wire n7000_1;
wire n7001;
wire n7002;
wire n7003;
wire n7004;
wire n7005;
wire n7005_1;
wire n7006;
wire n7007;
wire n7008;
wire n7009;
wire n7009_1;
wire n7010;
wire n7011;
wire n7012;
wire n7013;
wire n7013_1;
wire n7014;
wire n7015;
wire n7016;
wire n7017;
wire n7018;
wire n7018_1;
wire n7019;
wire n7020;
wire n7021;
wire n7022;
wire n7023;
wire n7023_1;
wire n7025;
wire n7026;
wire n7027;
wire n7027_1;
wire n7028;
wire n7029;
wire n703;
wire n7030;
wire n7031;
wire n7032;
wire n7032_1;
wire n7033;
wire n7034;
wire n7036;
wire n7036_1;
wire n7037;
wire n7038;
wire n7039;
wire n7040;
wire n7041;
wire n7041_1;
wire n7042;
wire n7043;
wire n7044;
wire n7045;
wire n7045_1;
wire n7046;
wire n7047;
wire n7048;
wire n7049;
wire n7049_1;
wire n7050;
wire n7051;
wire n7052;
wire n7053;
wire n7053_1;
wire n7054;
wire n7055;
wire n7056;
wire n7057;
wire n7058;
wire n7058_1;
wire n7059;
wire n7060;
wire n7061;
wire n7062;
wire n7062_1;
wire n7063;
wire n7064;
wire n7065;
wire n7067;
wire n7067_1;
wire n7069;
wire n7071;
wire n7072;
wire n7072_1;
wire n7073;
wire n7074;
wire n7075;
wire n7076;
wire n7077;
wire n7077_1;
wire n7078;
wire n7079;
wire n708;
wire n7080;
wire n7081;
wire n7082;
wire n7082_1;
wire n7083;
wire n7084;
wire n7085;
wire n7085_1;
wire n7086;
wire n7087;
wire n7088;
wire n7089;
wire n7089_1;
wire n7090;
wire n7091;
wire n7092;
wire n7093;
wire n7093_1;
wire n7094;
wire n7095;
wire n7096;
wire n7097;
wire n7098;
wire n7098_1;
wire n7099;
wire n7100;
wire n7101;
wire n7102;
wire n7102_1;
wire n7103;
wire n7105;
wire n7106;
wire n7107;
wire n7107_1;
wire n7108;
wire n7109;
wire n7110;
wire n7111;
wire n7111_1;
wire n7112;
wire n7113;
wire n7114;
wire n7116;
wire n7116_1;
wire n7117;
wire n7118;
wire n7119;
wire n7120;
wire n7120_1;
wire n7121;
wire n7122;
wire n7123;
wire n7124;
wire n7125;
wire n7125_1;
wire n7126;
wire n7127;
wire n7128;
wire n7128_1;
wire n7129;
wire n713;
wire n7130;
wire n7131;
wire n7132;
wire n7133;
wire n7133_1;
wire n7134;
wire n7135;
wire n7136;
wire n7137;
wire n7138;
wire n7138_1;
wire n7140;
wire n7141;
wire n7142;
wire n7142_1;
wire n7143;
wire n7144;
wire n7145;
wire n7147;
wire n7147_1;
wire n7148;
wire n7149;
wire n7150;
wire n7151;
wire n7151_1;
wire n7153;
wire n7154;
wire n7155;
wire n7155_1;
wire n7156;
wire n7158;
wire n7159;
wire n7160;
wire n7160_1;
wire n7161;
wire n7162;
wire n7163;
wire n7164;
wire n7164_1;
wire n7165;
wire n7166;
wire n7167;
wire n7167_1;
wire n7168;
wire n7169;
wire n7171;
wire n7172;
wire n7173;
wire n7175;
wire n7177;
wire n7177_1;
wire n7178;
wire n7179;
wire n718;
wire n7180;
wire n7181;
wire n7182;
wire n7182_1;
wire n7183;
wire n7184;
wire n7185;
wire n7186;
wire n7188;
wire n7190;
wire n7190_1;
wire n7191;
wire n7193;
wire n7194;
wire n7194_1;
wire n7195;
wire n7196;
wire n7197;
wire n7198;
wire n7199;
wire n7199_1;
wire n7200;
wire n7201;
wire n7203;
wire n7203_1;
wire n7205;
wire n7206;
wire n7207;
wire n7207_1;
wire n7208;
wire n7210;
wire n7211;
wire n7212;
wire n7212_1;
wire n7213;
wire n7214;
wire n7215;
wire n7216;
wire n7216_1;
wire n7217;
wire n7218;
wire n7219;
wire n722;
wire n7220;
wire n7221;
wire n7221_1;
wire n7223;
wire n7224;
wire n7225;
wire n7226;
wire n7226_1;
wire n7227;
wire n7228;
wire n7229;
wire n7230;
wire n7230_1;
wire n7232;
wire n7234;
wire n7235;
wire n7235_1;
wire n7237;
wire n7239;
wire n7240;
wire n7240_1;
wire n7241;
wire n7242;
wire n7243;
wire n7245;
wire n7245_1;
wire n7246;
wire n7248;
wire n7249;
wire n7250;
wire n7252;
wire n7252_1;
wire n7253;
wire n7254;
wire n7255;
wire n7256;
wire n7256_1;
wire n7257;
wire n7259;
wire n7260;
wire n7260_1;
wire n7261;
wire n7262;
wire n7263;
wire n7264;
wire n7265;
wire n7265_1;
wire n7266;
wire n7267;
wire n7268;
wire n7269;
wire n727;
wire n7270;
wire n7270_1;
wire n7271;
wire n7272;
wire n7273;
wire n7274;
wire n7275;
wire n7276;
wire n7278;
wire n7279;
wire n7280;
wire n7281;
wire n7282;
wire n7283;
wire n7284;
wire n7284_1;
wire n7285;
wire n7286;
wire n7287;
wire n7288;
wire n7288_1;
wire n7289;
wire n7290;
wire n7291;
wire n7292;
wire n7292_1;
wire n7293;
wire n7294;
wire n7295;
wire n7296;
wire n7297;
wire n7297_1;
wire n7298;
wire n7299;
wire n7300;
wire n7301;
wire n7302;
wire n7302_1;
wire n7303;
wire n7304;
wire n7305;
wire n7306;
wire n7307;
wire n7307_1;
wire n7308;
wire n7309;
wire n7310;
wire n7311;
wire n7312;
wire n7312_1;
wire n7313;
wire n7315;
wire n7316;
wire n7316_1;
wire n7318;
wire n7319;
wire n732;
wire n7321;
wire n7321_1;
wire n7322;
wire n7323;
wire n7324;
wire n7325;
wire n7326;
wire n7326_1;
wire n7327;
wire n7328;
wire n7330;
wire n7330_1;
wire n7331;
wire n7332;
wire n7334;
wire n7335;
wire n7335_1;
wire n7336;
wire n7337;
wire n7338;
wire n7339;
wire n7340;
wire n7340_1;
wire n7341;
wire n7342;
wire n7343;
wire n7344;
wire n7345;
wire n7346;
wire n7347;
wire n7348;
wire n7349;
wire n7349_1;
wire n7351;
wire n7353;
wire n7354;
wire n7354_1;
wire n7355;
wire n7356;
wire n7357;
wire n7358;
wire n7359;
wire n7359_1;
wire n736;
wire n7360;
wire n7361;
wire n7362;
wire n7363;
wire n7363_1;
wire n7365;
wire n7366;
wire n7368;
wire n7368_1;
wire n7369;
wire n7371;
wire n7372;
wire n7372_1;
wire n7374;
wire n7375;
wire n7376;
wire n7377;
wire n7378;
wire n7381;
wire n7381_1;
wire n7382;
wire n7384;
wire n7385;
wire n7386;
wire n7386_1;
wire n7387;
wire n7388;
wire n7390;
wire n7391;
wire n7391_1;
wire n7392;
wire n7393;
wire n7394;
wire n7395;
wire n7396;
wire n7397;
wire n7398;
wire n7399;
wire n7400;
wire n7400_1;
wire n7401;
wire n7402;
wire n7403;
wire n7404;
wire n7404_1;
wire n7406;
wire n7407;
wire n7408;
wire n7408_1;
wire n7409;
wire n741;
wire n7410;
wire n7411;
wire n7412;
wire n7413;
wire n7413_1;
wire n7414;
wire n7415;
wire n7416;
wire n7417;
wire n7417_1;
wire n7418;
wire n7419;
wire n7420;
wire n7421;
wire n7422;
wire n7422_1;
wire n7423;
wire n7425;
wire n7426;
wire n7427;
wire n7427_1;
wire n7428;
wire n7429;
wire n7431;
wire n7432;
wire n7432_1;
wire n7434;
wire n7435;
wire n7436;
wire n7437;
wire n7437_1;
wire n7438;
wire n7440;
wire n7441;
wire n7442;
wire n7443;
wire n7444;
wire n7445;
wire n7446;
wire n7446_1;
wire n7447;
wire n7448;
wire n7449;
wire n7450;
wire n7450_1;
wire n7452;
wire n7453;
wire n7454;
wire n7454_1;
wire n7456;
wire n7457;
wire n7459;
wire n7459_1;
wire n746;
wire n7460;
wire n7461;
wire n7462;
wire n7463;
wire n7463_1;
wire n7464;
wire n7465;
wire n7466;
wire n7467;
wire n7468;
wire n7468_1;
wire n7469;
wire n7470;
wire n7471;
wire n7472;
wire n7473;
wire n7473_1;
wire n7474;
wire n7475;
wire n7476;
wire n7477;
wire n7478;
wire n7478_1;
wire n7479;
wire n7480;
wire n7481;
wire n7482;
wire n7482_1;
wire n7483;
wire n7484;
wire n7485;
wire n7486;
wire n7487;
wire n7487_1;
wire n7488;
wire n7489;
wire n7490;
wire n7491;
wire n7492;
wire n7492_1;
wire n7493;
wire n7494;
wire n7495;
wire n7496;
wire n7496_1;
wire n7497;
wire n7498;
wire n7499;
wire n7501;
wire n7501_1;
wire n7502;
wire n7503;
wire n7504;
wire n7505;
wire n7505_1;
wire n7507;
wire n7509;
wire n7509_1;
wire n751;
wire n7511;
wire n7513;
wire n7513_1;
wire n7514;
wire n7516;
wire n7518;
wire n7518_1;
wire n7519;
wire n7520;
wire n7522;
wire n7522_1;
wire n7524;
wire n7525;
wire n7526;
wire n7527;
wire n7527_1;
wire n7528;
wire n7529;
wire n7530;
wire n7530_1;
wire n7531;
wire n7533;
wire n7534;
wire n7535;
wire n7535_1;
wire n7536;
wire n7537;
wire n7538;
wire n7539;
wire n7539_1;
wire n7540;
wire n7541;
wire n7542;
wire n7543;
wire n7543_1;
wire n7544;
wire n7545;
wire n7547;
wire n7548;
wire n7549;
wire n7550;
wire n7551;
wire n7552;
wire n7553;
wire n7553_1;
wire n7554;
wire n7556;
wire n7557;
wire n7558;
wire n7559;
wire n756;
wire n7560;
wire n7562;
wire n7563;
wire n7564;
wire n7565;
wire n7566;
wire n7567;
wire n7567_1;
wire n7568;
wire n7570;
wire n7571;
wire n7572;
wire n7572_1;
wire n7573;
wire n7574;
wire n7575;
wire n7576;
wire n7577;
wire n7577_1;
wire n7578;
wire n7579;
wire n7580;
wire n7581;
wire n7581_1;
wire n7582;
wire n7583;
wire n7584;
wire n7585;
wire n7586;
wire n7586_1;
wire n7587;
wire n7588;
wire n7589;
wire n7590;
wire n7591;
wire n7591_1;
wire n7592;
wire n7593;
wire n7594;
wire n7595;
wire n7596;
wire n7596_1;
wire n7597;
wire n7599;
wire n7599_1;
wire n7601;
wire n7603;
wire n7604;
wire n7604_1;
wire n7605;
wire n7606;
wire n7607;
wire n7608;
wire n7608_1;
wire n7609;
wire n761;
wire n7610;
wire n7611;
wire n7612;
wire n7613;
wire n7613_1;
wire n7614;
wire n7615;
wire n7616;
wire n7617;
wire n7618;
wire n7618_1;
wire n7619;
wire n7620;
wire n7621;
wire n7622;
wire n7623;
wire n7624;
wire n7625;
wire n7626;
wire n7626_1;
wire n7627;
wire n7629;
wire n7630;
wire n7631;
wire n7632;
wire n7633;
wire n7635;
wire n7635_1;
wire n7636;
wire n7637;
wire n7638;
wire n7639;
wire n7640;
wire n7641;
wire n7642;
wire n7643;
wire n7644;
wire n7644_1;
wire n7645;
wire n7647;
wire n7648;
wire n7649;
wire n765;
wire n7650;
wire n7652;
wire n7653;
wire n7654;
wire n7654_1;
wire n7656;
wire n7657;
wire n7658;
wire n7658_1;
wire n7659;
wire n7660;
wire n7661;
wire n7662;
wire n7663;
wire n7664;
wire n7665;
wire n7666;
wire n7666_1;
wire n7667;
wire n7668;
wire n7669;
wire n7670;
wire n7671;
wire n7671_1;
wire n7673;
wire n7674;
wire n7676;
wire n7676_1;
wire n7677;
wire n7679;
wire n7680;
wire n7681;
wire n7682;
wire n7684;
wire n7685;
wire n7686;
wire n7687;
wire n7688;
wire n7689;
wire n7690;
wire n7691;
wire n7691_1;
wire n7692;
wire n7693;
wire n7694;
wire n7695;
wire n7695_1;
wire n7696;
wire n7697;
wire n7698;
wire n7699;
wire n770;
wire n7700;
wire n7701;
wire n7702;
wire n7704;
wire n7704_1;
wire n7705;
wire n7706;
wire n7707;
wire n7708;
wire n7709;
wire n7710;
wire n7712;
wire n7713;
wire n7714;
wire n7714_1;
wire n7715;
wire n7716;
wire n7717;
wire n7718;
wire n7719;
wire n7719_1;
wire n7720;
wire n7721;
wire n7722;
wire n7723;
wire n7723_1;
wire n7724;
wire n7725;
wire n7726;
wire n7727;
wire n7728;
wire n7728_1;
wire n7729;
wire n7730;
wire n7731;
wire n7732;
wire n7732_1;
wire n7733;
wire n7734;
wire n7735;
wire n7736;
wire n7737;
wire n7737_1;
wire n7738;
wire n7739;
wire n774;
wire n7740;
wire n7741;
wire n7741_1;
wire n7742;
wire n7743;
wire n7744;
wire n7745;
wire n7746;
wire n7746_1;
wire n7747;
wire n7749;
wire n7750;
wire n7751;
wire n7751_1;
wire n7752;
wire n7753;
wire n7754;
wire n7755;
wire n7756;
wire n7756_1;
wire n7757;
wire n7758;
wire n7759;
wire n7760;
wire n7760_1;
wire n7761;
wire n7762;
wire n7763;
wire n7764;
wire n7764_1;
wire n7765;
wire n7766;
wire n7767;
wire n7768;
wire n7768_1;
wire n7769;
wire n7770;
wire n7771;
wire n7773;
wire n7773_1;
wire n7774;
wire n7776;
wire n7776_1;
wire n7777;
wire n7778;
wire n7779;
wire n7779_1;
wire n7780;
wire n7782;
wire n7784;
wire n7784_1;
wire n7785;
wire n7787;
wire n7788;
wire n7788_1;
wire n779;
wire n7790;
wire n7791;
wire n7793;
wire n7793_1;
wire n7794;
wire n7796;
wire n7797;
wire n7798;
wire n7799;
wire n7800;
wire n7801;
wire n7802;
wire n7802_1;
wire n7803;
wire n7804;
wire n7805;
wire n7806;
wire n7806_1;
wire n7807;
wire n7808;
wire n7809;
wire n7810;
wire n7810_1;
wire n7811;
wire n7812;
wire n7813;
wire n7814;
wire n7815;
wire n7815_1;
wire n7816;
wire n7817;
wire n7818;
wire n7818_1;
wire n7819;
wire n7820;
wire n7821;
wire n7822;
wire n7822_1;
wire n7823;
wire n7824;
wire n7825;
wire n7826;
wire n7826_1;
wire n7827;
wire n7828;
wire n7829;
wire n783;
wire n7830;
wire n7831;
wire n7831_1;
wire n7833;
wire n7834;
wire n7835;
wire n7836;
wire n7837;
wire n7838;
wire n7839;
wire n7840;
wire n7840_1;
wire n7841;
wire n7842;
wire n7844;
wire n7845;
wire n7845_1;
wire n7846;
wire n7847;
wire n7848;
wire n7848_1;
wire n7849;
wire n7850;
wire n7851;
wire n7852;
wire n7853;
wire n7853_1;
wire n7854;
wire n7855;
wire n7857;
wire n7858;
wire n7858_1;
wire n7859;
wire n7860;
wire n7861;
wire n7863;
wire n7863_1;
wire n7864;
wire n7866;
wire n7867;
wire n7867_1;
wire n7868;
wire n7869;
wire n7870;
wire n7871;
wire n7871_1;
wire n7872;
wire n7873;
wire n7874;
wire n7875;
wire n7877;
wire n7878;
wire n7878_1;
wire n788;
wire n7880;
wire n7881;
wire n7882;
wire n7883;
wire n7883_1;
wire n7884;
wire n7886;
wire n7887;
wire n7888;
wire n7889;
wire n7890;
wire n7891;
wire n7892;
wire n7893;
wire n7893_1;
wire n7895;
wire n7897;
wire n7897_1;
wire n7898;
wire n7900;
wire n7901;
wire n7902;
wire n7903;
wire n7904;
wire n7906;
wire n7906_1;
wire n7907;
wire n7908;
wire n7909;
wire n7910;
wire n7911;
wire n7911_1;
wire n7912;
wire n7913;
wire n7914;
wire n7915;
wire n7916;
wire n7916_1;
wire n7917;
wire n7918;
wire n7919;
wire n7920;
wire n7920_1;
wire n7921;
wire n7923;
wire n7924;
wire n7924_1;
wire n7925;
wire n7926;
wire n7927;
wire n7929;
wire n7929_1;
wire n793;
wire n7930;
wire n7931;
wire n7932;
wire n7933;
wire n7933_1;
wire n7934;
wire n7935;
wire n7936;
wire n7937;
wire n7937_1;
wire n7938;
wire n7939;
wire n7940;
wire n7941;
wire n7942;
wire n7942_1;
wire n7943;
wire n7944;
wire n7945;
wire n7945_1;
wire n7946;
wire n7947;
wire n7949;
wire n7950;
wire n7950_1;
wire n7951;
wire n7952;
wire n7953;
wire n7955;
wire n7955_1;
wire n7956;
wire n7958;
wire n7958_1;
wire n7959;
wire n7960;
wire n7961;
wire n7962;
wire n7962_1;
wire n7963;
wire n7964;
wire n7965;
wire n7966;
wire n7967;
wire n7967_1;
wire n7968;
wire n7969;
wire n7970;
wire n7970_1;
wire n7971;
wire n7972;
wire n7973;
wire n7974;
wire n7975;
wire n7975_1;
wire n7976;
wire n7978;
wire n798;
wire n7980;
wire n7980_1;
wire n7981;
wire n7983;
wire n7985;
wire n7986;
wire n7988;
wire n7989;
wire n7989_1;
wire n7991;
wire n7992;
wire n7993;
wire n7994;
wire n7994_1;
wire n7995;
wire n7997;
wire n7997_1;
wire n7998;
wire n7999;
wire n8000;
wire n8001;
wire n8002;
wire n8003;
wire n8004;
wire n8005;
wire n8005_1;
wire n8006;
wire n8007;
wire n8008;
wire n8009;
wire n8010;
wire n8010_1;
wire n8012;
wire n8014;
wire n8015;
wire n8016;
wire n8017;
wire n8019;
wire n8019_1;
wire n802;
wire n8020;
wire n8021;
wire n8022;
wire n8023;
wire n8024;
wire n8025;
wire n8026;
wire n8028;
wire n8028_1;
wire n8029;
wire n8030;
wire n8031;
wire n8032;
wire n8033;
wire n8033_1;
wire n8034;
wire n8035;
wire n8036;
wire n8037;
wire n8038;
wire n8038_1;
wire n8040;
wire n8041;
wire n8042;
wire n8042_1;
wire n8043;
wire n8044;
wire n8046;
wire n8047;
wire n8047_1;
wire n8048;
wire n8049;
wire n8050;
wire n8051;
wire n8051_1;
wire n8052;
wire n8053;
wire n8054;
wire n8055;
wire n8056;
wire n8056_1;
wire n8057;
wire n8058;
wire n8059;
wire n8059_1;
wire n806;
wire n8060;
wire n8061;
wire n8062;
wire n8063;
wire n8064;
wire n8064_1;
wire n8065;
wire n8066;
wire n8067;
wire n8067_1;
wire n8068;
wire n8069;
wire n8070;
wire n8071;
wire n8072;
wire n8072_1;
wire n8073;
wire n8074;
wire n8075;
wire n8075_1;
wire n8076;
wire n8077;
wire n8078;
wire n8079;
wire n8080;
wire n8080_1;
wire n8081;
wire n8082;
wire n8084;
wire n8085;
wire n8085_1;
wire n8086;
wire n8087;
wire n8088;
wire n8088_1;
wire n8089;
wire n8090;
wire n8092;
wire n8092_1;
wire n8093;
wire n8094;
wire n8096;
wire n8097;
wire n8097_1;
wire n8099;
wire n8100;
wire n8101;
wire n8102;
wire n8102_1;
wire n8103;
wire n8104;
wire n8105;
wire n8106;
wire n8107;
wire n8107_1;
wire n8108;
wire n8109;
wire n811;
wire n8110;
wire n8111;
wire n8112;
wire n8112_1;
wire n8113;
wire n8114;
wire n8115;
wire n8116;
wire n8116_1;
wire n8117;
wire n8119;
wire n8120;
wire n8121;
wire n8121_1;
wire n8122;
wire n8123;
wire n8124;
wire n8125;
wire n8125_1;
wire n8126;
wire n8127;
wire n8128;
wire n8129;
wire n8130;
wire n8130_1;
wire n8131;
wire n8132;
wire n8133;
wire n8135;
wire n8135_1;
wire n8136;
wire n8138;
wire n8139;
wire n8140;
wire n8140_1;
wire n8141;
wire n8142;
wire n8144;
wire n8144_1;
wire n8145;
wire n8146;
wire n8147;
wire n8147_1;
wire n8149;
wire n815;
wire n8150;
wire n8152;
wire n8152_1;
wire n8153;
wire n8155;
wire n8156;
wire n8156_1;
wire n8157;
wire n8158;
wire n8159;
wire n8160;
wire n8161;
wire n8161_1;
wire n8162;
wire n8163;
wire n8164;
wire n8165;
wire n8166;
wire n8166_1;
wire n8167;
wire n8168;
wire n8170;
wire n8170_1;
wire n8172;
wire n8173;
wire n8174;
wire n8175;
wire n8177;
wire n8178;
wire n8179;
wire n8179_1;
wire n8181;
wire n8182;
wire n8183;
wire n8183_1;
wire n8184;
wire n8185;
wire n8186;
wire n8187;
wire n8188;
wire n8188_1;
wire n8190;
wire n8191;
wire n8192;
wire n8192_1;
wire n8193;
wire n8194;
wire n8196;
wire n8197;
wire n8197_1;
wire n8198;
wire n8199;
wire n820;
wire n8200;
wire n8202;
wire n8202_1;
wire n8203;
wire n8205;
wire n8206;
wire n8206_1;
wire n8207;
wire n8208;
wire n8209;
wire n8211;
wire n8211_1;
wire n8212;
wire n8213;
wire n8214;
wire n8215;
wire n8216;
wire n8216_1;
wire n8217;
wire n8219;
wire n8220;
wire n8220_1;
wire n8221;
wire n8222;
wire n8223;
wire n8224;
wire n8224_1;
wire n8226;
wire n8227;
wire n8228;
wire n8229;
wire n8231;
wire n8232;
wire n8232_1;
wire n8233;
wire n8234;
wire n8235;
wire n8236;
wire n8237;
wire n8237_1;
wire n8238;
wire n8240;
wire n8241;
wire n8241_1;
wire n8243;
wire n8244;
wire n8245;
wire n8245_1;
wire n8246;
wire n8247;
wire n8249;
wire n8249_1;
wire n825;
wire n8250;
wire n8251;
wire n8252;
wire n8253;
wire n8253_1;
wire n8254;
wire n8255;
wire n8256;
wire n8258;
wire n8258_1;
wire n8259;
wire n8260;
wire n8261;
wire n8262;
wire n8262_1;
wire n8263;
wire n8264;
wire n8265;
wire n8266;
wire n8268;
wire n8269;
wire n8270;
wire n8271;
wire n8271_1;
wire n8272;
wire n8273;
wire n8274;
wire n8275;
wire n8276;
wire n8276_1;
wire n8277;
wire n8278;
wire n8279;
wire n8280;
wire n8280_1;
wire n8281;
wire n8282;
wire n8283;
wire n8284;
wire n8284_1;
wire n8285;
wire n8286;
wire n8287;
wire n8288;
wire n8289;
wire n8289_1;
wire n8290;
wire n8291;
wire n8292;
wire n8293;
wire n8294;
wire n8294_1;
wire n8295;
wire n8296;
wire n8297;
wire n8298;
wire n8299;
wire n8299_1;
wire n830;
wire n8300;
wire n8302;
wire n8303;
wire n8303_1;
wire n8304;
wire n8305;
wire n8306;
wire n8307;
wire n8307_1;
wire n8308;
wire n8309;
wire n8310;
wire n8311;
wire n8311_1;
wire n8312;
wire n8313;
wire n8315;
wire n8316;
wire n8316_1;
wire n8317;
wire n8319;
wire n8320;
wire n8320_1;
wire n8321;
wire n8322;
wire n8323;
wire n8324;
wire n8324_1;
wire n8325;
wire n8326;
wire n8328;
wire n8329;
wire n8330;
wire n8332;
wire n8333;
wire n8334;
wire n8334_1;
wire n8335;
wire n8336;
wire n8337;
wire n8337_1;
wire n8338;
wire n8339;
wire n834;
wire n8340;
wire n8340_1;
wire n8341;
wire n8342;
wire n8343;
wire n8344;
wire n8345;
wire n8345_1;
wire n8346;
wire n8348;
wire n8349;
wire n8350;
wire n8350_1;
wire n8351;
wire n8352;
wire n8353;
wire n8354;
wire n8354_1;
wire n8355;
wire n8356;
wire n8358;
wire n8359;
wire n8359_1;
wire n8360;
wire n8361;
wire n8362;
wire n8362_1;
wire n8365;
wire n8366;
wire n8367;
wire n8368;
wire n8369;
wire n8370;
wire n8371;
wire n8372;
wire n8372_1;
wire n8373;
wire n8374;
wire n8375;
wire n8377;
wire n8377_1;
wire n8378;
wire n8379;
wire n8380;
wire n8382;
wire n8382_1;
wire n8383;
wire n8385;
wire n8386;
wire n8387;
wire n8387_1;
wire n8388;
wire n839;
wire n8390;
wire n8391;
wire n8392;
wire n8392_1;
wire n8393;
wire n8394;
wire n8395;
wire n8396;
wire n8396_1;
wire n8397;
wire n8398;
wire n8399;
wire n8400;
wire n8401;
wire n8401_1;
wire n8402;
wire n8403;
wire n8404;
wire n8405;
wire n8405_1;
wire n8406;
wire n8407;
wire n8408;
wire n8409;
wire n8410;
wire n8410_1;
wire n8411;
wire n8412;
wire n8413;
wire n8414;
wire n8415;
wire n8415_1;
wire n8417;
wire n8418;
wire n8419;
wire n8421;
wire n8422;
wire n8423;
wire n8424;
wire n8425;
wire n8426;
wire n8426_1;
wire n8427;
wire n8429;
wire n8430;
wire n8430_1;
wire n8431;
wire n8432;
wire n8433;
wire n8434;
wire n8435;
wire n8435_1;
wire n8436;
wire n8437;
wire n8438;
wire n8438_1;
wire n8439;
wire n844;
wire n8440;
wire n8441;
wire n8442;
wire n8443;
wire n8443_1;
wire n8444;
wire n8445;
wire n8446;
wire n8447;
wire n8447_1;
wire n8448;
wire n8449;
wire n8450;
wire n8451;
wire n8451_1;
wire n8452;
wire n8453;
wire n8454;
wire n8455;
wire n8455_1;
wire n8456;
wire n8457;
wire n8458;
wire n8459;
wire n8459_1;
wire n8460;
wire n8461;
wire n8463;
wire n8464;
wire n8465;
wire n8466;
wire n8467;
wire n8467_1;
wire n8468;
wire n8469;
wire n8470;
wire n8471;
wire n8472;
wire n8472_1;
wire n8473;
wire n8474;
wire n8475;
wire n8476;
wire n8477;
wire n8477_1;
wire n8478;
wire n8479;
wire n8480;
wire n8481;
wire n8481_1;
wire n8482;
wire n8483;
wire n8484;
wire n8485;
wire n8486;
wire n8486_1;
wire n8487;
wire n8488;
wire n8489;
wire n849;
wire n8490;
wire n8491;
wire n8491_1;
wire n8492;
wire n8493;
wire n8494;
wire n8495;
wire n8497;
wire n8498;
wire n8499;
wire n8499_1;
wire n8500;
wire n8501;
wire n8502;
wire n8503;
wire n8504;
wire n8504_1;
wire n8505;
wire n8506;
wire n8507;
wire n8508;
wire n8508_1;
wire n8509;
wire n8511;
wire n8512;
wire n8513;
wire n8514;
wire n8516;
wire n8517;
wire n8517_1;
wire n8519;
wire n8520;
wire n8521;
wire n8522;
wire n8522_1;
wire n8523;
wire n8524;
wire n8525;
wire n8526;
wire n8526_1;
wire n8528;
wire n8529;
wire n8531;
wire n8531_1;
wire n8532;
wire n8534;
wire n8535;
wire n8535_1;
wire n8536;
wire n8537;
wire n8538;
wire n8539;
wire n854;
wire n8540;
wire n8540_1;
wire n8541;
wire n8542;
wire n8543;
wire n8544;
wire n8544_1;
wire n8545;
wire n8546;
wire n8547;
wire n8549;
wire n8549_1;
wire n8551;
wire n8552;
wire n8552_1;
wire n8553;
wire n8554;
wire n8555;
wire n8556;
wire n8557;
wire n8557_1;
wire n8558;
wire n8559;
wire n8560;
wire n8561;
wire n8561_1;
wire n8562;
wire n8563;
wire n8564;
wire n8565;
wire n8565_1;
wire n8566;
wire n8567;
wire n8568;
wire n8569;
wire n857;
wire n8570;
wire n8571;
wire n8572;
wire n8574;
wire n8575;
wire n8575_1;
wire n8577;
wire n8578;
wire n8578_1;
wire n8580;
wire n8581;
wire n8583;
wire n8583_1;
wire n8584;
wire n8585;
wire n8586;
wire n8587;
wire n8588;
wire n8588_1;
wire n8590;
wire n8591;
wire n8593;
wire n8593_1;
wire n8594;
wire n8596;
wire n8597;
wire n8598;
wire n8598_1;
wire n8599;
wire n8600;
wire n8601;
wire n8602;
wire n8602_1;
wire n8603;
wire n8604;
wire n8605;
wire n8606;
wire n8607;
wire n8607_1;
wire n8608;
wire n8609;
wire n8610;
wire n8611;
wire n8612;
wire n8612_1;
wire n8613;
wire n8614;
wire n8615;
wire n8616;
wire n8616_1;
wire n8617;
wire n8618;
wire n8619;
wire n862;
wire n8620;
wire n8621;
wire n8621_1;
wire n8622;
wire n8623;
wire n8624;
wire n8625;
wire n8625_1;
wire n8626;
wire n8627;
wire n8628;
wire n8628_1;
wire n8630;
wire n8631;
wire n8632;
wire n8632_1;
wire n8633;
wire n8634;
wire n8636;
wire n8637;
wire n8637_1;
wire n8638;
wire n8639;
wire n8640;
wire n8641;
wire n8642;
wire n8643;
wire n8645;
wire n8645_1;
wire n8646;
wire n8648;
wire n8650;
wire n8650_1;
wire n8653;
wire n8654;
wire n8654_1;
wire n8656;
wire n8657;
wire n8658;
wire n8659;
wire n8660;
wire n8661;
wire n8662;
wire n8662_1;
wire n8663;
wire n8664;
wire n8665;
wire n8666;
wire n8666_1;
wire n8667;
wire n8668;
wire n8669;
wire n867;
wire n8670;
wire n8671;
wire n8671_1;
wire n8672;
wire n8673;
wire n8674;
wire n8675;
wire n8676;
wire n8676_1;
wire n8677;
wire n8678;
wire n8679;
wire n8680;
wire n8681;
wire n8681_1;
wire n8682;
wire n8683;
wire n8684;
wire n8685;
wire n8685_1;
wire n8686;
wire n8687;
wire n8688;
wire n8689;
wire n8689_1;
wire n8690;
wire n8691;
wire n8693;
wire n8694;
wire n8694_1;
wire n8695;
wire n8696;
wire n8697;
wire n8698;
wire n8698_1;
wire n8699;
wire n870;
wire n8700;
wire n8701;
wire n8702;
wire n8703;
wire n8703_1;
wire n8704;
wire n8705;
wire n8706;
wire n8707;
wire n8708;
wire n8708_1;
wire n8710;
wire n8711;
wire n8711_1;
wire n8712;
wire n8713;
wire n8714;
wire n8715;
wire n8715_1;
wire n8716;
wire n8717;
wire n8719;
wire n8720;
wire n8720_1;
wire n8722;
wire n8723;
wire n8725;
wire n8725_1;
wire n8726;
wire n8728;
wire n8729;
wire n8730;
wire n8730_1;
wire n8731;
wire n8732;
wire n8734;
wire n8734_1;
wire n8735;
wire n8737;
wire n8738;
wire n8739;
wire n8739_1;
wire n8740;
wire n8741;
wire n8742;
wire n8743;
wire n8743_1;
wire n8744;
wire n8745;
wire n8746;
wire n8747;
wire n8748;
wire n8748_1;
wire n8749;
wire n875;
wire n8750;
wire n8751;
wire n8752;
wire n8753;
wire n8753_1;
wire n8754;
wire n8755;
wire n8757;
wire n8757_1;
wire n8759;
wire n8760;
wire n8761;
wire n8762;
wire n8762_1;
wire n8763;
wire n8764;
wire n8765;
wire n8766;
wire n8767;
wire n8767_1;
wire n8768;
wire n8770;
wire n8771;
wire n8771_1;
wire n8773;
wire n8774;
wire n8775;
wire n8776;
wire n8777;
wire n8778;
wire n8779;
wire n8780;
wire n8780_1;
wire n8781;
wire n8782;
wire n8783;
wire n8784;
wire n8784_1;
wire n8785;
wire n8786;
wire n8787;
wire n8788;
wire n8788_1;
wire n8789;
wire n8790;
wire n8791;
wire n8792;
wire n8793;
wire n8793_1;
wire n8794;
wire n8795;
wire n8796;
wire n8797;
wire n8797_1;
wire n8798;
wire n8799;
wire n880;
wire n8800;
wire n8800_1;
wire n8801;
wire n8803;
wire n8804;
wire n8805;
wire n8806;
wire n8807;
wire n8808;
wire n8809;
wire n8809_1;
wire n8810;
wire n8812;
wire n8813;
wire n8814;
wire n8815;
wire n8816;
wire n8817;
wire n8818;
wire n8818_1;
wire n8820;
wire n8821;
wire n8823;
wire n8823_1;
wire n8824;
wire n8826;
wire n8826_1;
wire n8828;
wire n8829;
wire n8830;
wire n8831;
wire n8831_1;
wire n8832;
wire n8833;
wire n8834;
wire n8835;
wire n8835_1;
wire n8837;
wire n8839;
wire n8840;
wire n8840_1;
wire n8841;
wire n8842;
wire n8843;
wire n8845;
wire n8845_1;
wire n8847;
wire n8848;
wire n8849;
wire n885;
wire n8850;
wire n8850_1;
wire n8851;
wire n8852;
wire n8853;
wire n8855;
wire n8855_1;
wire n8856;
wire n8857;
wire n8858;
wire n8859;
wire n8860;
wire n8860_1;
wire n8861;
wire n8862;
wire n8863;
wire n8864;
wire n8866;
wire n8867;
wire n8868;
wire n8869;
wire n8869_1;
wire n8870;
wire n8872;
wire n8873;
wire n8873_1;
wire n8875;
wire n8876;
wire n8877;
wire n8877_1;
wire n8878;
wire n8880;
wire n8881;
wire n8882;
wire n8882_1;
wire n8883;
wire n8884;
wire n8885;
wire n8886;
wire n8886_1;
wire n8887;
wire n8888;
wire n8889;
wire n8890;
wire n8891;
wire n8891_1;
wire n8892;
wire n8893;
wire n8894;
wire n8895;
wire n8895_1;
wire n8896;
wire n8899;
wire n8899_1;
wire n890;
wire n8901;
wire n8902;
wire n8903;
wire n8904;
wire n8905;
wire n8907;
wire n8908;
wire n8908_1;
wire n8910;
wire n8911;
wire n8912;
wire n8913;
wire n8914;
wire n8915;
wire n8916;
wire n8917;
wire n8917_1;
wire n8918;
wire n8919;
wire n8921;
wire n8922;
wire n8922_1;
wire n8923;
wire n8924;
wire n8925;
wire n8926;
wire n8927;
wire n8928;
wire n8930;
wire n8931;
wire n8931_1;
wire n8933;
wire n8934;
wire n8934_1;
wire n8935;
wire n8936;
wire n8937;
wire n8939;
wire n8939_1;
wire n894;
wire n8941;
wire n8942;
wire n8943;
wire n8944;
wire n8945;
wire n8947;
wire n8948;
wire n8948_1;
wire n8950;
wire n8951;
wire n8953;
wire n8954;
wire n8955;
wire n8957;
wire n8958;
wire n8958_1;
wire n8959;
wire n8960;
wire n8961;
wire n8963;
wire n8963_1;
wire n8964;
wire n8966;
wire n8967;
wire n8968;
wire n8969;
wire n8971;
wire n8971_1;
wire n8972;
wire n8974;
wire n8975;
wire n8976;
wire n8976_1;
wire n8977;
wire n8978;
wire n8979;
wire n8980;
wire n8981;
wire n8981_1;
wire n8982;
wire n8983;
wire n8984;
wire n8985;
wire n8986;
wire n8986_1;
wire n8987;
wire n8988;
wire n8989;
wire n899;
wire n8990;
wire n8991;
wire n8992;
wire n8993;
wire n8994;
wire n8995;
wire n8995_1;
wire n8997;
wire n8999;
wire n9000;
wire n9000_1;
wire n9001;
wire n9002;
wire n9003;
wire n9004;
wire n9005;
wire n9005_1;
wire n9006;
wire n9007;
wire n9008;
wire n9009;
wire n9010;
wire n9010_1;
wire n9011;
wire n9012;
wire n9013;
wire n9014;
wire n9014_1;
wire n9015;
wire n9016;
wire n9017;
wire n9017_1;
wire n9019;
wire n9020;
wire n9022;
wire n9022_1;
wire n9023;
wire n9025;
wire n9025_1;
wire n9026;
wire n9027;
wire n9028;
wire n9029;
wire n903;
wire n9030;
wire n9030_1;
wire n9031;
wire n9032;
wire n9033;
wire n9034;
wire n9034_1;
wire n9035;
wire n9036;
wire n9037;
wire n9038;
wire n9040;
wire n9041;
wire n9042;
wire n9042_1;
wire n9043;
wire n9044;
wire n9045;
wire n9046;
wire n9047;
wire n9047_1;
wire n9048;
wire n9049;
wire n9050;
wire n9051;
wire n9052;
wire n9052_1;
wire n9053;
wire n9054;
wire n9055;
wire n9056;
wire n9057;
wire n9057_1;
wire n9058;
wire n9059;
wire n9060;
wire n9060_1;
wire n9061;
wire n9063;
wire n9064;
wire n9065;
wire n9066;
wire n9067;
wire n9068;
wire n9069;
wire n9069_1;
wire n907;
wire n9070;
wire n9071;
wire n9072;
wire n9073;
wire n9074;
wire n9074_1;
wire n9075;
wire n9077;
wire n9078;
wire n9079;
wire n9079_1;
wire n9080;
wire n9081;
wire n9082;
wire n9082_1;
wire n9083;
wire n9084;
wire n9086;
wire n9086_1;
wire n9087;
wire n9089;
wire n9090;
wire n9091;
wire n9091_1;
wire n9092;
wire n9093;
wire n9094;
wire n9095;
wire n9096;
wire n9096_1;
wire n9098;
wire n9100;
wire n9101;
wire n9102;
wire n9103;
wire n9104;
wire n9105;
wire n9106;
wire n9106_1;
wire n9107;
wire n9108;
wire n9109;
wire n911;
wire n9110;
wire n9110_1;
wire n9111;
wire n9112;
wire n9113;
wire n9114;
wire n9115;
wire n9115_1;
wire n9116;
wire n9117;
wire n9118;
wire n9119;
wire n9120;
wire n9121;
wire n9122;
wire n9123;
wire n9124;
wire n9124_1;
wire n9125;
wire n9126;
wire n9127;
wire n9128;
wire n9129;
wire n9129_1;
wire n9130;
wire n9131;
wire n9132;
wire n9133;
wire n9134;
wire n9134_1;
wire n9135;
wire n9136;
wire n9137;
wire n9138;
wire n9138_1;
wire n9139;
wire n9140;
wire n9141;
wire n9142;
wire n9143;
wire n9143_1;
wire n9144;
wire n9145;
wire n9146;
wire n9146_1;
wire n9147;
wire n9148;
wire n9149;
wire n9151;
wire n9151_1;
wire n9152;
wire n9153;
wire n9154;
wire n9155;
wire n9156;
wire n9157;
wire n9158;
wire n916;
wire n9160;
wire n9160_1;
wire n9161;
wire n9163;
wire n9164;
wire n9164_1;
wire n9166;
wire n9167;
wire n9168;
wire n9169;
wire n9169_1;
wire n9170;
wire n9171;
wire n9172;
wire n9173;
wire n9173_1;
wire n9175;
wire n9176;
wire n9177;
wire n9178;
wire n9178_1;
wire n9179;
wire n9180;
wire n9181;
wire n9182;
wire n9182_1;
wire n9183;
wire n9184;
wire n9185;
wire n9186;
wire n9187;
wire n9187_1;
wire n9188;
wire n9189;
wire n9190;
wire n9191;
wire n9192;
wire n9192_1;
wire n9193;
wire n9195;
wire n9196;
wire n9196_1;
wire n9197;
wire n9199;
wire n920;
wire n9200;
wire n9201;
wire n9201_1;
wire n9202;
wire n9203;
wire n9204;
wire n9205;
wire n9206;
wire n9206_1;
wire n9207;
wire n9208;
wire n9209;
wire n9210;
wire n9211;
wire n9211_1;
wire n9212;
wire n9214;
wire n9215;
wire n9216;
wire n9217;
wire n9219;
wire n9220;
wire n9220_1;
wire n9221;
wire n9222;
wire n9223;
wire n9224;
wire n9225;
wire n9225_1;
wire n9226;
wire n9227;
wire n9228;
wire n9228_1;
wire n9229;
wire n9230;
wire n9231;
wire n9232;
wire n9233;
wire n9233_1;
wire n9234;
wire n9235;
wire n9236;
wire n9237;
wire n9238;
wire n9238_1;
wire n9239;
wire n9240;
wire n9241;
wire n9242;
wire n9242_1;
wire n9243;
wire n9244;
wire n9245;
wire n9246;
wire n9247;
wire n9248;
wire n9249;
wire n925;
wire n9250;
wire n9250_1;
wire n9251;
wire n9253;
wire n9254;
wire n9255;
wire n9256;
wire n9258;
wire n9258_1;
wire n9259;
wire n9260;
wire n9261;
wire n9262;
wire n9263;
wire n9264;
wire n9265;
wire n9267;
wire n9267_1;
wire n9268;
wire n9269;
wire n9270;
wire n9271;
wire n9272;
wire n9272_1;
wire n9273;
wire n9274;
wire n9275;
wire n9276;
wire n9277;
wire n9277_1;
wire n9279;
wire n9282;
wire n9282_1;
wire n9283;
wire n9284;
wire n9285;
wire n9286;
wire n9287;
wire n9287_1;
wire n9288;
wire n9289;
wire n9290;
wire n9290_1;
wire n9291;
wire n9292;
wire n9293;
wire n9294;
wire n9294_1;
wire n9295;
wire n9296;
wire n9297;
wire n9298;
wire n9298_1;
wire n9299;
wire n930;
wire n9300;
wire n9301;
wire n9302;
wire n9303;
wire n9305;
wire n9306;
wire n9307;
wire n9307_1;
wire n9308;
wire n9309;
wire n9310;
wire n9311;
wire n9312;
wire n9312_1;
wire n9313;
wire n9315;
wire n9316;
wire n9316_1;
wire n9317;
wire n9318;
wire n9319;
wire n9321;
wire n9321_1;
wire n9322;
wire n9323;
wire n9324;
wire n9326;
wire n9326_1;
wire n9327;
wire n9329;
wire n9330;
wire n9330_1;
wire n9332;
wire n9333;
wire n9334;
wire n9335;
wire n9335_1;
wire n9336;
wire n9337;
wire n9338;
wire n9339;
wire n9339_1;
wire n9340;
wire n9341;
wire n9342;
wire n9343;
wire n9343_1;
wire n9344;
wire n9345;
wire n9346;
wire n9347;
wire n9348;
wire n9348_1;
wire n935;
wire n9350;
wire n9351;
wire n9352;
wire n9353;
wire n9354;
wire n9355;
wire n9356;
wire n9357;
wire n9358;
wire n9359;
wire n9360;
wire n9361;
wire n9361_1;
wire n9362;
wire n9363;
wire n9364;
wire n9365;
wire n9365_1;
wire n9367;
wire n9368;
wire n9370;
wire n9370_1;
wire n9371;
wire n9372;
wire n9373;
wire n9373_1;
wire n9374;
wire n9376;
wire n9377;
wire n9377_1;
wire n9379;
wire n9380;
wire n9381;
wire n9382;
wire n9383;
wire n9384;
wire n9385;
wire n9385_1;
wire n9386;
wire n9387;
wire n9389;
wire n9390;
wire n9391;
wire n9392;
wire n9393;
wire n9394;
wire n9395;
wire n9396;
wire n9397;
wire n9398;
wire n9398_1;
wire n9399;
wire n940;
wire n9401;
wire n9402;
wire n9402_1;
wire n9403;
wire n9404;
wire n9405;
wire n9405_1;
wire n9406;
wire n9407;
wire n9409;
wire n9410;
wire n9410_1;
wire n9411;
wire n9412;
wire n9413;
wire n9414;
wire n9415;
wire n9416;
wire n9417;
wire n9419;
wire n9420;
wire n9420_1;
wire n9421;
wire n9422;
wire n9423;
wire n9424;
wire n9425;
wire n9425_1;
wire n9426;
wire n9427;
wire n9428;
wire n9428_1;
wire n9429;
wire n9430;
wire n9431;
wire n9432;
wire n9433;
wire n9435;
wire n9436;
wire n9436_1;
wire n9437;
wire n9438;
wire n9439;
wire n944;
wire n9440;
wire n9441;
wire n9441_1;
wire n9442;
wire n9443;
wire n9444;
wire n9445;
wire n9446;
wire n9447;
wire n9449;
wire n9449_1;
wire n9450;
wire n9452;
wire n9453;
wire n9454;
wire n9455;
wire n9456;
wire n9458;
wire n9459;
wire n9459_1;
wire n9461;
wire n9462;
wire n9462_1;
wire n9463;
wire n9464;
wire n9465;
wire n9466;
wire n9467;
wire n9467_1;
wire n9468;
wire n9469;
wire n9470;
wire n9470_1;
wire n9471;
wire n9472;
wire n9473;
wire n9474;
wire n9475;
wire n9475_1;
wire n9476;
wire n9477;
wire n9478;
wire n9478_1;
wire n9479;
wire n948;
wire n9481;
wire n9482;
wire n9483;
wire n9484;
wire n9485;
wire n9486;
wire n9487;
wire n9487_1;
wire n9488;
wire n9490;
wire n9491;
wire n9492;
wire n9492_1;
wire n9493;
wire n9494;
wire n9496;
wire n9497;
wire n9497_1;
wire n9499;
wire n9501;
wire n9502;
wire n9502_1;
wire n9503;
wire n9504;
wire n9505;
wire n9506;
wire n9507;
wire n9507_1;
wire n9508;
wire n9509;
wire n9510;
wire n9511;
wire n9512;
wire n9512_1;
wire n9513;
wire n9515;
wire n9516;
wire n9517;
wire n9517_1;
wire n9518;
wire n9519;
wire n9520;
wire n9520_1;
wire n9521;
wire n9522;
wire n9523;
wire n9525;
wire n9525_1;
wire n9526;
wire n9528;
wire n9528_1;
wire n9529;
wire n953;
wire n9531;
wire n9532;
wire n9533;
wire n9534;
wire n9535;
wire n9536;
wire n9537;
wire n9537_1;
wire n9538;
wire n9540;
wire n9541;
wire n9541_1;
wire n9543;
wire n9544;
wire n9545;
wire n9546;
wire n9546_1;
wire n9547;
wire n9549;
wire n9549_1;
wire n9550;
wire n9552;
wire n9553;
wire n9554;
wire n9555;
wire n9556;
wire n9558;
wire n9559;
wire n9559_1;
wire n956;
wire n9561;
wire n9562;
wire n9563;
wire n9564;
wire n9564_1;
wire n9565;
wire n9566;
wire n9568;
wire n9569;
wire n9569_1;
wire n9570;
wire n9571;
wire n9572;
wire n9574;
wire n9574_1;
wire n9575;
wire n9577;
wire n9578;
wire n9579;
wire n9581;
wire n9582;
wire n9583;
wire n9584;
wire n9585;
wire n9586;
wire n9587;
wire n9588;
wire n9588_1;
wire n9590;
wire n9591;
wire n9592;
wire n9592_1;
wire n9594;
wire n9595;
wire n9597;
wire n9597_1;
wire n9598;
wire n9600;
wire n9601;
wire n9602;
wire n9602_1;
wire n9603;
wire n9604;
wire n9605;
wire n9606;
wire n9606_1;
wire n9607;
wire n9608;
wire n9609;
wire n961;
wire n9610;
wire n9611;
wire n9611_1;
wire n9612;
wire n9613;
wire n9614;
wire n9615;
wire n9616;
wire n9616_1;
wire n9617;
wire n9618;
wire n9619;
wire n9620;
wire n9620_1;
wire n9622;
wire n9623;
wire n9624;
wire n9625;
wire n9626;
wire n9627;
wire n9628;
wire n9628_1;
wire n9629;
wire n9630;
wire n9631;
wire n9632;
wire n9633;
wire n9633_1;
wire n9634;
wire n9635;
wire n9636;
wire n9637;
wire n9638;
wire n9639;
wire n9640;
wire n9641;
wire n9642;
wire n9643;
wire n9644;
wire n9645;
wire n9646;
wire n9647;
wire n9647_1;
wire n9648;
wire n9649;
wire n9651;
wire n9651_1;
wire n9652;
wire n9654;
wire n9655;
wire n9655_1;
wire n9656;
wire n9657;
wire n9658;
wire n9659;
wire n966;
wire n9660;
wire n9660_1;
wire n9663;
wire n9664;
wire n9664_1;
wire n9665;
wire n9666;
wire n9667;
wire n9668;
wire n9668_1;
wire n9670;
wire n9671;
wire n9672;
wire n9673;
wire n9674;
wire n9675;
wire n9677;
wire n9678;
wire n9678_1;
wire n9680;
wire n9681;
wire n9683;
wire n9683_1;
wire n9684;
wire n9685;
wire n9686;
wire n9687;
wire n9688;
wire n9689;
wire n9691;
wire n9692;
wire n9692_1;
wire n9694;
wire n9695;
wire n9695_1;
wire n9697;
wire n9698;
wire n9699;
wire n9700;
wire n9700_1;
wire n9701;
wire n9703;
wire n9704;
wire n9705;
wire n9706;
wire n9707;
wire n9708;
wire n9709;
wire n9709_1;
wire n971;
wire n9710;
wire n9712;
wire n9713;
wire n9714;
wire n9715;
wire n9716;
wire n9717;
wire n9718;
wire n9719;
wire n9719_1;
wire n9720;
wire n9721;
wire n9723;
wire n9724;
wire n9724_1;
wire n9727;
wire n9728;
wire n9729;
wire n9730;
wire n9731;
wire n9732;
wire n9733;
wire n9733_1;
wire n9734;
wire n9735;
wire n9736;
wire n9737;
wire n9737_1;
wire n9738;
wire n9739;
wire n9740;
wire n9741;
wire n9742;
wire n9743;
wire n9744;
wire n9746;
wire n9746_1;
wire n9748;
wire n9750;
wire n9750_1;
wire n9751;
wire n9752;
wire n9753;
wire n9754;
wire n9754_1;
wire n9755;
wire n9756;
wire n9757;
wire n9758;
wire n9758_1;
wire n9759;
wire n976;
wire n9760;
wire n9761;
wire n9762;
wire n9763;
wire n9763_1;
wire n9764;
wire n9765;
wire n9766;
wire n9767;
wire n9768;
wire n9768_1;
wire n9769;
wire n9770;
wire n9771;
wire n9772;
wire n9773;
wire n9773_1;
wire n9774;
wire n9775;
wire n9777;
wire n9778;
wire n9778_1;
wire n9780;
wire n9781;
wire n9783;
wire n9783_1;
wire n9784;
wire n9785;
wire n9786;
wire n9787;
wire n9787_1;
wire n9789;
wire n9791;
wire n9792;
wire n9792_1;
wire n9793;
wire n9795;
wire n9796;
wire n9796_1;
wire n9798;
wire n9799;
wire n9801;
wire n9801_1;
wire n9802;
wire n9804;
wire n9805;
wire n9805_1;
wire n9807;
wire n9808;
wire n9809;
wire n9809_1;
wire n981;
wire n9810;
wire n9811;
wire n9813;
wire n9814;
wire n9814_1;
wire n9816;
wire n9817;
wire n9819;
wire n9819_1;
wire n9821;
wire n9822;
wire n9823;
wire n9824;
wire n9824_1;
wire n9825;
wire n9826;
wire n9827;
wire n9828;
wire n9828_1;
wire n9831;
wire n9832;
wire n9833;
wire n9833_1;
wire n9834;
wire n9835;
wire n9836;
wire n9837;
wire n9837_1;
wire n9838;
wire n9839;
wire n9840;
wire n9840_1;
wire n9841;
wire n9842;
wire n9843;
wire n9844;
wire n9844_1;
wire n9846;
wire n9847;
wire n9849;
wire n9849_1;
wire n985;
wire n9850;
wire n9852;
wire n9853;
wire n9853_1;
wire n9854;
wire n9855;
wire n9856;
wire n9857;
wire n9858;
wire n9858_1;
wire n9859;
wire n9860;
wire n9861;
wire n9863;
wire n9863_1;
wire n9864;
wire n9866;
wire n9867;
wire n9867_1;
wire n9869;
wire n9870;
wire n9871;
wire n9871_1;
wire n9872;
wire n9873;
wire n9875;
wire n9875_1;
wire n9876;
wire n9878;
wire n9879;
wire n9880;
wire n9880_1;
wire n9881;
wire n9882;
wire n9884;
wire n9885;
wire n9885_1;
wire n9886;
wire n9887;
wire n9889;
wire n9889_1;
wire n9890;
wire n9892;
wire n9893;
wire n9894;
wire n9895;
wire n9896;
wire n9898;
wire n9899;
wire n990;
wire n9900;
wire n9901;
wire n9902;
wire n9904;
wire n9906;
wire n9907;
wire n9907_1;
wire n9908;
wire n9909;
wire n9910;
wire n9911;
wire n9911_1;
wire n9913;
wire n9914;
wire n9914_1;
wire n9915;
wire n9916;
wire n9918;
wire n9918_1;
wire n9919;
wire n9921;
wire n9922;
wire n9923;
wire n9924;
wire n9925;
wire n9926;
wire n9927;
wire n9928;
wire n9929;
wire n9930;
wire n9930_1;
wire n9931;
wire n9932;
wire n9933;
wire n9934;
wire n9935;
wire n9935_1;
wire n9936;
wire n9937;
wire n9938;
wire n9939;
wire n9939_1;
wire n9940;
wire n9941;
wire n9942;
wire n9943;
wire n9944;
wire n9944_1;
wire n9945;
wire n9947;
wire n9948;
wire n9949;
wire n995;
wire n9950;
wire n9951;
wire n9952;
wire n9953;
wire n9953_1;
wire n9954;
wire n9955;
wire n9956;
wire n9957;
wire n9957_1;
wire n9958;
wire n9959;
wire n9960;
wire n9961;
wire n9961_1;
wire n9962;
wire n9963;
wire n9964;
wire n9965;
wire n9966;
wire n9966_1;
wire n9967;
wire n9968;
wire n9970;
wire n9971;
wire n9971_1;
wire n9973;
wire n9974;
wire n9975;
wire n9976;
wire n9976_1;
wire n9977;
wire n9978;
wire n9980;
wire n9981;
wire n9982;
wire n9983;
wire n9985;
wire n9985_1;
wire n9986;
wire n9988;
wire n9988_1;
wire n9989;
wire n9991;
wire n9992;
wire n9992_1;
wire n9994;
wire n9995;
wire n9997;
wire n9997_1;
wire n9998;
wire net_130;
wire net_131;
wire net_132;
wire net_133;
wire net_134;
wire net_135;
wire net_136;
wire net_137;
wire net_138;
wire net_139;
wire net_140;
wire net_141;
wire net_142;
wire net_143;
wire net_144;
wire net_145;
wire net_146;
wire net_147;
wire net_148;
wire net_149;
wire net_150;
wire net_151;
wire net_152;
wire net_153;
wire net_155;
wire net_156;
wire net_157;
wire net_158;
wire net_159;
wire net_160;
wire net_161;
wire net_162;
wire net_163;
wire net_164;
wire net_165;
wire net_166;
wire net_167;
wire net_168;
wire net_169;
wire net_170;
wire net_171;
wire net_179;
wire net_181;
wire net_182;
wire net_183;
wire net_185;
wire net_186;
wire net_187;
wire net_194;
wire net_195;
wire net_196;
wire net_197;
wire net_198;
wire net_199;
wire net_200;
wire net_202;
wire net_203;
wire net_204;
wire net_205;
wire net_206;
wire net_207;
wire net_208;
wire net_216;
wire net_218;
wire net_219;
wire net_220;
wire net_222;
wire net_223;
wire net_224;
wire net_230;
wire net_231;
wire net_232;
wire net_233;
wire net_234;
wire net_235;
wire net_236;
wire net_237;
wire net_238;
wire net_239;
wire net_240;
wire net_241;
wire net_242;
wire net_243;
wire net_244;
wire net_245;
wire net_246;
wire net_247;
wire net_248;
wire net_249;
wire net_250;
wire net_251;
wire net_252;
wire net_253;
wire net_254;
wire net_255;
wire net_256;
wire net_257;
wire net_258;
wire net_259;
wire net_260;
wire net_261;
wire net_274;
wire net_285;
wire net_296;
wire net_297;
wire net_303;
wire net_304;
wire net_305;
wire net_306;
wire net_307;
wire net_308;
wire net_309;
wire net_310;
wire net_311;
wire net_312;
wire net_313;
wire net_314;
wire net_315;
wire net_316;
wire net_317;
wire net_318;
wire net_319;
wire net_320;
wire net_321;
wire net_322;
wire net_323;
wire net_324;
wire net_325;
wire net_326;
wire net_327;
wire net_328;
wire net_329;
wire net_330;
wire net_331;
wire net_332;
wire net_333;
wire net_334;
wire net_335;
wire net_336;
wire net_337;
wire net_338;
wire net_339;
wire net_340;
wire net_341;
wire net_342;
wire net_343;
wire net_344;
wire net_345;
wire net_346;
wire net_347;
wire net_348;
wire net_349;
wire net_350;
wire net_351;
wire net_352;
wire net_353;
wire net_354;
wire net_355;
wire net_356;
wire net_357;
wire net_358;
wire net_359;
wire net_360;
wire net_361;
wire net_362;
wire net_363;
wire net_364;
wire net_365;
wire net_366;
wire net_367;
wire net_368;
wire net_369;
wire net_370;
wire net_371;
wire net_372;
wire net_373;
wire net_374;
wire net_375;
wire net_376;
wire net_377;
wire net_378;
wire net_379;
wire net_380;
wire net_381;
wire net_382;
wire net_383;
wire net_384;
wire net_385;
wire net_386;
wire net_387;
wire net_388;
wire net_389;
wire net_390;
wire net_391;
wire net_5858;
wire net_5860;
wire net_5861;
wire net_5992;
wire net_6003;
wire net_6013;
wire net_6014;
wire net_6024;
wire net_6025;
wire net_6035;
wire net_6036;
wire net_6046;
wire net_6056;
wire net_6057;
wire net_6058;
wire net_6059;
wire net_6060;
wire net_6061;
wire net_6380;
wire net_6381;
wire net_6382;
wire net_6383;
wire net_6384;
wire net_6385;
wire net_6386;
wire net_6387;
wire net_6388;
wire net_6389;
wire net_6390;
wire net_6391;
wire net_6392;
wire net_6393;
wire net_6394;
wire net_6395;
wire net_6396;
wire net_6397;
wire net_6398;
wire net_6399;
wire net_6400;
wire net_6403;
wire net_6412;
wire net_6416;
wire net_6417;
wire net_6424;
wire net_6425;
wire net_6426;
wire net_6427;
wire net_6428;
wire net_6429;
wire net_6430;
wire net_6431;
wire net_6432;
wire net_6433;
wire net_6434;
wire net_6435;
wire net_6436;
wire net_6437;
wire net_6438;
wire net_6439;
wire net_6440;
wire net_6441;
wire net_6442;
wire net_6443;
wire net_6444;
wire net_6445;
wire net_6446;
wire net_6447;
wire net_6448;
wire net_6449;
wire net_6450;
wire net_6451;
wire net_6452;
wire net_6453;
wire net_6454;
wire net_6455;
wire net_6456;
wire net_6457;
wire net_6458;
wire net_6459;
wire net_6460;
wire net_6461;
wire net_6462;
wire net_6463;
wire net_6464;
wire net_6465;
wire net_6466;
wire net_6467;
wire net_6468;
wire net_6469;
wire net_6470;
wire net_6471;
wire net_6472;
wire net_6473;
wire net_6474;
wire net_6475;
wire net_6476;
wire net_6477;
wire net_6478;
wire net_6479;
wire net_6480;
wire net_6481;
wire net_6482;
wire net_6483;
wire net_6484;
wire net_6485;
wire net_6486;
wire net_6487;
wire net_6488;
wire net_6489;
wire net_6490;
wire net_6491;
wire net_6492;
wire net_6493;
wire net_6494;
wire net_6495;
wire net_6496;
wire net_6497;
wire net_6498;
wire net_6499;
wire net_6500;
wire net_6501;
wire net_6502;
wire net_6503;
wire net_6504;
wire net_6505;
wire net_6506;
wire net_6507;
wire net_6508;
wire net_6509;
wire net_6510;
wire net_6511;
wire net_6512;
wire net_6513;
wire net_6514;
wire net_6515;
wire net_6516;
wire net_6517;
wire net_6518;
wire net_6519;
wire net_6520;
wire net_6521;
wire net_6522;
wire net_6523;
wire net_6524;
wire net_6525;
wire net_6526;
wire net_6527;
wire net_6528;
wire net_6529;
wire net_6530;
wire net_6531;
wire net_6532;
wire net_6533;
wire net_6534;
wire net_6535;
wire net_6536;
wire net_6537;
wire net_6538;
wire net_6539;
wire net_6540;
wire net_6541;
wire net_6542;
wire net_6543;
wire net_6544;
wire net_6545;
wire net_6546;
wire net_6547;
wire net_6548;
wire net_6549;
wire net_6550;
wire net_6551;
wire net_6556;
wire net_6559;
wire net_6560;
wire net_6561;
wire net_6562;
wire net_6563;
wire net_6564;
wire net_6565;
wire net_6566;
wire net_6567;
wire net_6568;
wire net_6569;
wire net_6570;
wire net_6571;
wire net_6572;
wire net_6573;
wire net_6574;
wire net_6575;
wire net_6576;
wire net_6577;
wire net_6578;
wire net_6579;
wire net_6580;
wire net_6581;
wire net_6582;
wire net_6583;
wire net_6584;
wire net_6585;
wire net_6586;
wire net_6587;
wire net_6588;
wire net_6589;
wire net_6590;
wire net_6591;
wire net_6592;
wire net_6593;
wire net_6594;
wire net_6595;
wire net_6596;
wire net_6597;
wire net_6598;
wire net_6599;
wire net_6600;
wire net_6601;
wire net_6602;
wire net_6603;
wire net_6604;
wire net_6605;
wire net_6606;
wire net_6607;
wire net_6608;
wire net_6609;
wire net_6610;
wire net_6611;
wire net_6612;
wire net_6613;
wire net_6614;
wire net_6615;
wire net_6616;
wire net_6617;
wire net_6618;
wire net_6619;
wire net_6620;
wire net_6621;
wire net_6622;
wire net_6623;
wire net_6624;
wire net_6625;
wire net_6626;
wire net_6627;
wire net_6628;
wire net_6629;
wire net_6630;
wire net_6631;
wire net_6632;
wire net_6633;
wire net_6634;
wire net_6635;
wire net_6636;
wire net_6637;
wire net_6638;
wire net_6639;
wire net_6640;
wire net_6641;
wire net_6642;
wire net_6643;
wire net_6644;
wire net_6645;
wire net_6646;
wire net_6647;
wire net_6648;
wire net_6649;
wire net_6650;
wire net_6651;
wire net_6652;
wire net_6653;
wire net_6654;
wire net_6655;
wire net_6656;
wire net_6657;
wire net_6658;
wire net_6659;
wire net_6660;
wire net_6661;
wire net_6662;
wire net_6663;
wire net_6664;
wire net_6665;
wire net_6666;
wire net_6667;
wire net_6668;
wire net_6669;
wire net_6670;
wire net_6671;
wire net_6672;
wire net_6673;
wire net_6674;
wire net_6675;
wire net_6676;
wire net_6677;
wire net_6678;
wire net_6679;
wire net_6680;
wire net_6681;
wire net_6682;
wire net_6683;
wire net_6684;
wire net_6685;
wire net_6686;
wire net_6691;
wire net_6694;
wire net_6695;
wire net_6696;
wire net_6697;
wire net_6698;
wire net_6699;
wire net_6700;
wire net_6701;
wire net_6702;
wire net_6703;
wire net_6704;
wire net_6705;
wire net_6706;
wire net_6707;
wire net_6708;
wire net_6709;
wire net_6710;
wire net_6711;
wire net_6712;
wire net_6713;
wire net_6714;
wire net_6715;
wire net_6716;
wire net_6717;
wire net_6718;
wire net_6719;
wire net_6720;
wire net_6721;
wire net_6722;
wire net_6723;
wire net_6724;
wire net_6725;
wire net_6726;
wire net_6727;
wire net_6728;
wire net_6729;
wire net_6730;
wire net_6731;
wire net_6732;
wire net_6733;
wire net_6734;
wire net_6735;
wire net_6736;
wire net_6737;
wire net_6738;
wire net_6739;
wire net_6740;
wire net_6741;
wire net_6742;
wire net_6743;
wire net_6744;
wire net_6745;
wire net_6746;
wire net_6747;
wire net_6748;
wire net_6749;
wire net_6750;
wire net_6751;
wire net_6752;
wire net_6753;
wire net_6754;
wire net_6755;
wire net_6756;
wire net_6757;
wire net_6758;
wire net_6759;
wire net_6760;
wire net_6761;
wire net_6762;
wire net_6763;
wire net_6764;
wire net_6765;
wire net_6766;
wire net_6767;
wire net_6768;
wire net_6769;
wire net_6770;
wire net_6771;
wire net_6772;
wire net_6773;
wire net_6774;
wire net_6775;
wire net_6776;
wire net_6777;
wire net_6778;
wire net_6779;
wire net_6780;
wire net_6781;
wire net_6782;
wire net_6783;
wire net_6784;
wire net_6785;
wire net_6786;
wire net_6787;
wire net_6788;
wire net_6789;
wire net_6790;
wire net_6791;
wire net_6792;
wire net_6793;
wire net_6794;
wire net_6795;
wire net_6796;
wire net_6797;
wire net_6798;
wire net_6799;
wire net_6800;
wire net_6801;
wire net_6802;
wire net_6803;
wire net_6804;
wire net_6805;
wire net_6806;
wire net_6807;
wire net_6808;
wire net_6809;
wire net_6810;
wire net_6811;
wire net_6812;
wire net_6813;
wire net_6814;
wire net_6815;
wire net_6816;
wire net_6817;
wire net_6818;
wire net_6819;
wire net_6820;
wire net_6821;
wire net_6826;
wire net_6829;
wire net_6830;
wire net_6831;
wire net_6832;
wire net_6833;
wire net_6834;
wire net_6835;
wire net_6836;
wire net_6837;
wire net_6838;
wire net_6839;
wire net_6840;
wire net_6841;
wire net_6842;
wire net_6843;
wire net_6844;
wire net_6845;
wire net_6846;
wire net_6847;
wire net_6848;
wire net_6849;
wire net_6850;
wire net_6851;
wire net_6852;
wire net_6853;
wire net_6854;
wire net_6855;
wire net_6856;
wire net_6857;
wire net_6858;
wire net_6859;
wire net_6860;
wire net_6861;
wire net_6862;
wire net_6863;
wire net_6864;
wire net_6865;
wire net_6866;
wire net_6867;
wire net_6868;
wire net_6869;
wire net_6870;
wire net_6871;
wire net_6872;
wire net_6873;
wire net_6874;
wire net_6875;
wire net_6876;
wire net_6877;
wire net_6878;
wire net_6879;
wire net_6880;
wire net_6881;
wire net_6882;
wire net_6883;
wire net_6884;
wire net_6885;
wire net_6886;
wire net_6887;
wire net_6888;
wire net_6889;
wire net_6890;
wire net_6891;
wire net_6892;
wire net_6893;
wire net_6894;
wire net_6895;
wire net_6896;
wire net_6897;
wire net_6898;
wire net_6899;
wire net_6900;
wire net_6901;
wire net_6902;
wire net_6903;
wire net_6904;
wire net_6905;
wire net_6906;
wire net_6907;
wire net_6908;
wire net_6909;
wire net_6910;
wire net_6911;
wire net_6912;
wire net_6913;
wire net_6914;
wire net_6915;
wire net_6916;
wire net_6917;
wire net_6918;
wire net_6919;
wire net_6920;
wire net_6921;
wire net_6922;
wire net_6923;
wire net_6924;
wire net_6925;
wire net_6926;
wire net_6927;
wire net_6928;
wire net_6929;
wire net_6930;
wire net_6931;
wire net_6932;
wire net_6933;
wire net_6934;
wire net_6935;
wire net_6936;
wire net_6937;
wire net_6938;
wire net_6939;
wire net_6940;
wire net_6941;
wire net_6942;
wire net_6943;
wire net_6944;
wire net_6945;
wire net_6946;
wire net_6947;
wire net_6948;
wire net_6949;
wire net_6950;
wire net_6951;
wire net_6952;
wire net_6953;
wire net_6954;
wire net_6955;
wire net_6956;
wire net_6961;
wire net_6964;
wire net_6965;
wire net_6966;
wire net_6967;
wire net_6968;
wire net_6969;
wire net_6970;
wire net_6971;
wire net_6972;
wire net_6973;
wire net_6974;
wire net_6975;
wire net_6976;
wire net_6977;
wire net_6978;
wire net_6979;
wire net_6980;
wire net_6981;
wire net_6982;
wire net_6983;
wire net_6984;
wire net_6985;
wire net_6986;
wire net_6987;
wire net_6988;
wire net_6989;
wire net_6990;
wire net_6991;
wire net_6992;
wire net_6993;
wire net_6994;
wire net_6995;
wire net_6996;
wire net_6997;
wire net_6998;
wire net_6999;
wire net_7000;
wire net_7001;
wire net_7002;
wire net_7003;
wire net_7004;
wire net_7005;
wire net_7006;
wire net_7007;
wire net_7008;
wire net_7009;
wire net_7010;
wire net_7011;
wire net_7012;
wire net_7013;
wire net_7014;
wire net_7015;
wire net_7016;
wire net_7017;
wire net_7018;
wire net_7019;
wire net_7020;
wire net_7021;
wire net_7022;
wire net_7023;
wire net_7024;
wire net_7025;
wire net_7026;
wire net_7027;
wire net_7028;
wire net_7029;
wire net_7030;
wire net_7031;
wire net_7032;
wire net_7033;
wire net_7034;
wire net_7035;
wire net_7036;
wire net_7037;
wire net_7038;
wire net_7039;
wire net_7040;
wire net_7041;
wire net_7042;
wire net_7043;
wire net_7044;
wire net_7045;
wire net_7046;
wire net_7047;
wire net_7048;
wire net_7049;
wire net_7050;
wire net_7051;
wire net_7052;
wire net_7053;
wire net_7054;
wire net_7055;
wire net_7056;
wire net_7057;
wire net_7058;
wire net_7059;
wire net_7060;
wire net_7061;
wire net_7062;
wire net_7063;
wire net_7064;
wire net_7065;
wire net_7066;
wire net_7067;
wire net_7068;
wire net_7069;
wire net_7070;
wire net_7071;
wire net_7072;
wire net_7073;
wire net_7074;
wire net_7075;
wire net_7076;
wire net_7077;
wire net_7078;
wire net_7079;
wire net_7080;
wire net_7081;
wire net_7082;
wire net_7083;
wire net_7084;
wire net_7085;
wire net_7086;
wire net_7087;
wire net_7088;
wire net_7089;
wire net_7090;
wire net_7091;
wire net_7096;
wire net_7099;
wire net_7100;
wire net_7101;
wire net_7102;
wire net_7103;
wire net_7104;
wire net_7105;
wire net_7106;
wire net_7107;
wire net_7108;
wire net_7109;
wire net_7110;
wire net_7111;
wire net_7112;
wire net_7113;
wire net_7114;
wire net_7115;
wire net_7116;
wire net_7117;
wire net_7118;
wire net_7119;
wire net_7120;
wire net_7121;
wire net_7122;
wire net_7123;
wire net_7124;
wire net_7125;
wire net_7126;
wire net_7127;
wire net_7128;
wire net_7129;
wire net_7130;
wire net_7131;
wire net_7132;
wire net_7133;
wire net_7134;
wire net_7135;
wire net_7136;
wire net_7137;
wire net_7138;
wire net_7139;
wire net_7140;
wire net_7141;
wire net_7142;
wire net_7143;
wire net_7144;
wire net_7145;
wire net_7146;
wire net_7147;
wire net_7148;
wire net_7149;
wire net_7150;
wire net_7151;
wire net_7152;
wire net_7153;
wire net_7154;
wire net_7155;
wire net_7156;
wire net_7157;
wire net_7158;
wire net_7159;
wire net_7160;
wire net_7161;
wire net_7162;
wire net_7163;
wire net_7164;
wire net_7165;
wire net_7166;
wire net_7167;
wire net_7168;
wire net_7169;
wire net_7170;
wire net_7171;
wire net_7172;
wire net_7173;
wire net_7174;
wire net_7175;
wire net_7176;
wire net_7177;
wire net_7178;
wire net_7179;
wire net_7180;
wire net_7181;
wire net_7182;
wire net_7183;
wire net_7184;
wire net_7185;
wire net_7186;
wire net_7187;
wire net_7188;
wire net_7189;
wire net_7190;
wire net_7191;
wire net_7192;
wire net_7193;
wire net_7194;
wire net_7195;
wire net_7196;
wire net_7197;
wire net_7198;
wire net_7199;
wire net_7200;
wire net_7201;
wire net_7202;
wire net_7203;
wire net_7204;
wire net_7205;
wire net_7206;
wire net_7207;
wire net_7208;
wire net_7209;
wire net_7210;
wire net_7211;
wire net_7212;
wire net_7213;
wire net_7214;
wire net_7215;
wire net_7216;
wire net_7217;
wire net_7218;
wire net_7219;
wire net_7220;
wire net_7221;
wire net_7222;
wire net_7223;
wire net_7224;
wire net_7225;
wire net_7226;
wire net_7231;
wire net_7234;
wire net_7235;
wire net_7236;
wire net_7237;
wire net_7238;
wire net_7239;
wire net_7240;
wire net_7241;
wire net_7242;
wire net_7243;
wire net_7244;
wire net_7245;
wire net_7246;
wire net_7247;
wire net_7248;
wire net_7249;
wire net_7302;
wire net_7303;
wire net_7304;
wire net_7305;
wire net_7306;
wire net_7307;
wire net_7308;
wire net_7309;
wire net_7310;
wire net_7311;
wire net_7312;
wire net_7313;
wire net_7334;
wire net_7335;
wire net_7336;
wire net_7337;
wire net_7338;
wire net_7339;
wire net_7340;
wire net_7341;
wire net_7342;
wire net_7343;
wire net_7344;
wire net_7345;
wire net_7366;
wire net_7367;
wire net_7368;
wire net_7369;
wire net_7370;
wire net_7371;
wire net_7372;
wire net_7373;
wire net_7374;
wire net_7375;
wire net_7376;
wire net_7377;
wire net_7378;
wire net_7385;
wire net_7386;
wire net_7387;
wire net_7388;
wire net_7389;
wire net_7390;
wire net_7391;
wire net_7392;
wire net_7393;
wire net_7394;
wire net_7395;
wire net_7396;
wire net_7397;
wire net_7398;
wire net_7399;
wire net_7400;
wire net_7453;
wire net_7454;
wire net_7455;
wire net_7456;
wire net_7457;
wire net_7458;
wire net_7459;
wire net_7460;
wire net_7461;
wire net_7462;
wire net_7463;
wire net_7464;
wire net_7485;
wire net_7486;
wire net_7487;
wire net_7488;
wire net_7489;
wire net_7490;
wire net_7491;
wire net_7492;
wire net_7493;
wire net_7494;
wire net_7495;
wire net_7496;
wire net_7517;
wire net_7518;
wire net_7519;
wire net_7520;
wire net_7521;
wire net_7522;
wire net_7523;
wire net_7524;
wire net_7525;
wire net_7526;
wire net_7527;
wire net_7528;
wire net_7529;
wire net_7536;
wire net_7537;
wire net_7538;
wire net_7539;
wire net_7540;
wire net_7541;
wire net_7542;
wire net_7543;
wire net_7544;
wire net_7545;
wire net_7546;
wire net_7547;
wire net_7548;
wire net_7549;
wire net_7550;
wire net_7551;
wire net_7604;
wire net_7605;
wire net_7606;
wire net_7607;
wire net_7608;
wire net_7609;
wire net_7610;
wire net_7611;
wire net_7612;
wire net_7613;
wire net_7614;
wire net_7615;
wire net_7636;
wire net_7637;
wire net_7638;
wire net_7639;
wire net_7640;
wire net_7641;
wire net_7642;
wire net_7643;
wire net_7644;
wire net_7645;
wire net_7646;
wire net_7647;
wire net_7668;
wire net_7669;
wire net_7670;
wire net_7671;
wire net_7672;
wire net_7673;
wire net_7674;
wire net_7675;
wire net_7676;
wire net_7677;
wire net_7678;
wire net_7679;
wire net_7680;
wire net_7691;
wire net_7708;
wire net_7709;
wire net_7710;
wire net_7711;
wire net_7712;
wire net_7713;
wire net_7714;
wire net_7715;
wire net_7737;
wire net_7738;
wire net_7739;
wire net_7740;
wire net_7741;
wire net_7742;
wire net_7743;
wire net_7744;
wire net_7750;
wire net_7752;
wire net_7754;
wire net_7756;
wire net_7758;
wire net_7760;
wire net_7767;
wire net_7769;
wire net_7770;
wire net_7771;
wire net_7772;
wire net_7773;
wire net_7774;
wire net_7775;
wire net_7776;
wire net_7777;
wire net_7778;
wire net_7779;
wire net_7780;
wire net_7790;
wire net_7792;
wire net_7799;
wire net_7802;
wire net_7807;
wire x130629;
wire x130630;
wire x130631;
wire x130632;
wire x130633;
wire x130634;
wire x130635;
wire x130636;
wire x130637;
wire x130638;
wire x130639;
wire x130640;
wire x130641;
wire x130642;
wire x130643;
wire x130644;
wire x130645;
wire x130646;
wire x130647;
wire x130648;
wire x130649;
wire x130650;
wire x130651;
wire x130652;
wire x130653;
wire x130654;
wire x130655;
wire x130656;
wire x1822;
wire x821;

// Start cells
in01f01  g0000 ( .o(n6730), .a(net_6416) );
in01f01  g0001 ( .o(n6731), .a(net_6417) );
na02f01  g0002 ( .o(x30), .a(n6731), .b(n6730) );
in01f01  g0003 ( .o(n6733), .a(net_7680) );
no02f01  g0004 ( .o(n6734), .a(n6733), .b(_net_7681) );
in01f01  g0005 ( .o(n6735), .a(_net_7681) );
no02f01  g0006 ( .o(n6736_1), .a(net_7680), .b(n6735) );
ao22f01  g0007 ( .o(n6737), .a(n6736_1), .b(_net_7635), .c(n6734), .d(_net_7603) );
no02f01  g0008 ( .o(n6738), .a(net_7680), .b(_net_7681) );
no02f01  g0009 ( .o(n6739), .a(n6733), .b(n6735) );
ao22f01  g0010 ( .o(n6740), .a(n6739), .b(_net_7667), .c(n6738), .d(_net_7571) );
na02f01  g0011 ( .o(n266), .a(n6740), .b(n6737) );
ao22f01  g0012 ( .o(n6742), .a(n6736_1), .b(net_7640), .c(n6734), .d(net_7608) );
ao22f01  g0013 ( .o(n6743), .a(n6739), .b(net_7672), .c(n6738), .d(_net_7576) );
na02f01  g0014 ( .o(n271), .a(n6743), .b(n6742) );
in01f01  g0015 ( .o(n6745), .a(net_6438) );
in01f01  g0016 ( .o(n6746_1), .a(net_6502) );
in01f01  g0017 ( .o(n6747), .a(_net_6553) );
na02f01  g0018 ( .o(n6748), .a(_net_6554), .b(n6747) );
in01f01  g0019 ( .o(n6749_1), .a(_net_6554) );
na02f01  g0020 ( .o(n6750), .a(n6749_1), .b(n6747) );
oa22f01  g0021 ( .o(n6751), .a(n6750), .b(n6745), .c(n6748), .d(n6746_1) );
in01f01  g0022 ( .o(n6752_1), .a(net_6470) );
in01f01  g0023 ( .o(n6753), .a(net_6534) );
na02f01  g0024 ( .o(n6754), .a(_net_6554), .b(_net_6553) );
na02f01  g0025 ( .o(n6755), .a(n6749_1), .b(_net_6553) );
oa22f01  g0026 ( .o(n6756_1), .a(n6755), .b(n6752_1), .c(n6754), .d(n6753) );
no02f01  g0027 ( .o(n6757), .a(n6756_1), .b(n6751) );
in01f01  g0028 ( .o(n6758), .a(_net_6552) );
in01f01  g0029 ( .o(n6759), .a(_net_5984) );
in01f01  g0030 ( .o(n6760), .a(_net_7749) );
na03f01  g0031 ( .o(n6761_1), .a(_net_7791), .b(net_6061), .c(n6760) );
no02f01  g0032 ( .o(n6762), .a(n6761_1), .b(n6759) );
no02f01  g0033 ( .o(n6763), .a(_net_5986), .b(_net_5987) );
na03f01  g0034 ( .o(n6764), .a(n6763), .b(n6762), .c(n6758) );
no02f01  g0035 ( .o(n6765_1), .a(n6764), .b(n6757) );
na02f01  g0036 ( .o(n6766), .a(n6762), .b(_net_5986) );
in01f01  g0037 ( .o(n6767), .a(net_6440) );
in01f01  g0038 ( .o(n6768), .a(net_6504) );
oa22f01  g0039 ( .o(n6769), .a(n6750), .b(n6767), .c(n6748), .d(n6768) );
in01f01  g0040 ( .o(n6770_1), .a(net_6536) );
in01f01  g0041 ( .o(n6771), .a(net_6472) );
oa22f01  g0042 ( .o(n6772), .a(n6755), .b(n6771), .c(n6754), .d(n6770_1) );
no02f01  g0043 ( .o(n6773), .a(n6772), .b(n6769) );
no02f01  g0044 ( .o(n6774_1), .a(n6773), .b(n6766) );
na02f01  g0045 ( .o(n6775), .a(n6762), .b(_net_5987) );
in01f01  g0046 ( .o(n6776), .a(n6748) );
in01f01  g0047 ( .o(n6777), .a(n6750) );
ao22f01  g0048 ( .o(n6778), .a(n6777), .b(net_6442), .c(n6776), .d(net_6506) );
in01f01  g0049 ( .o(n6779_1), .a(n6754) );
in01f01  g0050 ( .o(n6780), .a(n6755) );
ao22f01  g0051 ( .o(n6781), .a(n6780), .b(net_6474), .c(n6779_1), .d(net_6538) );
ao12f01  g0052 ( .o(n6782), .a(n6775), .b(n6781), .c(n6778) );
in01f01  g0053 ( .o(n6783_1), .a(_net_6082) );
na02f01  g0054 ( .o(n6784), .a(n6761_1), .b(_net_5984) );
no02f01  g0055 ( .o(n6785), .a(n6784), .b(n6783_1) );
no04f01  g0056 ( .o(n6786), .a(n6785), .b(n6782), .c(n6774_1), .d(n6765_1) );
in01f01  g0057 ( .o(n6787), .a(net_6486) );
in01f01  g0058 ( .o(n6788_1), .a(net_6454) );
na04f01  g0059 ( .o(n6789), .a(n6763), .b(n6762), .c(n6780), .d(_net_6552) );
na04f01  g0060 ( .o(n6790), .a(n6763), .b(n6762), .c(n6777), .d(_net_6552) );
oa22f01  g0061 ( .o(n6791), .a(n6790), .b(n6788_1), .c(n6789), .d(n6787) );
in01f01  g0062 ( .o(n6792), .a(net_6550) );
in01f01  g0063 ( .o(n6793_1), .a(net_6518) );
na04f01  g0064 ( .o(n6794), .a(n6763), .b(n6762), .c(n6776), .d(_net_6552) );
na04f01  g0065 ( .o(n6795), .a(n6763), .b(n6762), .c(n6779_1), .d(_net_6552) );
oa22f01  g0066 ( .o(n6796_1), .a(n6795), .b(n6792), .c(n6794), .d(n6793_1) );
no02f01  g0067 ( .o(n6797), .a(n6796_1), .b(n6791) );
na02f01  g0068 ( .o(n281), .a(n6797), .b(n6786) );
in01f01  g0069 ( .o(n6799), .a(_net_7797) );
in01f01  g0070 ( .o(n6800), .a(x1322) );
in01f01  g0071 ( .o(n6801_1), .a(x1286) );
no02f01  g0072 ( .o(n6802), .a(n6801_1), .b(x1261) );
na03f01  g0073 ( .o(n6803), .a(n6802), .b(_net_6184), .c(n6800) );
na02f01  g0074 ( .o(n6804), .a(n6803), .b(_net_6032) );
oa12f01  g0075 ( .o(n295), .a(n6804), .b(n6803), .c(n6799) );
in01f01  g0076 ( .o(n6806_1), .a(_net_6958) );
na02f01  g0077 ( .o(n6807), .a(n6806_1), .b(_net_6959) );
in01f01  g0078 ( .o(n6808), .a(n6807) );
in01f01  g0079 ( .o(n6809_1), .a(_net_6959) );
na02f01  g0080 ( .o(n6810), .a(n6806_1), .b(n6809_1) );
in01f01  g0081 ( .o(n6811), .a(n6810) );
ao22f01  g0082 ( .o(n6812), .a(n6811), .b(net_6834), .c(n6808), .d(net_6898) );
na02f01  g0083 ( .o(n6813_1), .a(_net_6958), .b(_net_6959) );
in01f01  g0084 ( .o(n6814), .a(n6813_1) );
na02f01  g0085 ( .o(n6815), .a(_net_6958), .b(n6809_1) );
in01f01  g0086 ( .o(n6816), .a(n6815) );
ao22f01  g0087 ( .o(n6817), .a(n6816), .b(net_6866), .c(n6814), .d(net_6930) );
in01f01  g0088 ( .o(n6818_1), .a(_net_6957) );
in01f01  g0089 ( .o(n6819), .a(_net_6017) );
in01f01  g0090 ( .o(n6820), .a(_net_7755) );
na03f01  g0091 ( .o(n6821), .a(net_6058), .b(n6820), .c(_net_7791) );
no02f01  g0092 ( .o(n6822_1), .a(n6821), .b(n6819) );
no02f01  g0093 ( .o(n6823), .a(_net_6020), .b(_net_6019) );
na03f01  g0094 ( .o(n6824), .a(n6823), .b(n6822_1), .c(n6818_1) );
ao12f01  g0095 ( .o(n6825), .a(n6824), .b(n6817), .c(n6812) );
na02f01  g0096 ( .o(n6826_1), .a(n6822_1), .b(_net_6019) );
in01f01  g0097 ( .o(n6827), .a(net_6900) );
in01f01  g0098 ( .o(n6828), .a(net_6836) );
oa22f01  g0099 ( .o(n6829), .a(n6810), .b(n6828), .c(n6807), .d(n6827) );
in01f01  g0100 ( .o(n6830), .a(net_6868) );
in01f01  g0101 ( .o(n6831_1), .a(net_6932) );
oa22f01  g0102 ( .o(n6832), .a(n6815), .b(n6830), .c(n6813_1), .d(n6831_1) );
no02f01  g0103 ( .o(n6833), .a(n6832), .b(n6829) );
no02f01  g0104 ( .o(n6834), .a(n6833), .b(n6826_1) );
in01f01  g0105 ( .o(n6835), .a(_net_6133) );
na02f01  g0106 ( .o(n6836_1), .a(n6822_1), .b(_net_6020) );
in01f01  g0107 ( .o(n6837), .a(net_6902) );
in01f01  g0108 ( .o(n6838), .a(net_6838) );
oa22f01  g0109 ( .o(n6839), .a(n6810), .b(n6838), .c(n6807), .d(n6837) );
in01f01  g0110 ( .o(n6840_1), .a(net_6870) );
in01f01  g0111 ( .o(n6841), .a(net_6934) );
oa22f01  g0112 ( .o(n6842), .a(n6815), .b(n6840_1), .c(n6813_1), .d(n6841) );
no02f01  g0113 ( .o(n6843), .a(n6842), .b(n6839) );
na02f01  g0114 ( .o(n6844), .a(n6821), .b(_net_6017) );
oa22f01  g0115 ( .o(n6845_1), .a(n6844), .b(n6835), .c(n6843), .d(n6836_1) );
no03f01  g0116 ( .o(n6846), .a(n6845_1), .b(n6834), .c(n6825) );
in01f01  g0117 ( .o(n6847), .a(net_6850) );
in01f01  g0118 ( .o(n6848), .a(net_6882) );
na04f01  g0119 ( .o(n6849), .a(n6823), .b(n6822_1), .c(n6816), .d(_net_6957) );
na04f01  g0120 ( .o(n6850_1), .a(n6823), .b(n6822_1), .c(n6811), .d(_net_6957) );
oa22f01  g0121 ( .o(n6851), .a(n6850_1), .b(n6847), .c(n6849), .d(n6848) );
in01f01  g0122 ( .o(n6852), .a(net_6914) );
in01f01  g0123 ( .o(n6853), .a(net_6946) );
na04f01  g0124 ( .o(n6854), .a(n6823), .b(n6822_1), .c(n6808), .d(_net_6957) );
na04f01  g0125 ( .o(n6855_1), .a(n6823), .b(n6822_1), .c(n6814), .d(_net_6957) );
oa22f01  g0126 ( .o(n6856), .a(n6855_1), .b(n6853), .c(n6854), .d(n6852) );
no02f01  g0127 ( .o(n6857), .a(n6856), .b(n6851) );
na02f01  g0128 ( .o(n300), .a(n6857), .b(n6846) );
in01f01  g0129 ( .o(n6859), .a(_net_7481) );
in01f01  g0130 ( .o(n6860_1), .a(_net_7534) );
no02f01  g0131 ( .o(n6861), .a(_net_7533), .b(n6860_1) );
in01f01  g0132 ( .o(n6862), .a(n6861) );
in01f01  g0133 ( .o(n6863_1), .a(_net_5920) );
in01f01  g0134 ( .o(n6864), .a(net_5860) );
no03f01  g0135 ( .o(n6865), .a(n6864), .b(n6863_1), .c(_net_7763) );
no02f01  g0136 ( .o(n6866), .a(_net_281), .b(_net_280) );
in01f01  g0137 ( .o(n6867_1), .a(n6866) );
oa12f01  g0138 ( .o(n6868), .a(n6865), .b(n6867_1), .c(_net_7532) );
no02f01  g0139 ( .o(n6869), .a(n6868), .b(n6862) );
na02f01  g0140 ( .o(n6870), .a(n6866), .b(net_350) );
ao22f01  g0141 ( .o(n6871), .a(_net_281), .b(net_362), .c(net_364), .d(_net_280) );
na02f01  g0142 ( .o(n6872_1), .a(n6871), .b(n6870) );
na02f01  g0143 ( .o(n6873), .a(n6872_1), .b(n6869) );
oa12f01  g0144 ( .o(n314), .a(n6873), .b(n6869), .c(n6859) );
in01f01  g0145 ( .o(n6875), .a(_net_7379) );
no02f01  g0146 ( .o(n6876_1), .a(net_7378), .b(n6875) );
no02f01  g0147 ( .o(n6877), .a(net_7378), .b(_net_7379) );
ao22f01  g0148 ( .o(n6878), .a(n6877), .b(_net_7269), .c(n6876_1), .d(_net_7333) );
in01f01  g0149 ( .o(n6879), .a(net_7378) );
no02f01  g0150 ( .o(n6880), .a(n6879), .b(n6875) );
no02f01  g0151 ( .o(n6881_1), .a(n6879), .b(_net_7379) );
ao22f01  g0152 ( .o(n6882), .a(n6881_1), .b(_net_7301), .c(n6880), .d(_net_7365) );
na02f01  g0153 ( .o(n319), .a(n6882), .b(n6878) );
in01f01  g0154 ( .o(n6884), .a(_net_6062) );
in01f01  g0155 ( .o(n6885), .a(net_155) );
oa12f01  g0156 ( .o(n6886_1), .a(_net_7791), .b(net_155), .c(net_7767) );
oa22f01  g0157 ( .o(n329), .a(n6886_1), .b(n6885), .c(_net_7791), .d(n6884) );
in01f01  g0158 ( .o(n6888), .a(_net_7474) );
na02f01  g0159 ( .o(n6889), .a(n6866), .b(net_7394) );
ao22f01  g0160 ( .o(n6890_1), .a(_net_281), .b(net_355), .c(_net_280), .d(net_357) );
na02f01  g0161 ( .o(n6891), .a(n6890_1), .b(n6889) );
na02f01  g0162 ( .o(n6892), .a(n6891), .b(n6869) );
oa12f01  g0163 ( .o(n370), .a(n6892), .b(n6869), .c(n6888) );
in01f01  g0164 ( .o(n6894), .a(_net_7252) );
in01f01  g0165 ( .o(n6895_1), .a(net_5861) );
in01f01  g0166 ( .o(n6896), .a(_net_5922) );
no03f01  g0167 ( .o(n6897), .a(_net_7761), .b(n6896), .c(n6895_1) );
no02f01  g0168 ( .o(n6898), .a(_net_269), .b(_net_270) );
in01f01  g0169 ( .o(n6899_1), .a(n6898) );
oa12f01  g0170 ( .o(n6900), .a(n6897), .b(n6899_1), .c(_net_7381) );
no03f01  g0171 ( .o(n6901), .a(n6900), .b(_net_7383), .c(_net_7382) );
na02f01  g0172 ( .o(n6902_1), .a(n6898), .b(net_7236) );
ao22f01  g0173 ( .o(n6903), .a(net_328), .b(_net_270), .c(net_330), .d(_net_269) );
na02f01  g0174 ( .o(n6904), .a(n6903), .b(n6902_1) );
na02f01  g0175 ( .o(n6905), .a(n6904), .b(n6901) );
oa12f01  g0176 ( .o(n375), .a(n6905), .b(n6901), .c(n6894) );
in01f01  g0177 ( .o(n6907), .a(_net_298) );
na02f01  g0178 ( .o(n6908), .a(_net_262), .b(_net_264) );
na02f01  g0179 ( .o(n380), .a(n6908), .b(n6907) );
in01f01  g0180 ( .o(n6910_1), .a(x38) );
na02f01  g0181 ( .o(n385), .a(n6910_1), .b(_net_6404) );
in01f01  g0182 ( .o(n6912), .a(_net_5995) );
in01f01  g0183 ( .o(n6913), .a(_net_7751) );
na03f01  g0184 ( .o(n6914), .a(_net_7791), .b(n6913), .c(net_6060) );
no02f01  g0185 ( .o(n6915_1), .a(n6914), .b(n6912) );
na02f01  g0186 ( .o(n6916), .a(n6915_1), .b(_net_5998) );
in01f01  g0187 ( .o(n6917), .a(n6916) );
in01f01  g0188 ( .o(n6918), .a(_net_6688) );
na02f01  g0189 ( .o(n6919_1), .a(_net_6689), .b(n6918) );
in01f01  g0190 ( .o(n6920), .a(n6919_1) );
in01f01  g0191 ( .o(n6921), .a(_net_6689) );
na02f01  g0192 ( .o(n6922), .a(n6921), .b(n6918) );
in01f01  g0193 ( .o(n6923), .a(n6922) );
ao22f01  g0194 ( .o(n6924_1), .a(n6923), .b(net_6563), .c(n6920), .d(net_6627) );
na02f01  g0195 ( .o(n6925), .a(_net_6689), .b(_net_6688) );
in01f01  g0196 ( .o(n6926), .a(n6925) );
na02f01  g0197 ( .o(n6927), .a(n6921), .b(_net_6688) );
in01f01  g0198 ( .o(n6928), .a(n6927) );
ao22f01  g0199 ( .o(n6929_1), .a(n6928), .b(net_6595), .c(n6926), .d(net_6659) );
na02f01  g0200 ( .o(n6930), .a(n6929_1), .b(n6924_1) );
na02f01  g0201 ( .o(n6931), .a(n6930), .b(n6917) );
na02f01  g0202 ( .o(n6932), .a(n6914), .b(_net_5995) );
in01f01  g0203 ( .o(n6933), .a(n6932) );
na02f01  g0204 ( .o(n6934_1), .a(n6915_1), .b(_net_5997) );
in01f01  g0205 ( .o(n6935), .a(n6934_1) );
ao22f01  g0206 ( .o(n6936), .a(n6923), .b(net_6561), .c(n6920), .d(net_6625) );
ao22f01  g0207 ( .o(n6937), .a(n6928), .b(net_6593), .c(n6926), .d(net_6657) );
na02f01  g0208 ( .o(n6938_1), .a(n6937), .b(n6936) );
ao22f01  g0209 ( .o(n6939), .a(n6938_1), .b(n6935), .c(n6933), .d(_net_6088) );
ao22f01  g0210 ( .o(n6940), .a(n6923), .b(net_6559), .c(n6920), .d(net_6623) );
ao22f01  g0211 ( .o(n6941), .a(n6928), .b(net_6591), .c(n6926), .d(net_6655) );
na02f01  g0212 ( .o(n6942), .a(n6941), .b(n6940) );
in01f01  g0213 ( .o(n6943_1), .a(_net_6687) );
no02f01  g0214 ( .o(n6944), .a(_net_5998), .b(_net_5997) );
na03f01  g0215 ( .o(n6945), .a(n6944), .b(n6915_1), .c(n6943_1) );
in01f01  g0216 ( .o(n6946), .a(n6945) );
na02f01  g0217 ( .o(n6947_1), .a(n6944), .b(n6915_1) );
in01f01  g0218 ( .o(n6948), .a(net_6639) );
in01f01  g0219 ( .o(n6949), .a(net_6575) );
oa22f01  g0220 ( .o(n6950), .a(n6922), .b(n6949), .c(n6919_1), .d(n6948) );
in01f01  g0221 ( .o(n6951), .a(net_6671) );
in01f01  g0222 ( .o(n6952_1), .a(net_6607) );
oa22f01  g0223 ( .o(n6953), .a(n6927), .b(n6952_1), .c(n6925), .d(n6951) );
no02f01  g0224 ( .o(n6954), .a(n6953), .b(n6950) );
no03f01  g0225 ( .o(n6955), .a(n6954), .b(n6947_1), .c(n6943_1) );
ao12f01  g0226 ( .o(n6956), .a(n6955), .b(n6946), .c(n6942) );
na03f01  g0227 ( .o(n390), .a(n6956), .b(n6939), .c(n6931) );
in01f01  g0228 ( .o(n6958), .a(_net_7595) );
in01f01  g0229 ( .o(n6959), .a(_net_7684) );
no02f01  g0230 ( .o(n6960_1), .a(_net_7685), .b(n6959) );
in01f01  g0231 ( .o(n6961), .a(n6960_1) );
in01f01  g0232 ( .o(n6962), .a(net_5858) );
in01f01  g0233 ( .o(n6963), .a(_net_5924) );
no03f01  g0234 ( .o(n6964_1), .a(n6963), .b(n6962), .c(_net_7765) );
no02f01  g0235 ( .o(n6965), .a(_net_292), .b(_net_291) );
in01f01  g0236 ( .o(n6966), .a(n6965) );
oa12f01  g0237 ( .o(n6967), .a(n6964_1), .b(n6966), .c(_net_7683) );
no02f01  g0238 ( .o(n6968), .a(n6967), .b(n6961) );
na02f01  g0239 ( .o(n6969_1), .a(n6965), .b(net_7547) );
ao22f01  g0240 ( .o(n6970), .a(_net_292), .b(net_377), .c(_net_291), .d(net_379) );
na02f01  g0241 ( .o(n6971), .a(n6970), .b(n6969_1) );
na02f01  g0242 ( .o(n6972), .a(n6971), .b(n6968) );
oa12f01  g0243 ( .o(n400), .a(n6972), .b(n6968), .c(n6958) );
in01f01  g0244 ( .o(n6974_1), .a(net_362) );
no02f01  g0245 ( .o(n420), .a(n6867_1), .b(n6974_1) );
in01f01  g0246 ( .o(n6976), .a(_net_6028) );
in01f01  g0247 ( .o(n6977_1), .a(_net_7757) );
na03f01  g0248 ( .o(n6978), .a(n6977_1), .b(_net_7791), .c(net_6057) );
no02f01  g0249 ( .o(n6979), .a(n6978), .b(n6976) );
na02f01  g0250 ( .o(n6980), .a(n6979), .b(_net_6031) );
in01f01  g0251 ( .o(n6981), .a(n6980) );
in01f01  g0252 ( .o(n6982_1), .a(net_7034) );
in01f01  g0253 ( .o(n6983), .a(net_6970) );
in01f01  g0254 ( .o(n6984), .a(_net_7093) );
na02f01  g0255 ( .o(n6985), .a(n6984), .b(_net_7094) );
in01f01  g0256 ( .o(n6986_1), .a(_net_7094) );
na02f01  g0257 ( .o(n6987), .a(n6984), .b(n6986_1) );
oa22f01  g0258 ( .o(n6988), .a(n6987), .b(n6983), .c(n6985), .d(n6982_1) );
in01f01  g0259 ( .o(n6989), .a(net_7066) );
in01f01  g0260 ( .o(n6990_1), .a(net_7002) );
na02f01  g0261 ( .o(n6991), .a(_net_7093), .b(_net_7094) );
na02f01  g0262 ( .o(n6992), .a(_net_7093), .b(n6986_1) );
oa22f01  g0263 ( .o(n6993), .a(n6992), .b(n6990_1), .c(n6991), .d(n6989) );
oa12f01  g0264 ( .o(n6994), .a(n6981), .b(n6993), .c(n6988) );
na02f01  g0265 ( .o(n6995_1), .a(n6978), .b(_net_6028) );
in01f01  g0266 ( .o(n6996), .a(n6995_1) );
na02f01  g0267 ( .o(n6997), .a(n6979), .b(_net_6030) );
in01f01  g0268 ( .o(n6998), .a(n6997) );
in01f01  g0269 ( .o(n6999), .a(n6985) );
in01f01  g0270 ( .o(n7000_1), .a(n6987) );
ao22f01  g0271 ( .o(n7001), .a(n7000_1), .b(net_6968), .c(n6999), .d(net_7032) );
in01f01  g0272 ( .o(n7002), .a(n6991) );
in01f01  g0273 ( .o(n7003), .a(n6992) );
ao22f01  g0274 ( .o(n7004), .a(n7003), .b(net_7000), .c(n7002), .d(net_7064) );
na02f01  g0275 ( .o(n7005_1), .a(n7004), .b(n7001) );
ao22f01  g0276 ( .o(n7006), .a(n7005_1), .b(n6998), .c(n6996), .d(_net_6150) );
ao22f01  g0277 ( .o(n7007), .a(n7000_1), .b(net_6966), .c(n6999), .d(net_7030) );
ao22f01  g0278 ( .o(n7008), .a(n7003), .b(net_6998), .c(n7002), .d(net_7062) );
na02f01  g0279 ( .o(n7009_1), .a(n7008), .b(n7007) );
in01f01  g0280 ( .o(n7010), .a(_net_7092) );
no02f01  g0281 ( .o(n7011), .a(_net_6031), .b(_net_6030) );
na03f01  g0282 ( .o(n7012), .a(n7011), .b(n6979), .c(n7010) );
in01f01  g0283 ( .o(n7013_1), .a(n7012) );
na02f01  g0284 ( .o(n7014), .a(n7013_1), .b(n7009_1) );
in01f01  g0285 ( .o(n7015), .a(net_6982) );
in01f01  g0286 ( .o(n7016), .a(net_7046) );
oa22f01  g0287 ( .o(n7017), .a(n6987), .b(n7015), .c(n6985), .d(n7016) );
in01f01  g0288 ( .o(n7018_1), .a(net_7014) );
in01f01  g0289 ( .o(n7019), .a(net_7078) );
oa22f01  g0290 ( .o(n7020), .a(n6992), .b(n7018_1), .c(n6991), .d(n7019) );
na02f01  g0291 ( .o(n7021), .a(n7011), .b(n6979) );
no02f01  g0292 ( .o(n7022), .a(n7021), .b(n7010) );
oa12f01  g0293 ( .o(n7023_1), .a(n7022), .b(n7020), .c(n7017) );
na04f01  g0294 ( .o(n447), .a(n7023_1), .b(n7014), .c(n7006), .d(n6994) );
in01f01  g0295 ( .o(n7025), .a(_net_7355) );
in01f01  g0296 ( .o(n7026), .a(_net_7382) );
in01f01  g0297 ( .o(n7027_1), .a(_net_7383) );
no02f01  g0298 ( .o(n7028), .a(n7027_1), .b(n7026) );
in01f01  g0299 ( .o(n7029), .a(n7028) );
no02f01  g0300 ( .o(n7030), .a(n7029), .b(n6900) );
na02f01  g0301 ( .o(n7031), .a(n6898), .b(net_7243) );
ao22f01  g0302 ( .o(n7032_1), .a(net_335), .b(_net_270), .c(_net_269), .d(net_337) );
na02f01  g0303 ( .o(n7033), .a(n7032_1), .b(n7031) );
na02f01  g0304 ( .o(n7034), .a(n7033), .b(n7030) );
oa12f01  g0305 ( .o(n460), .a(n7034), .b(n7030), .c(n7025) );
in01f01  g0306 ( .o(n7036_1), .a(net_6635) );
in01f01  g0307 ( .o(n7037), .a(net_6571) );
oa22f01  g0308 ( .o(n7038), .a(n6922), .b(n7037), .c(n6919_1), .d(n7036_1) );
in01f01  g0309 ( .o(n7039), .a(net_6603) );
in01f01  g0310 ( .o(n7040), .a(net_6667) );
oa22f01  g0311 ( .o(n7041_1), .a(n6927), .b(n7039), .c(n6925), .d(n7040) );
no02f01  g0312 ( .o(n7042), .a(n7041_1), .b(n7038) );
no02f01  g0313 ( .o(n7043), .a(n7042), .b(n6945) );
in01f01  g0314 ( .o(n7044), .a(net_6637) );
in01f01  g0315 ( .o(n7045_1), .a(net_6573) );
oa22f01  g0316 ( .o(n7046), .a(n6922), .b(n7045_1), .c(n6919_1), .d(n7044) );
in01f01  g0317 ( .o(n7047), .a(net_6605) );
in01f01  g0318 ( .o(n7048), .a(net_6669) );
oa22f01  g0319 ( .o(n7049_1), .a(n6927), .b(n7047), .c(n6925), .d(n7048) );
no02f01  g0320 ( .o(n7050), .a(n7049_1), .b(n7046) );
no02f01  g0321 ( .o(n7051), .a(n7050), .b(n6934_1) );
in01f01  g0322 ( .o(n7052), .a(_net_6100) );
oa22f01  g0323 ( .o(n7053_1), .a(n6954), .b(n6916), .c(n6932), .d(n7052) );
no03f01  g0324 ( .o(n7054), .a(n7053_1), .b(n7051), .c(n7043) );
in01f01  g0325 ( .o(n7055), .a(net_6619) );
in01f01  g0326 ( .o(n7056), .a(net_6587) );
na04f01  g0327 ( .o(n7057), .a(n6944), .b(n6928), .c(n6915_1), .d(_net_6687) );
na04f01  g0328 ( .o(n7058_1), .a(n6944), .b(n6923), .c(n6915_1), .d(_net_6687) );
oa22f01  g0329 ( .o(n7059), .a(n7058_1), .b(n7056), .c(n7057), .d(n7055) );
in01f01  g0330 ( .o(n7060), .a(net_6651) );
in01f01  g0331 ( .o(n7061), .a(net_6683) );
na04f01  g0332 ( .o(n7062_1), .a(n6944), .b(n6920), .c(n6915_1), .d(_net_6687) );
na04f01  g0333 ( .o(n7063), .a(n6944), .b(n6926), .c(n6915_1), .d(_net_6687) );
oa22f01  g0334 ( .o(n7064), .a(n7063), .b(n7061), .c(n7062_1), .d(n7060) );
no02f01  g0335 ( .o(n7065), .a(n7064), .b(n7059) );
na02f01  g0336 ( .o(n465), .a(n7065), .b(n7054) );
in01f01  g0337 ( .o(n7067_1), .a(_net_5967) );
no02f01  g0338 ( .o(n513), .a(n6912), .b(n7067_1) );
in01f01  g0339 ( .o(n7069), .a(net_337) );
no02f01  g0340 ( .o(n518), .a(n6899_1), .b(n7069) );
in01f01  g0341 ( .o(n7071), .a(net_6435) );
in01f01  g0342 ( .o(n7072_1), .a(net_6499) );
oa22f01  g0343 ( .o(n7073), .a(n6750), .b(n7071), .c(n6748), .d(n7072_1) );
in01f01  g0344 ( .o(n7074), .a(net_6467) );
in01f01  g0345 ( .o(n7075), .a(net_6531) );
oa22f01  g0346 ( .o(n7076), .a(n6755), .b(n7074), .c(n6754), .d(n7075) );
no02f01  g0347 ( .o(n7077_1), .a(n7076), .b(n7073) );
no02f01  g0348 ( .o(n7078), .a(n7077_1), .b(n6764) );
in01f01  g0349 ( .o(n7079), .a(net_6501) );
in01f01  g0350 ( .o(n7080), .a(net_6437) );
oa22f01  g0351 ( .o(n7081), .a(n6750), .b(n7080), .c(n6748), .d(n7079) );
in01f01  g0352 ( .o(n7082_1), .a(net_6469) );
in01f01  g0353 ( .o(n7083), .a(net_6533) );
oa22f01  g0354 ( .o(n7084), .a(n6755), .b(n7082_1), .c(n6754), .d(n7083) );
no02f01  g0355 ( .o(n7085_1), .a(n7084), .b(n7081) );
no02f01  g0356 ( .o(n7086), .a(n7085_1), .b(n6766) );
in01f01  g0357 ( .o(n7087), .a(_net_6079) );
in01f01  g0358 ( .o(n7088), .a(net_6439) );
in01f01  g0359 ( .o(n7089_1), .a(net_6503) );
oa22f01  g0360 ( .o(n7090), .a(n6750), .b(n7088), .c(n6748), .d(n7089_1) );
in01f01  g0361 ( .o(n7091), .a(net_6471) );
in01f01  g0362 ( .o(n7092), .a(net_6535) );
oa22f01  g0363 ( .o(n7093_1), .a(n6755), .b(n7091), .c(n6754), .d(n7092) );
no02f01  g0364 ( .o(n7094), .a(n7093_1), .b(n7090) );
oa22f01  g0365 ( .o(n7095), .a(n7094), .b(n6775), .c(n6784), .d(n7087) );
no03f01  g0366 ( .o(n7096), .a(n7095), .b(n7086), .c(n7078) );
in01f01  g0367 ( .o(n7097), .a(net_6451) );
in01f01  g0368 ( .o(n7098_1), .a(net_6483) );
oa22f01  g0369 ( .o(n7099), .a(n6790), .b(n7097), .c(n6789), .d(n7098_1) );
in01f01  g0370 ( .o(n7100), .a(net_6515) );
in01f01  g0371 ( .o(n7101), .a(net_6547) );
oa22f01  g0372 ( .o(n7102_1), .a(n6795), .b(n7101), .c(n6794), .d(n7100) );
no02f01  g0373 ( .o(n7103), .a(n7102_1), .b(n7099) );
na02f01  g0374 ( .o(n523), .a(n7103), .b(n7096) );
in01f01  g0375 ( .o(n7105), .a(x1155) );
in01f01  g0376 ( .o(n7106), .a(x1101) );
in01f01  g0377 ( .o(n7107_1), .a(x1126) );
no02f01  g0378 ( .o(n7108), .a(n7107_1), .b(n7106) );
in01f01  g0379 ( .o(n7109), .a(_net_7689) );
no03f01  g0380 ( .o(n7110), .a(_net_7690), .b(n7109), .c(n7105) );
na02f01  g0381 ( .o(n7111_1), .a(n7110), .b(n7108) );
in01f01  g0382 ( .o(n7112), .a(n7111_1) );
no03f01  g0383 ( .o(n7113), .a(x1193), .b(x1209), .c(x1203) );
na02f01  g0384 ( .o(n7114), .a(n7113), .b(n7108) );
no03f01  g0385 ( .o(n528), .a(n7114), .b(n7112), .c(n7105) );
in01f01  g0386 ( .o(n7116_1), .a(_net_7753) );
na03f01  g0387 ( .o(n7117), .a(_net_7791), .b(net_6059), .c(n7116_1) );
na02f01  g0388 ( .o(n7118), .a(n7117), .b(_net_6006) );
in01f01  g0389 ( .o(n7119), .a(n7118) );
na02f01  g0390 ( .o(n7120_1), .a(n7119), .b(_net_6104) );
in01f01  g0391 ( .o(n7121), .a(_net_6006) );
no02f01  g0392 ( .o(n7122), .a(n7117), .b(n7121) );
na02f01  g0393 ( .o(n7123), .a(n7122), .b(_net_6009) );
in01f01  g0394 ( .o(n7124), .a(n7123) );
in01f01  g0395 ( .o(n7125_1), .a(_net_6823) );
na02f01  g0396 ( .o(n7126), .a(_net_6824), .b(n7125_1) );
in01f01  g0397 ( .o(n7127), .a(n7126) );
in01f01  g0398 ( .o(n7128_1), .a(_net_6824) );
na02f01  g0399 ( .o(n7129), .a(n7128_1), .b(n7125_1) );
in01f01  g0400 ( .o(n7130), .a(n7129) );
ao22f01  g0401 ( .o(n7131), .a(n7130), .b(net_6694), .c(n7127), .d(net_6758) );
na02f01  g0402 ( .o(n7132), .a(_net_6824), .b(_net_6823) );
in01f01  g0403 ( .o(n7133_1), .a(n7132) );
na02f01  g0404 ( .o(n7134), .a(n7128_1), .b(_net_6823) );
in01f01  g0405 ( .o(n7135), .a(n7134) );
ao22f01  g0406 ( .o(n7136), .a(n7135), .b(net_6726), .c(n7133_1), .d(net_6790) );
na02f01  g0407 ( .o(n7137), .a(n7136), .b(n7131) );
na02f01  g0408 ( .o(n7138_1), .a(n7137), .b(n7124) );
na02f01  g0409 ( .o(n533), .a(n7138_1), .b(n7120_1) );
in01f01  g0410 ( .o(n7140), .a(_net_7603) );
in01f01  g0411 ( .o(n7141), .a(net_373) );
in01f01  g0412 ( .o(n7142_1), .a(net_385) );
in01f01  g0413 ( .o(n7143), .a(_net_292) );
oa22f01  g0414 ( .o(n7144), .a(n6966), .b(n7141), .c(n7143), .d(n7142_1) );
na02f01  g0415 ( .o(n7145), .a(n7144), .b(n6968) );
oa12f01  g0416 ( .o(n538), .a(n7145), .b(n6968), .c(n7140) );
in01f01  g0417 ( .o(n7147_1), .a(_net_7316) );
no02f01  g0418 ( .o(n7148), .a(n7027_1), .b(_net_7382) );
in01f01  g0419 ( .o(n7149), .a(n7148) );
no02f01  g0420 ( .o(n7150), .a(n7149), .b(n6900) );
na02f01  g0421 ( .o(n7151_1), .a(n7150), .b(n6904) );
oa12f01  g0422 ( .o(n543), .a(n7151_1), .b(n7150), .c(n7147_1) );
in01f01  g0423 ( .o(n7153), .a(net_6691) );
no02f01  g0424 ( .o(n7154), .a(n6918), .b(n7153) );
no02f01  g0425 ( .o(n7155_1), .a(_net_6688), .b(net_6691) );
no02f01  g0426 ( .o(n7156), .a(n7155_1), .b(n7154) );
in01f01  g0427 ( .o(n548), .a(n7156) );
in01f01  g0428 ( .o(n7158), .a(net_6057) );
in01f01  g0429 ( .o(n7159), .a(net_6061) );
in01f01  g0430 ( .o(n7160_1), .a(net_6056) );
in01f01  g0431 ( .o(n7161), .a(net_6058) );
na04f01  g0432 ( .o(n7162), .a(n7161), .b(n7160_1), .c(n7159), .d(n7158) );
in01f01  g0433 ( .o(n7163), .a(net_6060) );
in01f01  g0434 ( .o(n7164_1), .a(net_6059) );
in01f01  g0435 ( .o(n7165), .a(_net_6063) );
na04f01  g0436 ( .o(n7166), .a(n7165), .b(n7164_1), .c(n7163), .d(n6884) );
oa12f01  g0437 ( .o(n7167_1), .a(_net_392), .b(n7166), .c(n7162) );
in01f01  g0438 ( .o(n7168), .a(_net_392) );
na02f01  g0439 ( .o(n7169), .a(n7168), .b(_net_6199) );
na02f01  g0440 ( .o(n553), .a(n7169), .b(n7167_1) );
in01f01  g0441 ( .o(n7171), .a(_net_6293) );
no02f01  g0442 ( .o(n561), .a(_net_392), .b(n7171) );
in01f01  g0443 ( .o(n7173), .a(net_342) );
no02f01  g0444 ( .o(n576), .a(n6899_1), .b(n7173) );
in01f01  g0445 ( .o(n7175), .a(net_361) );
no02f01  g0446 ( .o(n595), .a(n6867_1), .b(n7175) );
in01f01  g0447 ( .o(n7177_1), .a(_net_7285) );
no02f01  g0448 ( .o(n7178), .a(_net_7383), .b(n7026) );
in01f01  g0449 ( .o(n7179), .a(n7178) );
no02f01  g0450 ( .o(n7180), .a(n7179), .b(n6900) );
na02f01  g0451 ( .o(n7181), .a(n6898), .b(net_7237) );
ao22f01  g0452 ( .o(n7182_1), .a(_net_269), .b(net_331), .c(_net_270), .d(net_329) );
na02f01  g0453 ( .o(n7183), .a(n7182_1), .b(n7181) );
na02f01  g0454 ( .o(n7184), .a(n7183), .b(n7180) );
oa12f01  g0455 ( .o(n600), .a(n7184), .b(n7180), .c(n7177_1) );
in01f01  g0456 ( .o(n7186), .a(_net_6209) );
no02f01  g0457 ( .o(n605), .a(_net_392), .b(n7186) );
in01f01  g0458 ( .o(n7188), .a(net_374) );
no02f01  g0459 ( .o(n615), .a(n6966), .b(n7188) );
in01f01  g0460 ( .o(n7190_1), .a(_net_6004) );
in01f01  g0461 ( .o(n7191), .a(_net_5964) );
oa12f01  g0462 ( .o(n620), .a(n7190_1), .b(n6914), .c(n7191) );
in01f01  g0463 ( .o(n7193), .a(_net_7441) );
in01f01  g0464 ( .o(n7194_1), .a(_net_7533) );
no02f01  g0465 ( .o(n7195), .a(n7194_1), .b(_net_7534) );
in01f01  g0466 ( .o(n7196), .a(n7195) );
no02f01  g0467 ( .o(n7197), .a(n7196), .b(n6868) );
na02f01  g0468 ( .o(n7198), .a(n6866), .b(net_7393) );
ao22f01  g0469 ( .o(n7199_1), .a(net_354), .b(_net_281), .c(net_356), .d(_net_280) );
na02f01  g0470 ( .o(n7200), .a(n7199_1), .b(n7198) );
na02f01  g0471 ( .o(n7201), .a(n7200), .b(n7197) );
oa12f01  g0472 ( .o(n629), .a(n7201), .b(n7197), .c(n7193) );
in01f01  g0473 ( .o(n7203_1), .a(net_356) );
no02f01  g0474 ( .o(n634), .a(n6867_1), .b(n7203_1) );
in01f01  g0475 ( .o(n7205), .a(_net_7694) );
na02f01  g0476 ( .o(n7206), .a(_net_6184), .b(x1261) );
no03f01  g0477 ( .o(n7207_1), .a(n7206), .b(x1286), .c(n6800) );
na02f01  g0478 ( .o(n7208), .a(n7207_1), .b(_net_7796) );
oa12f01  g0479 ( .o(n639), .a(n7208), .b(n7207_1), .c(n7205) );
no02f01  g0480 ( .o(n7210), .a(n7010), .b(n6984) );
na02f01  g0481 ( .o(n7211), .a(n7210), .b(n6986_1) );
in01f01  g0482 ( .o(n7212_1), .a(n7210) );
na02f01  g0483 ( .o(n7213), .a(n7212_1), .b(_net_7094) );
na02f01  g0484 ( .o(n7214), .a(n7213), .b(n7211) );
no04f01  g0485 ( .o(n7215), .a(n6978), .b(_net_6031), .c(n6976), .d(_net_6030) );
na02f01  g0486 ( .o(n7216_1), .a(n7215), .b(n7214) );
na02f01  g0487 ( .o(n7217), .a(n6992), .b(n6985) );
no03f01  g0488 ( .o(n7218), .a(n7011), .b(n6978), .c(n6976) );
in01f01  g0489 ( .o(n7219), .a(n6978) );
no02f01  g0490 ( .o(n7220), .a(n7219), .b(n6976) );
ao22f01  g0491 ( .o(n7221_1), .a(n7220), .b(_net_7094), .c(n7218), .d(n7217) );
na02f01  g0492 ( .o(n644), .a(n7221_1), .b(n7216_1) );
in01f01  g0493 ( .o(n7223), .a(net_7529) );
no02f01  g0494 ( .o(n7224), .a(_net_7530), .b(n7223) );
no02f01  g0495 ( .o(n7225), .a(_net_7530), .b(net_7529) );
ao22f01  g0496 ( .o(n7226_1), .a(n7225), .b(_net_7420), .c(n7224), .d(_net_7452) );
in01f01  g0497 ( .o(n7227), .a(_net_7530) );
no02f01  g0498 ( .o(n7228), .a(n7227), .b(net_7529) );
no02f01  g0499 ( .o(n7229), .a(n7227), .b(n7223) );
ao22f01  g0500 ( .o(n7230_1), .a(n7229), .b(_net_7516), .c(n7228), .d(_net_7484) );
na02f01  g0501 ( .o(n649), .a(n7230_1), .b(n7226_1) );
in01f01  g0502 ( .o(n7232), .a(_net_7791) );
no02f01  g0503 ( .o(n654), .a(n7232), .b(n7164_1) );
ao22f01  g0504 ( .o(n7234), .a(n6877), .b(_net_7254), .c(n6876_1), .d(_net_7318) );
ao22f01  g0505 ( .o(n7235_1), .a(n6881_1), .b(_net_7286), .c(n6880), .d(_net_7350) );
na02f01  g0506 ( .o(n659), .a(n7235_1), .b(n7234) );
in01f01  g0507 ( .o(n7237), .a(_net_6207) );
no02f01  g0508 ( .o(n673), .a(_net_392), .b(n7237) );
in01f01  g0509 ( .o(n7239), .a(_net_7330) );
na02f01  g0510 ( .o(n7240_1), .a(n6898), .b(net_330) );
ao22f01  g0511 ( .o(n7241), .a(net_344), .b(_net_269), .c(net_342), .d(_net_270) );
na02f01  g0512 ( .o(n7242), .a(n7241), .b(n7240_1) );
na02f01  g0513 ( .o(n7243), .a(n7242), .b(n7150) );
oa12f01  g0514 ( .o(n688), .a(n7243), .b(n7150), .c(n7239) );
in01f01  g0515 ( .o(n7245_1), .a(_net_7271) );
in01f01  g0516 ( .o(n7246), .a(net_335) );
no02f01  g0517 ( .o(n1350), .a(n6899_1), .b(n7246) );
na02f01  g0518 ( .o(n7248), .a(n1350), .b(n6901) );
oa12f01  g0519 ( .o(n693), .a(n7248), .b(n6901), .c(n7245_1) );
in01f01  g0520 ( .o(n7250), .a(net_383) );
no02f01  g0521 ( .o(n698), .a(n6966), .b(n7250) );
in01f01  g0522 ( .o(n7252_1), .a(_net_7300) );
in01f01  g0523 ( .o(n7253), .a(_net_270) );
in01f01  g0524 ( .o(n7254), .a(net_344) );
in01f01  g0525 ( .o(n7255), .a(net_332) );
oa22f01  g0526 ( .o(n7256_1), .a(n6899_1), .b(n7255), .c(n7254), .d(n7253) );
na02f01  g0527 ( .o(n7257), .a(n7256_1), .b(n7180) );
oa12f01  g0528 ( .o(n708), .a(n7257), .b(n7180), .c(n7252_1) );
in01f01  g0529 ( .o(n7259), .a(_net_6010) );
no02f01  g0530 ( .o(n7260_1), .a(n7259), .b(_net_6011) );
in01f01  g0531 ( .o(n7261), .a(_net_5968) );
na02f01  g0532 ( .o(n7262), .a(_net_6006), .b(_net_6012) );
ao12f01  g0533 ( .o(n7263), .a(n7262), .b(_net_5970), .c(n7261) );
na02f01  g0534 ( .o(n7264), .a(n7263), .b(n7260_1) );
in01f01  g0535 ( .o(n7265_1), .a(_net_6011) );
in01f01  g0536 ( .o(n7266), .a(n7262) );
na03f01  g0537 ( .o(n7267), .a(_net_5970), .b(n7261), .c(_net_5969) );
na04f01  g0538 ( .o(n7268), .a(n7267), .b(n7266), .c(n7259), .d(n7265_1) );
oa12f01  g0539 ( .o(n7269), .a(n7261), .b(_net_5970), .c(_net_5969) );
na04f01  g0540 ( .o(n7270_1), .a(n7269), .b(n7266), .c(n7259), .d(_net_6011) );
no02f01  g0541 ( .o(n7271), .a(n7259), .b(n7265_1) );
na03f01  g0542 ( .o(n7272), .a(n7271), .b(n7266), .c(_net_5968) );
na04f01  g0543 ( .o(n7273), .a(n7272), .b(n7270_1), .c(n7268), .d(n7264) );
in01f01  g0544 ( .o(n7274), .a(n7273) );
no02f01  g0545 ( .o(n713), .a(n7274), .b(x1006) );
in01f01  g0546 ( .o(n7276), .a(net_375) );
no02f01  g0547 ( .o(n718), .a(n6966), .b(n7276) );
ao22f01  g0548 ( .o(n7278), .a(n6738), .b(_net_7558), .c(n6736_1), .d(_net_7622) );
ao22f01  g0549 ( .o(n7279), .a(n6739), .b(_net_7654), .c(n6734), .d(_net_7590) );
na02f01  g0550 ( .o(n727), .a(n7279), .b(n7278) );
in01f01  g0551 ( .o(n7281), .a(x1215) );
na04f01  g0552 ( .o(n7282), .a(x1231), .b(x1286), .c(x1261), .d(n7281) );
no02f01  g0553 ( .o(n7283), .a(x1231), .b(x1261) );
na04f01  g0554 ( .o(n7284_1), .a(n7283), .b(n6801_1), .c(x1215), .d(n6800) );
na04f01  g0555 ( .o(n7285), .a(n7284_1), .b(n7282), .c(x1286), .d(x1322) );
in01f01  g0556 ( .o(n7286), .a(n7285) );
na04f01  g0557 ( .o(n7287), .a(n7284_1), .b(n7282), .c(n6802), .d(n6800) );
in01f01  g0558 ( .o(n7288_1), .a(n7287) );
ao22f01  g0559 ( .o(n7289), .a(n7288_1), .b(_net_6041), .c(n7286), .d(_net_280) );
na04f01  g0560 ( .o(n7290), .a(n7284_1), .b(n7282), .c(x1261), .d(x1322) );
in01f01  g0561 ( .o(n7291), .a(n7290) );
na02f01  g0562 ( .o(n7292_1), .a(x1286), .b(x1261) );
no02f01  g0563 ( .o(n7293), .a(n7282), .b(n6800) );
in01f01  g0564 ( .o(n7294), .a(n7283) );
na03f01  g0565 ( .o(n7295), .a(n6801_1), .b(x1215), .c(n6800) );
no02f01  g0566 ( .o(n7296), .a(n7295), .b(n7294) );
no02f01  g0567 ( .o(n7297_1), .a(n7282), .b(x1322) );
no04f01  g0568 ( .o(n7298), .a(n7297_1), .b(n7296), .c(n7293), .d(n7292_1) );
ao22f01  g0569 ( .o(n7299), .a(n7298), .b(_net_7730), .c(n7291), .d(_net_7701) );
in01f01  g0570 ( .o(n7300), .a(x1261) );
na04f01  g0571 ( .o(n7301), .a(n7284_1), .b(n7282), .c(n6801_1), .d(n6800) );
no02f01  g0572 ( .o(n7302_1), .a(n7301), .b(n7300) );
na02f01  g0573 ( .o(n7303), .a(n7302_1), .b(_net_124) );
no02f01  g0574 ( .o(n7304), .a(x1286), .b(x1261) );
na04f01  g0575 ( .o(n7305), .a(n7304), .b(n7284_1), .c(n7282), .d(x1322) );
in01f01  g0576 ( .o(n7306), .a(n7305) );
na02f01  g0577 ( .o(n7307_1), .a(x1231), .b(n7281) );
no02f01  g0578 ( .o(n7308), .a(n7307_1), .b(n7292_1) );
na03f01  g0579 ( .o(n7309), .a(n7308), .b(net_203), .c(x1322) );
na02f01  g0580 ( .o(n7310), .a(n7296), .b(net_240) );
na03f01  g0581 ( .o(n7311), .a(n7308), .b(net_166), .c(n6800) );
na03f01  g0582 ( .o(n7312_1), .a(n7311), .b(n7310), .c(n7309) );
ao12f01  g0583 ( .o(n7313), .a(n7312_1), .b(n7306), .c(_net_5997) );
na04f01  g0584 ( .o(n732), .a(n7313), .b(n7303), .c(n7299), .d(n7289) );
in01f01  g0585 ( .o(n7315), .a(_net_6037) );
in01f01  g0586 ( .o(n7316_1), .a(_net_5976) );
oa12f01  g0587 ( .o(n736), .a(n7315), .b(n6978), .c(n7316_1) );
ao22f01  g0588 ( .o(n7318), .a(n6738), .b(_net_7557), .c(n6736_1), .d(_net_7621) );
ao22f01  g0589 ( .o(n7319), .a(n6739), .b(_net_7653), .c(n6734), .d(_net_7589) );
na02f01  g0590 ( .o(n746), .a(n7319), .b(n7318) );
ao22f01  g0591 ( .o(n7321_1), .a(n7000_1), .b(net_6967), .c(n6999), .d(net_7031) );
ao22f01  g0592 ( .o(n7322), .a(n7003), .b(net_6999), .c(n7002), .d(net_7063) );
na02f01  g0593 ( .o(n7323), .a(n7322), .b(n7321_1) );
na02f01  g0594 ( .o(n7324), .a(n7323), .b(n6981) );
ao22f01  g0595 ( .o(n7325), .a(n7000_1), .b(net_6965), .c(n6999), .d(net_7029) );
ao22f01  g0596 ( .o(n7326_1), .a(n7003), .b(net_6997), .c(n7002), .d(net_7061) );
na02f01  g0597 ( .o(n7327), .a(n7326_1), .b(n7325) );
ao22f01  g0598 ( .o(n7328), .a(n7327), .b(n6998), .c(n6996), .d(_net_6147) );
na02f01  g0599 ( .o(n756), .a(n7328), .b(n7324) );
in01f01  g0600 ( .o(n7330_1), .a(_net_7793) );
no02f01  g0601 ( .o(n7331), .a(x1286), .b(x1322) );
na03f01  g0602 ( .o(n7332), .a(n7331), .b(_net_6184), .c(n7300) );
no02f01  g0603 ( .o(n765), .a(n7332), .b(n7330_1) );
in01f01  g0604 ( .o(n7334), .a(_net_7732) );
in01f01  g0605 ( .o(n7335_1), .a(_net_6026) );
in01f01  g0606 ( .o(n7336), .a(n7108) );
in01f01  g0607 ( .o(n7337), .a(_net_7688) );
na03f01  g0608 ( .o(n7338), .a(_net_7687), .b(n7337), .c(n7105) );
no02f01  g0609 ( .o(n7339), .a(n7338), .b(n7336) );
in01f01  g0610 ( .o(n7340_1), .a(n7339) );
in01f01  g0611 ( .o(n7341), .a(x1231) );
na02f01  g0612 ( .o(n7342), .a(n7341), .b(n7281) );
no04f01  g0613 ( .o(n7343), .a(n7342), .b(n7340_1), .c(n7292_1), .d(x1322) );
ao12f01  g0614 ( .o(n770), .a(n7343), .b(n7335_1), .c(n7334) );
in01f01  g0615 ( .o(n7345), .a(_net_6012) );
in01f01  g0616 ( .o(n7346), .a(_net_6184) );
na02f01  g0617 ( .o(n7347), .a(n7304), .b(x1322) );
no02f01  g0618 ( .o(n7348), .a(n7347), .b(n7346) );
na02f01  g0619 ( .o(n7349_1), .a(n7348), .b(_net_7815) );
oa12f01  g0620 ( .o(n788), .a(n7349_1), .b(n7348), .c(n7345) );
in01f01  g0621 ( .o(n7351), .a(net_377) );
no02f01  g0622 ( .o(n793), .a(n6966), .b(n7351) );
in01f01  g0623 ( .o(n7353), .a(_net_113) );
no02f01  g0624 ( .o(n7354_1), .a(_net_7785), .b(_net_7786) );
in01f01  g0625 ( .o(n7355), .a(_net_7788) );
no02f01  g0626 ( .o(n7356), .a(n7355), .b(_net_7787) );
na04f01  g0627 ( .o(n7357), .a(n7356), .b(n7354_1), .c(_net_7789), .d(_net_7784) );
na02f01  g0628 ( .o(n7358), .a(n7357), .b(n7353) );
in01f01  g0629 ( .o(n7359_1), .a(_net_7786) );
na02f01  g0630 ( .o(n7360), .a(_net_7784), .b(_net_7785) );
no02f01  g0631 ( .o(n7361), .a(n7360), .b(n7359_1) );
in01f01  g0632 ( .o(n7362), .a(n7360) );
no02f01  g0633 ( .o(n7363_1), .a(n7362), .b(_net_7786) );
no03f01  g0634 ( .o(n806), .a(n7363_1), .b(n7361), .c(n7358) );
in01f01  g0635 ( .o(n7365), .a(_net_121) );
na02f01  g0636 ( .o(n7366), .a(net_317), .b(_net_154) );
oa12f01  g0637 ( .o(n820), .a(n7366), .b(_net_154), .c(n7365) );
in01f01  g0638 ( .o(n7368_1), .a(_net_120) );
na02f01  g0639 ( .o(n7369), .a(net_316), .b(_net_154) );
oa12f01  g0640 ( .o(n825), .a(n7369), .b(_net_154), .c(n7368_1) );
ao22f01  g0641 ( .o(n7371), .a(n7225), .b(_net_7428), .c(n7224), .d(net_7460) );
ao22f01  g0642 ( .o(n7372_1), .a(n7229), .b(net_7524), .c(n7228), .d(net_7492) );
na02f01  g0643 ( .o(n834), .a(n7372_1), .b(n7371) );
ao22f01  g0644 ( .o(n7374), .a(n6877), .b(_net_7265), .c(n6876_1), .d(_net_7329) );
ao22f01  g0645 ( .o(n7375), .a(n6881_1), .b(_net_7297), .c(n6880), .d(_net_7361) );
na02f01  g0646 ( .o(n849), .a(n7375), .b(n7374) );
na02f01  g0647 ( .o(n7377), .a(n6938_1), .b(n6917) );
ao22f01  g0648 ( .o(n7378), .a(n6942), .b(n6935), .c(n6933), .d(_net_6086) );
na02f01  g0649 ( .o(n862), .a(n7378), .b(n7377) );
no02f01  g0650 ( .o(n875), .a(n6899_1), .b(n7254) );
in01f01  g0651 ( .o(n7381_1), .a(_net_6008) );
na02f01  g0652 ( .o(n7382), .a(n7348), .b(_net_7811) );
oa12f01  g0653 ( .o(n885), .a(n7382), .b(n7348), .c(n7381_1) );
in01f01  g0654 ( .o(n7384), .a(_net_7439) );
na02f01  g0655 ( .o(n7385), .a(n6866), .b(net_7391) );
ao22f01  g0656 ( .o(n7386_1), .a(net_354), .b(_net_280), .c(_net_281), .d(net_352) );
na02f01  g0657 ( .o(n7387), .a(n7386_1), .b(n7385) );
na02f01  g0658 ( .o(n7388), .a(n7387), .b(n7197) );
oa12f01  g0659 ( .o(n903), .a(n7388), .b(n7197), .c(n7384) );
in01f01  g0660 ( .o(n7390), .a(_net_7354) );
na02f01  g0661 ( .o(n7391_1), .a(n6898), .b(net_7242) );
ao22f01  g0662 ( .o(n7392), .a(_net_269), .b(net_336), .c(_net_270), .d(net_334) );
na02f01  g0663 ( .o(n7393), .a(n7392), .b(n7391_1) );
na02f01  g0664 ( .o(n7394), .a(n7393), .b(n7030) );
oa12f01  g0665 ( .o(n925), .a(n7394), .b(n7030), .c(n7390) );
in01f01  g0666 ( .o(n7396), .a(_net_7632) );
in01f01  g0667 ( .o(n7397), .a(_net_7685) );
no02f01  g0668 ( .o(n7398), .a(n7397), .b(_net_7684) );
in01f01  g0669 ( .o(n7399), .a(n7398) );
no02f01  g0670 ( .o(n7400_1), .a(n7399), .b(n6967) );
na02f01  g0671 ( .o(n7401), .a(n6965), .b(net_370) );
ao22f01  g0672 ( .o(n7402), .a(net_384), .b(_net_291), .c(_net_292), .d(net_382) );
na02f01  g0673 ( .o(n7403), .a(n7402), .b(n7401) );
na02f01  g0674 ( .o(n7404_1), .a(n7403), .b(n7400_1) );
oa12f01  g0675 ( .o(n930), .a(n7404_1), .b(n7400_1), .c(n7396) );
in01f01  g0676 ( .o(n7406), .a(_net_5851) );
in01f01  g0677 ( .o(n7407), .a(x868) );
in01f01  g0678 ( .o(n7408_1), .a(_net_282) );
no02f01  g0679 ( .o(n7409), .a(_net_283), .b(n7408_1) );
in01f01  g0680 ( .o(n7410), .a(_net_226) );
na02f01  g0681 ( .o(n7411), .a(_net_278), .b(_net_284) );
ao12f01  g0682 ( .o(n7412), .a(n7411), .b(_net_229), .c(n7410) );
na02f01  g0683 ( .o(n7413_1), .a(n7412), .b(n7409) );
in01f01  g0684 ( .o(n7414), .a(n7411) );
in01f01  g0685 ( .o(n7415), .a(_net_283) );
no02f01  g0686 ( .o(n7416), .a(n7415), .b(n7408_1) );
na03f01  g0687 ( .o(n7417_1), .a(n7416), .b(n7414), .c(_net_226) );
na03f01  g0688 ( .o(n7418), .a(_net_228), .b(_net_229), .c(n7410) );
na04f01  g0689 ( .o(n7419), .a(n7418), .b(n7414), .c(n7415), .d(n7408_1) );
oa12f01  g0690 ( .o(n7420), .a(n7410), .b(_net_228), .c(_net_229) );
na04f01  g0691 ( .o(n7421), .a(n7420), .b(n7414), .c(_net_283), .d(n7408_1) );
na04f01  g0692 ( .o(n7422_1), .a(n7421), .b(n7419), .c(n7417_1), .d(n7413_1) );
na03f01  g0693 ( .o(n7423), .a(n7422_1), .b(net_7779), .c(n7407) );
oa12f01  g0694 ( .o(n944), .a(n7423), .b(n7406), .c(x868) );
in01f01  g0695 ( .o(n7425), .a(_net_7629) );
na02f01  g0696 ( .o(n7426), .a(n6965), .b(net_7549) );
ao22f01  g0697 ( .o(n7427_1), .a(_net_292), .b(net_379), .c(_net_291), .d(net_381) );
na02f01  g0698 ( .o(n7428), .a(n7427_1), .b(n7426) );
na02f01  g0699 ( .o(n7429), .a(n7428), .b(n7400_1) );
oa12f01  g0700 ( .o(n961), .a(n7429), .b(n7400_1), .c(n7425) );
ao22f01  g0701 ( .o(n7431), .a(n7225), .b(_net_7412), .c(n7224), .d(_net_7444) );
ao22f01  g0702 ( .o(n7432_1), .a(n7229), .b(_net_7508), .c(n7228), .d(_net_7476) );
na02f01  g0703 ( .o(n966), .a(n7432_1), .b(n7431) );
in01f01  g0704 ( .o(n7434), .a(_net_7296) );
na02f01  g0705 ( .o(n7435), .a(n6898), .b(net_7248) );
ao22f01  g0706 ( .o(n7436), .a(net_342), .b(_net_269), .c(net_340), .d(_net_270) );
na02f01  g0707 ( .o(n7437_1), .a(n7436), .b(n7435) );
na02f01  g0708 ( .o(n7438), .a(n7437_1), .b(n7180) );
oa12f01  g0709 ( .o(n971), .a(n7438), .b(n7180), .c(n7434) );
no04f01  g0710 ( .o(n7440), .a(n7346), .b(n6801_1), .c(x1261), .d(n6800) );
na02f01  g0711 ( .o(n7441), .a(n7440), .b(_net_7805) );
oa12f01  g0712 ( .o(n985), .a(n7441), .b(n7440), .c(n7408_1) );
in01f01  g0713 ( .o(n7443), .a(_net_7653) );
no02f01  g0714 ( .o(n7444), .a(n7397), .b(n6959) );
in01f01  g0715 ( .o(n7445), .a(n7444) );
no02f01  g0716 ( .o(n7446_1), .a(n7445), .b(n6967) );
na02f01  g0717 ( .o(n7447), .a(n6965), .b(net_7541) );
ao22f01  g0718 ( .o(n7448), .a(_net_292), .b(net_371), .c(_net_291), .d(net_373) );
na02f01  g0719 ( .o(n7449), .a(n7448), .b(n7447) );
na02f01  g0720 ( .o(n7450_1), .a(n7449), .b(n7446_1) );
oa12f01  g0721 ( .o(n990), .a(n7450_1), .b(n7446_1), .c(n7443) );
in01f01  g0722 ( .o(n7452), .a(_net_5856) );
in01f01  g0723 ( .o(n7453), .a(x1006) );
na03f01  g0724 ( .o(n7454_1), .a(n7273), .b(net_7774), .c(n7453) );
oa12f01  g0725 ( .o(n995), .a(n7454_1), .b(n7452), .c(x1006) );
in01f01  g0726 ( .o(n7456), .a(_net_7621) );
na02f01  g0727 ( .o(n7457), .a(n7449), .b(n7400_1) );
oa12f01  g0728 ( .o(n1010), .a(n7457), .b(n7400_1), .c(n7456) );
in01f01  g0729 ( .o(n7459_1), .a(net_6770) );
in01f01  g0730 ( .o(n7460), .a(net_6706) );
oa22f01  g0731 ( .o(n7461), .a(n7129), .b(n7460), .c(n7126), .d(n7459_1) );
in01f01  g0732 ( .o(n7462), .a(net_6802) );
in01f01  g0733 ( .o(n7463_1), .a(net_6738) );
oa22f01  g0734 ( .o(n7464), .a(n7134), .b(n7463_1), .c(n7132), .d(n7462) );
no02f01  g0735 ( .o(n7465), .a(n7464), .b(n7461) );
in01f01  g0736 ( .o(n7466), .a(_net_6822) );
no02f01  g0737 ( .o(n7467), .a(_net_6009), .b(_net_6008) );
na03f01  g0738 ( .o(n7468_1), .a(n7467), .b(n7122), .c(n7466) );
no02f01  g0739 ( .o(n7469), .a(n7468_1), .b(n7465) );
na02f01  g0740 ( .o(n7470), .a(n7122), .b(_net_6008) );
in01f01  g0741 ( .o(n7471), .a(net_6708) );
in01f01  g0742 ( .o(n7472), .a(net_6772) );
oa22f01  g0743 ( .o(n7473_1), .a(n7129), .b(n7471), .c(n7126), .d(n7472) );
in01f01  g0744 ( .o(n7474), .a(net_6804) );
in01f01  g0745 ( .o(n7475), .a(net_6740) );
oa22f01  g0746 ( .o(n7476), .a(n7134), .b(n7475), .c(n7132), .d(n7474) );
no02f01  g0747 ( .o(n7477), .a(n7476), .b(n7473_1) );
no02f01  g0748 ( .o(n7478_1), .a(n7477), .b(n7470) );
in01f01  g0749 ( .o(n7479), .a(_net_6120) );
in01f01  g0750 ( .o(n7480), .a(net_6774) );
in01f01  g0751 ( .o(n7481), .a(net_6710) );
oa22f01  g0752 ( .o(n7482_1), .a(n7129), .b(n7481), .c(n7126), .d(n7480) );
in01f01  g0753 ( .o(n7483), .a(net_6806) );
in01f01  g0754 ( .o(n7484), .a(net_6742) );
oa22f01  g0755 ( .o(n7485), .a(n7134), .b(n7484), .c(n7132), .d(n7483) );
no02f01  g0756 ( .o(n7486), .a(n7485), .b(n7482_1) );
oa22f01  g0757 ( .o(n7487_1), .a(n7486), .b(n7123), .c(n7118), .d(n7479) );
no03f01  g0758 ( .o(n7488), .a(n7487_1), .b(n7478_1), .c(n7469) );
in01f01  g0759 ( .o(n7489), .a(net_6754) );
in01f01  g0760 ( .o(n7490), .a(net_6722) );
na04f01  g0761 ( .o(n7491), .a(n7467), .b(n7135), .c(n7122), .d(_net_6822) );
na04f01  g0762 ( .o(n7492_1), .a(n7467), .b(n7130), .c(n7122), .d(_net_6822) );
oa22f01  g0763 ( .o(n7493), .a(n7492_1), .b(n7490), .c(n7491), .d(n7489) );
in01f01  g0764 ( .o(n7494), .a(net_6786) );
in01f01  g0765 ( .o(n7495), .a(net_6818) );
na04f01  g0766 ( .o(n7496_1), .a(n7467), .b(n7127), .c(n7122), .d(_net_6822) );
na04f01  g0767 ( .o(n7497), .a(n7467), .b(n7133_1), .c(n7122), .d(_net_6822) );
oa22f01  g0768 ( .o(n7498), .a(n7497), .b(n7495), .c(n7496_1), .d(n7494) );
no02f01  g0769 ( .o(n7499), .a(n7498), .b(n7493) );
na02f01  g0770 ( .o(n1015), .a(n7499), .b(n7488) );
in01f01  g0771 ( .o(n7501_1), .a(_net_7447) );
na02f01  g0772 ( .o(n7502), .a(n6866), .b(net_7399) );
ao22f01  g0773 ( .o(n7503), .a(_net_281), .b(net_360), .c(_net_280), .d(net_362) );
na02f01  g0774 ( .o(n7504), .a(n7503), .b(n7502) );
na02f01  g0775 ( .o(n7505_1), .a(n7504), .b(n7197) );
oa12f01  g0776 ( .o(n1024), .a(n7505_1), .b(n7197), .c(n7501_1) );
in01f01  g0777 ( .o(n7507), .a(net_334) );
no02f01  g0778 ( .o(n1029), .a(n6899_1), .b(n7507) );
in01f01  g0779 ( .o(n7509_1), .a(net_343) );
no02f01  g0780 ( .o(n1034), .a(n6899_1), .b(n7509_1) );
in01f01  g0781 ( .o(n7511), .a(_net_6259) );
no02f01  g0782 ( .o(n1039), .a(_net_392), .b(n7511) );
in01f01  g0783 ( .o(n7513_1), .a(_net_7281) );
in01f01  g0784 ( .o(n7514), .a(net_345) );
no02f01  g0785 ( .o(n6722), .a(n6899_1), .b(n7514) );
na02f01  g0786 ( .o(n7516), .a(n6722), .b(n6901) );
oa12f01  g0787 ( .o(n1044), .a(n7516), .b(n6901), .c(n7513_1) );
in01f01  g0788 ( .o(n7518_1), .a(_net_7578) );
no03f01  g0789 ( .o(n7519), .a(n6967), .b(_net_7685), .c(_net_7684) );
in01f01  g0790 ( .o(n7520), .a(net_380) );
no02f01  g0791 ( .o(n3546), .a(n6966), .b(n7520) );
na02f01  g0792 ( .o(n7522_1), .a(n3546), .b(n7519) );
oa12f01  g0793 ( .o(n1049), .a(n7522_1), .b(n7519), .c(n7518_1) );
ao22f01  g0794 ( .o(n7524), .a(n7288_1), .b(_net_6034), .c(n7286), .d(_net_273) );
ao22f01  g0795 ( .o(n7525), .a(n7298), .b(_net_7726), .c(n7291), .d(_net_7697) );
na02f01  g0796 ( .o(n7526), .a(n7302_1), .b(_net_120) );
na03f01  g0797 ( .o(n7527_1), .a(n7308), .b(net_199), .c(x1322) );
na02f01  g0798 ( .o(n7528), .a(n7296), .b(net_236) );
na03f01  g0799 ( .o(n7529), .a(n7308), .b(net_162), .c(n6800) );
na03f01  g0800 ( .o(n7530_1), .a(n7529), .b(n7528), .c(n7527_1) );
ao12f01  g0801 ( .o(n7531), .a(n7530_1), .b(n7306), .c(_net_5990) );
na04f01  g0802 ( .o(n1058), .a(n7531), .b(n7526), .c(n7525), .d(n7524) );
in01f01  g0803 ( .o(n7533), .a(_net_5960) );
oa12f01  g0804 ( .o(n7534), .a(n7533), .b(_net_5961), .c(_net_5962) );
in01f01  g0805 ( .o(n7535_1), .a(_net_5989) );
no03f01  g0806 ( .o(n7536), .a(n7535_1), .b(_net_5988), .c(n6759) );
no02f01  g0807 ( .o(n7537), .a(n6759), .b(n7533) );
in01f01  g0808 ( .o(n7538), .a(_net_5988) );
no02f01  g0809 ( .o(n7539_1), .a(n7535_1), .b(n7538) );
ao22f01  g0810 ( .o(n7540), .a(n7539_1), .b(n7537), .c(n7536), .d(n7534) );
no02f01  g0811 ( .o(n7541), .a(_net_5989), .b(n7538) );
ao12f01  g0812 ( .o(n7542), .a(n6759), .b(_net_5962), .c(n7533) );
na03f01  g0813 ( .o(n7543_1), .a(_net_5961), .b(_net_5962), .c(n7533) );
no03f01  g0814 ( .o(n7544), .a(_net_5989), .b(_net_5988), .c(n6759) );
ao22f01  g0815 ( .o(n7545), .a(n7544), .b(n7543_1), .c(n7542), .d(n7541) );
na02f01  g0816 ( .o(n1067), .a(n7545), .b(n7540) );
in01f01  g0817 ( .o(n7547), .a(_net_6285) );
no02f01  g0818 ( .o(n1072), .a(_net_392), .b(n7547) );
in01f01  g0819 ( .o(n7549), .a(_net_7412) );
no03f01  g0820 ( .o(n7550), .a(n6868), .b(_net_7533), .c(_net_7534) );
na02f01  g0821 ( .o(n7551), .a(n6866), .b(net_7396) );
ao22f01  g0822 ( .o(n7552), .a(net_359), .b(_net_280), .c(_net_281), .d(net_357) );
na02f01  g0823 ( .o(n7553_1), .a(n7552), .b(n7551) );
na02f01  g0824 ( .o(n7554), .a(n7553_1), .b(n7550) );
oa12f01  g0825 ( .o(n1106), .a(n7554), .b(n7550), .c(n7549) );
in01f01  g0826 ( .o(n7556), .a(net_7752) );
na04f01  g0827 ( .o(n7557), .a(_net_5995), .b(_net_7791), .c(n7556), .d(net_303) );
ao12f01  g0828 ( .o(n1116), .a(n7557), .b(net_308), .c(_net_5996) );
in01f01  g0829 ( .o(n7559), .a(_net_7274) );
in01f01  g0830 ( .o(n7560), .a(net_338) );
no02f01  g0831 ( .o(n4263), .a(n6899_1), .b(n7560) );
na02f01  g0832 ( .o(n7562), .a(n4263), .b(n6901) );
oa12f01  g0833 ( .o(n1125), .a(n7562), .b(n6901), .c(n7559) );
in01f01  g0834 ( .o(n7564), .a(_net_7299) );
na02f01  g0835 ( .o(n7565), .a(n6898), .b(net_331) );
ao22f01  g0836 ( .o(n7566), .a(_net_269), .b(net_345), .c(net_343), .d(_net_270) );
na02f01  g0837 ( .o(n7567_1), .a(n7566), .b(n7565) );
na02f01  g0838 ( .o(n7568), .a(n7567_1), .b(n7180) );
oa12f01  g0839 ( .o(n1135), .a(n7568), .b(n7180), .c(n7564) );
in01f01  g0840 ( .o(n7570), .a(_net_6039) );
in01f01  g0841 ( .o(n7571), .a(_net_7759) );
na03f01  g0842 ( .o(n7572_1), .a(net_6056), .b(_net_7791), .c(n7571) );
no02f01  g0843 ( .o(n7573), .a(n7572_1), .b(n7570) );
na02f01  g0844 ( .o(n7574), .a(n7573), .b(_net_6042) );
in01f01  g0845 ( .o(n7575), .a(n7574) );
in01f01  g0846 ( .o(n7576), .a(_net_7228) );
na02f01  g0847 ( .o(n7577_1), .a(n7576), .b(_net_7229) );
in01f01  g0848 ( .o(n7578), .a(n7577_1) );
in01f01  g0849 ( .o(n7579), .a(_net_7229) );
na02f01  g0850 ( .o(n7580), .a(n7576), .b(n7579) );
in01f01  g0851 ( .o(n7581_1), .a(n7580) );
ao22f01  g0852 ( .o(n7582), .a(n7581_1), .b(net_7102), .c(n7578), .d(net_7166) );
na02f01  g0853 ( .o(n7583), .a(_net_7228), .b(_net_7229) );
in01f01  g0854 ( .o(n7584), .a(n7583) );
na02f01  g0855 ( .o(n7585), .a(_net_7228), .b(n7579) );
in01f01  g0856 ( .o(n7586_1), .a(n7585) );
ao22f01  g0857 ( .o(n7587), .a(n7586_1), .b(net_7134), .c(n7584), .d(net_7198) );
na02f01  g0858 ( .o(n7588), .a(n7587), .b(n7582) );
na02f01  g0859 ( .o(n7589), .a(n7588), .b(n7575) );
na02f01  g0860 ( .o(n7590), .a(n7572_1), .b(_net_6039) );
in01f01  g0861 ( .o(n7591_1), .a(n7590) );
na02f01  g0862 ( .o(n7592), .a(n7573), .b(_net_6041) );
in01f01  g0863 ( .o(n7593), .a(n7592) );
ao22f01  g0864 ( .o(n7594), .a(n7581_1), .b(net_7100), .c(n7578), .d(net_7164) );
ao22f01  g0865 ( .o(n7595), .a(n7586_1), .b(net_7132), .c(n7584), .d(net_7196) );
na02f01  g0866 ( .o(n7596_1), .a(n7595), .b(n7594) );
ao22f01  g0867 ( .o(n7597), .a(n7596_1), .b(n7593), .c(n7591_1), .d(_net_6167) );
na02f01  g0868 ( .o(n1153), .a(n7597), .b(n7589) );
in01f01  g0869 ( .o(n7599_1), .a(net_381) );
no02f01  g0870 ( .o(n1163), .a(n6966), .b(n7599_1) );
in01f01  g0871 ( .o(n7601), .a(net_360) );
no02f01  g0872 ( .o(n1173), .a(n6867_1), .b(n7601) );
no02f01  g0873 ( .o(n7603), .a(n6833), .b(n6824) );
no02f01  g0874 ( .o(n7604_1), .a(n6843), .b(n6826_1) );
in01f01  g0875 ( .o(n7605), .a(_net_6135) );
in01f01  g0876 ( .o(n7606), .a(net_6904) );
in01f01  g0877 ( .o(n7607), .a(net_6840) );
oa22f01  g0878 ( .o(n7608_1), .a(n6810), .b(n7607), .c(n6807), .d(n7606) );
in01f01  g0879 ( .o(n7609), .a(net_6872) );
in01f01  g0880 ( .o(n7610), .a(net_6936) );
oa22f01  g0881 ( .o(n7611), .a(n6815), .b(n7609), .c(n6813_1), .d(n7610) );
no02f01  g0882 ( .o(n7612), .a(n7611), .b(n7608_1) );
oa22f01  g0883 ( .o(n7613_1), .a(n7612), .b(n6836_1), .c(n6844), .d(n7605) );
no03f01  g0884 ( .o(n7614), .a(n7613_1), .b(n7604_1), .c(n7603) );
in01f01  g0885 ( .o(n7615), .a(net_6852) );
in01f01  g0886 ( .o(n7616), .a(net_6884) );
oa22f01  g0887 ( .o(n7617), .a(n6850_1), .b(n7615), .c(n6849), .d(n7616) );
in01f01  g0888 ( .o(n7618_1), .a(net_6948) );
in01f01  g0889 ( .o(n7619), .a(net_6916) );
oa22f01  g0890 ( .o(n7620), .a(n6855_1), .b(n7618_1), .c(n6854), .d(n7619) );
no02f01  g0891 ( .o(n7621), .a(n7620), .b(n7617) );
na02f01  g0892 ( .o(n1178), .a(n7621), .b(n7614) );
in01f01  g0893 ( .o(n7623), .a(_net_7503) );
no02f01  g0894 ( .o(n7624), .a(n7194_1), .b(n6860_1) );
in01f01  g0895 ( .o(n7625), .a(n7624) );
no02f01  g0896 ( .o(n7626_1), .a(n7625), .b(n6868) );
na02f01  g0897 ( .o(n7627), .a(n7626_1), .b(n7387) );
oa12f01  g0898 ( .o(n1214), .a(n7627), .b(n7626_1), .c(n7623) );
in01f01  g0899 ( .o(n7629), .a(_net_7428) );
na02f01  g0900 ( .o(n7630), .a(n7550), .b(n595) );
oa12f01  g0901 ( .o(n1219), .a(n7630), .b(n7550), .c(n7629) );
in01f01  g0902 ( .o(n7632), .a(_net_7730) );
in01f01  g0903 ( .o(n7633), .a(_net_6016) );
ao12f01  g0904 ( .o(n1228), .a(n7343), .b(n7633), .c(n7632) );
in01f01  g0905 ( .o(n7635_1), .a(_net_7512) );
na02f01  g0906 ( .o(n7636), .a(n6866), .b(net_7400) );
ao22f01  g0907 ( .o(n7637), .a(_net_281), .b(net_361), .c(_net_280), .d(net_363) );
na02f01  g0908 ( .o(n7638), .a(n7637), .b(n7636) );
na02f01  g0909 ( .o(n7639), .a(n7638), .b(n7626_1) );
oa12f01  g0910 ( .o(n1253), .a(n7639), .b(n7626_1), .c(n7635_1) );
in01f01  g0911 ( .o(n7641), .a(_net_7590) );
na02f01  g0912 ( .o(n7642), .a(n6965), .b(net_7542) );
ao22f01  g0913 ( .o(n7643), .a(net_374), .b(_net_291), .c(_net_292), .d(net_372) );
na02f01  g0914 ( .o(n7644_1), .a(n7643), .b(n7642) );
na02f01  g0915 ( .o(n7645), .a(n7644_1), .b(n6968) );
oa12f01  g0916 ( .o(n1267), .a(n7645), .b(n6968), .c(n7641) );
in01f01  g0917 ( .o(n7647), .a(_net_273) );
na02f01  g0918 ( .o(n7648), .a(n7440), .b(net_7799) );
oa12f01  g0919 ( .o(n1272), .a(n7648), .b(n7440), .c(n7647) );
in01f01  g0920 ( .o(n7650), .a(net_354) );
no02f01  g0921 ( .o(n1277), .a(n6867_1), .b(n7650) );
in01f01  g0922 ( .o(n7652), .a(_net_299) );
in01f01  g0923 ( .o(n7653), .a(_net_263) );
in01f01  g0924 ( .o(n7654_1), .a(n6964_1) );
oa12f01  g0925 ( .o(n1282), .a(n7652), .b(n7654_1), .c(n7653) );
in01f01  g0926 ( .o(n7656), .a(_net_7315) );
na02f01  g0927 ( .o(n7657), .a(n6898), .b(net_7235) );
ao22f01  g0928 ( .o(n7658_1), .a(net_327), .b(_net_270), .c(_net_269), .d(net_329) );
na02f01  g0929 ( .o(n7659), .a(n7658_1), .b(n7657) );
na02f01  g0930 ( .o(n7660), .a(n7659), .b(n7150) );
oa12f01  g0931 ( .o(n1295), .a(n7660), .b(n7150), .c(n7656) );
no02f01  g0932 ( .o(n7662), .a(_net_6692), .b(n6921) );
in01f01  g0933 ( .o(n7663), .a(_net_6692) );
no02f01  g0934 ( .o(n7664), .a(n7663), .b(_net_6689) );
no02f01  g0935 ( .o(n7665), .a(n7664), .b(n7662) );
no02f01  g0936 ( .o(n7666_1), .a(n6918), .b(net_6691) );
no02f01  g0937 ( .o(n7667), .a(n7666_1), .b(n7665) );
no04f01  g0938 ( .o(n7668), .a(n7664), .b(n7662), .c(n6918), .d(net_6691) );
oa12f01  g0939 ( .o(n7669), .a(n7156), .b(n7668), .c(n7667) );
no02f01  g0940 ( .o(n7670), .a(n7668), .b(n7667) );
na02f01  g0941 ( .o(n7671_1), .a(n7670), .b(n548) );
na02f01  g0942 ( .o(n1309), .a(n7671_1), .b(n7669) );
in01f01  g0943 ( .o(n7673), .a(_net_6000) );
na02f01  g0944 ( .o(n7674), .a(n7348), .b(_net_7806) );
oa12f01  g0945 ( .o(n1314), .a(n7674), .b(n7348), .c(n7673) );
in01f01  g0946 ( .o(n7676_1), .a(_net_5991) );
na02f01  g0947 ( .o(n7677), .a(n7348), .b(_net_7800) );
oa12f01  g0948 ( .o(n1335), .a(n7677), .b(n7348), .c(n7676_1) );
in01f01  g0949 ( .o(n7679), .a(_net_7707) );
na02f01  g0950 ( .o(n7680), .a(n7207_1), .b(_net_7809) );
oa12f01  g0951 ( .o(n1340), .a(n7680), .b(n7207_1), .c(n7679) );
in01f01  g0952 ( .o(n7682), .a(_net_5975) );
no02f01  g0953 ( .o(n1345), .a(n6819), .b(n7682) );
ao22f01  g0954 ( .o(n7684), .a(n7225), .b(_net_7421), .c(n7224), .d(net_7453) );
ao22f01  g0955 ( .o(n7685), .a(n7229), .b(net_7517), .c(n7228), .d(net_7485) );
na02f01  g0956 ( .o(n1363), .a(n7685), .b(n7684) );
in01f01  g0957 ( .o(n7687), .a(_net_5972) );
oa12f01  g0958 ( .o(n7688), .a(n7687), .b(_net_5973), .c(_net_5974) );
in01f01  g0959 ( .o(n7689), .a(_net_6022) );
no03f01  g0960 ( .o(n7690), .a(n6819), .b(_net_6021), .c(n7689) );
no02f01  g0961 ( .o(n7691_1), .a(n6819), .b(n7687) );
in01f01  g0962 ( .o(n7692), .a(_net_6021) );
no02f01  g0963 ( .o(n7693), .a(n7692), .b(n7689) );
ao22f01  g0964 ( .o(n7694), .a(n7693), .b(n7691_1), .c(n7690), .d(n7688) );
no02f01  g0965 ( .o(n7695_1), .a(n7692), .b(_net_6022) );
ao12f01  g0966 ( .o(n7696), .a(n6819), .b(_net_5974), .c(n7687) );
na03f01  g0967 ( .o(n7697), .a(_net_5973), .b(_net_5974), .c(n7687) );
no03f01  g0968 ( .o(n7698), .a(n6819), .b(_net_6021), .c(_net_6022) );
ao22f01  g0969 ( .o(n7699), .a(n7698), .b(n7697), .c(n7696), .d(n7695_1) );
na02f01  g0970 ( .o(n1368), .a(n7699), .b(n7694) );
in01f01  g0971 ( .o(n7701), .a(_net_5997) );
na02f01  g0972 ( .o(n7702), .a(n7348), .b(_net_7803) );
oa12f01  g0973 ( .o(n1373), .a(n7702), .b(n7348), .c(n7701) );
in01f01  g0974 ( .o(n7704_1), .a(_net_7658) );
na02f01  g0975 ( .o(n7705), .a(n6965), .b(net_7546) );
ao22f01  g0976 ( .o(n7706), .a(_net_292), .b(net_376), .c(_net_291), .d(net_378) );
na02f01  g0977 ( .o(n7707), .a(n7706), .b(n7705) );
na02f01  g0978 ( .o(n7708), .a(n7707), .b(n7446_1) );
oa12f01  g0979 ( .o(n1391), .a(n7708), .b(n7446_1), .c(n7704_1) );
in01f01  g0980 ( .o(n7710), .a(_net_6189) );
no02f01  g0981 ( .o(n1396), .a(_net_392), .b(n7710) );
in01f01  g0982 ( .o(n7712), .a(net_7113) );
in01f01  g0983 ( .o(n7713), .a(net_7177) );
oa22f01  g0984 ( .o(n7714_1), .a(n7580), .b(n7712), .c(n7577_1), .d(n7713) );
in01f01  g0985 ( .o(n7715), .a(net_7145) );
in01f01  g0986 ( .o(n7716), .a(net_7209) );
oa22f01  g0987 ( .o(n7717), .a(n7585), .b(n7715), .c(n7583), .d(n7716) );
no02f01  g0988 ( .o(n7718), .a(n7717), .b(n7714_1) );
in01f01  g0989 ( .o(n7719_1), .a(_net_7227) );
no02f01  g0990 ( .o(n7720), .a(_net_6041), .b(_net_6042) );
na03f01  g0991 ( .o(n7721), .a(n7720), .b(n7573), .c(n7719_1) );
no02f01  g0992 ( .o(n7722), .a(n7721), .b(n7718) );
in01f01  g0993 ( .o(n7723_1), .a(net_7179) );
in01f01  g0994 ( .o(n7724), .a(net_7115) );
oa22f01  g0995 ( .o(n7725), .a(n7580), .b(n7724), .c(n7577_1), .d(n7723_1) );
in01f01  g0996 ( .o(n7726), .a(net_7147) );
in01f01  g0997 ( .o(n7727), .a(net_7211) );
oa22f01  g0998 ( .o(n7728_1), .a(n7585), .b(n7726), .c(n7583), .d(n7727) );
no02f01  g0999 ( .o(n7729), .a(n7728_1), .b(n7725) );
no02f01  g1000 ( .o(n7730), .a(n7729), .b(n7592) );
ao22f01  g1001 ( .o(n7731), .a(n7581_1), .b(net_7117), .c(n7578), .d(net_7181) );
ao22f01  g1002 ( .o(n7732_1), .a(n7586_1), .b(net_7149), .c(n7584), .d(net_7213) );
ao12f01  g1003 ( .o(n7733), .a(n7574), .b(n7732_1), .c(n7731) );
in01f01  g1004 ( .o(n7734), .a(_net_6182) );
no02f01  g1005 ( .o(n7735), .a(n7590), .b(n7734) );
no04f01  g1006 ( .o(n7736), .a(n7735), .b(n7733), .c(n7730), .d(n7722) );
in01f01  g1007 ( .o(n7737_1), .a(net_7129) );
in01f01  g1008 ( .o(n7738), .a(net_7161) );
na04f01  g1009 ( .o(n7739), .a(n7720), .b(n7586_1), .c(n7573), .d(_net_7227) );
na04f01  g1010 ( .o(n7740), .a(n7720), .b(n7581_1), .c(n7573), .d(_net_7227) );
oa22f01  g1011 ( .o(n7741_1), .a(n7740), .b(n7737_1), .c(n7739), .d(n7738) );
in01f01  g1012 ( .o(n7742), .a(net_7225) );
in01f01  g1013 ( .o(n7743), .a(net_7193) );
na04f01  g1014 ( .o(n7744), .a(n7720), .b(n7578), .c(n7573), .d(_net_7227) );
na04f01  g1015 ( .o(n7745), .a(n7720), .b(n7584), .c(n7573), .d(_net_7227) );
oa22f01  g1016 ( .o(n7746_1), .a(n7745), .b(n7742), .c(n7744), .d(n7743) );
no02f01  g1017 ( .o(n7747), .a(n7746_1), .b(n7741_1) );
na02f01  g1018 ( .o(n1405), .a(n7747), .b(n7736) );
in01f01  g1019 ( .o(n7749), .a(_net_6555) );
no02f01  g1020 ( .o(n7750), .a(n6758), .b(n6747) );
na03f01  g1021 ( .o(n7751_1), .a(n7750), .b(n7749), .c(_net_6554) );
in01f01  g1022 ( .o(n7752), .a(n7750) );
oa12f01  g1023 ( .o(n7753), .a(_net_6555), .b(n7752), .c(n6749_1) );
na02f01  g1024 ( .o(n7754), .a(n7753), .b(n7751_1) );
na02f01  g1025 ( .o(n7755), .a(n7754), .b(_net_6558) );
in01f01  g1026 ( .o(n7756_1), .a(_net_6558) );
na03f01  g1027 ( .o(n7757), .a(n7753), .b(n7751_1), .c(n7756_1) );
na02f01  g1028 ( .o(n7758), .a(n6758), .b(_net_6553) );
na02f01  g1029 ( .o(n7759), .a(_net_6552), .b(n6747) );
na02f01  g1030 ( .o(n7760_1), .a(n7759), .b(n7758) );
na02f01  g1031 ( .o(n7761), .a(n7760_1), .b(net_6556) );
in01f01  g1032 ( .o(n7762), .a(net_6556) );
na03f01  g1033 ( .o(n7763), .a(n7759), .b(n7758), .c(n7762) );
ao22f01  g1034 ( .o(n7764_1), .a(n7763), .b(n7761), .c(n6763), .d(_net_6552) );
in01f01  g1035 ( .o(n7765), .a(_net_6557) );
na02f01  g1036 ( .o(n7766), .a(n7750), .b(n6749_1) );
na02f01  g1037 ( .o(n7767), .a(n7752), .b(_net_6554) );
na02f01  g1038 ( .o(n7768_1), .a(n7767), .b(n7766) );
na02f01  g1039 ( .o(n7769), .a(n7768_1), .b(n7765) );
na03f01  g1040 ( .o(n7770), .a(n7767), .b(n7766), .c(_net_6557) );
na03f01  g1041 ( .o(n7771), .a(n7770), .b(n7769), .c(n7764_1) );
ao12f01  g1042 ( .o(n1410), .a(n7771), .b(n7757), .c(n7755) );
in01f01  g1043 ( .o(n7773_1), .a(_net_7253) );
na02f01  g1044 ( .o(n7774), .a(n7183), .b(n6901) );
oa12f01  g1045 ( .o(n1419), .a(n7774), .b(n6901), .c(n7773_1) );
in01f01  g1046 ( .o(n7776_1), .a(_net_7497) );
na02f01  g1047 ( .o(n7777), .a(n6866), .b(net_7385) );
ao22f01  g1048 ( .o(n7778), .a(net_348), .b(_net_280), .c(_net_281), .d(net_346) );
na02f01  g1049 ( .o(n7779_1), .a(n7778), .b(n7777) );
na02f01  g1050 ( .o(n7780), .a(n7779_1), .b(n7626_1) );
oa12f01  g1051 ( .o(n1428), .a(n7780), .b(n7626_1), .c(n7776_1) );
in01f01  g1052 ( .o(n7782), .a(n7331) );
no02f01  g1053 ( .o(n1433), .a(n7782), .b(n7206) );
in01f01  g1054 ( .o(n7784_1), .a(_net_7565) );
na02f01  g1055 ( .o(n7785), .a(n7519), .b(n7428) );
oa12f01  g1056 ( .o(n1442), .a(n7785), .b(n7519), .c(n7784_1) );
in01f01  g1057 ( .o(n7787), .a(_net_7806) );
na02f01  g1058 ( .o(n7788_1), .a(n6803), .b(_net_6044) );
oa12f01  g1059 ( .o(n1451), .a(n7788_1), .b(n6803), .c(n7787) );
in01f01  g1060 ( .o(n7790), .a(_net_7746) );
in01f01  g1061 ( .o(n7791), .a(net_297) );
ao12f01  g1062 ( .o(n1487), .a(n7343), .b(n7791), .c(n7790) );
in01f01  g1063 ( .o(n7793_1), .a(net_7754) );
na04f01  g1064 ( .o(n7794), .a(_net_7791), .b(_net_6006), .c(net_303), .d(n7793_1) );
ao12f01  g1065 ( .o(n1496), .a(n7794), .b(net_307), .c(_net_6007) );
in01f01  g1066 ( .o(n7796), .a(_net_7698) );
na02f01  g1067 ( .o(n7797), .a(n7207_1), .b(_net_7800) );
oa12f01  g1068 ( .o(n1501), .a(n7797), .b(n7207_1), .c(n7796) );
in01f01  g1069 ( .o(n7799), .a(net_6630) );
in01f01  g1070 ( .o(n7800), .a(net_6566) );
oa22f01  g1071 ( .o(n7801), .a(n6922), .b(n7800), .c(n6919_1), .d(n7799) );
in01f01  g1072 ( .o(n7802_1), .a(net_6598) );
in01f01  g1073 ( .o(n7803), .a(net_6662) );
oa22f01  g1074 ( .o(n7804), .a(n6927), .b(n7802_1), .c(n6925), .d(n7803) );
no02f01  g1075 ( .o(n7805), .a(n7804), .b(n7801) );
no02f01  g1076 ( .o(n7806_1), .a(n7805), .b(n6945) );
in01f01  g1077 ( .o(n7807), .a(net_6632) );
in01f01  g1078 ( .o(n7808), .a(net_6568) );
oa22f01  g1079 ( .o(n7809), .a(n6922), .b(n7808), .c(n6919_1), .d(n7807) );
in01f01  g1080 ( .o(n7810_1), .a(net_6664) );
in01f01  g1081 ( .o(n7811), .a(net_6600) );
oa22f01  g1082 ( .o(n7812), .a(n6927), .b(n7811), .c(n6925), .d(n7810_1) );
no02f01  g1083 ( .o(n7813), .a(n7812), .b(n7809) );
no02f01  g1084 ( .o(n7814), .a(n7813), .b(n6934_1) );
in01f01  g1085 ( .o(n7815_1), .a(_net_6095) );
in01f01  g1086 ( .o(n7816), .a(net_6570) );
in01f01  g1087 ( .o(n7817), .a(net_6634) );
oa22f01  g1088 ( .o(n7818_1), .a(n6922), .b(n7816), .c(n6919_1), .d(n7817) );
in01f01  g1089 ( .o(n7819), .a(net_6602) );
in01f01  g1090 ( .o(n7820), .a(net_6666) );
oa22f01  g1091 ( .o(n7821), .a(n6927), .b(n7819), .c(n6925), .d(n7820) );
no02f01  g1092 ( .o(n7822_1), .a(n7821), .b(n7818_1) );
oa22f01  g1093 ( .o(n7823), .a(n7822_1), .b(n6916), .c(n6932), .d(n7815_1) );
no03f01  g1094 ( .o(n7824), .a(n7823), .b(n7814), .c(n7806_1) );
in01f01  g1095 ( .o(n7825), .a(net_6614) );
in01f01  g1096 ( .o(n7826_1), .a(net_6582) );
oa22f01  g1097 ( .o(n7827), .a(n7058_1), .b(n7826_1), .c(n7057), .d(n7825) );
in01f01  g1098 ( .o(n7828), .a(net_6646) );
in01f01  g1099 ( .o(n7829), .a(net_6678) );
oa22f01  g1100 ( .o(n7830), .a(n7063), .b(n7829), .c(n7062_1), .d(n7828) );
no02f01  g1101 ( .o(n7831_1), .a(n7830), .b(n7827) );
na02f01  g1102 ( .o(n1519), .a(n7831_1), .b(n7824) );
ao22f01  g1103 ( .o(n7833), .a(n7225), .b(_net_7411), .c(n7224), .d(_net_7443) );
ao22f01  g1104 ( .o(n7834), .a(n7229), .b(_net_7507), .c(n7228), .d(_net_7475) );
na02f01  g1105 ( .o(n1533), .a(n7834), .b(n7833) );
na02f01  g1106 ( .o(n7836), .a(n7293), .b(net_216) );
na02f01  g1107 ( .o(n7837), .a(n7296), .b(net_253) );
na02f01  g1108 ( .o(n7838), .a(n7297_1), .b(net_179) );
na03f01  g1109 ( .o(n7839), .a(n7838), .b(n7837), .c(n7836) );
ao12f01  g1110 ( .o(n7840_1), .a(n7839), .b(n7291), .c(net_7714) );
na02f01  g1111 ( .o(n7841), .a(n7298), .b(net_7743) );
ao22f01  g1112 ( .o(n7842), .a(n7306), .b(net_6013), .c(n7286), .d(net_296) );
na03f01  g1113 ( .o(n1542), .a(n7842), .b(n7841), .c(n7840_1) );
na02f01  g1114 ( .o(n7844), .a(n6865), .b(_net_278) );
no02f01  g1115 ( .o(n7845_1), .a(n7844), .b(n6867_1) );
in01f01  g1116 ( .o(n7846), .a(_net_7532) );
oa12f01  g1117 ( .o(n7847), .a(n6860_1), .b(n7194_1), .c(n7846) );
na03f01  g1118 ( .o(n7848_1), .a(_net_7533), .b(_net_7532), .c(_net_7534) );
na03f01  g1119 ( .o(n7849), .a(n7848_1), .b(n7847), .c(n7845_1) );
in01f01  g1120 ( .o(n7850), .a(_net_278) );
in01f01  g1121 ( .o(n7851), .a(n6865) );
no03f01  g1122 ( .o(n7852), .a(n6866), .b(n7851), .c(n7850) );
na02f01  g1123 ( .o(n7853_1), .a(n7196), .b(n6862) );
no02f01  g1124 ( .o(n7854), .a(n6865), .b(n7850) );
ao22f01  g1125 ( .o(n7855), .a(n7854), .b(_net_7534), .c(n7853_1), .d(n7852) );
na02f01  g1126 ( .o(n1546), .a(n7855), .b(n7849) );
in01f01  g1127 ( .o(n7857), .a(_net_7406) );
na02f01  g1128 ( .o(n7858_1), .a(n6866), .b(net_7390) );
ao22f01  g1129 ( .o(n7859), .a(_net_281), .b(net_351), .c(_net_280), .d(net_353) );
na02f01  g1130 ( .o(n7860), .a(n7859), .b(n7858_1) );
na02f01  g1131 ( .o(n7861), .a(n7860), .b(n7550) );
oa12f01  g1132 ( .o(n1555), .a(n7861), .b(n7550), .c(n7857) );
ao22f01  g1133 ( .o(n7863_1), .a(n6736_1), .b(net_7644), .c(n6734), .d(net_7612) );
ao22f01  g1134 ( .o(n7864), .a(n6739), .b(net_7676), .c(n6738), .d(_net_7580) );
na02f01  g1135 ( .o(n1572), .a(n7864), .b(n7863_1) );
na02f01  g1136 ( .o(n7866), .a(n7624), .b(_net_7535) );
in01f01  g1137 ( .o(n7867_1), .a(_net_7535) );
na02f01  g1138 ( .o(n7868), .a(n7625), .b(n7867_1) );
na03f01  g1139 ( .o(n7869), .a(n7868), .b(n7866), .c(n7852) );
na02f01  g1140 ( .o(n7870), .a(n7848_1), .b(n7867_1) );
in01f01  g1141 ( .o(n7871_1), .a(n7848_1) );
na02f01  g1142 ( .o(n7872), .a(n7871_1), .b(_net_7535) );
na03f01  g1143 ( .o(n7873), .a(n7872), .b(n7870), .c(n7845_1) );
na02f01  g1144 ( .o(n7874), .a(n7854), .b(_net_7535) );
na03f01  g1145 ( .o(n1582), .a(n7874), .b(n7873), .c(n7869) );
no02f01  g1146 ( .o(n1600), .a(n7160_1), .b(n7232) );
ao22f01  g1147 ( .o(n7877), .a(n6877), .b(_net_7259), .c(n6876_1), .d(_net_7323) );
ao22f01  g1148 ( .o(n7878_1), .a(n6881_1), .b(_net_7291), .c(n6880), .d(_net_7355) );
na02f01  g1149 ( .o(n1605), .a(n7878_1), .b(n7877) );
in01f01  g1150 ( .o(n7880), .a(_net_7498) );
na02f01  g1151 ( .o(n7881), .a(n6866), .b(net_7386) );
ao22f01  g1152 ( .o(n7882), .a(_net_281), .b(net_347), .c(net_349), .d(_net_280) );
na02f01  g1153 ( .o(n7883_1), .a(n7882), .b(n7881) );
na02f01  g1154 ( .o(n7884), .a(n7883_1), .b(n7626_1) );
oa12f01  g1155 ( .o(n1610), .a(n7884), .b(n7626_1), .c(n7880) );
in01f01  g1156 ( .o(n7886), .a(_net_7696) );
na02f01  g1157 ( .o(n7887), .a(n7207_1), .b(_net_7798) );
oa12f01  g1158 ( .o(n1624), .a(n7887), .b(n7207_1), .c(n7886) );
in01f01  g1159 ( .o(n7889), .a(_net_7570) );
in01f01  g1160 ( .o(n7890), .a(net_372) );
in01f01  g1161 ( .o(n7891), .a(net_384) );
oa22f01  g1162 ( .o(n7892), .a(n6966), .b(n7890), .c(n7891), .d(n7143) );
na02f01  g1163 ( .o(n7893_1), .a(n7892), .b(n7519) );
oa12f01  g1164 ( .o(n1634), .a(n7893_1), .b(n7519), .c(n7889) );
in01f01  g1165 ( .o(n7895), .a(net_340) );
no02f01  g1166 ( .o(n1639), .a(n6899_1), .b(n7895) );
ao22f01  g1167 ( .o(n7897_1), .a(n6736_1), .b(net_7646), .c(n6734), .d(net_7614) );
ao22f01  g1168 ( .o(n7898), .a(n6739), .b(net_7678), .c(n6738), .d(_net_7582) );
na02f01  g1169 ( .o(n1644), .a(n7898), .b(n7897_1) );
ao22f01  g1170 ( .o(n7900), .a(n6736_1), .b(_net_7631), .c(n6734), .d(_net_7599) );
ao22f01  g1171 ( .o(n7901), .a(n6739), .b(_net_7663), .c(n6738), .d(_net_7567) );
na02f01  g1172 ( .o(n1658), .a(n7901), .b(n7900) );
in01f01  g1173 ( .o(n7903), .a(_net_7804) );
na02f01  g1174 ( .o(n7904), .a(n6803), .b(_net_6042) );
oa12f01  g1175 ( .o(n1677), .a(n7904), .b(n6803), .c(n7903) );
ao22f01  g1176 ( .o(n7906_1), .a(n7581_1), .b(net_7103), .c(n7578), .d(net_7167) );
ao22f01  g1177 ( .o(n7907), .a(n7586_1), .b(net_7135), .c(n7584), .d(net_7199) );
na02f01  g1178 ( .o(n7908), .a(n7907), .b(n7906_1) );
na02f01  g1179 ( .o(n7909), .a(n7908), .b(n7575) );
ao22f01  g1180 ( .o(n7910), .a(n7581_1), .b(net_7101), .c(n7578), .d(net_7165) );
ao22f01  g1181 ( .o(n7911_1), .a(n7586_1), .b(net_7133), .c(n7584), .d(net_7197) );
na02f01  g1182 ( .o(n7912), .a(n7911_1), .b(n7910) );
ao22f01  g1183 ( .o(n7913), .a(n7912), .b(n7593), .c(n7591_1), .d(_net_6168) );
in01f01  g1184 ( .o(n7914), .a(n7721) );
ao22f01  g1185 ( .o(n7915), .a(n7581_1), .b(net_7099), .c(n7578), .d(net_7163) );
ao22f01  g1186 ( .o(n7916_1), .a(n7586_1), .b(net_7131), .c(n7584), .d(net_7195) );
na02f01  g1187 ( .o(n7917), .a(n7916_1), .b(n7915) );
na02f01  g1188 ( .o(n7918), .a(n7917), .b(n7914) );
na02f01  g1189 ( .o(n7919), .a(n7720), .b(n7573) );
no02f01  g1190 ( .o(n7920_1), .a(n7919), .b(n7719_1) );
oa12f01  g1191 ( .o(n7921), .a(n7920_1), .b(n7728_1), .c(n7725) );
na04f01  g1192 ( .o(n1696), .a(n7921), .b(n7918), .c(n7913), .d(n7909) );
in01f01  g1193 ( .o(n7923), .a(_net_7358) );
na02f01  g1194 ( .o(n7924_1), .a(n6898), .b(net_7246) );
ao22f01  g1195 ( .o(n7925), .a(net_338), .b(_net_270), .c(net_340), .d(_net_269) );
na02f01  g1196 ( .o(n7926), .a(n7925), .b(n7924_1) );
na02f01  g1197 ( .o(n7927), .a(n7926), .b(n7030) );
oa12f01  g1198 ( .o(n1714), .a(n7927), .b(n7030), .c(n7923) );
in01f01  g1199 ( .o(n7929_1), .a(net_7111) );
in01f01  g1200 ( .o(n7930), .a(net_7175) );
oa22f01  g1201 ( .o(n7931), .a(n7580), .b(n7929_1), .c(n7577_1), .d(n7930) );
in01f01  g1202 ( .o(n7932), .a(net_7207) );
in01f01  g1203 ( .o(n7933_1), .a(net_7143) );
oa22f01  g1204 ( .o(n7934), .a(n7585), .b(n7933_1), .c(n7583), .d(n7932) );
no02f01  g1205 ( .o(n7935), .a(n7934), .b(n7931) );
no02f01  g1206 ( .o(n7936), .a(n7935), .b(n7721) );
no02f01  g1207 ( .o(n7937_1), .a(n7718), .b(n7592) );
in01f01  g1208 ( .o(n7938), .a(_net_6180) );
oa22f01  g1209 ( .o(n7939), .a(n7729), .b(n7574), .c(n7590), .d(n7938) );
no03f01  g1210 ( .o(n7940), .a(n7939), .b(n7937_1), .c(n7936) );
in01f01  g1211 ( .o(n7941), .a(net_7159) );
in01f01  g1212 ( .o(n7942_1), .a(net_7127) );
oa22f01  g1213 ( .o(n7943), .a(n7740), .b(n7942_1), .c(n7739), .d(n7941) );
in01f01  g1214 ( .o(n7944), .a(net_7223) );
in01f01  g1215 ( .o(n7945_1), .a(net_7191) );
oa22f01  g1216 ( .o(n7946), .a(n7745), .b(n7944), .c(n7744), .d(n7945_1) );
no02f01  g1217 ( .o(n7947), .a(n7946), .b(n7943) );
na02f01  g1218 ( .o(n1727), .a(n7947), .b(n7940) );
in01f01  g1219 ( .o(n7949), .a(_net_7468) );
na02f01  g1220 ( .o(n7950_1), .a(n6866), .b(net_7388) );
ao22f01  g1221 ( .o(n7951), .a(_net_281), .b(net_349), .c(_net_280), .d(net_351) );
na02f01  g1222 ( .o(n7952), .a(n7951), .b(n7950_1) );
na02f01  g1223 ( .o(n7953), .a(n7952), .b(n6869) );
oa12f01  g1224 ( .o(n1737), .a(n7953), .b(n6869), .c(n7949) );
in01f01  g1225 ( .o(n7955_1), .a(_net_5996) );
na02f01  g1226 ( .o(n7956), .a(n7348), .b(net_7802) );
oa12f01  g1227 ( .o(n1742), .a(n7956), .b(n7348), .c(n7955_1) );
in01f01  g1228 ( .o(n7958_1), .a(net_6433) );
in01f01  g1229 ( .o(n7959), .a(net_6497) );
oa22f01  g1230 ( .o(n7960), .a(n6750), .b(n7958_1), .c(n6748), .d(n7959) );
in01f01  g1231 ( .o(n7961), .a(net_6465) );
in01f01  g1232 ( .o(n7962_1), .a(net_6529) );
oa22f01  g1233 ( .o(n7963), .a(n6755), .b(n7961), .c(n6754), .d(n7962_1) );
no02f01  g1234 ( .o(n7964), .a(n7963), .b(n7960) );
no02f01  g1235 ( .o(n7965), .a(n7964), .b(n6764) );
no02f01  g1236 ( .o(n7966), .a(n7077_1), .b(n6766) );
in01f01  g1237 ( .o(n7967_1), .a(_net_6077) );
oa22f01  g1238 ( .o(n7968), .a(n7085_1), .b(n6775), .c(n6784), .d(n7967_1) );
no03f01  g1239 ( .o(n7969), .a(n7968), .b(n7966), .c(n7965) );
in01f01  g1240 ( .o(n7970_1), .a(net_6449) );
in01f01  g1241 ( .o(n7971), .a(net_6481) );
oa22f01  g1242 ( .o(n7972), .a(n6790), .b(n7970_1), .c(n6789), .d(n7971) );
in01f01  g1243 ( .o(n7973), .a(net_6545) );
in01f01  g1244 ( .o(n7974), .a(net_6513) );
oa22f01  g1245 ( .o(n7975_1), .a(n6795), .b(n7973), .c(n6794), .d(n7974) );
no02f01  g1246 ( .o(n7976), .a(n7975_1), .b(n7972) );
na02f01  g1247 ( .o(n1747), .a(n7976), .b(n7969) );
in01f01  g1248 ( .o(n7978), .a(net_364) );
no02f01  g1249 ( .o(n1752), .a(n6867_1), .b(n7978) );
in01f01  g1250 ( .o(n7980_1), .a(_net_5985) );
na02f01  g1251 ( .o(n7981), .a(n7348), .b(_net_7794) );
oa12f01  g1252 ( .o(n1770), .a(n7981), .b(n7348), .c(n7980_1) );
in01f01  g1253 ( .o(n7983), .a(_net_6295) );
no02f01  g1254 ( .o(n1787), .a(_net_392), .b(n7983) );
in01f01  g1255 ( .o(n1792), .a(n7343) );
in01f01  g1256 ( .o(n7986), .a(_net_6219) );
no02f01  g1257 ( .o(n1802), .a(n7986), .b(_net_392) );
in01f01  g1258 ( .o(n7988), .a(_net_7328) );
na02f01  g1259 ( .o(n7989_1), .a(n7437_1), .b(n7150) );
oa12f01  g1260 ( .o(n1807), .a(n7989_1), .b(n7150), .c(n7988) );
in01f01  g1261 ( .o(n7991), .a(_net_7359) );
na02f01  g1262 ( .o(n7992), .a(n6898), .b(net_7247) );
ao22f01  g1263 ( .o(n7993), .a(net_341), .b(_net_269), .c(_net_270), .d(net_339) );
na02f01  g1264 ( .o(n7994_1), .a(n7993), .b(n7992) );
na02f01  g1265 ( .o(n7995), .a(n7994_1), .b(n7030) );
oa12f01  g1266 ( .o(n1812), .a(n7995), .b(n7030), .c(n7991) );
in01f01  g1267 ( .o(n7997_1), .a(_net_7650) );
na02f01  g1268 ( .o(n7998), .a(n6965), .b(net_7538) );
ao22f01  g1269 ( .o(n7999), .a(net_368), .b(_net_292), .c(net_370), .d(_net_291) );
na02f01  g1270 ( .o(n8000), .a(n7999), .b(n7998) );
na02f01  g1271 ( .o(n8001), .a(n8000), .b(n7446_1) );
oa12f01  g1272 ( .o(n1832), .a(n8001), .b(n7446_1), .c(n7997_1) );
ao22f01  g1273 ( .o(n8003), .a(n6923), .b(net_6562), .c(n6920), .d(net_6626) );
ao22f01  g1274 ( .o(n8004), .a(n6928), .b(net_6594), .c(n6926), .d(net_6658) );
na02f01  g1275 ( .o(n8005_1), .a(n8004), .b(n8003) );
na02f01  g1276 ( .o(n8006), .a(n8005_1), .b(n6917) );
ao22f01  g1277 ( .o(n8007), .a(n6923), .b(net_6560), .c(n6920), .d(net_6624) );
ao22f01  g1278 ( .o(n8008), .a(n6928), .b(net_6592), .c(n6926), .d(net_6656) );
na02f01  g1279 ( .o(n8009), .a(n8008), .b(n8007) );
ao22f01  g1280 ( .o(n8010_1), .a(n8009), .b(n6935), .c(n6933), .d(_net_6087) );
na02f01  g1281 ( .o(n1841), .a(n8010_1), .b(n8006) );
in01f01  g1282 ( .o(n8012), .a(_net_6291) );
no02f01  g1283 ( .o(n1846), .a(_net_392), .b(n8012) );
in01f01  g1284 ( .o(n8014), .a(_net_6222) );
no02f01  g1285 ( .o(n1851), .a(_net_392), .b(n8014) );
in01f01  g1286 ( .o(n8016), .a(_net_7768) );
in01f01  g1287 ( .o(n8017), .a(net_153) );
no02f01  g1288 ( .o(n1860), .a(n8017), .b(n8016) );
in01f01  g1289 ( .o(n8019_1), .a(_net_7255) );
na02f01  g1290 ( .o(n8020), .a(n6898), .b(net_7239) );
ao22f01  g1291 ( .o(n8021), .a(net_333), .b(_net_269), .c(_net_270), .d(net_331) );
na02f01  g1292 ( .o(n8022), .a(n8021), .b(n8020) );
na02f01  g1293 ( .o(n8023), .a(n8022), .b(n6901) );
oa12f01  g1294 ( .o(n1869), .a(n8023), .b(n6901), .c(n8019_1) );
in01f01  g1295 ( .o(n8025), .a(_net_7600) );
na02f01  g1296 ( .o(n8026), .a(n7403), .b(n6968) );
oa12f01  g1297 ( .o(n1878), .a(n8026), .b(n6968), .c(n8025) );
in01f01  g1298 ( .o(n8028_1), .a(n6775) );
ao22f01  g1299 ( .o(n8029), .a(n6777), .b(net_6427), .c(n6776), .d(net_6491) );
ao22f01  g1300 ( .o(n8030), .a(n6780), .b(net_6459), .c(n6779_1), .d(net_6523) );
na02f01  g1301 ( .o(n8031), .a(n8030), .b(n8029) );
na02f01  g1302 ( .o(n8032), .a(n8031), .b(n8028_1) );
in01f01  g1303 ( .o(n8033_1), .a(n6766) );
in01f01  g1304 ( .o(n8034), .a(n6784) );
ao22f01  g1305 ( .o(n8035), .a(n6777), .b(net_6425), .c(n6776), .d(net_6489) );
ao22f01  g1306 ( .o(n8036), .a(n6780), .b(net_6457), .c(n6779_1), .d(net_6521) );
na02f01  g1307 ( .o(n8037), .a(n8036), .b(n8035) );
ao22f01  g1308 ( .o(n8038_1), .a(n8037), .b(n8033_1), .c(n8034), .d(_net_6067) );
na02f01  g1309 ( .o(n1883), .a(n8038_1), .b(n8032) );
in01f01  g1310 ( .o(n8040), .a(_net_7628) );
na02f01  g1311 ( .o(n8041), .a(n6965), .b(net_7548) );
ao22f01  g1312 ( .o(n8042_1), .a(_net_292), .b(net_378), .c(_net_291), .d(net_380) );
na02f01  g1313 ( .o(n8043), .a(n8042_1), .b(n8041) );
na02f01  g1314 ( .o(n8044), .a(n8043), .b(n7400_1) );
oa12f01  g1315 ( .o(n1888), .a(n8044), .b(n7400_1), .c(n8040) );
in01f01  g1316 ( .o(n8046), .a(net_7035) );
in01f01  g1317 ( .o(n8047_1), .a(net_6971) );
oa22f01  g1318 ( .o(n8048), .a(n6987), .b(n8047_1), .c(n6985), .d(n8046) );
in01f01  g1319 ( .o(n8049), .a(net_7067) );
in01f01  g1320 ( .o(n8050), .a(net_7003) );
oa22f01  g1321 ( .o(n8051_1), .a(n6992), .b(n8050), .c(n6991), .d(n8049) );
no02f01  g1322 ( .o(n8052), .a(n8051_1), .b(n8048) );
no02f01  g1323 ( .o(n8053), .a(n8052), .b(n7012) );
in01f01  g1324 ( .o(n8054), .a(net_7037) );
in01f01  g1325 ( .o(n8055), .a(net_6973) );
oa22f01  g1326 ( .o(n8056_1), .a(n6987), .b(n8055), .c(n6985), .d(n8054) );
in01f01  g1327 ( .o(n8057), .a(net_7069) );
in01f01  g1328 ( .o(n8058), .a(net_7005) );
oa22f01  g1329 ( .o(n8059_1), .a(n6992), .b(n8058), .c(n6991), .d(n8057) );
no02f01  g1330 ( .o(n8060), .a(n8059_1), .b(n8056_1) );
no02f01  g1331 ( .o(n8061), .a(n8060), .b(n6997) );
in01f01  g1332 ( .o(n8062), .a(_net_6155) );
in01f01  g1333 ( .o(n8063), .a(net_6975) );
in01f01  g1334 ( .o(n8064_1), .a(net_7039) );
oa22f01  g1335 ( .o(n8065), .a(n6987), .b(n8063), .c(n6985), .d(n8064_1) );
in01f01  g1336 ( .o(n8066), .a(net_7007) );
in01f01  g1337 ( .o(n8067_1), .a(net_7071) );
oa22f01  g1338 ( .o(n8068), .a(n6992), .b(n8066), .c(n6991), .d(n8067_1) );
no02f01  g1339 ( .o(n8069), .a(n8068), .b(n8065) );
oa22f01  g1340 ( .o(n8070), .a(n8069), .b(n6980), .c(n6995_1), .d(n8062) );
no03f01  g1341 ( .o(n8071), .a(n8070), .b(n8061), .c(n8053) );
in01f01  g1342 ( .o(n8072_1), .a(net_7019) );
in01f01  g1343 ( .o(n8073), .a(net_6987) );
na04f01  g1344 ( .o(n8074), .a(n7011), .b(n7003), .c(n6979), .d(_net_7092) );
na04f01  g1345 ( .o(n8075_1), .a(n7011), .b(n7000_1), .c(n6979), .d(_net_7092) );
oa22f01  g1346 ( .o(n8076), .a(n8075_1), .b(n8073), .c(n8074), .d(n8072_1) );
in01f01  g1347 ( .o(n8077), .a(net_7083) );
in01f01  g1348 ( .o(n8078), .a(net_7051) );
na04f01  g1349 ( .o(n8079), .a(n7011), .b(n6999), .c(n6979), .d(_net_7092) );
na04f01  g1350 ( .o(n8080_1), .a(n7011), .b(n7002), .c(n6979), .d(_net_7092) );
oa22f01  g1351 ( .o(n8081), .a(n8080_1), .b(n8077), .c(n8079), .d(n8078) );
no02f01  g1352 ( .o(n8082), .a(n8081), .b(n8076) );
na02f01  g1353 ( .o(n1893), .a(n8082), .b(n8071) );
in01f01  g1354 ( .o(n8084), .a(_net_6411) );
na04f01  g1355 ( .o(n8085_1), .a(_net_6407), .b(_net_6410), .c(_net_6406), .d(n8084) );
no02f01  g1356 ( .o(n8086), .a(_net_6409), .b(_net_6408) );
in01f01  g1357 ( .o(n8087), .a(n8086) );
in01f01  g1358 ( .o(n8088_1), .a(_net_6404) );
no02f01  g1359 ( .o(n8089), .a(_net_6405), .b(n8088_1) );
in01f01  g1360 ( .o(n8090), .a(n8089) );
no03f01  g1361 ( .o(n1898), .a(n8090), .b(n8087), .c(n8085_1) );
no02f01  g1362 ( .o(n8092_1), .a(n6881_1), .b(n6876_1) );
in01f01  g1363 ( .o(n8093), .a(_net_190) );
in01f01  g1364 ( .o(n8094), .a(_net_267) );
no02f01  g1365 ( .o(n3638), .a(n8094), .b(n8093) );
in01f01  g1366 ( .o(n8096), .a(n3638) );
na02f01  g1367 ( .o(n8097_1), .a(_net_267), .b(n8093) );
oa22f01  g1368 ( .o(n1908), .a(n8097_1), .b(n6875), .c(n8096), .d(n8092_1) );
in01f01  g1369 ( .o(n8099), .a(net_6430) );
in01f01  g1370 ( .o(n8100), .a(net_6494) );
oa22f01  g1371 ( .o(n8101), .a(n6750), .b(n8099), .c(n6748), .d(n8100) );
in01f01  g1372 ( .o(n8102_1), .a(net_6462) );
in01f01  g1373 ( .o(n8103), .a(net_6526) );
oa22f01  g1374 ( .o(n8104), .a(n6755), .b(n8102_1), .c(n6754), .d(n8103) );
oa12f01  g1375 ( .o(n8105), .a(n8028_1), .b(n8104), .c(n8101) );
ao22f01  g1376 ( .o(n8106), .a(n6777), .b(net_6428), .c(n6776), .d(net_6492) );
ao22f01  g1377 ( .o(n8107_1), .a(n6780), .b(net_6460), .c(n6779_1), .d(net_6524) );
na02f01  g1378 ( .o(n8108), .a(n8107_1), .b(n8106) );
ao22f01  g1379 ( .o(n8109), .a(n8108), .b(n8033_1), .c(n8034), .d(_net_6070) );
in01f01  g1380 ( .o(n8110), .a(n6764) );
na02f01  g1381 ( .o(n8111), .a(n6781), .b(n6778) );
na02f01  g1382 ( .o(n8112_1), .a(n6763), .b(n6762) );
no02f01  g1383 ( .o(n8113), .a(n8112_1), .b(n6758) );
ao22f01  g1384 ( .o(n8114), .a(n6777), .b(net_6426), .c(n6776), .d(net_6490) );
ao22f01  g1385 ( .o(n8115), .a(n6780), .b(net_6458), .c(n6779_1), .d(net_6522) );
na02f01  g1386 ( .o(n8116_1), .a(n8115), .b(n8114) );
ao22f01  g1387 ( .o(n8117), .a(n8116_1), .b(n8110), .c(n8113), .d(n8111) );
na03f01  g1388 ( .o(n1922), .a(n8117), .b(n8109), .c(n8105) );
in01f01  g1389 ( .o(n8119), .a(_net_6690) );
no02f01  g1390 ( .o(n8120), .a(n6943_1), .b(n6918) );
na03f01  g1391 ( .o(n8121_1), .a(n8120), .b(_net_6689), .c(n8119) );
in01f01  g1392 ( .o(n8122), .a(n8120) );
oa12f01  g1393 ( .o(n8123), .a(_net_6690), .b(n8122), .c(n6921) );
na02f01  g1394 ( .o(n8124), .a(n8123), .b(n8121_1) );
no04f01  g1395 ( .o(n8125_1), .a(n6914), .b(n6912), .c(_net_5998), .d(_net_5997) );
na02f01  g1396 ( .o(n8126), .a(n8125_1), .b(n8124) );
no03f01  g1397 ( .o(n8127), .a(n6944), .b(n6914), .c(n6912) );
no02f01  g1398 ( .o(n8128), .a(n6925), .b(n8119) );
no02f01  g1399 ( .o(n8129), .a(n6926), .b(_net_6690) );
no02f01  g1400 ( .o(n8130_1), .a(n8129), .b(n8128) );
in01f01  g1401 ( .o(n8131), .a(n6914) );
no02f01  g1402 ( .o(n8132), .a(n8131), .b(n6912) );
ao22f01  g1403 ( .o(n8133), .a(n8132), .b(_net_6690), .c(n8130_1), .d(n8127) );
na02f01  g1404 ( .o(n1927), .a(n8133), .b(n8126) );
ao22f01  g1405 ( .o(n8135_1), .a(n6736_1), .b(_net_7627), .c(n6734), .d(_net_7595) );
ao22f01  g1406 ( .o(n8136), .a(n6739), .b(_net_7659), .c(n6738), .d(_net_7563) );
na02f01  g1407 ( .o(n1936), .a(n8136), .b(n8135_1) );
in01f01  g1408 ( .o(n8138), .a(_net_7472) );
na02f01  g1409 ( .o(n8139), .a(n6866), .b(net_7392) );
ao22f01  g1410 ( .o(n8140_1), .a(_net_281), .b(net_353), .c(net_355), .d(_net_280) );
na02f01  g1411 ( .o(n8141), .a(n8140_1), .b(n8139) );
na02f01  g1412 ( .o(n8142), .a(n8141), .b(n6869) );
oa12f01  g1413 ( .o(n1945), .a(n8142), .b(n6869), .c(n8138) );
in01f01  g1414 ( .o(n8144_1), .a(n7854) );
na02f01  g1415 ( .o(n8145), .a(n6867_1), .b(n7846) );
na02f01  g1416 ( .o(n8146), .a(n6866), .b(_net_7532) );
na02f01  g1417 ( .o(n8147_1), .a(n8146), .b(n8145) );
oa22f01  g1418 ( .o(n1950), .a(n8147_1), .b(n7844), .c(n8144_1), .d(n7846) );
in01f01  g1419 ( .o(n8149), .a(_net_129) );
na02f01  g1420 ( .o(n8150), .a(_net_154), .b(net_325) );
oa12f01  g1421 ( .o(n1959), .a(n8150), .b(_net_154), .c(n8149) );
in01f01  g1422 ( .o(n8152_1), .a(_net_7594) );
na02f01  g1423 ( .o(n8153), .a(n7707), .b(n6968) );
oa12f01  g1424 ( .o(n1969), .a(n8153), .b(n6968), .c(n8152_1) );
ao22f01  g1425 ( .o(n8155), .a(n7130), .b(net_6698), .c(n7127), .d(net_6762) );
ao22f01  g1426 ( .o(n8156_1), .a(n7135), .b(net_6730), .c(n7133_1), .d(net_6794) );
na02f01  g1427 ( .o(n8157), .a(n8156_1), .b(n8155) );
na02f01  g1428 ( .o(n8158), .a(n8157), .b(n7124) );
in01f01  g1429 ( .o(n8159), .a(n7470) );
ao22f01  g1430 ( .o(n8160), .a(n7130), .b(net_6696), .c(n7127), .d(net_6760) );
ao22f01  g1431 ( .o(n8161_1), .a(n7135), .b(net_6728), .c(n7133_1), .d(net_6792) );
na02f01  g1432 ( .o(n8162), .a(n8161_1), .b(n8160) );
ao22f01  g1433 ( .o(n8163), .a(n8162), .b(n8159), .c(n7119), .d(_net_6108) );
in01f01  g1434 ( .o(n8164), .a(n7468_1) );
na02f01  g1435 ( .o(n8165), .a(n8164), .b(n7137) );
na02f01  g1436 ( .o(n8166_1), .a(n7467), .b(n7122) );
no02f01  g1437 ( .o(n8167), .a(n8166_1), .b(n7466) );
oa12f01  g1438 ( .o(n8168), .a(n8167), .b(n7485), .c(n7482_1) );
na04f01  g1439 ( .o(n1988), .a(n8168), .b(n8165), .c(n8163), .d(n8158) );
in01f01  g1440 ( .o(n8170_1), .a(net_357) );
no02f01  g1441 ( .o(n1993), .a(n6867_1), .b(n8170_1) );
in01f01  g1442 ( .o(n8172), .a(_net_7426) );
in01f01  g1443 ( .o(n8173), .a(net_359) );
no02f01  g1444 ( .o(n2256), .a(n6867_1), .b(n8173) );
na02f01  g1445 ( .o(n8175), .a(n2256), .b(n7550) );
oa12f01  g1446 ( .o(n2016), .a(n8175), .b(n7550), .c(n8172) );
no02f01  g1447 ( .o(n8177), .a(_net_6410), .b(_net_6411) );
na02f01  g1448 ( .o(n8178), .a(_net_6409), .b(_net_6408) );
oa12f01  g1449 ( .o(n8179_1), .a(_net_6407), .b(_net_6405), .c(_net_6406) );
oa12f01  g1450 ( .o(n2021), .a(n8177), .b(n8179_1), .c(n8178) );
ao22f01  g1451 ( .o(n8181), .a(n7130), .b(net_6697), .c(n7127), .d(net_6761) );
ao22f01  g1452 ( .o(n8182), .a(n7135), .b(net_6729), .c(n7133_1), .d(net_6793) );
na02f01  g1453 ( .o(n8183_1), .a(n8182), .b(n8181) );
na02f01  g1454 ( .o(n8184), .a(n8183_1), .b(n7124) );
ao22f01  g1455 ( .o(n8185), .a(n7130), .b(net_6695), .c(n7127), .d(net_6759) );
ao22f01  g1456 ( .o(n8186), .a(n7135), .b(net_6727), .c(n7133_1), .d(net_6791) );
na02f01  g1457 ( .o(n8187), .a(n8186), .b(n8185) );
ao22f01  g1458 ( .o(n8188_1), .a(n8187), .b(n8159), .c(n7119), .d(_net_6107) );
na02f01  g1459 ( .o(n2026), .a(n8188_1), .b(n8184) );
in01f01  g1460 ( .o(n8190), .a(_net_7483) );
in01f01  g1461 ( .o(n8191), .a(net_352) );
in01f01  g1462 ( .o(n8192_1), .a(_net_281) );
oa22f01  g1463 ( .o(n8193), .a(n6867_1), .b(n8191), .c(n8192_1), .d(n7978) );
na02f01  g1464 ( .o(n8194), .a(n8193), .b(n6869) );
oa12f01  g1465 ( .o(n2041), .a(n8194), .b(n6869), .c(n8190) );
na02f01  g1466 ( .o(n8196), .a(n7218), .b(n6984) );
na02f01  g1467 ( .o(n8197_1), .a(n7010), .b(_net_7093) );
na02f01  g1468 ( .o(n8198), .a(_net_7092), .b(n6984) );
na02f01  g1469 ( .o(n8199), .a(n8198), .b(n8197_1) );
ao22f01  g1470 ( .o(n8200), .a(n8199), .b(n7215), .c(n7220), .d(_net_7093) );
na02f01  g1471 ( .o(n2046), .a(n8200), .b(n8196) );
in01f01  g1472 ( .o(n8202_1), .a(_net_7465) );
na02f01  g1473 ( .o(n8203), .a(n7779_1), .b(n6869) );
oa12f01  g1474 ( .o(n2055), .a(n8203), .b(n6869), .c(n8202_1) );
in01f01  g1475 ( .o(n8205), .a(_net_7352) );
na02f01  g1476 ( .o(n8206_1), .a(n6898), .b(net_7240) );
ao22f01  g1477 ( .o(n8207), .a(net_332), .b(_net_270), .c(_net_269), .d(net_334) );
na02f01  g1478 ( .o(n8208), .a(n8207), .b(n8206_1) );
na02f01  g1479 ( .o(n8209), .a(n8208), .b(n7030) );
oa12f01  g1480 ( .o(n2060), .a(n8209), .b(n7030), .c(n8205) );
in01f01  g1481 ( .o(n8211_1), .a(n6844) );
na02f01  g1482 ( .o(n8212), .a(n8211_1), .b(_net_6125) );
in01f01  g1483 ( .o(n8213), .a(n6836_1) );
ao22f01  g1484 ( .o(n8214), .a(n6811), .b(net_6830), .c(n6808), .d(net_6894) );
ao22f01  g1485 ( .o(n8215), .a(n6816), .b(net_6862), .c(n6814), .d(net_6926) );
na02f01  g1486 ( .o(n8216_1), .a(n8215), .b(n8214) );
na02f01  g1487 ( .o(n8217), .a(n8216_1), .b(n8213) );
na02f01  g1488 ( .o(n2065), .a(n8217), .b(n8212) );
in01f01  g1489 ( .o(n8219), .a(_net_6827) );
in01f01  g1490 ( .o(n8220_1), .a(net_6826) );
no02f01  g1491 ( .o(n8221), .a(n8220_1), .b(_net_6827) );
no02f01  g1492 ( .o(n8222), .a(net_6826), .b(n8219) );
no02f01  g1493 ( .o(n8223), .a(n8222), .b(n8221) );
in01f01  g1494 ( .o(n8224_1), .a(_net_5971) );
no02f01  g1495 ( .o(n6427), .a(n8224_1), .b(n7121) );
in01f01  g1496 ( .o(n8226), .a(n6427) );
na02f01  g1497 ( .o(n8227), .a(n8224_1), .b(_net_6006) );
oa22f01  g1498 ( .o(n2070), .a(n8227), .b(n8219), .c(n8226), .d(n8223) );
in01f01  g1499 ( .o(n8229), .a(net_339) );
no02f01  g1500 ( .o(n2084), .a(n6899_1), .b(n8229) );
in01f01  g1501 ( .o(n8231), .a(_net_7683) );
na02f01  g1502 ( .o(n8232_1), .a(n6964_1), .b(_net_289) );
na02f01  g1503 ( .o(n8233), .a(n6966), .b(n8231) );
na02f01  g1504 ( .o(n8234), .a(n6965), .b(_net_7683) );
na02f01  g1505 ( .o(n8235), .a(n8234), .b(n8233) );
in01f01  g1506 ( .o(n8236), .a(_net_289) );
no02f01  g1507 ( .o(n8237_1), .a(n6964_1), .b(n8236) );
in01f01  g1508 ( .o(n8238), .a(n8237_1) );
oa22f01  g1509 ( .o(n2140), .a(n8238), .b(n8231), .c(n8235), .d(n8232_1) );
in01f01  g1510 ( .o(n8240), .a(_net_7554) );
na02f01  g1511 ( .o(n8241_1), .a(n8000), .b(n7519) );
oa12f01  g1512 ( .o(n2162), .a(n8241_1), .b(n7519), .c(n8240) );
in01f01  g1513 ( .o(n8243), .a(_net_7649) );
na02f01  g1514 ( .o(n8244), .a(n6965), .b(net_7537) );
ao22f01  g1515 ( .o(n8245_1), .a(_net_292), .b(net_367), .c(_net_291), .d(net_369) );
na02f01  g1516 ( .o(n8246), .a(n8245_1), .b(n8244) );
na02f01  g1517 ( .o(n8247), .a(n8246), .b(n7446_1) );
oa12f01  g1518 ( .o(n2167), .a(n8247), .b(n7446_1), .c(n8243) );
in01f01  g1519 ( .o(n8249_1), .a(_net_6963) );
in01f01  g1520 ( .o(n8250), .a(n1345) );
ao12f01  g1521 ( .o(n8251), .a(n8249_1), .b(_net_6962), .c(net_6961) );
in01f01  g1522 ( .o(n8252), .a(net_6961) );
in01f01  g1523 ( .o(n8253_1), .a(_net_6962) );
no03f01  g1524 ( .o(n8254), .a(n8253_1), .b(_net_6963), .c(n8252) );
no02f01  g1525 ( .o(n8255), .a(n8254), .b(n8251) );
na02f01  g1526 ( .o(n8256), .a(_net_6017), .b(n7682) );
oa22f01  g1527 ( .o(n2172), .a(n8256), .b(n8249_1), .c(n8255), .d(n8250) );
na02f01  g1528 ( .o(n8258_1), .a(n7298), .b(net_7737) );
ao22f01  g1529 ( .o(n8259), .a(n7306), .b(_net_6007), .c(n7291), .d(net_7708) );
na02f01  g1530 ( .o(n8260), .a(n7302_1), .b(net_147) );
na02f01  g1531 ( .o(n8261), .a(n7296), .b(net_247) );
na03f01  g1532 ( .o(n8262_1), .a(n7308), .b(_net_173), .c(n6800) );
na03f01  g1533 ( .o(n8263), .a(n7308), .b(_net_210), .c(x1322) );
na03f01  g1534 ( .o(n8264), .a(n8263), .b(n8262_1), .c(n8261) );
ao12f01  g1535 ( .o(n8265), .a(n8264), .b(n7286), .c(_net_290) );
na04f01  g1536 ( .o(n2177), .a(n8265), .b(n8260), .c(n8259), .d(n8258_1) );
no02f01  g1537 ( .o(n2181), .a(n6864), .b(n6863_1) );
in01f01  g1538 ( .o(n8268), .a(net_7108) );
in01f01  g1539 ( .o(n8269), .a(net_7172) );
oa22f01  g1540 ( .o(n8270), .a(n7580), .b(n8268), .c(n7577_1), .d(n8269) );
in01f01  g1541 ( .o(n8271_1), .a(net_7204) );
in01f01  g1542 ( .o(n8272), .a(net_7140) );
oa22f01  g1543 ( .o(n8273), .a(n7585), .b(n8272), .c(n7583), .d(n8271_1) );
no02f01  g1544 ( .o(n8274), .a(n8273), .b(n8270) );
no02f01  g1545 ( .o(n8275), .a(n8274), .b(n7721) );
in01f01  g1546 ( .o(n8276_1), .a(net_7174) );
in01f01  g1547 ( .o(n8277), .a(net_7110) );
oa22f01  g1548 ( .o(n8278), .a(n7580), .b(n8277), .c(n7577_1), .d(n8276_1) );
in01f01  g1549 ( .o(n8279), .a(net_7142) );
in01f01  g1550 ( .o(n8280_1), .a(net_7206) );
oa22f01  g1551 ( .o(n8281), .a(n7585), .b(n8279), .c(n7583), .d(n8280_1) );
no02f01  g1552 ( .o(n8282), .a(n8281), .b(n8278) );
no02f01  g1553 ( .o(n8283), .a(n8282), .b(n7592) );
in01f01  g1554 ( .o(n8284_1), .a(_net_6177) );
in01f01  g1555 ( .o(n8285), .a(net_7176) );
in01f01  g1556 ( .o(n8286), .a(net_7112) );
oa22f01  g1557 ( .o(n8287), .a(n7580), .b(n8286), .c(n7577_1), .d(n8285) );
in01f01  g1558 ( .o(n8288), .a(net_7144) );
in01f01  g1559 ( .o(n8289_1), .a(net_7208) );
oa22f01  g1560 ( .o(n8290), .a(n7585), .b(n8288), .c(n7583), .d(n8289_1) );
no02f01  g1561 ( .o(n8291), .a(n8290), .b(n8287) );
oa22f01  g1562 ( .o(n8292), .a(n8291), .b(n7574), .c(n7590), .d(n8284_1) );
no03f01  g1563 ( .o(n8293), .a(n8292), .b(n8283), .c(n8275) );
in01f01  g1564 ( .o(n8294_1), .a(net_7124) );
in01f01  g1565 ( .o(n8295), .a(net_7156) );
oa22f01  g1566 ( .o(n8296), .a(n7740), .b(n8294_1), .c(n7739), .d(n8295) );
in01f01  g1567 ( .o(n8297), .a(net_7220) );
in01f01  g1568 ( .o(n8298), .a(net_7188) );
oa22f01  g1569 ( .o(n8299_1), .a(n7745), .b(n8297), .c(n7744), .d(n8298) );
no02f01  g1570 ( .o(n8300), .a(n8299_1), .b(n8296) );
na02f01  g1571 ( .o(n2194), .a(n8300), .b(n8293) );
no02f01  g1572 ( .o(n8302), .a(n7576), .b(n7719_1) );
na02f01  g1573 ( .o(n8303_1), .a(n8302), .b(n7579) );
in01f01  g1574 ( .o(n8304), .a(n8302) );
na02f01  g1575 ( .o(n8305), .a(n8304), .b(_net_7229) );
na02f01  g1576 ( .o(n8306), .a(n8305), .b(n8303_1) );
no04f01  g1577 ( .o(n8307_1), .a(n7572_1), .b(n7570), .c(_net_6041), .d(_net_6042) );
na02f01  g1578 ( .o(n8308), .a(n8307_1), .b(n8306) );
na02f01  g1579 ( .o(n8309), .a(n7585), .b(n7577_1) );
no03f01  g1580 ( .o(n8310), .a(n7720), .b(n7572_1), .c(n7570) );
in01f01  g1581 ( .o(n8311_1), .a(n7572_1) );
no02f01  g1582 ( .o(n8312), .a(n8311_1), .b(n7570) );
ao22f01  g1583 ( .o(n8313), .a(n8312), .b(_net_7229), .c(n8310), .d(n8309) );
na02f01  g1584 ( .o(n2199), .a(n8313), .b(n8308) );
in01f01  g1585 ( .o(n8315), .a(n7304) );
no02f01  g1586 ( .o(n8316_1), .a(n7111_1), .b(n7341) );
na03f01  g1587 ( .o(n8317), .a(n8316_1), .b(n7281), .c(n6800) );
no02f01  g1588 ( .o(n2208), .a(n8317), .b(n8315) );
ao12f01  g1589 ( .o(n8319), .a(n8224_1), .b(_net_6828), .c(_net_6825) );
oa12f01  g1590 ( .o(n8320_1), .a(n8319), .b(_net_6828), .c(_net_6825) );
no02f01  g1591 ( .o(n8321), .a(n7128_1), .b(_net_6827) );
no02f01  g1592 ( .o(n8322), .a(_net_6824), .b(n8219) );
no02f01  g1593 ( .o(n8323), .a(n8322), .b(n8321) );
no02f01  g1594 ( .o(n8324_1), .a(n7125_1), .b(n8220_1) );
no02f01  g1595 ( .o(n8325), .a(_net_6823), .b(net_6826) );
no02f01  g1596 ( .o(n8326), .a(n8325), .b(n8324_1) );
in01f01  g1597 ( .o(n2948), .a(n8326) );
na02f01  g1598 ( .o(n8328), .a(n2948), .b(n8323) );
oa12f01  g1599 ( .o(n2213), .a(n7633), .b(n8328), .c(n8320_1) );
in01f01  g1600 ( .o(n8330), .a(_net_5963) );
no02f01  g1601 ( .o(n2222), .a(n6759), .b(n8330) );
in01f01  g1602 ( .o(n8332), .a(_net_6960) );
no02f01  g1603 ( .o(n8333), .a(n6806_1), .b(n6818_1) );
na03f01  g1604 ( .o(n8334_1), .a(n8333), .b(_net_6959), .c(n8332) );
in01f01  g1605 ( .o(n8335), .a(n8333) );
oa12f01  g1606 ( .o(n8336), .a(_net_6960), .b(n8335), .c(n6809_1) );
na02f01  g1607 ( .o(n8337_1), .a(n8336), .b(n8334_1) );
no04f01  g1608 ( .o(n8338), .a(n6821), .b(n6819), .c(_net_6020), .d(_net_6019) );
na02f01  g1609 ( .o(n8339), .a(n8338), .b(n8337_1) );
no03f01  g1610 ( .o(n8340_1), .a(n6823), .b(n6821), .c(n6819) );
no02f01  g1611 ( .o(n8341), .a(n6813_1), .b(n8332) );
no02f01  g1612 ( .o(n8342), .a(n6814), .b(_net_6960) );
no02f01  g1613 ( .o(n8343), .a(n8342), .b(n8341) );
in01f01  g1614 ( .o(n8344), .a(n6821) );
no02f01  g1615 ( .o(n8345_1), .a(n8344), .b(n6819) );
ao22f01  g1616 ( .o(n8346), .a(n8345_1), .b(_net_6960), .c(n8343), .d(n8340_1) );
na02f01  g1617 ( .o(n2227), .a(n8346), .b(n8339) );
in01f01  g1618 ( .o(n8348), .a(_net_7686) );
in01f01  g1619 ( .o(n8349), .a(_net_7682) );
no02f01  g1620 ( .o(n8350_1), .a(n8349), .b(n8348) );
no02f01  g1621 ( .o(n8351), .a(_net_7682), .b(_net_7686) );
no02f01  g1622 ( .o(n8352), .a(n8351), .b(n8350_1) );
in01f01  g1623 ( .o(n8353), .a(n8352) );
no02f01  g1624 ( .o(n8354_1), .a(n6733), .b(n6959) );
no02f01  g1625 ( .o(n8355), .a(net_7680), .b(_net_7684) );
no02f01  g1626 ( .o(n8356), .a(n8355), .b(n8354_1) );
in01f01  g1627 ( .o(n4405), .a(n8356) );
no02f01  g1628 ( .o(n8358), .a(n7397), .b(n6735) );
no02f01  g1629 ( .o(n8359_1), .a(_net_7685), .b(_net_7681) );
no02f01  g1630 ( .o(n8360), .a(n8359_1), .b(n8358) );
in01f01  g1631 ( .o(n8361), .a(n8360) );
na02f01  g1632 ( .o(n8362_1), .a(n8361), .b(n4405) );
no02f01  g1633 ( .o(n2232), .a(n8362_1), .b(n8353) );
no02f01  g1634 ( .o(n2237), .a(n7342), .b(n7111_1) );
in01f01  g1635 ( .o(n8365), .a(_net_7724) );
in01f01  g1636 ( .o(n8366), .a(_net_5994) );
ao12f01  g1637 ( .o(n2242), .a(n7343), .b(n8366), .c(n8365) );
ao22f01  g1638 ( .o(n8368), .a(n7288_1), .b(_net_6044), .c(n7286), .d(_net_283) );
ao22f01  g1639 ( .o(n8369), .a(n7298), .b(_net_7733), .c(n7291), .d(_net_7704) );
na02f01  g1640 ( .o(n8370), .a(n7302_1), .b(_net_127) );
na03f01  g1641 ( .o(n8371), .a(n7308), .b(net_206), .c(x1322) );
na02f01  g1642 ( .o(n8372_1), .a(n7296), .b(net_243) );
na03f01  g1643 ( .o(n8373), .a(n7308), .b(net_169), .c(n6800) );
na03f01  g1644 ( .o(n8374), .a(n8373), .b(n8372_1), .c(n8371) );
ao12f01  g1645 ( .o(n8375), .a(n8374), .b(n7306), .c(_net_6000) );
na04f01  g1646 ( .o(n2247), .a(n8375), .b(n8370), .c(n8369), .d(n8368) );
in01f01  g1647 ( .o(n8377_1), .a(_net_6402) );
na02f01  g1648 ( .o(n8378), .a(n8377_1), .b(net_6403) );
in01f01  g1649 ( .o(n8379), .a(net_6403) );
na02f01  g1650 ( .o(n8380), .a(_net_6402), .b(n8379) );
na02f01  g1651 ( .o(n2251), .a(n8380), .b(n8378) );
in01f01  g1652 ( .o(n8382_1), .a(_net_7401) );
na02f01  g1653 ( .o(n8383), .a(n7779_1), .b(n7550) );
oa12f01  g1654 ( .o(n2265), .a(n8383), .b(n7550), .c(n8382_1) );
in01f01  g1655 ( .o(n8385), .a(net_7096) );
no02f01  g1656 ( .o(n8386), .a(n8385), .b(n6984) );
no02f01  g1657 ( .o(n8387_1), .a(net_7096), .b(_net_7093) );
no02f01  g1658 ( .o(n8388), .a(n8387_1), .b(n8386) );
in01f01  g1659 ( .o(n2270), .a(n8388) );
no02f01  g1660 ( .o(n8390), .a(n7612), .b(n6824) );
in01f01  g1661 ( .o(n8391), .a(net_6906) );
in01f01  g1662 ( .o(n8392_1), .a(net_6842) );
oa22f01  g1663 ( .o(n8393), .a(n6810), .b(n8392_1), .c(n6807), .d(n8391) );
in01f01  g1664 ( .o(n8394), .a(net_6938) );
in01f01  g1665 ( .o(n8395), .a(net_6874) );
oa22f01  g1666 ( .o(n8396_1), .a(n6815), .b(n8395), .c(n6813_1), .d(n8394) );
no02f01  g1667 ( .o(n8397), .a(n8396_1), .b(n8393) );
no02f01  g1668 ( .o(n8398), .a(n8397), .b(n6826_1) );
in01f01  g1669 ( .o(n8399), .a(_net_6139) );
in01f01  g1670 ( .o(n8400), .a(net_6844) );
in01f01  g1671 ( .o(n8401_1), .a(net_6908) );
oa22f01  g1672 ( .o(n8402), .a(n6810), .b(n8400), .c(n6807), .d(n8401_1) );
in01f01  g1673 ( .o(n8403), .a(net_6940) );
in01f01  g1674 ( .o(n8404), .a(net_6876) );
oa22f01  g1675 ( .o(n8405_1), .a(n6815), .b(n8404), .c(n6813_1), .d(n8403) );
no02f01  g1676 ( .o(n8406), .a(n8405_1), .b(n8402) );
oa22f01  g1677 ( .o(n8407), .a(n8406), .b(n6836_1), .c(n6844), .d(n8399) );
no03f01  g1678 ( .o(n8408), .a(n8407), .b(n8398), .c(n8390) );
in01f01  g1679 ( .o(n8409), .a(net_6856) );
in01f01  g1680 ( .o(n8410_1), .a(net_6888) );
oa22f01  g1681 ( .o(n8411), .a(n6850_1), .b(n8409), .c(n6849), .d(n8410_1) );
in01f01  g1682 ( .o(n8412), .a(net_6952) );
in01f01  g1683 ( .o(n8413), .a(net_6920) );
oa22f01  g1684 ( .o(n8414), .a(n6855_1), .b(n8412), .c(n6854), .d(n8413) );
no02f01  g1685 ( .o(n8415_1), .a(n8414), .b(n8411) );
na02f01  g1686 ( .o(n2275), .a(n8415_1), .b(n8408) );
in01f01  g1687 ( .o(n8417), .a(_net_7748) );
ao12f01  g1688 ( .o(n2280), .a(n7343), .b(n8417), .c(n7652) );
in01f01  g1689 ( .o(n8419), .a(_net_6015) );
oa12f01  g1690 ( .o(n2298), .a(n8419), .b(n7117), .c(n7261) );
in01f01  g1691 ( .o(n8421), .a(_net_6186) );
no02f01  g1692 ( .o(n2303), .a(n8421), .b(_net_392) );
in01f01  g1693 ( .o(n8423), .a(_net_7556) );
na02f01  g1694 ( .o(n8424), .a(n6965), .b(net_7540) );
ao22f01  g1695 ( .o(n8425), .a(_net_292), .b(net_370), .c(_net_291), .d(net_372) );
na02f01  g1696 ( .o(n8426_1), .a(n8425), .b(n8424) );
na02f01  g1697 ( .o(n8427), .a(n8426_1), .b(n7519) );
oa12f01  g1698 ( .o(n2312), .a(n8427), .b(n7519), .c(n8423) );
in01f01  g1699 ( .o(n8429), .a(net_6899) );
in01f01  g1700 ( .o(n8430_1), .a(net_6835) );
oa22f01  g1701 ( .o(n8431), .a(n6810), .b(n8430_1), .c(n6807), .d(n8429) );
in01f01  g1702 ( .o(n8432), .a(net_6867) );
in01f01  g1703 ( .o(n8433), .a(net_6931) );
oa22f01  g1704 ( .o(n8434), .a(n6815), .b(n8432), .c(n6813_1), .d(n8433) );
no02f01  g1705 ( .o(n8435_1), .a(n8434), .b(n8431) );
no02f01  g1706 ( .o(n8436), .a(n8435_1), .b(n6824) );
in01f01  g1707 ( .o(n8437), .a(net_6901) );
in01f01  g1708 ( .o(n8438_1), .a(net_6837) );
oa22f01  g1709 ( .o(n8439), .a(n6810), .b(n8438_1), .c(n6807), .d(n8437) );
in01f01  g1710 ( .o(n8440), .a(net_6933) );
in01f01  g1711 ( .o(n8441), .a(net_6869) );
oa22f01  g1712 ( .o(n8442), .a(n6815), .b(n8441), .c(n6813_1), .d(n8440) );
no02f01  g1713 ( .o(n8443_1), .a(n8442), .b(n8439) );
no02f01  g1714 ( .o(n8444), .a(n8443_1), .b(n6826_1) );
in01f01  g1715 ( .o(n8445), .a(_net_6134) );
in01f01  g1716 ( .o(n8446), .a(net_6903) );
in01f01  g1717 ( .o(n8447_1), .a(net_6839) );
oa22f01  g1718 ( .o(n8448), .a(n6810), .b(n8447_1), .c(n6807), .d(n8446) );
in01f01  g1719 ( .o(n8449), .a(net_6935) );
in01f01  g1720 ( .o(n8450), .a(net_6871) );
oa22f01  g1721 ( .o(n8451_1), .a(n6815), .b(n8450), .c(n6813_1), .d(n8449) );
no02f01  g1722 ( .o(n8452), .a(n8451_1), .b(n8448) );
oa22f01  g1723 ( .o(n8453), .a(n8452), .b(n6836_1), .c(n6844), .d(n8445) );
no03f01  g1724 ( .o(n8454), .a(n8453), .b(n8444), .c(n8436) );
in01f01  g1725 ( .o(n8455_1), .a(net_6883) );
in01f01  g1726 ( .o(n8456), .a(net_6851) );
oa22f01  g1727 ( .o(n8457), .a(n6850_1), .b(n8456), .c(n6849), .d(n8455_1) );
in01f01  g1728 ( .o(n8458), .a(net_6915) );
in01f01  g1729 ( .o(n8459_1), .a(net_6947) );
oa22f01  g1730 ( .o(n8460), .a(n6855_1), .b(n8459_1), .c(n6854), .d(n8458) );
no02f01  g1731 ( .o(n8461), .a(n8460), .b(n8457) );
na02f01  g1732 ( .o(n2329), .a(n8461), .b(n8454) );
in01f01  g1733 ( .o(n8463), .a(_net_7747) );
ao12f01  g1734 ( .o(n2334), .a(n7343), .b(n8463), .c(n6907) );
in01f01  g1735 ( .o(n8465), .a(net_6979) );
in01f01  g1736 ( .o(n8466), .a(net_7043) );
oa22f01  g1737 ( .o(n8467_1), .a(n6987), .b(n8465), .c(n6985), .d(n8466) );
in01f01  g1738 ( .o(n8468), .a(net_7075) );
in01f01  g1739 ( .o(n8469), .a(net_7011) );
oa22f01  g1740 ( .o(n8470), .a(n6992), .b(n8469), .c(n6991), .d(n8468) );
no02f01  g1741 ( .o(n8471), .a(n8470), .b(n8467_1) );
no02f01  g1742 ( .o(n8472_1), .a(n8471), .b(n7012) );
in01f01  g1743 ( .o(n8473), .a(net_6981) );
in01f01  g1744 ( .o(n8474), .a(net_7045) );
oa22f01  g1745 ( .o(n8475), .a(n6987), .b(n8473), .c(n6985), .d(n8474) );
in01f01  g1746 ( .o(n8476), .a(net_7013) );
in01f01  g1747 ( .o(n8477_1), .a(net_7077) );
oa22f01  g1748 ( .o(n8478), .a(n6992), .b(n8476), .c(n6991), .d(n8477_1) );
no02f01  g1749 ( .o(n8479), .a(n8478), .b(n8475) );
no02f01  g1750 ( .o(n8480), .a(n8479), .b(n6997) );
ao22f01  g1751 ( .o(n8481_1), .a(n7000_1), .b(net_6983), .c(n6999), .d(net_7047) );
ao22f01  g1752 ( .o(n8482), .a(n7003), .b(net_7015), .c(n7002), .d(net_7079) );
ao12f01  g1753 ( .o(n8483), .a(n6980), .b(n8482), .c(n8481_1) );
in01f01  g1754 ( .o(n8484), .a(_net_6163) );
no02f01  g1755 ( .o(n8485), .a(n6995_1), .b(n8484) );
no04f01  g1756 ( .o(n8486_1), .a(n8485), .b(n8483), .c(n8480), .d(n8472_1) );
in01f01  g1757 ( .o(n8487), .a(net_6995) );
in01f01  g1758 ( .o(n8488), .a(net_7027) );
oa22f01  g1759 ( .o(n8489), .a(n8075_1), .b(n8487), .c(n8074), .d(n8488) );
in01f01  g1760 ( .o(n8490), .a(net_7091) );
in01f01  g1761 ( .o(n8491_1), .a(net_7059) );
oa22f01  g1762 ( .o(n8492), .a(n8080_1), .b(n8490), .c(n8079), .d(n8491_1) );
no02f01  g1763 ( .o(n8493), .a(n8492), .b(n8489) );
na02f01  g1764 ( .o(n2365), .a(n8493), .b(n8486_1) );
no02f01  g1765 ( .o(n8495), .a(_net_154), .b(_net_7720) );
no02f01  g1766 ( .o(n2377), .a(n8495), .b(n7343) );
ao22f01  g1767 ( .o(n8497), .a(n7581_1), .b(net_7104), .c(n7578), .d(net_7168) );
ao22f01  g1768 ( .o(n8498), .a(n7586_1), .b(net_7136), .c(n7584), .d(net_7200) );
na02f01  g1769 ( .o(n8499_1), .a(n8498), .b(n8497) );
na02f01  g1770 ( .o(n8500), .a(n8499_1), .b(n7575) );
ao22f01  g1771 ( .o(n8501), .a(n7593), .b(n7588), .c(n7591_1), .d(_net_6169) );
na02f01  g1772 ( .o(n8502), .a(n7914), .b(n7596_1) );
in01f01  g1773 ( .o(n8503), .a(net_7116) );
in01f01  g1774 ( .o(n8504_1), .a(net_7180) );
oa22f01  g1775 ( .o(n8505), .a(n7580), .b(n8503), .c(n7577_1), .d(n8504_1) );
in01f01  g1776 ( .o(n8506), .a(net_7148) );
in01f01  g1777 ( .o(n8507), .a(net_7212) );
oa22f01  g1778 ( .o(n8508_1), .a(n7585), .b(n8506), .c(n7583), .d(n8507) );
oa12f01  g1779 ( .o(n8509), .a(n7920_1), .b(n8508_1), .c(n8505) );
na04f01  g1780 ( .o(n2386), .a(n8509), .b(n8502), .c(n8501), .d(n8500) );
ao22f01  g1781 ( .o(n8511), .a(n6877), .b(_net_7277), .c(n6876_1), .d(net_7341) );
ao22f01  g1782 ( .o(n8512), .a(n6881_1), .b(net_7309), .c(n6880), .d(net_7373) );
na02f01  g1783 ( .o(n2395), .a(n8512), .b(n8511) );
in01f01  g1784 ( .o(n8514), .a(net_378) );
no02f01  g1785 ( .o(n2404), .a(n6966), .b(n8514) );
in01f01  g1786 ( .o(n8516), .a(_net_7511) );
na02f01  g1787 ( .o(n8517_1), .a(n7626_1), .b(n7504) );
oa12f01  g1788 ( .o(n2409), .a(n8517_1), .b(n7626_1), .c(n8516) );
ao22f01  g1789 ( .o(n8519), .a(n7288_1), .b(_net_6032), .c(n7286), .d(_net_271) );
ao22f01  g1790 ( .o(n8520), .a(n7298), .b(_net_7724), .c(n7291), .d(_net_7695) );
na02f01  g1791 ( .o(n8521), .a(n7302_1), .b(_net_118) );
na03f01  g1792 ( .o(n8522_1), .a(n7308), .b(net_197), .c(x1322) );
na02f01  g1793 ( .o(n8523), .a(n7296), .b(net_234) );
na03f01  g1794 ( .o(n8524), .a(n7308), .b(net_160), .c(n6800) );
na03f01  g1795 ( .o(n8525), .a(n8524), .b(n8523), .c(n8522_1) );
ao12f01  g1796 ( .o(n8526_1), .a(n8525), .b(n7306), .c(_net_5988) );
na04f01  g1797 ( .o(n2414), .a(n8526_1), .b(n8521), .c(n8520), .d(n8519) );
in01f01  g1798 ( .o(n8528), .a(_net_7431) );
na02f01  g1799 ( .o(n8529), .a(n1752), .b(n7550) );
oa12f01  g1800 ( .o(n2430), .a(n8529), .b(n7550), .c(n8528) );
in01f01  g1801 ( .o(n8531_1), .a(_net_279) );
na02f01  g1802 ( .o(n8532), .a(n7440), .b(net_7802) );
oa12f01  g1803 ( .o(n2435), .a(n8532), .b(n7440), .c(n8531_1) );
na02f01  g1804 ( .o(n8534), .a(n8337_1), .b(_net_6963) );
na03f01  g1805 ( .o(n8535_1), .a(n8336), .b(n8334_1), .c(n8249_1) );
na02f01  g1806 ( .o(n8536), .a(_net_6958), .b(n6818_1) );
na02f01  g1807 ( .o(n8537), .a(n6806_1), .b(_net_6957) );
na02f01  g1808 ( .o(n8538), .a(n8537), .b(n8536) );
na02f01  g1809 ( .o(n8539), .a(n8538), .b(net_6961) );
na03f01  g1810 ( .o(n8540_1), .a(n8537), .b(n8536), .c(n8252) );
ao22f01  g1811 ( .o(n8541), .a(n8540_1), .b(n8539), .c(n6823), .d(_net_6957) );
na02f01  g1812 ( .o(n8542), .a(n8333), .b(n6809_1) );
na02f01  g1813 ( .o(n8543), .a(n8335), .b(_net_6959) );
na02f01  g1814 ( .o(n8544_1), .a(n8543), .b(n8542) );
na02f01  g1815 ( .o(n8545), .a(n8544_1), .b(n8253_1) );
na03f01  g1816 ( .o(n8546), .a(n8543), .b(n8542), .c(_net_6962) );
na03f01  g1817 ( .o(n8547), .a(n8546), .b(n8545), .c(n8541) );
ao12f01  g1818 ( .o(n2444), .a(n8547), .b(n8535_1), .c(n8534) );
na02f01  g1819 ( .o(n8549_1), .a(n7348), .b(_net_7793) );
oa12f01  g1820 ( .o(n2457), .a(n8549_1), .b(n7348), .c(n6759) );
in01f01  g1821 ( .o(n8551), .a(net_6704) );
in01f01  g1822 ( .o(n8552_1), .a(net_6768) );
oa22f01  g1823 ( .o(n8553), .a(n7129), .b(n8551), .c(n7126), .d(n8552_1) );
in01f01  g1824 ( .o(n8554), .a(net_6800) );
in01f01  g1825 ( .o(n8555), .a(net_6736) );
oa22f01  g1826 ( .o(n8556), .a(n7134), .b(n8555), .c(n7132), .d(n8554) );
no02f01  g1827 ( .o(n8557_1), .a(n8556), .b(n8553) );
no02f01  g1828 ( .o(n8558), .a(n8557_1), .b(n7468_1) );
no02f01  g1829 ( .o(n8559), .a(n7470), .b(n7465) );
in01f01  g1830 ( .o(n8560), .a(_net_6118) );
oa22f01  g1831 ( .o(n8561_1), .a(n7477), .b(n7123), .c(n7118), .d(n8560) );
no03f01  g1832 ( .o(n8562), .a(n8561_1), .b(n8559), .c(n8558) );
in01f01  g1833 ( .o(n8563), .a(net_6720) );
in01f01  g1834 ( .o(n8564), .a(net_6752) );
oa22f01  g1835 ( .o(n8565_1), .a(n7492_1), .b(n8563), .c(n7491), .d(n8564) );
in01f01  g1836 ( .o(n8566), .a(net_6784) );
in01f01  g1837 ( .o(n8567), .a(net_6816) );
oa22f01  g1838 ( .o(n8568), .a(n7497), .b(n8567), .c(n7496_1), .d(n8566) );
no02f01  g1839 ( .o(n8569), .a(n8568), .b(n8565_1) );
na02f01  g1840 ( .o(n2470), .a(n8569), .b(n8562) );
in01f01  g1841 ( .o(n8571), .a(_net_7294) );
na02f01  g1842 ( .o(n8572), .a(n7926), .b(n7180) );
oa12f01  g1843 ( .o(n2479), .a(n8572), .b(n7180), .c(n8571) );
ao22f01  g1844 ( .o(n8574), .a(n7225), .b(_net_7432), .c(n7224), .d(net_7464) );
ao22f01  g1845 ( .o(n8575_1), .a(n7229), .b(net_7528), .c(n7228), .d(net_7496) );
na02f01  g1846 ( .o(n2484), .a(n8575_1), .b(n8574) );
in01f01  g1847 ( .o(n8577), .a(_net_7704) );
na02f01  g1848 ( .o(n8578_1), .a(n7207_1), .b(_net_7806) );
oa12f01  g1849 ( .o(n2505), .a(n8578_1), .b(n7207_1), .c(n8577) );
ao22f01  g1850 ( .o(n8580), .a(n6736_1), .b(net_7638), .c(n6734), .d(net_7606) );
ao22f01  g1851 ( .o(n8581), .a(n6739), .b(net_7670), .c(n6738), .d(_net_7574) );
na02f01  g1852 ( .o(n2510), .a(n8581), .b(n8580) );
no03f01  g1853 ( .o(n8583_1), .a(_net_6010), .b(n7121), .c(n7265_1) );
no02f01  g1854 ( .o(n8584), .a(n7121), .b(n7261) );
ao22f01  g1855 ( .o(n8585), .a(n8584), .b(n7271), .c(n8583_1), .d(n7269) );
ao12f01  g1856 ( .o(n8586), .a(n7121), .b(_net_5970), .c(n7261) );
no03f01  g1857 ( .o(n8587), .a(_net_6010), .b(n7121), .c(_net_6011) );
ao22f01  g1858 ( .o(n8588_1), .a(n8587), .b(n7267), .c(n8586), .d(n7260_1) );
na02f01  g1859 ( .o(n2515), .a(n8588_1), .b(n8585) );
ao22f01  g1860 ( .o(n8590), .a(n6877), .b(_net_7273), .c(n6876_1), .d(net_7337) );
ao22f01  g1861 ( .o(n8591), .a(n6881_1), .b(net_7305), .c(n6880), .d(net_7369) );
na02f01  g1862 ( .o(n2524), .a(n8591), .b(n8590) );
in01f01  g1863 ( .o(n8593_1), .a(_net_7419) );
na02f01  g1864 ( .o(n8594), .a(n8193), .b(n7550) );
oa12f01  g1865 ( .o(n2529), .a(n8594), .b(n7550), .c(n8593_1) );
in01f01  g1866 ( .o(n8596), .a(net_7040) );
in01f01  g1867 ( .o(n8597), .a(net_6976) );
oa22f01  g1868 ( .o(n8598_1), .a(n6987), .b(n8597), .c(n6985), .d(n8596) );
in01f01  g1869 ( .o(n8599), .a(net_7008) );
in01f01  g1870 ( .o(n8600), .a(net_7072) );
oa22f01  g1871 ( .o(n8601), .a(n6992), .b(n8599), .c(n6991), .d(n8600) );
no02f01  g1872 ( .o(n8602_1), .a(n8601), .b(n8598_1) );
no02f01  g1873 ( .o(n8603), .a(n8602_1), .b(n7012) );
in01f01  g1874 ( .o(n8604), .a(net_7042) );
in01f01  g1875 ( .o(n8605), .a(net_6978) );
oa22f01  g1876 ( .o(n8606), .a(n6987), .b(n8605), .c(n6985), .d(n8604) );
in01f01  g1877 ( .o(n8607_1), .a(net_7010) );
in01f01  g1878 ( .o(n8608), .a(net_7074) );
oa22f01  g1879 ( .o(n8609), .a(n6992), .b(n8607_1), .c(n6991), .d(n8608) );
no02f01  g1880 ( .o(n8610), .a(n8609), .b(n8606) );
no02f01  g1881 ( .o(n8611), .a(n8610), .b(n6997) );
in01f01  g1882 ( .o(n8612_1), .a(_net_6160) );
in01f01  g1883 ( .o(n8613), .a(net_6980) );
in01f01  g1884 ( .o(n8614), .a(net_7044) );
oa22f01  g1885 ( .o(n8615), .a(n6987), .b(n8613), .c(n6985), .d(n8614) );
in01f01  g1886 ( .o(n8616_1), .a(net_7076) );
in01f01  g1887 ( .o(n8617), .a(net_7012) );
oa22f01  g1888 ( .o(n8618), .a(n6992), .b(n8617), .c(n6991), .d(n8616_1) );
no02f01  g1889 ( .o(n8619), .a(n8618), .b(n8615) );
oa22f01  g1890 ( .o(n8620), .a(n8619), .b(n6980), .c(n6995_1), .d(n8612_1) );
no03f01  g1891 ( .o(n8621_1), .a(n8620), .b(n8611), .c(n8603) );
in01f01  g1892 ( .o(n8622), .a(net_7024) );
in01f01  g1893 ( .o(n8623), .a(net_6992) );
oa22f01  g1894 ( .o(n8624), .a(n8075_1), .b(n8623), .c(n8074), .d(n8622) );
in01f01  g1895 ( .o(n8625_1), .a(net_7056) );
in01f01  g1896 ( .o(n8626), .a(net_7088) );
oa22f01  g1897 ( .o(n8627), .a(n8080_1), .b(n8626), .c(n8079), .d(n8625_1) );
no02f01  g1898 ( .o(n8628_1), .a(n8627), .b(n8624) );
na02f01  g1899 ( .o(n2534), .a(n8628_1), .b(n8621_1) );
in01f01  g1900 ( .o(n8630), .a(_net_7445) );
na02f01  g1901 ( .o(n8631), .a(n6866), .b(net_7397) );
ao22f01  g1902 ( .o(n8632_1), .a(net_358), .b(_net_281), .c(_net_280), .d(net_360) );
na02f01  g1903 ( .o(n8633), .a(n8632_1), .b(n8631) );
na02f01  g1904 ( .o(n8634), .a(n8633), .b(n7197) );
oa12f01  g1905 ( .o(n2552), .a(n8634), .b(n7197), .c(n8630) );
in01f01  g1906 ( .o(n8636), .a(_net_7663) );
na02f01  g1907 ( .o(n8637_1), .a(n6965), .b(net_7551) );
ao22f01  g1908 ( .o(n8638), .a(_net_292), .b(net_381), .c(_net_291), .d(net_383) );
na02f01  g1909 ( .o(n8639), .a(n8638), .b(n8637_1) );
na02f01  g1910 ( .o(n8640), .a(n8639), .b(n7446_1) );
oa12f01  g1911 ( .o(n2566), .a(n8640), .b(n7446_1), .c(n8636) );
ao22f01  g1912 ( .o(n8642), .a(n6877), .b(_net_7270), .c(n6876_1), .d(net_7334) );
ao22f01  g1913 ( .o(n8643), .a(n6881_1), .b(net_7302), .c(n6880), .d(net_7366) );
na02f01  g1914 ( .o(n2575), .a(n8643), .b(n8642) );
ao22f01  g1915 ( .o(n8645_1), .a(n7225), .b(_net_7415), .c(n7224), .d(_net_7447) );
ao22f01  g1916 ( .o(n8646), .a(n7229), .b(_net_7511), .c(n7228), .d(_net_7479) );
na02f01  g1917 ( .o(n2580), .a(n8646), .b(n8645_1) );
in01f01  g1918 ( .o(n8648), .a(n7422_1) );
no02f01  g1919 ( .o(n2585), .a(n8648), .b(x868) );
in01f01  g1920 ( .o(n8650_1), .a(_net_5979) );
no02f01  g1921 ( .o(n2590), .a(n6976), .b(n8650_1) );
no02f01  g1922 ( .o(n2632), .a(n6963), .b(n6962) );
ao22f01  g1923 ( .o(n8653), .a(n6736_1), .b(net_7643), .c(n6734), .d(net_7611) );
ao22f01  g1924 ( .o(n8654_1), .a(n6739), .b(net_7675), .c(n6738), .d(_net_7579) );
na02f01  g1925 ( .o(n2637), .a(n8654_1), .b(n8653) );
ao22f01  g1926 ( .o(n8656), .a(n6877), .b(_net_7281), .c(n6876_1), .d(net_7345) );
ao22f01  g1927 ( .o(n8657), .a(n6881_1), .b(net_7313), .c(n6880), .d(net_7377) );
na02f01  g1928 ( .o(n2651), .a(n8657), .b(n8656) );
in01f01  g1929 ( .o(n8659), .a(net_6771) );
in01f01  g1930 ( .o(n8660), .a(net_6707) );
oa22f01  g1931 ( .o(n8661), .a(n7129), .b(n8660), .c(n7126), .d(n8659) );
in01f01  g1932 ( .o(n8662_1), .a(net_6803) );
in01f01  g1933 ( .o(n8663), .a(net_6739) );
oa22f01  g1934 ( .o(n8664), .a(n7134), .b(n8663), .c(n7132), .d(n8662_1) );
no02f01  g1935 ( .o(n8665), .a(n8664), .b(n8661) );
no02f01  g1936 ( .o(n8666_1), .a(n8665), .b(n7468_1) );
in01f01  g1937 ( .o(n8667), .a(net_6773) );
in01f01  g1938 ( .o(n8668), .a(net_6709) );
oa22f01  g1939 ( .o(n8669), .a(n7129), .b(n8668), .c(n7126), .d(n8667) );
in01f01  g1940 ( .o(n8670), .a(net_6741) );
in01f01  g1941 ( .o(n8671_1), .a(net_6805) );
oa22f01  g1942 ( .o(n8672), .a(n7134), .b(n8670), .c(n7132), .d(n8671_1) );
no02f01  g1943 ( .o(n8673), .a(n8672), .b(n8669) );
no02f01  g1944 ( .o(n8674), .a(n8673), .b(n7470) );
in01f01  g1945 ( .o(n8675), .a(_net_6121) );
in01f01  g1946 ( .o(n8676_1), .a(net_6711) );
in01f01  g1947 ( .o(n8677), .a(net_6775) );
oa22f01  g1948 ( .o(n8678), .a(n7129), .b(n8676_1), .c(n7126), .d(n8677) );
in01f01  g1949 ( .o(n8679), .a(net_6743) );
in01f01  g1950 ( .o(n8680), .a(net_6807) );
oa22f01  g1951 ( .o(n8681_1), .a(n7134), .b(n8679), .c(n7132), .d(n8680) );
no02f01  g1952 ( .o(n8682), .a(n8681_1), .b(n8678) );
oa22f01  g1953 ( .o(n8683), .a(n8682), .b(n7123), .c(n7118), .d(n8675) );
no03f01  g1954 ( .o(n8684), .a(n8683), .b(n8674), .c(n8666_1) );
in01f01  g1955 ( .o(n8685_1), .a(net_6723) );
in01f01  g1956 ( .o(n8686), .a(net_6755) );
oa22f01  g1957 ( .o(n8687), .a(n7492_1), .b(n8685_1), .c(n7491), .d(n8686) );
in01f01  g1958 ( .o(n8688), .a(net_6819) );
in01f01  g1959 ( .o(n8689_1), .a(net_6787) );
oa22f01  g1960 ( .o(n8690), .a(n7497), .b(n8688), .c(n7496_1), .d(n8689_1) );
no02f01  g1961 ( .o(n8691), .a(n8690), .b(n8687) );
na02f01  g1962 ( .o(n2665), .a(n8691), .b(n8684) );
in01f01  g1963 ( .o(n8693), .a(_net_6043) );
no02f01  g1964 ( .o(n8694_1), .a(n8693), .b(_net_6044) );
in01f01  g1965 ( .o(n8695), .a(_net_5980) );
na02f01  g1966 ( .o(n8696), .a(_net_6039), .b(_net_6045) );
ao12f01  g1967 ( .o(n8697), .a(n8696), .b(_net_5982), .c(n8695) );
na02f01  g1968 ( .o(n8698_1), .a(n8697), .b(n8694_1) );
in01f01  g1969 ( .o(n8699), .a(_net_6044) );
in01f01  g1970 ( .o(n8700), .a(n8696) );
na03f01  g1971 ( .o(n8701), .a(_net_5982), .b(_net_5981), .c(n8695) );
na04f01  g1972 ( .o(n8702), .a(n8701), .b(n8700), .c(n8693), .d(n8699) );
oa12f01  g1973 ( .o(n8703_1), .a(n8695), .b(_net_5982), .c(_net_5981) );
na04f01  g1974 ( .o(n8704), .a(n8703_1), .b(n8700), .c(n8693), .d(_net_6044) );
no02f01  g1975 ( .o(n8705), .a(n8693), .b(n8699) );
na03f01  g1976 ( .o(n8706), .a(n8705), .b(n8700), .c(_net_5980) );
na04f01  g1977 ( .o(n8707), .a(n8706), .b(n8704), .c(n8702), .d(n8698_1) );
in01f01  g1978 ( .o(n8708_1), .a(n8707) );
no02f01  g1979 ( .o(n2687), .a(n8708_1), .b(x906) );
in01f01  g1980 ( .o(n8710), .a(n7117) );
na02f01  g1981 ( .o(n8711_1), .a(n8710), .b(_net_6006) );
na03f01  g1982 ( .o(n8712), .a(n7467), .b(n8710), .c(_net_6822) );
na02f01  g1983 ( .o(n8713), .a(n7467), .b(n8710) );
na02f01  g1984 ( .o(n8714), .a(n8713), .b(n7466) );
na02f01  g1985 ( .o(n8715_1), .a(n8714), .b(n8712) );
no02f01  g1986 ( .o(n8716), .a(n8710), .b(n7121) );
na02f01  g1987 ( .o(n8717), .a(n8716), .b(_net_6822) );
oa12f01  g1988 ( .o(n2696), .a(n8717), .b(n8715_1), .c(n8711_1) );
in01f01  g1989 ( .o(n8719), .a(_net_126) );
na02f01  g1990 ( .o(n8720_1), .a(_net_154), .b(net_322) );
oa12f01  g1991 ( .o(n2713), .a(n8720_1), .b(_net_154), .c(n8719) );
ao22f01  g1992 ( .o(n8722), .a(n6736_1), .b(_net_7624), .c(n6734), .d(_net_7592) );
ao22f01  g1993 ( .o(n8723), .a(n6739), .b(_net_7656), .c(n6738), .d(_net_7560) );
na02f01  g1994 ( .o(n2718), .a(n8723), .b(n8722) );
in01f01  g1995 ( .o(n8725_1), .a(_net_280) );
na02f01  g1996 ( .o(n8726), .a(n7440), .b(_net_7803) );
oa12f01  g1997 ( .o(n2723), .a(n8726), .b(n7440), .c(n8725_1) );
in01f01  g1998 ( .o(n8728), .a(_net_7314) );
na02f01  g1999 ( .o(n8729), .a(n6898), .b(net_7234) );
ao22f01  g2000 ( .o(n8730_1), .a(net_328), .b(_net_269), .c(_net_270), .d(net_326) );
na02f01  g2001 ( .o(n8731), .a(n8730_1), .b(n8729) );
na02f01  g2002 ( .o(n8732), .a(n8731), .b(n7150) );
oa12f01  g2003 ( .o(n2732), .a(n8732), .b(n7150), .c(n8728) );
ao22f01  g2004 ( .o(n8734_1), .a(n6877), .b(_net_7257), .c(n6876_1), .d(_net_7321) );
ao22f01  g2005 ( .o(n8735), .a(n6881_1), .b(_net_7289), .c(n6880), .d(_net_7353) );
na02f01  g2006 ( .o(n2753), .a(n8735), .b(n8734_1) );
no02f01  g2007 ( .o(n8737), .a(n7813), .b(n6945) );
no02f01  g2008 ( .o(n8738), .a(n7822_1), .b(n6934_1) );
in01f01  g2009 ( .o(n8739_1), .a(_net_6097) );
in01f01  g2010 ( .o(n8740), .a(net_6636) );
in01f01  g2011 ( .o(n8741), .a(net_6572) );
oa22f01  g2012 ( .o(n8742), .a(n6922), .b(n8741), .c(n6919_1), .d(n8740) );
in01f01  g2013 ( .o(n8743_1), .a(net_6668) );
in01f01  g2014 ( .o(n8744), .a(net_6604) );
oa22f01  g2015 ( .o(n8745), .a(n6927), .b(n8744), .c(n6925), .d(n8743_1) );
no02f01  g2016 ( .o(n8746), .a(n8745), .b(n8742) );
oa22f01  g2017 ( .o(n8747), .a(n8746), .b(n6916), .c(n6932), .d(n8739_1) );
no03f01  g2018 ( .o(n8748_1), .a(n8747), .b(n8738), .c(n8737) );
in01f01  g2019 ( .o(n8749), .a(net_6616) );
in01f01  g2020 ( .o(n8750), .a(net_6584) );
oa22f01  g2021 ( .o(n8751), .a(n7058_1), .b(n8750), .c(n7057), .d(n8749) );
in01f01  g2022 ( .o(n8752), .a(net_6680) );
in01f01  g2023 ( .o(n8753_1), .a(net_6648) );
oa22f01  g2024 ( .o(n8754), .a(n7063), .b(n8752), .c(n7062_1), .d(n8753_1) );
no02f01  g2025 ( .o(n8755), .a(n8754), .b(n8751) );
na02f01  g2026 ( .o(n2758), .a(n8755), .b(n8748_1) );
na02f01  g2027 ( .o(n8757_1), .a(n7348), .b(_net_7822) );
oa12f01  g2028 ( .o(n2771), .a(n8757_1), .b(n7348), .c(n7689) );
no02f01  g2029 ( .o(n8759), .a(_net_7097), .b(n6986_1) );
in01f01  g2030 ( .o(n8760), .a(_net_7097) );
no02f01  g2031 ( .o(n8761), .a(n8760), .b(_net_7094) );
no02f01  g2032 ( .o(n8762_1), .a(n8761), .b(n8759) );
no02f01  g2033 ( .o(n8763), .a(net_7096), .b(n6984) );
no02f01  g2034 ( .o(n8764), .a(n8763), .b(n8762_1) );
no04f01  g2035 ( .o(n8765), .a(n8761), .b(n8759), .c(net_7096), .d(n6984) );
oa12f01  g2036 ( .o(n8766), .a(n8388), .b(n8765), .c(n8764) );
no02f01  g2037 ( .o(n8767_1), .a(n8765), .b(n8764) );
na02f01  g2038 ( .o(n8768), .a(n8767_1), .b(n2270) );
na02f01  g2039 ( .o(n2776), .a(n8768), .b(n8766) );
ao22f01  g2040 ( .o(n8770), .a(n6738), .b(_net_7554), .c(n6736_1), .d(_net_7618) );
ao22f01  g2041 ( .o(n8771_1), .a(n6739), .b(_net_7650), .c(n6734), .d(_net_7586) );
na02f01  g2042 ( .o(n2797), .a(n8771_1), .b(n8770) );
ao22f01  g2043 ( .o(n8773), .a(n7225), .b(_net_7422), .c(n7224), .d(net_7454) );
ao22f01  g2044 ( .o(n8774), .a(n7229), .b(net_7518), .c(n7228), .d(net_7486) );
na02f01  g2045 ( .o(n2810), .a(n8774), .b(n8773) );
in01f01  g2046 ( .o(n8776), .a(net_7036) );
in01f01  g2047 ( .o(n8777), .a(net_6972) );
oa22f01  g2048 ( .o(n8778), .a(n6987), .b(n8777), .c(n6985), .d(n8776) );
in01f01  g2049 ( .o(n8779), .a(net_7004) );
in01f01  g2050 ( .o(n8780_1), .a(net_7068) );
oa22f01  g2051 ( .o(n8781), .a(n6992), .b(n8779), .c(n6991), .d(n8780_1) );
no02f01  g2052 ( .o(n8782), .a(n8781), .b(n8778) );
no02f01  g2053 ( .o(n8783), .a(n8782), .b(n7012) );
in01f01  g2054 ( .o(n8784_1), .a(net_6974) );
in01f01  g2055 ( .o(n8785), .a(net_7038) );
oa22f01  g2056 ( .o(n8786), .a(n6987), .b(n8784_1), .c(n6985), .d(n8785) );
in01f01  g2057 ( .o(n8787), .a(net_7070) );
in01f01  g2058 ( .o(n8788_1), .a(net_7006) );
oa22f01  g2059 ( .o(n8789), .a(n6992), .b(n8788_1), .c(n6991), .d(n8787) );
no02f01  g2060 ( .o(n8790), .a(n8789), .b(n8786) );
no02f01  g2061 ( .o(n8791), .a(n8790), .b(n6997) );
in01f01  g2062 ( .o(n8792), .a(_net_6156) );
oa22f01  g2063 ( .o(n8793_1), .a(n8602_1), .b(n6980), .c(n6995_1), .d(n8792) );
no03f01  g2064 ( .o(n8794), .a(n8793_1), .b(n8791), .c(n8783) );
in01f01  g2065 ( .o(n8795), .a(net_6988) );
in01f01  g2066 ( .o(n8796), .a(net_7020) );
oa22f01  g2067 ( .o(n8797_1), .a(n8075_1), .b(n8795), .c(n8074), .d(n8796) );
in01f01  g2068 ( .o(n8798), .a(net_7052) );
in01f01  g2069 ( .o(n8799), .a(net_7084) );
oa22f01  g2070 ( .o(n8800_1), .a(n8080_1), .b(n8799), .c(n8079), .d(n8798) );
no02f01  g2071 ( .o(n8801), .a(n8800_1), .b(n8797_1) );
na02f01  g2072 ( .o(n2831), .a(n8801), .b(n8794) );
in01f01  g2073 ( .o(n8803), .a(_net_7794) );
na02f01  g2074 ( .o(n8804), .a(n6803), .b(_net_6029) );
oa12f01  g2075 ( .o(n2836), .a(n8804), .b(n6803), .c(n8803) );
in01f01  g2076 ( .o(n8806), .a(_net_7261) );
na02f01  g2077 ( .o(n8807), .a(n6898), .b(net_7245) );
ao22f01  g2078 ( .o(n8808), .a(_net_269), .b(net_339), .c(_net_270), .d(net_337) );
na02f01  g2079 ( .o(n8809_1), .a(n8808), .b(n8807) );
na02f01  g2080 ( .o(n8810), .a(n8809_1), .b(n6901) );
oa12f01  g2081 ( .o(n2845), .a(n8810), .b(n6901), .c(n8806) );
in01f01  g2082 ( .o(n8812), .a(net_376) );
no02f01  g2083 ( .o(n2850), .a(n6966), .b(n8812) );
in01f01  g2084 ( .o(n8814), .a(_net_7501) );
na02f01  g2085 ( .o(n8815), .a(n6866), .b(net_7389) );
ao22f01  g2086 ( .o(n8816), .a(net_350), .b(_net_281), .c(_net_280), .d(net_352) );
na02f01  g2087 ( .o(n8817), .a(n8816), .b(n8815) );
na02f01  g2088 ( .o(n8818_1), .a(n8817), .b(n7626_1) );
oa12f01  g2089 ( .o(n2855), .a(n8818_1), .b(n7626_1), .c(n8814) );
in01f01  g2090 ( .o(n8820), .a(_net_7572) );
na02f01  g2091 ( .o(n8821), .a(n7519), .b(n615) );
oa12f01  g2092 ( .o(n2890), .a(n8821), .b(n7519), .c(n8820) );
in01f01  g2093 ( .o(n8823_1), .a(net_5992) );
in01f01  g2094 ( .o(n8824), .a(_net_7722) );
ao12f01  g2095 ( .o(n2900), .a(n7343), .b(n8824), .c(n8823_1) );
in01f01  g2096 ( .o(n8826_1), .a(net_336) );
no02f01  g2097 ( .o(n2913), .a(n6899_1), .b(n8826_1) );
na02f01  g2098 ( .o(n8828), .a(n7298), .b(net_7742) );
ao22f01  g2099 ( .o(n8829), .a(n7306), .b(_net_6012), .c(n7291), .d(net_7713) );
na02f01  g2100 ( .o(n8830), .a(n7302_1), .b(net_152) );
na02f01  g2101 ( .o(n8831_1), .a(n7296), .b(net_252) );
na03f01  g2102 ( .o(n8832), .a(n7308), .b(_net_178), .c(n6800) );
na03f01  g2103 ( .o(n8833), .a(n7308), .b(_net_215), .c(x1322) );
na03f01  g2104 ( .o(n8834), .a(n8833), .b(n8832), .c(n8831_1) );
ao12f01  g2105 ( .o(n8835_1), .a(n8834), .b(n7286), .c(_net_295) );
na04f01  g2106 ( .o(n2918), .a(n8835_1), .b(n8830), .c(n8829), .d(n8828) );
in01f01  g2107 ( .o(n8837), .a(_net_6220) );
no02f01  g2108 ( .o(n2930), .a(_net_392), .b(n8837) );
in01f01  g2109 ( .o(n8839), .a(_net_7552) );
na02f01  g2110 ( .o(n8840_1), .a(n6965), .b(net_7536) );
ao22f01  g2111 ( .o(n8841), .a(net_366), .b(_net_292), .c(net_368), .d(_net_291) );
na02f01  g2112 ( .o(n8842), .a(n8841), .b(n8840_1) );
na02f01  g2113 ( .o(n8843), .a(n8842), .b(n7519) );
oa12f01  g2114 ( .o(n2953), .a(n8843), .b(n7519), .c(n8839) );
in01f01  g2115 ( .o(n8845_1), .a(net_358) );
no02f01  g2116 ( .o(n2958), .a(n6867_1), .b(n8845_1) );
no02f01  g2117 ( .o(n8847), .a(net_7680), .b(n6959) );
in01f01  g2118 ( .o(n8848), .a(n8847) );
no02f01  g2119 ( .o(n8849), .a(n8848), .b(n8360) );
no02f01  g2120 ( .o(n8850_1), .a(n8847), .b(n8361) );
oa12f01  g2121 ( .o(n8851), .a(n8356), .b(n8850_1), .c(n8849) );
no02f01  g2122 ( .o(n8852), .a(n8850_1), .b(n8849) );
na02f01  g2123 ( .o(n8853), .a(n8852), .b(n4405) );
na02f01  g2124 ( .o(n2976), .a(n8853), .b(n8851) );
in01f01  g2125 ( .o(n8855_1), .a(n6761_1) );
na02f01  g2126 ( .o(n8856), .a(n6763), .b(n8855_1) );
in01f01  g2127 ( .o(n8857), .a(n8856) );
na02f01  g2128 ( .o(n8858), .a(n8855_1), .b(_net_5984) );
no02f01  g2129 ( .o(n8859), .a(n8858), .b(n8857) );
na02f01  g2130 ( .o(n8860_1), .a(n8859), .b(n6747) );
no02f01  g2131 ( .o(n8861), .a(n8858), .b(n8856) );
no02f01  g2132 ( .o(n8862), .a(n8855_1), .b(n6759) );
ao22f01  g2133 ( .o(n8863), .a(n8862), .b(_net_6553), .c(n8861), .d(n7760_1) );
na02f01  g2134 ( .o(n2981), .a(n8863), .b(n8860_1) );
oa12f01  g2135 ( .o(n2986), .a(n6886_1), .b(_net_7791), .c(n7165) );
in01f01  g2136 ( .o(n8866), .a(_net_7531) );
no02f01  g2137 ( .o(n8867), .a(n7229), .b(n8866) );
no03f01  g2138 ( .o(n8868), .a(n7227), .b(n7223), .c(_net_7531) );
no02f01  g2139 ( .o(n8869_1), .a(n8868), .b(n8867) );
in01f01  g2140 ( .o(n8870), .a(_net_227) );
no02f01  g2141 ( .o(n5792), .a(n7850), .b(n8870) );
in01f01  g2142 ( .o(n8872), .a(n5792) );
na02f01  g2143 ( .o(n8873_1), .a(_net_278), .b(n8870) );
oa22f01  g2144 ( .o(n2991), .a(n8873_1), .b(n8866), .c(n8872), .d(n8869_1) );
in01f01  g2145 ( .o(n8875), .a(_net_6038) );
ao12f01  g2146 ( .o(n8876), .a(n8650_1), .b(_net_7098), .c(_net_7095) );
oa12f01  g2147 ( .o(n8877_1), .a(n8876), .b(_net_7098), .c(_net_7095) );
na02f01  g2148 ( .o(n8878), .a(n8762_1), .b(n2270) );
oa12f01  g2149 ( .o(n3000), .a(n8875), .b(n8878), .c(n8877_1) );
in01f01  g2150 ( .o(n8880), .a(net_6629) );
in01f01  g2151 ( .o(n8881), .a(net_6565) );
oa22f01  g2152 ( .o(n8882_1), .a(n6922), .b(n8881), .c(n6919_1), .d(n8880) );
in01f01  g2153 ( .o(n8883), .a(net_6661) );
in01f01  g2154 ( .o(n8884), .a(net_6597) );
oa22f01  g2155 ( .o(n8885), .a(n6927), .b(n8884), .c(n6925), .d(n8883) );
oa12f01  g2156 ( .o(n8886_1), .a(n6917), .b(n8885), .c(n8882_1) );
ao22f01  g2157 ( .o(n8887), .a(n6935), .b(n6930), .c(n6933), .d(_net_6090) );
in01f01  g2158 ( .o(n8888), .a(net_6641) );
in01f01  g2159 ( .o(n8889), .a(net_6577) );
oa22f01  g2160 ( .o(n8890), .a(n6922), .b(n8889), .c(n6919_1), .d(n8888) );
in01f01  g2161 ( .o(n8891_1), .a(net_6609) );
in01f01  g2162 ( .o(n8892), .a(net_6673) );
oa22f01  g2163 ( .o(n8893), .a(n6927), .b(n8891_1), .c(n6925), .d(n8892) );
no02f01  g2164 ( .o(n8894), .a(n8893), .b(n8890) );
no03f01  g2165 ( .o(n8895_1), .a(n8894), .b(n6947_1), .c(n6943_1) );
ao12f01  g2166 ( .o(n8896), .a(n8895_1), .b(n6946), .c(n6938_1) );
na03f01  g2167 ( .o(n3005), .a(n8896), .b(n8887), .c(n8886_1) );
no02f01  g2168 ( .o(n3010), .a(n7232), .b(n7163) );
in01f01  g2169 ( .o(n8899_1), .a(net_379) );
no02f01  g2170 ( .o(n3015), .a(n6966), .b(n8899_1) );
in01f01  g2171 ( .o(n8901), .a(_net_7320) );
na02f01  g2172 ( .o(n8902), .a(n8208), .b(n7150) );
oa12f01  g2173 ( .o(n3020), .a(n8902), .b(n7150), .c(n8901) );
ao22f01  g2174 ( .o(n8904), .a(n6877), .b(_net_7267), .c(n6876_1), .d(_net_7331) );
ao22f01  g2175 ( .o(n8905), .a(n6881_1), .b(_net_7299), .c(n6880), .d(_net_7363) );
na02f01  g2176 ( .o(n3025), .a(n8905), .b(n8904) );
in01f01  g2177 ( .o(n8907), .a(_net_6023) );
na02f01  g2178 ( .o(n8908_1), .a(n7348), .b(_net_7823) );
oa12f01  g2179 ( .o(n3042), .a(n8908_1), .b(n7348), .c(n8907) );
in01f01  g2180 ( .o(n8910), .a(_net_7667) );
na02f01  g2181 ( .o(n8911), .a(n7446_1), .b(n7144) );
oa12f01  g2182 ( .o(n3047), .a(n8911), .b(n7446_1), .c(n8910) );
no02f01  g2183 ( .o(n8913), .a(n8866), .b(n7867_1) );
no02f01  g2184 ( .o(n8914), .a(_net_7531), .b(_net_7535) );
no02f01  g2185 ( .o(n8915), .a(n8914), .b(n8913) );
in01f01  g2186 ( .o(n8916), .a(n8915) );
no02f01  g2187 ( .o(n8917_1), .a(n7194_1), .b(n7223) );
no02f01  g2188 ( .o(n8918), .a(_net_7533), .b(net_7529) );
no02f01  g2189 ( .o(n8919), .a(n8918), .b(n8917_1) );
in01f01  g2190 ( .o(n8850), .a(n8919) );
no02f01  g2191 ( .o(n8921), .a(n7227), .b(n6860_1) );
no02f01  g2192 ( .o(n8922_1), .a(_net_7530), .b(_net_7534) );
no02f01  g2193 ( .o(n8923), .a(n8922_1), .b(n8921) );
in01f01  g2194 ( .o(n8924), .a(n8923) );
na02f01  g2195 ( .o(n8925), .a(n8924), .b(n8850) );
no02f01  g2196 ( .o(n3056), .a(n8925), .b(n8916) );
ao22f01  g2197 ( .o(n8927), .a(n6877), .b(_net_7278), .c(n6876_1), .d(net_7342) );
ao22f01  g2198 ( .o(n8928), .a(n6881_1), .b(net_7310), .c(n6880), .d(net_7374) );
na02f01  g2199 ( .o(n3065), .a(n8928), .b(n8927) );
ao22f01  g2200 ( .o(n8930), .a(n6738), .b(_net_7555), .c(n6736_1), .d(_net_7619) );
ao22f01  g2201 ( .o(n8931_1), .a(n6739), .b(_net_7651), .c(n6734), .d(_net_7587) );
na02f01  g2202 ( .o(n3078), .a(n8931_1), .b(n8930) );
na02f01  g2203 ( .o(n8933), .a(n8127), .b(n6918) );
na02f01  g2204 ( .o(n8934_1), .a(n6943_1), .b(_net_6688) );
na02f01  g2205 ( .o(n8935), .a(_net_6687), .b(n6918) );
na02f01  g2206 ( .o(n8936), .a(n8935), .b(n8934_1) );
ao22f01  g2207 ( .o(n8937), .a(n8936), .b(n8125_1), .c(n8132), .d(_net_6688) );
na02f01  g2208 ( .o(n3087), .a(n8937), .b(n8933) );
in01f01  g2209 ( .o(n8939_1), .a(_net_6280) );
no02f01  g2210 ( .o(n3092), .a(n8939_1), .b(_net_392) );
in01f01  g2211 ( .o(n8941), .a(_net_128) );
na02f01  g2212 ( .o(n8942), .a(net_324), .b(_net_154) );
oa12f01  g2213 ( .o(n3097), .a(n8942), .b(_net_154), .c(n8941) );
in01f01  g2214 ( .o(n8944), .a(_net_7410) );
na02f01  g2215 ( .o(n8945), .a(n7550), .b(n6891) );
oa12f01  g2216 ( .o(n3130), .a(n8945), .b(n7550), .c(n8944) );
in01f01  g2217 ( .o(n8947), .a(_net_7557) );
na02f01  g2218 ( .o(n8948_1), .a(n7519), .b(n7449) );
oa12f01  g2219 ( .o(n3139), .a(n8948_1), .b(n7519), .c(n8947) );
in01f01  g2220 ( .o(n8950), .a(_net_7449) );
na02f01  g2221 ( .o(n8951), .a(n7197), .b(n6872_1) );
oa12f01  g2222 ( .o(n3148), .a(n8951), .b(n7197), .c(n8950) );
no03f01  g2223 ( .o(n3157), .a(n7336), .b(n7109), .c(n7105) );
in01f01  g2224 ( .o(n8954), .a(_net_7470) );
na02f01  g2225 ( .o(n8955), .a(n7860), .b(n6869) );
oa12f01  g2226 ( .o(n3170), .a(n8955), .b(n6869), .c(n8954) );
in01f01  g2227 ( .o(n8957), .a(_net_7350) );
na02f01  g2228 ( .o(n8958_1), .a(n6898), .b(net_7238) );
ao22f01  g2229 ( .o(n8959), .a(net_332), .b(_net_269), .c(net_330), .d(_net_270) );
na02f01  g2230 ( .o(n8960), .a(n8959), .b(n8958_1) );
na02f01  g2231 ( .o(n8961), .a(n8960), .b(n7030) );
oa12f01  g2232 ( .o(n3182), .a(n8961), .b(n7030), .c(n8957) );
in01f01  g2233 ( .o(n8963_1), .a(_net_7277) );
in01f01  g2234 ( .o(n8964), .a(net_341) );
no02f01  g2235 ( .o(n6376), .a(n6899_1), .b(n8964) );
na02f01  g2236 ( .o(n8966), .a(n6376), .b(n6901) );
oa12f01  g2237 ( .o(n3194), .a(n8966), .b(n6901), .c(n8963_1) );
ao22f01  g2238 ( .o(n8968), .a(n6877), .b(_net_7272), .c(n6876_1), .d(net_7336) );
ao22f01  g2239 ( .o(n8969), .a(n6881_1), .b(net_7304), .c(n6880), .d(net_7368) );
na02f01  g2240 ( .o(n3203), .a(n8969), .b(n8968) );
in01f01  g2241 ( .o(n8971_1), .a(_net_7326) );
na02f01  g2242 ( .o(n8972), .a(n7926), .b(n7150) );
oa12f01  g2243 ( .o(n3212), .a(n8972), .b(n7150), .c(n8971_1) );
in01f01  g2244 ( .o(n8974), .a(net_6764) );
in01f01  g2245 ( .o(n8975), .a(net_6700) );
oa22f01  g2246 ( .o(n8976_1), .a(n7129), .b(n8975), .c(n7126), .d(n8974) );
in01f01  g2247 ( .o(n8977), .a(net_6732) );
in01f01  g2248 ( .o(n8978), .a(net_6796) );
oa22f01  g2249 ( .o(n8979), .a(n7134), .b(n8977), .c(n7132), .d(n8978) );
oa12f01  g2250 ( .o(n8980), .a(n7124), .b(n8979), .c(n8976_1) );
ao22f01  g2251 ( .o(n8981_1), .a(n8157), .b(n8159), .c(n7119), .d(_net_6110) );
na02f01  g2252 ( .o(n8982), .a(n8162), .b(n8164) );
in01f01  g2253 ( .o(n8983), .a(net_6776) );
in01f01  g2254 ( .o(n8984), .a(net_6712) );
oa22f01  g2255 ( .o(n8985), .a(n7129), .b(n8984), .c(n7126), .d(n8983) );
in01f01  g2256 ( .o(n8986_1), .a(net_6808) );
in01f01  g2257 ( .o(n8987), .a(net_6744) );
oa22f01  g2258 ( .o(n8988), .a(n7134), .b(n8987), .c(n7132), .d(n8986_1) );
oa12f01  g2259 ( .o(n8989), .a(n8167), .b(n8988), .c(n8985) );
na04f01  g2260 ( .o(n3217), .a(n8989), .b(n8982), .c(n8981_1), .d(n8980) );
in01f01  g2261 ( .o(n8991), .a(_net_7478) );
na02f01  g2262 ( .o(n8992), .a(n6866), .b(net_7398) );
ao22f01  g2263 ( .o(n8993), .a(net_359), .b(_net_281), .c(_net_280), .d(net_361) );
na02f01  g2264 ( .o(n8994), .a(n8993), .b(n8992) );
na02f01  g2265 ( .o(n8995_1), .a(n8994), .b(n6869) );
oa12f01  g2266 ( .o(n3222), .a(n8995_1), .b(n6869), .c(n8991) );
in01f01  g2267 ( .o(n8997), .a(net_7770) );
no03f01  g2268 ( .o(n3231), .a(n7232), .b(n8997), .c(net_7771) );
in01f01  g2269 ( .o(n8999), .a(net_7106) );
in01f01  g2270 ( .o(n9000_1), .a(net_7170) );
oa22f01  g2271 ( .o(n9001), .a(n7580), .b(n8999), .c(n7577_1), .d(n9000_1) );
in01f01  g2272 ( .o(n9002), .a(net_7202) );
in01f01  g2273 ( .o(n9003), .a(net_7138) );
oa22f01  g2274 ( .o(n9004), .a(n7585), .b(n9003), .c(n7583), .d(n9002) );
no02f01  g2275 ( .o(n9005_1), .a(n9004), .b(n9001) );
no02f01  g2276 ( .o(n9006), .a(n9005_1), .b(n7721) );
no02f01  g2277 ( .o(n9007), .a(n8274), .b(n7592) );
in01f01  g2278 ( .o(n9008), .a(_net_6175) );
oa22f01  g2279 ( .o(n9009), .a(n8282), .b(n7574), .c(n7590), .d(n9008) );
no03f01  g2280 ( .o(n9010_1), .a(n9009), .b(n9007), .c(n9006) );
in01f01  g2281 ( .o(n9011), .a(net_7154) );
in01f01  g2282 ( .o(n9012), .a(net_7122) );
oa22f01  g2283 ( .o(n9013), .a(n7740), .b(n9012), .c(n7739), .d(n9011) );
in01f01  g2284 ( .o(n9014_1), .a(net_7186) );
in01f01  g2285 ( .o(n9015), .a(net_7218) );
oa22f01  g2286 ( .o(n9016), .a(n7745), .b(n9015), .c(n7744), .d(n9014_1) );
no02f01  g2287 ( .o(n9017_1), .a(n9016), .b(n9013) );
na02f01  g2288 ( .o(n3240), .a(n9017_1), .b(n9010_1) );
in01f01  g2289 ( .o(n9019), .a(_net_272) );
na02f01  g2290 ( .o(n9020), .a(n7440), .b(_net_7798) );
oa12f01  g2291 ( .o(n3254), .a(n9020), .b(n7440), .c(n9019) );
in01f01  g2292 ( .o(n9022_1), .a(_net_116) );
na02f01  g2293 ( .o(n9023), .a(net_312), .b(_net_154) );
oa12f01  g2294 ( .o(n3263), .a(n9023), .b(n9022_1), .c(_net_154) );
no02f01  g2295 ( .o(n9025_1), .a(n7050), .b(n6945) );
no02f01  g2296 ( .o(n9026), .a(n6954), .b(n6934_1) );
in01f01  g2297 ( .o(n9027), .a(_net_6102) );
oa22f01  g2298 ( .o(n9028), .a(n8894), .b(n6916), .c(n6932), .d(n9027) );
no03f01  g2299 ( .o(n9029), .a(n9028), .b(n9026), .c(n9025_1) );
in01f01  g2300 ( .o(n9030_1), .a(net_6589) );
in01f01  g2301 ( .o(n9031), .a(net_6621) );
oa22f01  g2302 ( .o(n9032), .a(n7058_1), .b(n9030_1), .c(n7057), .d(n9031) );
in01f01  g2303 ( .o(n9033), .a(net_6653) );
in01f01  g2304 ( .o(n9034_1), .a(net_6685) );
oa22f01  g2305 ( .o(n9035), .a(n7063), .b(n9034_1), .c(n7062_1), .d(n9033) );
no02f01  g2306 ( .o(n9036), .a(n9035), .b(n9032) );
na02f01  g2307 ( .o(n3268), .a(n9036), .b(n9029) );
in01f01  g2308 ( .o(n9038), .a(_net_6203) );
no02f01  g2309 ( .o(n3285), .a(n9038), .b(_net_392) );
no02f01  g2310 ( .o(n9040), .a(n7094), .b(n6764) );
in01f01  g2311 ( .o(n9041), .a(net_6505) );
in01f01  g2312 ( .o(n9042_1), .a(net_6441) );
oa22f01  g2313 ( .o(n9043), .a(n6750), .b(n9042_1), .c(n6748), .d(n9041) );
in01f01  g2314 ( .o(n9044), .a(net_6537) );
in01f01  g2315 ( .o(n9045), .a(net_6473) );
oa22f01  g2316 ( .o(n9046), .a(n6755), .b(n9045), .c(n6754), .d(n9044) );
no02f01  g2317 ( .o(n9047_1), .a(n9046), .b(n9043) );
no02f01  g2318 ( .o(n9048), .a(n9047_1), .b(n6766) );
ao22f01  g2319 ( .o(n9049), .a(n6777), .b(net_6443), .c(n6776), .d(net_6507) );
ao22f01  g2320 ( .o(n9050), .a(n6780), .b(net_6475), .c(n6779_1), .d(net_6539) );
ao12f01  g2321 ( .o(n9051), .a(n6775), .b(n9050), .c(n9049) );
in01f01  g2322 ( .o(n9052_1), .a(_net_6083) );
no02f01  g2323 ( .o(n9053), .a(n6784), .b(n9052_1) );
no04f01  g2324 ( .o(n9054), .a(n9053), .b(n9051), .c(n9048), .d(n9040) );
in01f01  g2325 ( .o(n9055), .a(net_6487) );
in01f01  g2326 ( .o(n9056), .a(net_6455) );
oa22f01  g2327 ( .o(n9057_1), .a(n6790), .b(n9056), .c(n6789), .d(n9055) );
in01f01  g2328 ( .o(n9058), .a(net_6551) );
in01f01  g2329 ( .o(n9059), .a(net_6519) );
oa22f01  g2330 ( .o(n9060_1), .a(n6795), .b(n9058), .c(n6794), .d(n9059) );
no02f01  g2331 ( .o(n9061), .a(n9060_1), .b(n9057_1) );
na02f01  g2332 ( .o(n3294), .a(n9061), .b(n9054) );
in01f01  g2333 ( .o(n9063), .a(_net_7266) );
na02f01  g2334 ( .o(n9064), .a(n7242), .b(n6901) );
oa12f01  g2335 ( .o(n3308), .a(n9064), .b(n6901), .c(n9063) );
oa12f01  g2336 ( .o(n9066), .a(n7575), .b(n9004), .c(n9001) );
ao22f01  g2337 ( .o(n9067), .a(n8499_1), .b(n7593), .c(n7591_1), .d(_net_6171) );
na02f01  g2338 ( .o(n9068), .a(n7914), .b(n7588) );
in01f01  g2339 ( .o(n9069_1), .a(net_7182) );
in01f01  g2340 ( .o(n9070), .a(net_7118) );
oa22f01  g2341 ( .o(n9071), .a(n7580), .b(n9070), .c(n7577_1), .d(n9069_1) );
in01f01  g2342 ( .o(n9072), .a(net_7150) );
in01f01  g2343 ( .o(n9073), .a(net_7214) );
oa22f01  g2344 ( .o(n9074_1), .a(n7585), .b(n9072), .c(n7583), .d(n9073) );
oa12f01  g2345 ( .o(n9075), .a(n7920_1), .b(n9074_1), .c(n9071) );
na04f01  g2346 ( .o(n3313), .a(n9075), .b(n9068), .c(n9067), .d(n9066) );
ao22f01  g2347 ( .o(n9077), .a(n7288_1), .b(net_6046), .c(n7286), .d(net_285) );
ao22f01  g2348 ( .o(n9078), .a(n7298), .b(_net_7735), .c(n7291), .d(_net_7706) );
na02f01  g2349 ( .o(n9079_1), .a(n7302_1), .b(_net_129) );
na03f01  g2350 ( .o(n9080), .a(n7308), .b(net_208), .c(x1322) );
na02f01  g2351 ( .o(n9081), .a(n7296), .b(net_245) );
na03f01  g2352 ( .o(n9082_1), .a(n7308), .b(net_171), .c(n6800) );
na03f01  g2353 ( .o(n9083), .a(n9082_1), .b(n9081), .c(n9080) );
ao12f01  g2354 ( .o(n9084), .a(n9083), .b(n7306), .c(_net_6002) );
na04f01  g2355 ( .o(n3322), .a(n9084), .b(n9079_1), .c(n9078), .d(n9077) );
in01f01  g2356 ( .o(n9086_1), .a(_net_7803) );
na02f01  g2357 ( .o(n9087), .a(n6803), .b(_net_6041) );
oa12f01  g2358 ( .o(n3338), .a(n9087), .b(n6803), .c(n9086_1) );
ao22f01  g2359 ( .o(n9089), .a(n7288_1), .b(_net_6040), .c(n7286), .d(_net_279) );
ao22f01  g2360 ( .o(n9090), .a(n7298), .b(_net_7729), .c(n7291), .d(_net_7700) );
na02f01  g2361 ( .o(n9091_1), .a(n7302_1), .b(_net_123) );
na03f01  g2362 ( .o(n9092), .a(n7308), .b(net_202), .c(x1322) );
na02f01  g2363 ( .o(n9093), .a(n7296), .b(net_239) );
na03f01  g2364 ( .o(n9094), .a(n7308), .b(net_165), .c(n6800) );
na03f01  g2365 ( .o(n9095), .a(n9094), .b(n9093), .c(n9092) );
ao12f01  g2366 ( .o(n9096_1), .a(n9095), .b(n7306), .c(_net_5996) );
na04f01  g2367 ( .o(n3352), .a(n9096_1), .b(n9091_1), .c(n9090), .d(n9089) );
in01f01  g2368 ( .o(n9098), .a(_net_7583) );
no02f01  g2369 ( .o(n5628), .a(n6966), .b(n7142_1) );
na02f01  g2370 ( .o(n9100), .a(n5628), .b(n7519) );
oa12f01  g2371 ( .o(n3356), .a(n9100), .b(n7519), .c(n9098) );
in01f01  g2372 ( .o(n9102), .a(_net_7230) );
na03f01  g2373 ( .o(n9103), .a(n8302), .b(n9102), .c(_net_7229) );
oa12f01  g2374 ( .o(n9104), .a(_net_7230), .b(n8304), .c(n7579) );
na02f01  g2375 ( .o(n9105), .a(n9104), .b(n9103) );
na02f01  g2376 ( .o(n9106_1), .a(n9105), .b(_net_7233) );
in01f01  g2377 ( .o(n9107), .a(_net_7233) );
na03f01  g2378 ( .o(n9108), .a(n9104), .b(n9103), .c(n9107) );
na02f01  g2379 ( .o(n9109), .a(_net_7228), .b(n7719_1) );
na02f01  g2380 ( .o(n9110_1), .a(n7576), .b(_net_7227) );
na02f01  g2381 ( .o(n9111), .a(n9110_1), .b(n9109) );
na02f01  g2382 ( .o(n9112), .a(n9111), .b(net_7231) );
in01f01  g2383 ( .o(n9113), .a(net_7231) );
na03f01  g2384 ( .o(n9114), .a(n9110_1), .b(n9109), .c(n9113) );
ao22f01  g2385 ( .o(n9115_1), .a(n9114), .b(n9112), .c(n7720), .d(_net_7227) );
in01f01  g2386 ( .o(n9116), .a(_net_7232) );
na02f01  g2387 ( .o(n9117), .a(n8306), .b(n9116) );
na03f01  g2388 ( .o(n9118), .a(n8305), .b(n8303_1), .c(_net_7232) );
na03f01  g2389 ( .o(n9119), .a(n9118), .b(n9117), .c(n9115_1) );
ao12f01  g2390 ( .o(n3370), .a(n9119), .b(n9108), .c(n9106_1) );
in01f01  g2391 ( .o(n9121), .a(net_6907) );
in01f01  g2392 ( .o(n9122), .a(net_6843) );
oa22f01  g2393 ( .o(n9123), .a(n6810), .b(n9122), .c(n6807), .d(n9121) );
in01f01  g2394 ( .o(n9124_1), .a(net_6939) );
in01f01  g2395 ( .o(n9125), .a(net_6875) );
oa22f01  g2396 ( .o(n9126), .a(n6815), .b(n9125), .c(n6813_1), .d(n9124_1) );
no02f01  g2397 ( .o(n9127), .a(n9126), .b(n9123) );
no02f01  g2398 ( .o(n9128), .a(n9127), .b(n6824) );
in01f01  g2399 ( .o(n9129_1), .a(net_6845) );
in01f01  g2400 ( .o(n9130), .a(net_6909) );
oa22f01  g2401 ( .o(n9131), .a(n6810), .b(n9129_1), .c(n6807), .d(n9130) );
in01f01  g2402 ( .o(n9132), .a(net_6877) );
in01f01  g2403 ( .o(n9133), .a(net_6941) );
oa22f01  g2404 ( .o(n9134_1), .a(n6815), .b(n9132), .c(n6813_1), .d(n9133) );
no02f01  g2405 ( .o(n9135), .a(n9134_1), .b(n9131) );
no02f01  g2406 ( .o(n9136), .a(n9135), .b(n6826_1) );
ao22f01  g2407 ( .o(n9137), .a(n6811), .b(net_6847), .c(n6808), .d(net_6911) );
ao22f01  g2408 ( .o(n9138_1), .a(n6816), .b(net_6879), .c(n6814), .d(net_6943) );
ao12f01  g2409 ( .o(n9139), .a(n6836_1), .b(n9138_1), .c(n9137) );
in01f01  g2410 ( .o(n9140), .a(_net_6142) );
no02f01  g2411 ( .o(n9141), .a(n6844), .b(n9140) );
no04f01  g2412 ( .o(n9142), .a(n9141), .b(n9139), .c(n9136), .d(n9128) );
in01f01  g2413 ( .o(n9143_1), .a(net_6859) );
in01f01  g2414 ( .o(n9144), .a(net_6891) );
oa22f01  g2415 ( .o(n9145), .a(n6850_1), .b(n9143_1), .c(n6849), .d(n9144) );
in01f01  g2416 ( .o(n9146_1), .a(net_6955) );
in01f01  g2417 ( .o(n9147), .a(net_6923) );
oa22f01  g2418 ( .o(n9148), .a(n6855_1), .b(n9146_1), .c(n6854), .d(n9147) );
no02f01  g2419 ( .o(n9149), .a(n9148), .b(n9145) );
na02f01  g2420 ( .o(n3395), .a(n9149), .b(n9142) );
in01f01  g2421 ( .o(n9151_1), .a(_net_7619) );
na02f01  g2422 ( .o(n9152), .a(n6965), .b(net_7539) );
ao22f01  g2423 ( .o(n9153), .a(_net_292), .b(net_369), .c(_net_291), .d(net_371) );
na02f01  g2424 ( .o(n9154), .a(n9153), .b(n9152) );
na02f01  g2425 ( .o(n9155), .a(n9154), .b(n7400_1) );
oa12f01  g2426 ( .o(n3400), .a(n9155), .b(n7400_1), .c(n9151_1) );
ao22f01  g2427 ( .o(n9157), .a(n7225), .b(_net_7405), .c(n7224), .d(_net_7437) );
ao22f01  g2428 ( .o(n9158), .a(n7229), .b(_net_7501), .c(n7228), .d(_net_7469) );
na02f01  g2429 ( .o(n3422), .a(n9158), .b(n9157) );
in01f01  g2430 ( .o(n9160_1), .a(_net_7618) );
na02f01  g2431 ( .o(n9161), .a(n8000), .b(n7400_1) );
oa12f01  g2432 ( .o(n3427), .a(n9161), .b(n7400_1), .c(n9160_1) );
ao22f01  g2433 ( .o(n9163), .a(n7225), .b(_net_7419), .c(n7224), .d(_net_7451) );
ao22f01  g2434 ( .o(n9164_1), .a(n7229), .b(_net_7515), .c(n7228), .d(_net_7483) );
na02f01  g2435 ( .o(n3440), .a(n9164_1), .b(n9163) );
ao22f01  g2436 ( .o(n9166), .a(n7306), .b(_net_5984), .c(n7298), .d(_net_7720) );
ao22f01  g2437 ( .o(n9167), .a(n7288_1), .b(_net_6028), .c(n7286), .d(_net_267) );
na02f01  g2438 ( .o(n9168), .a(n7302_1), .b(_net_114) );
na03f01  g2439 ( .o(n9169_1), .a(n7308), .b(_net_193), .c(x1322) );
na02f01  g2440 ( .o(n9170), .a(n7296), .b(net_230) );
na03f01  g2441 ( .o(n9171), .a(n7308), .b(net_156), .c(n6800) );
na03f01  g2442 ( .o(n9172), .a(n9171), .b(n9170), .c(n9169_1) );
ao12f01  g2443 ( .o(n9173_1), .a(n9172), .b(n7291), .c(net_7691) );
na04f01  g2444 ( .o(n3455), .a(n9173_1), .b(n9168), .c(n9167), .d(n9166) );
in01f01  g2445 ( .o(n9175), .a(net_6431) );
in01f01  g2446 ( .o(n9176), .a(net_6495) );
oa22f01  g2447 ( .o(n9177), .a(n6750), .b(n9175), .c(n6748), .d(n9176) );
in01f01  g2448 ( .o(n9178_1), .a(net_6463) );
in01f01  g2449 ( .o(n9179), .a(net_6527) );
oa22f01  g2450 ( .o(n9180), .a(n6755), .b(n9178_1), .c(n6754), .d(n9179) );
no02f01  g2451 ( .o(n9181), .a(n9180), .b(n9177) );
no02f01  g2452 ( .o(n9182_1), .a(n9181), .b(n6764) );
no02f01  g2453 ( .o(n9183), .a(n7964), .b(n6766) );
in01f01  g2454 ( .o(n9184), .a(_net_6075) );
oa22f01  g2455 ( .o(n9185), .a(n7077_1), .b(n6775), .c(n6784), .d(n9184) );
no03f01  g2456 ( .o(n9186), .a(n9185), .b(n9183), .c(n9182_1) );
in01f01  g2457 ( .o(n9187_1), .a(net_6447) );
in01f01  g2458 ( .o(n9188), .a(net_6479) );
oa22f01  g2459 ( .o(n9189), .a(n6790), .b(n9187_1), .c(n6789), .d(n9188) );
in01f01  g2460 ( .o(n9190), .a(net_6543) );
in01f01  g2461 ( .o(n9191), .a(net_6511) );
oa22f01  g2462 ( .o(n9192_1), .a(n6795), .b(n9190), .c(n6794), .d(n9191) );
no02f01  g2463 ( .o(n9193), .a(n9192_1), .b(n9189) );
na02f01  g2464 ( .o(n3459), .a(n9193), .b(n9186) );
no02f01  g2465 ( .o(n9195), .a(n7026), .b(n6879) );
no02f01  g2466 ( .o(n9196_1), .a(_net_7382), .b(net_7378) );
no02f01  g2467 ( .o(n9197), .a(n9196_1), .b(n9195) );
in01f01  g2468 ( .o(n3464), .a(n9197) );
oa12f01  g2469 ( .o(n9199), .a(n8213), .b(n8434), .c(n8431) );
in01f01  g2470 ( .o(n9200), .a(n6826_1) );
ao22f01  g2471 ( .o(n9201_1), .a(n6811), .b(net_6833), .c(n6808), .d(net_6897) );
ao22f01  g2472 ( .o(n9202), .a(n6816), .b(net_6865), .c(n6814), .d(net_6929) );
na02f01  g2473 ( .o(n9203), .a(n9202), .b(n9201_1) );
ao22f01  g2474 ( .o(n9204), .a(n9203), .b(n9200), .c(n8211_1), .d(_net_6130) );
in01f01  g2475 ( .o(n9205), .a(n6824) );
na02f01  g2476 ( .o(n9206_1), .a(n6823), .b(n6822_1) );
no02f01  g2477 ( .o(n9207), .a(n9206_1), .b(n6818_1) );
na02f01  g2478 ( .o(n9208), .a(n9138_1), .b(n9137) );
ao22f01  g2479 ( .o(n9209), .a(n6811), .b(net_6831), .c(n6808), .d(net_6895) );
ao22f01  g2480 ( .o(n9210), .a(n6816), .b(net_6863), .c(n6814), .d(net_6927) );
na02f01  g2481 ( .o(n9211_1), .a(n9210), .b(n9209) );
ao22f01  g2482 ( .o(n9212), .a(n9211_1), .b(n9205), .c(n9208), .d(n9207) );
na03f01  g2483 ( .o(n3474), .a(n9212), .b(n9204), .c(n9199) );
in01f01  g2484 ( .o(n9214), .a(_net_6289) );
no02f01  g2485 ( .o(n3484), .a(n9214), .b(_net_392) );
in01f01  g2486 ( .o(n9216), .a(_net_7362) );
na02f01  g2487 ( .o(n9217), .a(n7242), .b(n7030) );
oa12f01  g2488 ( .o(n3489), .a(n9217), .b(n7030), .c(n9216) );
in01f01  g2489 ( .o(n9219), .a(net_6434) );
in01f01  g2490 ( .o(n9220_1), .a(net_6498) );
oa22f01  g2491 ( .o(n9221), .a(n6750), .b(n9219), .c(n6748), .d(n9220_1) );
in01f01  g2492 ( .o(n9222), .a(net_6530) );
in01f01  g2493 ( .o(n9223), .a(net_6466) );
oa22f01  g2494 ( .o(n9224), .a(n6755), .b(n9223), .c(n6754), .d(n9222) );
no02f01  g2495 ( .o(n9225_1), .a(n9224), .b(n9221) );
no02f01  g2496 ( .o(n9226), .a(n9225_1), .b(n6764) );
in01f01  g2497 ( .o(n9227), .a(net_6500) );
in01f01  g2498 ( .o(n9228_1), .a(net_6436) );
oa22f01  g2499 ( .o(n9229), .a(n6750), .b(n9228_1), .c(n6748), .d(n9227) );
in01f01  g2500 ( .o(n9230), .a(net_6468) );
in01f01  g2501 ( .o(n9231), .a(net_6532) );
oa22f01  g2502 ( .o(n9232), .a(n6755), .b(n9230), .c(n6754), .d(n9231) );
no02f01  g2503 ( .o(n9233_1), .a(n9232), .b(n9229) );
no02f01  g2504 ( .o(n9234), .a(n9233_1), .b(n6766) );
in01f01  g2505 ( .o(n9235), .a(_net_6078) );
oa22f01  g2506 ( .o(n9236), .a(n6784), .b(n9235), .c(n6775), .d(n6757) );
no03f01  g2507 ( .o(n9237), .a(n9236), .b(n9234), .c(n9226) );
in01f01  g2508 ( .o(n9238_1), .a(net_6482) );
in01f01  g2509 ( .o(n9239), .a(net_6450) );
oa22f01  g2510 ( .o(n9240), .a(n6790), .b(n9239), .c(n6789), .d(n9238_1) );
in01f01  g2511 ( .o(n9241), .a(net_6514) );
in01f01  g2512 ( .o(n9242_1), .a(net_6546) );
oa22f01  g2513 ( .o(n9243), .a(n6795), .b(n9242_1), .c(n6794), .d(n9241) );
no02f01  g2514 ( .o(n9244), .a(n9243), .b(n9240) );
na02f01  g2515 ( .o(n3507), .a(n9244), .b(n9237) );
no02f01  g2516 ( .o(n9246), .a(n6914), .b(n6912) );
na03f01  g2517 ( .o(n9247), .a(n6944), .b(n8131), .c(_net_6687) );
na02f01  g2518 ( .o(n9248), .a(n6944), .b(n8131) );
na02f01  g2519 ( .o(n9249), .a(n9248), .b(n6943_1) );
na03f01  g2520 ( .o(n9250_1), .a(n9249), .b(n9247), .c(n9246) );
na02f01  g2521 ( .o(n9251), .a(n8132), .b(_net_6687) );
na02f01  g2522 ( .o(n3516), .a(n9251), .b(n9250_1) );
in01f01  g2523 ( .o(n9253), .a(_net_5983) );
no02f01  g2524 ( .o(n3551), .a(n9253), .b(n7570) );
in01f01  g2525 ( .o(n9255), .a(_net_7703) );
na02f01  g2526 ( .o(n9256), .a(n7207_1), .b(_net_7805) );
oa12f01  g2527 ( .o(n3572), .a(n9256), .b(n7207_1), .c(n9255) );
in01f01  g2528 ( .o(n9258_1), .a(_net_6406) );
na02f01  g2529 ( .o(n9259), .a(_net_6405), .b(_net_6404) );
no02f01  g2530 ( .o(n9260), .a(n9259), .b(n9258_1) );
na02f01  g2531 ( .o(n9261), .a(n9260), .b(_net_6407) );
ao12f01  g2532 ( .o(n9262), .a(x38), .b(n9261), .c(_net_6408) );
oa12f01  g2533 ( .o(n3577), .a(n9262), .b(n9261), .c(_net_6408) );
ao22f01  g2534 ( .o(n9264), .a(n6736_1), .b(net_7641), .c(n6734), .d(net_7609) );
ao22f01  g2535 ( .o(n9265), .a(n6739), .b(net_7673), .c(n6738), .d(_net_7577) );
na02f01  g2536 ( .o(n3582), .a(n9265), .b(n9264) );
no02f01  g2537 ( .o(n9267_1), .a(_net_6557), .b(n6749_1) );
no02f01  g2538 ( .o(n9268), .a(n7765), .b(_net_6554) );
no02f01  g2539 ( .o(n9269), .a(n9268), .b(n9267_1) );
no02f01  g2540 ( .o(n9270), .a(n6747), .b(net_6556) );
no02f01  g2541 ( .o(n9271), .a(n9270), .b(n9269) );
no04f01  g2542 ( .o(n9272_1), .a(n9268), .b(n9267_1), .c(n6747), .d(net_6556) );
no02f01  g2543 ( .o(n9273), .a(n6747), .b(n7762) );
no02f01  g2544 ( .o(n9274), .a(_net_6553), .b(net_6556) );
no02f01  g2545 ( .o(n9275), .a(n9274), .b(n9273) );
oa12f01  g2546 ( .o(n9276), .a(n9275), .b(n9272_1), .c(n9271) );
no02f01  g2547 ( .o(n9277_1), .a(n9272_1), .b(n9271) );
in01f01  g2548 ( .o(n8472), .a(n9275) );
na02f01  g2549 ( .o(n9279), .a(n8472), .b(n9277_1) );
na02f01  g2550 ( .o(n3595), .a(n9279), .b(n9276) );
no02f01  g2551 ( .o(n3604), .a(n6966), .b(n7891) );
ao12f01  g2552 ( .o(n9282_1), .a(n6945), .b(n6929_1), .c(n6924_1) );
no02f01  g2553 ( .o(n9283), .a(n8885), .b(n8882_1) );
no02f01  g2554 ( .o(n9284), .a(n9283), .b(n6934_1) );
in01f01  g2555 ( .o(n9285), .a(_net_6092) );
in01f01  g2556 ( .o(n9286), .a(net_6631) );
in01f01  g2557 ( .o(n9287_1), .a(net_6567) );
oa22f01  g2558 ( .o(n9288), .a(n6922), .b(n9287_1), .c(n6919_1), .d(n9286) );
in01f01  g2559 ( .o(n9289), .a(net_6599) );
in01f01  g2560 ( .o(n9290_1), .a(net_6663) );
oa22f01  g2561 ( .o(n9291), .a(n6927), .b(n9289), .c(n6925), .d(n9290_1) );
no02f01  g2562 ( .o(n9292), .a(n9291), .b(n9288) );
oa22f01  g2563 ( .o(n9293), .a(n9292), .b(n6916), .c(n6932), .d(n9285) );
no03f01  g2564 ( .o(n9294_1), .a(n9293), .b(n9284), .c(n9282_1) );
in01f01  g2565 ( .o(n9295), .a(net_6579) );
in01f01  g2566 ( .o(n9296), .a(net_6611) );
oa22f01  g2567 ( .o(n9297), .a(n7058_1), .b(n9295), .c(n7057), .d(n9296) );
in01f01  g2568 ( .o(n9298_1), .a(net_6643) );
in01f01  g2569 ( .o(n9299), .a(net_6675) );
oa22f01  g2570 ( .o(n9300), .a(n7063), .b(n9299), .c(n7062_1), .d(n9298_1) );
no02f01  g2571 ( .o(n9301), .a(n9300), .b(n9297) );
na02f01  g2572 ( .o(n3609), .a(n9301), .b(n9294_1) );
na02f01  g2573 ( .o(n9303), .a(n7348), .b(_net_7797) );
oa12f01  g2574 ( .o(n3614), .a(n9303), .b(n7348), .c(n7538) );
in01f01  g2575 ( .o(n9305), .a(n7357) );
in01f01  g2576 ( .o(n9306), .a(_net_7783) );
in01f01  g2577 ( .o(n9307_1), .a(_net_7781) );
in01f01  g2578 ( .o(n9308), .a(_net_7782) );
na02f01  g2579 ( .o(n9309), .a(n9308), .b(n9307_1) );
no02f01  g2580 ( .o(n9310), .a(n9309), .b(n9306) );
no02f01  g2581 ( .o(n9311), .a(n9310), .b(_net_113) );
ao12f01  g2582 ( .o(n9312_1), .a(_net_7781), .b(n9311), .c(n9305) );
oa12f01  g2583 ( .o(n9313), .a(n7353), .b(n9310), .c(n7357) );
ao12f01  g2584 ( .o(n3628), .a(n9312_1), .b(n9313), .c(_net_7781) );
in01f01  g2585 ( .o(n9315), .a(_net_7665) );
na02f01  g2586 ( .o(n9316_1), .a(n6965), .b(net_371) );
ao22f01  g2587 ( .o(n9317), .a(_net_292), .b(net_383), .c(_net_291), .d(net_385) );
na02f01  g2588 ( .o(n9318), .a(n9317), .b(n9316_1) );
na02f01  g2589 ( .o(n9319), .a(n9318), .b(n7446_1) );
oa12f01  g2590 ( .o(n3633), .a(n9319), .b(n7446_1), .c(n9315) );
na02f01  g2591 ( .o(n9321_1), .a(n7306), .b(_net_6020) );
na02f01  g2592 ( .o(n9322), .a(n7293), .b(net_220) );
ao22f01  g2593 ( .o(n9323), .a(n7297_1), .b(net_183), .c(n7296), .d(net_257) );
ao22f01  g2594 ( .o(n9324), .a(n7298), .b(_net_7747), .c(n7291), .d(_net_7718) );
na04f01  g2595 ( .o(n3647), .a(n9324), .b(n9323), .c(n9322), .d(n9321_1) );
in01f01  g2596 ( .o(n9326_1), .a(_net_7424) );
na02f01  g2597 ( .o(n9327), .a(n1993), .b(n7550) );
oa12f01  g2598 ( .o(n3666), .a(n9327), .b(n7550), .c(n9326_1) );
in01f01  g2599 ( .o(n9329), .a(net_6014) );
in01f01  g2600 ( .o(n9330_1), .a(_net_7728) );
ao12f01  g2601 ( .o(n3675), .a(n7343), .b(n9330_1), .c(n9329) );
in01f01  g2602 ( .o(n9332), .a(_net_5854) );
in01f01  g2603 ( .o(n9333), .a(x940) );
in01f01  g2604 ( .o(n9334), .a(_net_6032) );
no02f01  g2605 ( .o(n9335_1), .a(_net_6033), .b(n9334) );
na02f01  g2606 ( .o(n9336), .a(_net_6028), .b(_net_6034) );
ao12f01  g2607 ( .o(n9337), .a(n9336), .b(n7316_1), .c(_net_5978) );
na02f01  g2608 ( .o(n9338), .a(n9337), .b(n9335_1) );
in01f01  g2609 ( .o(n9339_1), .a(_net_6033) );
in01f01  g2610 ( .o(n9340), .a(n9336) );
na03f01  g2611 ( .o(n9341), .a(n7316_1), .b(_net_5978), .c(_net_5977) );
na04f01  g2612 ( .o(n9342), .a(n9341), .b(n9340), .c(n9339_1), .d(n9334) );
oa12f01  g2613 ( .o(n9343_1), .a(n7316_1), .b(_net_5978), .c(_net_5977) );
na04f01  g2614 ( .o(n9344), .a(n9343_1), .b(n9340), .c(_net_6033), .d(n9334) );
no02f01  g2615 ( .o(n9345), .a(n9339_1), .b(n9334) );
na03f01  g2616 ( .o(n9346), .a(n9345), .b(n9340), .c(_net_5976) );
na04f01  g2617 ( .o(n9347), .a(n9346), .b(n9344), .c(n9342), .d(n9338) );
na03f01  g2618 ( .o(n9348_1), .a(n9347), .b(net_7776), .c(n9333) );
oa12f01  g2619 ( .o(n3684), .a(n9348_1), .b(n9332), .c(x940) );
in01f01  g2620 ( .o(n9350), .a(_net_7250) );
na02f01  g2621 ( .o(n9351), .a(n8731), .b(n6901) );
oa12f01  g2622 ( .o(n3693), .a(n9351), .b(n6901), .c(n9350) );
in01f01  g2623 ( .o(n9353), .a(_net_5853) );
in01f01  g2624 ( .o(n9354), .a(x906) );
na03f01  g2625 ( .o(n9355), .a(n8707), .b(net_7777), .c(n9354) );
oa12f01  g2626 ( .o(n3698), .a(n9355), .b(n9353), .c(x906) );
na02f01  g2627 ( .o(n9357), .a(_net_6017), .b(_net_6023) );
ao12f01  g2628 ( .o(n9358), .a(n9357), .b(_net_5974), .c(n7687) );
na02f01  g2629 ( .o(n9359), .a(n9358), .b(n7695_1) );
in01f01  g2630 ( .o(n9360), .a(n9357) );
na04f01  g2631 ( .o(n9361_1), .a(n9360), .b(n7697), .c(n7692), .d(n7689) );
na04f01  g2632 ( .o(n9362), .a(n9360), .b(n7688), .c(n7692), .d(_net_6022) );
na03f01  g2633 ( .o(n9363), .a(n9360), .b(n7693), .c(_net_5972) );
na04f01  g2634 ( .o(n9364), .a(n9363), .b(n9362), .c(n9361_1), .d(n9359) );
in01f01  g2635 ( .o(n9365_1), .a(n9364) );
no02f01  g2636 ( .o(n3711), .a(n9365_1), .b(x977) );
in01f01  g2637 ( .o(n9367), .a(_net_7444) );
na02f01  g2638 ( .o(n9368), .a(n7553_1), .b(n7197) );
oa12f01  g2639 ( .o(n3737), .a(n9368), .b(n7197), .c(n9367) );
in01f01  g2640 ( .o(n9370_1), .a(_net_7598) );
na02f01  g2641 ( .o(n9371), .a(n6965), .b(net_7550) );
ao22f01  g2642 ( .o(n9372), .a(_net_292), .b(net_380), .c(_net_291), .d(net_382) );
na02f01  g2643 ( .o(n9373_1), .a(n9372), .b(n9371) );
na02f01  g2644 ( .o(n9374), .a(n9373_1), .b(n6968) );
oa12f01  g2645 ( .o(n3742), .a(n9374), .b(n6968), .c(n9370_1) );
in01f01  g2646 ( .o(n9376), .a(_net_290) );
na02f01  g2647 ( .o(n9377_1), .a(n7440), .b(_net_7810) );
oa12f01  g2648 ( .o(n3765), .a(n9377_1), .b(n7440), .c(n9376) );
in01f01  g2649 ( .o(n9379), .a(_net_7626) );
na02f01  g2650 ( .o(n9380), .a(n7707), .b(n7400_1) );
oa12f01  g2651 ( .o(n3782), .a(n9380), .b(n7400_1), .c(n9379) );
no02f01  g2652 ( .o(n9382), .a(n6978), .b(n6976) );
na03f01  g2653 ( .o(n9383), .a(n7011), .b(n7219), .c(_net_7092) );
na02f01  g2654 ( .o(n9384), .a(n7011), .b(n7219) );
na02f01  g2655 ( .o(n9385_1), .a(n9384), .b(n7010) );
na03f01  g2656 ( .o(n9386), .a(n9385_1), .b(n9383), .c(n9382) );
na02f01  g2657 ( .o(n9387), .a(n7220), .b(_net_7092) );
na02f01  g2658 ( .o(n3787), .a(n9387), .b(n9386) );
no02f01  g2659 ( .o(n9389), .a(_net_7784), .b(_net_7785) );
no03f01  g2660 ( .o(n3796), .a(n9389), .b(n7362), .c(n7358) );
ao22f01  g2661 ( .o(n9391), .a(n6877), .b(_net_7276), .c(n6876_1), .d(net_7340) );
ao22f01  g2662 ( .o(n9392), .a(n6881_1), .b(net_7308), .c(n6880), .d(net_7372) );
na02f01  g2663 ( .o(n3813), .a(n9392), .b(n9391) );
no03f01  g2664 ( .o(n9394), .a(n7850), .b(n7415), .c(_net_282) );
no02f01  g2665 ( .o(n9395), .a(n7850), .b(n7410) );
ao22f01  g2666 ( .o(n9396), .a(n9395), .b(n7416), .c(n9394), .d(n7420) );
ao12f01  g2667 ( .o(n9397), .a(n7850), .b(_net_229), .c(n7410) );
no03f01  g2668 ( .o(n9398_1), .a(n7850), .b(_net_283), .c(_net_282) );
ao22f01  g2669 ( .o(n9399), .a(n9398_1), .b(n7418), .c(n9397), .d(n7409) );
na02f01  g2670 ( .o(n3827), .a(n9399), .b(n9396) );
in01f01  g2671 ( .o(n9401), .a(_net_6419) );
in01f01  g2672 ( .o(n9402_1), .a(_net_6401) );
in01f01  g2673 ( .o(n9403), .a(_net_6422) );
in01f01  g2674 ( .o(n9404), .a(_net_6423) );
in01f01  g2675 ( .o(n9405_1), .a(_net_6418) );
no04f01  g2676 ( .o(n9406), .a(_net_6421), .b(n9405_1), .c(n9404), .d(_net_6420) );
na03f01  g2677 ( .o(n9407), .a(n9406), .b(n9403), .c(n9401) );
in01f01  g2678 ( .o(n7691), .a(n9407) );
na02f01  g2679 ( .o(n9409), .a(n7691), .b(n9402_1) );
no02f01  g2680 ( .o(n9410_1), .a(n7691), .b(_net_6401) );
in01f01  g2681 ( .o(n9411), .a(n9410_1) );
na02f01  g2682 ( .o(n9412), .a(_net_6418), .b(_net_6419) );
na02f01  g2683 ( .o(n9413), .a(n9405_1), .b(n9401) );
na02f01  g2684 ( .o(n9414), .a(n9413), .b(n9412) );
oa22f01  g2685 ( .o(n3836), .a(n9414), .b(n9411), .c(n9409), .d(n9401) );
in01f01  g2686 ( .o(n9416), .a(_net_7652) );
na02f01  g2687 ( .o(n9417), .a(n8426_1), .b(n7446_1) );
oa12f01  g2688 ( .o(n3841), .a(n9417), .b(n7446_1), .c(n9416) );
no02f01  g2689 ( .o(n9419), .a(n8790), .b(n7012) );
no02f01  g2690 ( .o(n9420_1), .a(n8602_1), .b(n6997) );
in01f01  g2691 ( .o(n9421), .a(_net_6158) );
oa22f01  g2692 ( .o(n9422), .a(n8610), .b(n6980), .c(n6995_1), .d(n9421) );
no03f01  g2693 ( .o(n9423), .a(n9422), .b(n9420_1), .c(n9419) );
in01f01  g2694 ( .o(n9424), .a(net_7022) );
in01f01  g2695 ( .o(n9425_1), .a(net_6990) );
oa22f01  g2696 ( .o(n9426), .a(n8075_1), .b(n9425_1), .c(n8074), .d(n9424) );
in01f01  g2697 ( .o(n9427), .a(net_7054) );
in01f01  g2698 ( .o(n9428_1), .a(net_7086) );
oa22f01  g2699 ( .o(n9429), .a(n8080_1), .b(n9428_1), .c(n8079), .d(n9427) );
no02f01  g2700 ( .o(n9430), .a(n9429), .b(n9426) );
na02f01  g2701 ( .o(n3846), .a(n9430), .b(n9423) );
in01f01  g2702 ( .o(n9432), .a(_net_7290) );
na02f01  g2703 ( .o(n9433), .a(n7393), .b(n7180) );
oa12f01  g2704 ( .o(n3859), .a(n9433), .b(n7180), .c(n9432) );
no02f01  g2705 ( .o(n9435), .a(n7027_1), .b(n6875) );
no02f01  g2706 ( .o(n9436_1), .a(_net_7383), .b(_net_7379) );
no02f01  g2707 ( .o(n9437), .a(n9436_1), .b(n9435) );
in01f01  g2708 ( .o(n9438), .a(n9437) );
na02f01  g2709 ( .o(n9439), .a(n9438), .b(n3464) );
in01f01  g2710 ( .o(n9440), .a(_net_7380) );
in01f01  g2711 ( .o(n9441_1), .a(_net_7384) );
no02f01  g2712 ( .o(n9442), .a(n9441_1), .b(n9440) );
no02f01  g2713 ( .o(n9443), .a(_net_7384), .b(_net_7380) );
no02f01  g2714 ( .o(n9444), .a(n9443), .b(n9442) );
no04f01  g2715 ( .o(n3872), .a(n9444), .b(n9439), .c(n6899_1), .d(_net_7381) );
na02f01  g2716 ( .o(n9446), .a(n8034), .b(_net_6065) );
na02f01  g2717 ( .o(n9447), .a(n8037), .b(n8028_1) );
na02f01  g2718 ( .o(n3877), .a(n9447), .b(n9446) );
in01f01  g2719 ( .o(n9449_1), .a(_net_7574) );
na02f01  g2720 ( .o(n9450), .a(n2850), .b(n7519) );
oa12f01  g2721 ( .o(n3886), .a(n9450), .b(n7519), .c(n9449_1) );
in01f01  g2722 ( .o(n9452), .a(_net_123) );
na02f01  g2723 ( .o(n9453), .a(_net_154), .b(net_319) );
oa12f01  g2724 ( .o(n3891), .a(n9453), .b(n9452), .c(_net_154) );
ao22f01  g2725 ( .o(n9455), .a(n7225), .b(_net_7431), .c(n7224), .d(net_7463) );
ao22f01  g2726 ( .o(n9456), .a(n7229), .b(net_7527), .c(n7228), .d(net_7495) );
na02f01  g2727 ( .o(n3908), .a(n9456), .b(n9455) );
in01f01  g2728 ( .o(n9458), .a(_net_7270) );
na02f01  g2729 ( .o(n9459_1), .a(n1029), .b(n6901) );
oa12f01  g2730 ( .o(n3913), .a(n9459_1), .b(n6901), .c(n9458) );
in01f01  g2731 ( .o(n9461), .a(net_6766) );
in01f01  g2732 ( .o(n9462_1), .a(net_6702) );
oa22f01  g2733 ( .o(n9463), .a(n7129), .b(n9462_1), .c(n7126), .d(n9461) );
in01f01  g2734 ( .o(n9464), .a(net_6734) );
in01f01  g2735 ( .o(n9465), .a(net_6798) );
oa22f01  g2736 ( .o(n9466), .a(n7134), .b(n9464), .c(n7132), .d(n9465) );
no02f01  g2737 ( .o(n9467_1), .a(n9466), .b(n9463) );
no02f01  g2738 ( .o(n9468), .a(n9467_1), .b(n7468_1) );
no02f01  g2739 ( .o(n9469), .a(n8557_1), .b(n7470) );
in01f01  g2740 ( .o(n9470_1), .a(_net_6116) );
oa22f01  g2741 ( .o(n9471), .a(n7465), .b(n7123), .c(n7118), .d(n9470_1) );
no03f01  g2742 ( .o(n9472), .a(n9471), .b(n9469), .c(n9468) );
in01f01  g2743 ( .o(n9473), .a(net_6718) );
in01f01  g2744 ( .o(n9474), .a(net_6750) );
oa22f01  g2745 ( .o(n9475_1), .a(n7492_1), .b(n9473), .c(n7491), .d(n9474) );
in01f01  g2746 ( .o(n9476), .a(net_6814) );
in01f01  g2747 ( .o(n9477), .a(net_6782) );
oa22f01  g2748 ( .o(n9478_1), .a(n7497), .b(n9476), .c(n7496_1), .d(n9477) );
no02f01  g2749 ( .o(n9479), .a(n9478_1), .b(n9475_1) );
na02f01  g2750 ( .o(n3922), .a(n9479), .b(n9472) );
in01f01  g2751 ( .o(n9481), .a(_net_7563) );
na02f01  g2752 ( .o(n9482), .a(n7519), .b(n6971) );
oa12f01  g2753 ( .o(n3927), .a(n9482), .b(n7519), .c(n9481) );
in01f01  g2754 ( .o(n9484), .a(_net_7418) );
na02f01  g2755 ( .o(n9485), .a(n6866), .b(net_351) );
ao22f01  g2756 ( .o(n9486), .a(_net_281), .b(net_363), .c(_net_280), .d(net_365) );
na02f01  g2757 ( .o(n9487_1), .a(n9486), .b(n9485) );
na02f01  g2758 ( .o(n9488), .a(n9487_1), .b(n7550) );
oa12f01  g2759 ( .o(n3932), .a(n9488), .b(n7550), .c(n9484) );
in01f01  g2760 ( .o(n9490), .a(_net_7591) );
na02f01  g2761 ( .o(n9491), .a(n6965), .b(net_7543) );
ao22f01  g2762 ( .o(n9492_1), .a(_net_292), .b(net_373), .c(_net_291), .d(net_375) );
na02f01  g2763 ( .o(n9493), .a(n9492_1), .b(n9491) );
na02f01  g2764 ( .o(n9494), .a(n9493), .b(n6968) );
oa12f01  g2765 ( .o(n3941), .a(n9494), .b(n6968), .c(n9490) );
in01f01  g2766 ( .o(n9496), .a(_net_7510) );
na02f01  g2767 ( .o(n9497_1), .a(n8994), .b(n7626_1) );
oa12f01  g2768 ( .o(n3967), .a(n9497_1), .b(n7626_1), .c(n9496) );
in01f01  g2769 ( .o(n9499), .a(_net_6201) );
no02f01  g2770 ( .o(n3976), .a(n9499), .b(_net_392) );
ao12f01  g2771 ( .o(n9501), .a(n7468_1), .b(n8156_1), .c(n8155) );
no02f01  g2772 ( .o(n9502_1), .a(n8979), .b(n8976_1) );
no02f01  g2773 ( .o(n9503), .a(n9502_1), .b(n7470) );
in01f01  g2774 ( .o(n9504), .a(_net_6112) );
oa22f01  g2775 ( .o(n9505), .a(n9467_1), .b(n7123), .c(n7118), .d(n9504) );
no03f01  g2776 ( .o(n9506), .a(n9505), .b(n9503), .c(n9501) );
in01f01  g2777 ( .o(n9507_1), .a(net_6746) );
in01f01  g2778 ( .o(n9508), .a(net_6714) );
oa22f01  g2779 ( .o(n9509), .a(n7492_1), .b(n9508), .c(n7491), .d(n9507_1) );
in01f01  g2780 ( .o(n9510), .a(net_6810) );
in01f01  g2781 ( .o(n9511), .a(net_6778) );
oa22f01  g2782 ( .o(n9512_1), .a(n7497), .b(n9510), .c(n7496_1), .d(n9511) );
no02f01  g2783 ( .o(n9513), .a(n9512_1), .b(n9509) );
na02f01  g2784 ( .o(n3981), .a(n9513), .b(n9506) );
in01f01  g2785 ( .o(n9515), .a(_net_7095) );
na03f01  g2786 ( .o(n9516), .a(n7210), .b(n9515), .c(_net_7094) );
oa12f01  g2787 ( .o(n9517_1), .a(_net_7095), .b(n7212_1), .c(n6986_1) );
na02f01  g2788 ( .o(n9518), .a(n9517_1), .b(n9516) );
na02f01  g2789 ( .o(n9519), .a(n9518), .b(n7215) );
no02f01  g2790 ( .o(n9520_1), .a(n6991), .b(n9515) );
no02f01  g2791 ( .o(n9521), .a(n7002), .b(_net_7095) );
no02f01  g2792 ( .o(n9522), .a(n9521), .b(n9520_1) );
ao22f01  g2793 ( .o(n9523), .a(n9522), .b(n7218), .c(n7220), .d(_net_7095) );
na02f01  g2794 ( .o(n3998), .a(n9523), .b(n9519) );
in01f01  g2795 ( .o(n9525_1), .a(_net_7733) );
in01f01  g2796 ( .o(n9526), .a(_net_6027) );
ao12f01  g2797 ( .o(n4016), .a(n7343), .b(n9526), .c(n9525_1) );
in01f01  g2798 ( .o(n9528_1), .a(_net_7601) );
na02f01  g2799 ( .o(n9529), .a(n9318), .b(n6968) );
oa12f01  g2800 ( .o(n4029), .a(n9529), .b(n6968), .c(n9528_1) );
in01f01  g2801 ( .o(n9531), .a(_net_7633) );
na02f01  g2802 ( .o(n9532), .a(n9318), .b(n7400_1) );
oa12f01  g2803 ( .o(n4042), .a(n9532), .b(n7400_1), .c(n9531) );
in01f01  g2804 ( .o(n9534), .a(_net_7329) );
na02f01  g2805 ( .o(n9535), .a(n6898), .b(net_7249) );
ao22f01  g2806 ( .o(n9536), .a(net_341), .b(_net_270), .c(_net_269), .d(net_343) );
na02f01  g2807 ( .o(n9537_1), .a(n9536), .b(n9535) );
na02f01  g2808 ( .o(n9538), .a(n9537_1), .b(n7150) );
oa12f01  g2809 ( .o(n4063), .a(n9538), .b(n7150), .c(n9534) );
in01f01  g2810 ( .o(n9540), .a(_net_294) );
na02f01  g2811 ( .o(n9541_1), .a(n7440), .b(_net_7814) );
oa12f01  g2812 ( .o(n4084), .a(n9541_1), .b(n7440), .c(n9540) );
no02f01  g2813 ( .o(n9543), .a(n9261), .b(n8178) );
na03f01  g2814 ( .o(n9544), .a(n9543), .b(_net_6410), .c(n8084) );
in01f01  g2815 ( .o(n9545), .a(_net_6410) );
in01f01  g2816 ( .o(n9546_1), .a(n9543) );
oa12f01  g2817 ( .o(n9547), .a(_net_6411), .b(n9546_1), .c(n9545) );
na03f01  g2818 ( .o(n4089), .a(n9547), .b(n9544), .c(n6910_1) );
in01f01  g2819 ( .o(n9549_1), .a(_net_7404) );
na02f01  g2820 ( .o(n9550), .a(n7952), .b(n7550) );
oa12f01  g2821 ( .o(n4094), .a(n9550), .b(n7550), .c(n9549_1) );
in01f01  g2822 ( .o(n9552), .a(_net_7719) );
na02f01  g2823 ( .o(n9553), .a(n7207_1), .b(_net_7821) );
oa12f01  g2824 ( .o(n4107), .a(n9553), .b(n7207_1), .c(n9552) );
in01f01  g2825 ( .o(n9555), .a(_net_7364) );
na02f01  g2826 ( .o(n9556), .a(n7256_1), .b(n7030) );
oa12f01  g2827 ( .o(n4116), .a(n9556), .b(n7030), .c(n9555) );
in01f01  g2828 ( .o(n9558), .a(_net_276) );
na02f01  g2829 ( .o(n9559_1), .a(_net_190), .b(_net_188) );
na02f01  g2830 ( .o(n4121), .a(n9559_1), .b(n9558) );
no02f01  g2831 ( .o(n9561), .a(n7572_1), .b(n7570) );
na03f01  g2832 ( .o(n9562), .a(n7720), .b(n8311_1), .c(_net_7227) );
na02f01  g2833 ( .o(n9563), .a(n7720), .b(n8311_1) );
na02f01  g2834 ( .o(n9564_1), .a(n9563), .b(n7719_1) );
na03f01  g2835 ( .o(n9565), .a(n9564_1), .b(n9562), .c(n9561) );
na02f01  g2836 ( .o(n9566), .a(n8312), .b(_net_7227) );
na02f01  g2837 ( .o(n4126), .a(n9566), .b(n9565) );
in01f01  g2838 ( .o(n9568), .a(n3551) );
no02f01  g2839 ( .o(n9569_1), .a(_net_7232), .b(n9113) );
no02f01  g2840 ( .o(n9570), .a(n9116), .b(net_7231) );
no02f01  g2841 ( .o(n9571), .a(n9570), .b(n9569_1) );
na02f01  g2842 ( .o(n9572), .a(n9253), .b(_net_6039) );
oa22f01  g2843 ( .o(n4135), .a(n9572), .b(n9116), .c(n9571), .d(n9568) );
in01f01  g2844 ( .o(n9574_1), .a(_net_7347) );
na02f01  g2845 ( .o(n9575), .a(n7659), .b(n7030) );
oa12f01  g2846 ( .o(n4140), .a(n9575), .b(n7030), .c(n9574_1) );
in01f01  g2847 ( .o(n9577), .a(_net_7437) );
na02f01  g2848 ( .o(n9578), .a(n8817), .b(n7197) );
oa12f01  g2849 ( .o(n4166), .a(n9578), .b(n7197), .c(n9577) );
no02f01  g2850 ( .o(n4171), .a(_net_7784), .b(_net_113) );
ao22f01  g2851 ( .o(n9581), .a(n6738), .b(_net_7556), .c(n6736_1), .d(_net_7620) );
ao22f01  g2852 ( .o(n9582), .a(n6739), .b(_net_7652), .c(n6734), .d(_net_7588) );
na02f01  g2853 ( .o(n4181), .a(n9582), .b(n9581) );
in01f01  g2854 ( .o(n9584), .a(_net_7321) );
na02f01  g2855 ( .o(n9585), .a(n6898), .b(net_7241) );
ao22f01  g2856 ( .o(n9586), .a(net_333), .b(_net_270), .c(net_335), .d(_net_269) );
na02f01  g2857 ( .o(n9587), .a(n9586), .b(n9585) );
na02f01  g2858 ( .o(n9588_1), .a(n9587), .b(n7150) );
oa12f01  g2859 ( .o(n4186), .a(n9588_1), .b(n7150), .c(n9584) );
in01f01  g2860 ( .o(n9590), .a(_net_277) );
in01f01  g2861 ( .o(n9591), .a(_net_189) );
in01f01  g2862 ( .o(n9592_1), .a(n6897) );
oa12f01  g2863 ( .o(n4203), .a(n9590), .b(n9592_1), .c(n9591) );
ao22f01  g2864 ( .o(n9594), .a(n7225), .b(_net_7414), .c(n7224), .d(_net_7446) );
ao22f01  g2865 ( .o(n9595), .a(n7229), .b(_net_7510), .c(n7228), .d(_net_7478) );
na02f01  g2866 ( .o(n4212), .a(n9595), .b(n9594) );
in01f01  g2867 ( .o(n9597_1), .a(_net_7630) );
na02f01  g2868 ( .o(n9598), .a(n9373_1), .b(n7400_1) );
oa12f01  g2869 ( .o(n4217), .a(n9598), .b(n7400_1), .c(n9597_1) );
in01f01  g2870 ( .o(n9600), .a(_net_6825) );
no02f01  g2871 ( .o(n9601), .a(n7125_1), .b(n7466) );
na03f01  g2872 ( .o(n9602_1), .a(n9601), .b(_net_6824), .c(n9600) );
in01f01  g2873 ( .o(n9603), .a(n9601) );
oa12f01  g2874 ( .o(n9604), .a(_net_6825), .b(n9603), .c(n7128_1) );
na02f01  g2875 ( .o(n9605), .a(n9604), .b(n9602_1) );
na02f01  g2876 ( .o(n9606_1), .a(n9605), .b(_net_6828) );
in01f01  g2877 ( .o(n9607), .a(_net_6828) );
na03f01  g2878 ( .o(n9608), .a(n9604), .b(n9602_1), .c(n9607) );
na02f01  g2879 ( .o(n9609), .a(_net_6823), .b(n7466) );
na02f01  g2880 ( .o(n9610), .a(n7125_1), .b(_net_6822) );
na02f01  g2881 ( .o(n9611_1), .a(n9610), .b(n9609) );
na02f01  g2882 ( .o(n9612), .a(n9611_1), .b(net_6826) );
na03f01  g2883 ( .o(n9613), .a(n9610), .b(n9609), .c(n8220_1) );
ao22f01  g2884 ( .o(n9614), .a(n9613), .b(n9612), .c(n7467), .d(_net_6822) );
na02f01  g2885 ( .o(n9615), .a(n9601), .b(n7128_1) );
na02f01  g2886 ( .o(n9616_1), .a(n9603), .b(_net_6824) );
na02f01  g2887 ( .o(n9617), .a(n9616_1), .b(n9615) );
na02f01  g2888 ( .o(n9618), .a(n9617), .b(n8219) );
na03f01  g2889 ( .o(n9619), .a(n9616_1), .b(n9615), .c(_net_6827) );
na03f01  g2890 ( .o(n9620_1), .a(n9619), .b(n9618), .c(n9614) );
ao12f01  g2891 ( .o(n4226), .a(n9620_1), .b(n9608), .c(n9606_1) );
in01f01  g2892 ( .o(n9622), .a(_net_7635) );
na02f01  g2893 ( .o(n9623), .a(n7400_1), .b(n7144) );
oa12f01  g2894 ( .o(n4240), .a(n9623), .b(n7400_1), .c(n9622) );
ao12f01  g2895 ( .o(n9625), .a(n7012), .b(n7004), .c(n7001) );
no02f01  g2896 ( .o(n9626), .a(n6993), .b(n6988) );
no02f01  g2897 ( .o(n9627), .a(n6997), .b(n9626) );
in01f01  g2898 ( .o(n9628_1), .a(_net_6152) );
oa22f01  g2899 ( .o(n9629), .a(n8782), .b(n6980), .c(n6995_1), .d(n9628_1) );
no03f01  g2900 ( .o(n9630), .a(n9629), .b(n9627), .c(n9625) );
in01f01  g2901 ( .o(n9631), .a(net_7016) );
in01f01  g2902 ( .o(n9632), .a(net_6984) );
oa22f01  g2903 ( .o(n9633_1), .a(n8075_1), .b(n9632), .c(n8074), .d(n9631) );
in01f01  g2904 ( .o(n9634), .a(net_7048) );
in01f01  g2905 ( .o(n9635), .a(net_7080) );
oa22f01  g2906 ( .o(n9636), .a(n8080_1), .b(n9635), .c(n8079), .d(n9634) );
no02f01  g2907 ( .o(n9637), .a(n9636), .b(n9633_1) );
na02f01  g2908 ( .o(n4249), .a(n9637), .b(n9630) );
no02f01  g2909 ( .o(n9639), .a(n7576), .b(n9113) );
no02f01  g2910 ( .o(n9640), .a(_net_7228), .b(net_7231) );
no02f01  g2911 ( .o(n9641), .a(n9640), .b(n9639) );
in01f01  g2912 ( .o(n4276), .a(n9641) );
no02f01  g2913 ( .o(n9643), .a(n7194_1), .b(net_7529) );
in01f01  g2914 ( .o(n9644), .a(n9643) );
no02f01  g2915 ( .o(n9645), .a(n9644), .b(n8923) );
no02f01  g2916 ( .o(n9646), .a(n9643), .b(n8924) );
oa12f01  g2917 ( .o(n9647_1), .a(n8919), .b(n9646), .c(n9645) );
no02f01  g2918 ( .o(n9648), .a(n9646), .b(n9645) );
na02f01  g2919 ( .o(n9649), .a(n9648), .b(n8850) );
na02f01  g2920 ( .o(n4289), .a(n9649), .b(n9647_1) );
in01f01  g2921 ( .o(n9651_1), .a(_net_7318) );
na02f01  g2922 ( .o(n9652), .a(n8960), .b(n7150) );
oa12f01  g2923 ( .o(n4294), .a(n9652), .b(n7150), .c(n9651_1) );
na02f01  g2924 ( .o(n9654), .a(n9203), .b(n8213) );
ao22f01  g2925 ( .o(n9655_1), .a(n9211_1), .b(n9200), .c(n8211_1), .d(_net_6128) );
ao22f01  g2926 ( .o(n9656), .a(n6811), .b(net_6829), .c(n6808), .d(net_6893) );
ao22f01  g2927 ( .o(n9657), .a(n6816), .b(net_6861), .c(n6814), .d(net_6925) );
na02f01  g2928 ( .o(n9658), .a(n9657), .b(n9656) );
na02f01  g2929 ( .o(n9659), .a(n9658), .b(n9205) );
oa12f01  g2930 ( .o(n9660_1), .a(n9207), .b(n9134_1), .c(n9131) );
na04f01  g2931 ( .o(n4299), .a(n9660_1), .b(n9659), .c(n9655_1), .d(n9654) );
no04f01  g2932 ( .o(n4304), .a(n7338), .b(n7107_1), .c(n7106), .d(x1155) );
in01f01  g2933 ( .o(n9663), .a(_net_6421) );
na03f01  g2934 ( .o(n9664_1), .a(_net_6418), .b(_net_6420), .c(_net_6419) );
no02f01  g2935 ( .o(n9665), .a(n9664_1), .b(n9663) );
no02f01  g2936 ( .o(n9666), .a(n9665), .b(_net_6422) );
na02f01  g2937 ( .o(n9667), .a(n9665), .b(_net_6422) );
na02f01  g2938 ( .o(n9668_1), .a(n9667), .b(n9410_1) );
oa22f01  g2939 ( .o(n4313), .a(n9668_1), .b(n9666), .c(n9409), .d(n9403) );
na03f01  g2940 ( .o(n9670), .a(n8089), .b(n8084), .c(_net_6408) );
in01f01  g2941 ( .o(n9671), .a(_net_6409) );
na02f01  g2942 ( .o(n9672), .a(n9671), .b(n9545) );
no04f01  g2943 ( .o(n4322), .a(n9672), .b(n9670), .c(_net_6407), .d(_net_6406) );
in01f01  g2944 ( .o(n9674), .a(_net_7505) );
na02f01  g2945 ( .o(n9675), .a(n7626_1), .b(n7200) );
oa12f01  g2946 ( .o(n4348), .a(n9675), .b(n7626_1), .c(n9674) );
in01f01  g2947 ( .o(n9677), .a(_net_6009) );
na02f01  g2948 ( .o(n9678_1), .a(n7348), .b(_net_7812) );
oa12f01  g2949 ( .o(n4357), .a(n9678_1), .b(n7348), .c(n9677) );
in01f01  g2950 ( .o(n9680), .a(_net_7278) );
na02f01  g2951 ( .o(n9681), .a(n576), .b(n6901) );
oa12f01  g2952 ( .o(n4379), .a(n9681), .b(n6901), .c(n9680) );
in01f01  g2953 ( .o(n9683_1), .a(_net_7301) );
in01f01  g2954 ( .o(n9684), .a(net_333) );
oa22f01  g2955 ( .o(n9685), .a(n6899_1), .b(n9684), .c(n7253), .d(n7514) );
na02f01  g2956 ( .o(n9686), .a(n9685), .b(n7180) );
oa12f01  g2957 ( .o(n4392), .a(n9686), .b(n7180), .c(n9683_1) );
in01f01  g2958 ( .o(n9688), .a(_net_7718) );
na02f01  g2959 ( .o(n9689), .a(n7207_1), .b(_net_7820) );
oa12f01  g2960 ( .o(n4414), .a(n9689), .b(n7207_1), .c(n9688) );
in01f01  g2961 ( .o(n9691), .a(net_7807) );
na02f01  g2962 ( .o(n9692_1), .a(n6803), .b(_net_6045) );
oa12f01  g2963 ( .o(n4424), .a(n9692_1), .b(n6803), .c(n9691) );
in01f01  g2964 ( .o(n9694), .a(_net_7332) );
na02f01  g2965 ( .o(n9695_1), .a(n7256_1), .b(n7150) );
oa12f01  g2966 ( .o(n4433), .a(n9695_1), .b(n7150), .c(n9694) );
in01f01  g2967 ( .o(n9697), .a(_net_7403) );
na02f01  g2968 ( .o(n9698), .a(n6866), .b(net_7387) );
ao22f01  g2969 ( .o(n9699), .a(net_350), .b(_net_280), .c(net_348), .d(_net_281) );
na02f01  g2970 ( .o(n9700_1), .a(n9699), .b(n9698) );
na02f01  g2971 ( .o(n9701), .a(n9700_1), .b(n7550) );
oa12f01  g2972 ( .o(n4438), .a(n9701), .b(n7550), .c(n9697) );
in01f01  g2973 ( .o(n9703), .a(_net_6205) );
no02f01  g2974 ( .o(n4443), .a(_net_392), .b(n9703) );
oa12f01  g2975 ( .o(n9705), .a(n7284_1), .b(n7282), .c(x1322) );
no02f01  g2976 ( .o(n9706), .a(n9705), .b(n7293) );
in01f01  g2977 ( .o(n9707), .a(n7347) );
na03f01  g2978 ( .o(n9708), .a(n9707), .b(n9706), .c(_net_6023) );
na02f01  g2979 ( .o(n9709_1), .a(n7293), .b(net_223) );
ao22f01  g2980 ( .o(n9710), .a(n7297_1), .b(net_186), .c(n7296), .d(net_260) );
na03f01  g2981 ( .o(n4456), .a(n9710), .b(n9709_1), .c(n9708) );
in01f01  g2982 ( .o(n9712), .a(_net_7323) );
na02f01  g2983 ( .o(n9713), .a(n7150), .b(n7033) );
oa12f01  g2984 ( .o(n4464), .a(n9713), .b(n7150), .c(n9712) );
na02f01  g2985 ( .o(n9715), .a(n7005_1), .b(n6981) );
ao22f01  g2986 ( .o(n9716), .a(n7009_1), .b(n6998), .c(n6996), .d(_net_6148) );
ao22f01  g2987 ( .o(n9717), .a(n7000_1), .b(net_6964), .c(n6999), .d(net_7028) );
ao22f01  g2988 ( .o(n9718), .a(n7003), .b(net_6996), .c(n7002), .d(net_7060) );
na02f01  g2989 ( .o(n9719_1), .a(n9718), .b(n9717) );
na02f01  g2990 ( .o(n9720), .a(n9719_1), .b(n7013_1) );
oa12f01  g2991 ( .o(n9721), .a(n7022), .b(n8618), .c(n8615) );
na04f01  g2992 ( .o(n4482), .a(n9721), .b(n9720), .c(n9716), .d(n9715) );
in01f01  g2993 ( .o(n9723), .a(_net_6018) );
na02f01  g2994 ( .o(n9724_1), .a(n7348), .b(_net_7818) );
oa12f01  g2995 ( .o(n4491), .a(n9724_1), .b(n7348), .c(n9723) );
no02f01  g2996 ( .o(n4501), .a(net_153), .b(n8016) );
in01f01  g2997 ( .o(n9727), .a(_net_7469) );
na02f01  g2998 ( .o(n9728), .a(n8817), .b(n6869) );
oa12f01  g2999 ( .o(n4510), .a(n9728), .b(n6869), .c(n9727) );
ao12f01  g3000 ( .o(n9730), .a(n7721), .b(n8498), .c(n8497) );
no02f01  g3001 ( .o(n9731), .a(n9005_1), .b(n7592) );
in01f01  g3002 ( .o(n9732), .a(_net_6173) );
oa22f01  g3003 ( .o(n9733_1), .a(n8274), .b(n7574), .c(n7590), .d(n9732) );
no03f01  g3004 ( .o(n9734), .a(n9733_1), .b(n9731), .c(n9730) );
in01f01  g3005 ( .o(n9735), .a(net_7120) );
in01f01  g3006 ( .o(n9736), .a(net_7152) );
oa22f01  g3007 ( .o(n9737_1), .a(n7740), .b(n9735), .c(n7739), .d(n9736) );
in01f01  g3008 ( .o(n9738), .a(net_7184) );
in01f01  g3009 ( .o(n9739), .a(net_7216) );
oa22f01  g3010 ( .o(n9740), .a(n7745), .b(n9739), .c(n7744), .d(n9738) );
no02f01  g3011 ( .o(n9741), .a(n9740), .b(n9737_1) );
na02f01  g3012 ( .o(n4515), .a(n9741), .b(n9734) );
ao22f01  g3013 ( .o(n9743), .a(n6736_1), .b(_net_7632), .c(n6734), .d(_net_7600) );
ao22f01  g3014 ( .o(n9744), .a(n6739), .b(_net_7664), .c(n6738), .d(_net_7568) );
na02f01  g3015 ( .o(n4520), .a(n9744), .b(n9743) );
in01f01  g3016 ( .o(n9746_1), .a(_net_6188) );
no02f01  g3017 ( .o(n4529), .a(n9746_1), .b(_net_392) );
in01f01  g3018 ( .o(n9748), .a(_net_6194) );
no02f01  g3019 ( .o(n4534), .a(_net_392), .b(n9748) );
ao12f01  g3020 ( .o(n9750_1), .a(n7721), .b(n7907), .c(n7906_1) );
in01f01  g3021 ( .o(n9751), .a(net_7105) );
in01f01  g3022 ( .o(n9752), .a(net_7169) );
oa22f01  g3023 ( .o(n9753), .a(n7580), .b(n9751), .c(n7577_1), .d(n9752) );
in01f01  g3024 ( .o(n9754_1), .a(net_7201) );
in01f01  g3025 ( .o(n9755), .a(net_7137) );
oa22f01  g3026 ( .o(n9756), .a(n7585), .b(n9755), .c(n7583), .d(n9754_1) );
no02f01  g3027 ( .o(n9757), .a(n9756), .b(n9753) );
no02f01  g3028 ( .o(n9758_1), .a(n9757), .b(n7592) );
in01f01  g3029 ( .o(n9759), .a(_net_6172) );
in01f01  g3030 ( .o(n9760), .a(net_7171) );
in01f01  g3031 ( .o(n9761), .a(net_7107) );
oa22f01  g3032 ( .o(n9762), .a(n7580), .b(n9761), .c(n7577_1), .d(n9760) );
in01f01  g3033 ( .o(n9763_1), .a(net_7203) );
in01f01  g3034 ( .o(n9764), .a(net_7139) );
oa22f01  g3035 ( .o(n9765), .a(n7585), .b(n9764), .c(n7583), .d(n9763_1) );
no02f01  g3036 ( .o(n9766), .a(n9765), .b(n9762) );
oa22f01  g3037 ( .o(n9767), .a(n9766), .b(n7574), .c(n7590), .d(n9759) );
no03f01  g3038 ( .o(n9768_1), .a(n9767), .b(n9758_1), .c(n9750_1) );
in01f01  g3039 ( .o(n9769), .a(net_7119) );
in01f01  g3040 ( .o(n9770), .a(net_7151) );
oa22f01  g3041 ( .o(n9771), .a(n7740), .b(n9769), .c(n7739), .d(n9770) );
in01f01  g3042 ( .o(n9772), .a(net_7215) );
in01f01  g3043 ( .o(n9773_1), .a(net_7183) );
oa22f01  g3044 ( .o(n9774), .a(n7745), .b(n9772), .c(n7744), .d(n9773_1) );
no02f01  g3045 ( .o(n9775), .a(n9774), .b(n9771) );
na02f01  g3046 ( .o(n4539), .a(n9775), .b(n9768_1) );
in01f01  g3047 ( .o(n9777), .a(_net_7480) );
na02f01  g3048 ( .o(n9778_1), .a(n7638), .b(n6869) );
oa12f01  g3049 ( .o(n4544), .a(n9778_1), .b(n6869), .c(n9777) );
na02f01  g3050 ( .o(n9780), .a(n7591_1), .b(_net_6165) );
na02f01  g3051 ( .o(n9781), .a(n7596_1), .b(n7575) );
na02f01  g3052 ( .o(n4553), .a(n9781), .b(n9780) );
in01f01  g3053 ( .o(n9783_1), .a(_net_7475) );
na02f01  g3054 ( .o(n9784), .a(n6866), .b(net_7395) );
ao22f01  g3055 ( .o(n9785), .a(net_358), .b(_net_280), .c(_net_281), .d(net_356) );
na02f01  g3056 ( .o(n9786), .a(n9785), .b(n9784) );
na02f01  g3057 ( .o(n9787_1), .a(n9786), .b(n6869) );
oa12f01  g3058 ( .o(n4572), .a(n9787_1), .b(n6869), .c(n9783_1) );
in01f01  g3059 ( .o(n9789), .a(_net_6296) );
no02f01  g3060 ( .o(n4586), .a(_net_392), .b(n9789) );
ao12f01  g3061 ( .o(n9791), .a(n9107), .b(_net_7232), .c(net_7231) );
no03f01  g3062 ( .o(n9792_1), .a(_net_7233), .b(n9116), .c(n9113) );
no02f01  g3063 ( .o(n9793), .a(n9792_1), .b(n9791) );
oa22f01  g3064 ( .o(n4591), .a(n9793), .b(n9568), .c(n9572), .d(n9107) );
in01f01  g3065 ( .o(n9795), .a(_net_7413) );
na02f01  g3066 ( .o(n9796_1), .a(n8633), .b(n7550) );
oa12f01  g3067 ( .o(n4596), .a(n9796_1), .b(n7550), .c(n9795) );
in01f01  g3068 ( .o(n9798), .a(_net_7586) );
na02f01  g3069 ( .o(n9799), .a(n8000), .b(n6968) );
oa12f01  g3070 ( .o(n4609), .a(n9799), .b(n6968), .c(n9798) );
in01f01  g3071 ( .o(n9801_1), .a(_net_7346) );
na02f01  g3072 ( .o(n9802), .a(n8731), .b(n7030) );
oa12f01  g3073 ( .o(n4627), .a(n9802), .b(n7030), .c(n9801_1) );
ao22f01  g3074 ( .o(n9804), .a(n6736_1), .b(net_7639), .c(n6734), .d(net_7607) );
ao22f01  g3075 ( .o(n9805_1), .a(n6739), .b(net_7671), .c(n6738), .d(_net_7575) );
na02f01  g3076 ( .o(n4636), .a(n9805_1), .b(n9804) );
na02f01  g3077 ( .o(n9807), .a(n8034), .b(_net_6064) );
ao22f01  g3078 ( .o(n9808), .a(n6777), .b(net_6424), .c(n6776), .d(net_6488) );
ao22f01  g3079 ( .o(n9809_1), .a(n6780), .b(net_6456), .c(n6779_1), .d(net_6520) );
na02f01  g3080 ( .o(n9810), .a(n9809_1), .b(n9808) );
na02f01  g3081 ( .o(n9811), .a(n9810), .b(n8028_1) );
na02f01  g3082 ( .o(n4641), .a(n9811), .b(n9807) );
in01f01  g3083 ( .o(n9813), .a(_net_7269) );
na02f01  g3084 ( .o(n9814_1), .a(n9685), .b(n6901) );
oa12f01  g3085 ( .o(n4646), .a(n9814_1), .b(n6901), .c(n9813) );
in01f01  g3086 ( .o(n9816), .a(_net_7288) );
na02f01  g3087 ( .o(n9817), .a(n8208), .b(n7180) );
oa12f01  g3088 ( .o(n4656), .a(n9817), .b(n7180), .c(n9816) );
na03f01  g3089 ( .o(n9819_1), .a(n8089), .b(_net_6407), .c(n9258_1) );
no04f01  g3090 ( .o(n4673), .a(n9819_1), .b(n9672), .c(n8084), .d(_net_6408) );
ao22f01  g3091 ( .o(n9821), .a(n7288_1), .b(_net_6030), .c(n7286), .d(_net_269) );
ao22f01  g3092 ( .o(n9822), .a(n7298), .b(_net_7722), .c(n7291), .d(_net_7693) );
na02f01  g3093 ( .o(n9823), .a(n7302_1), .b(_net_116) );
na03f01  g3094 ( .o(n9824_1), .a(n7308), .b(net_195), .c(x1322) );
na02f01  g3095 ( .o(n9825), .a(n7296), .b(net_232) );
na03f01  g3096 ( .o(n9826), .a(n7308), .b(net_158), .c(n6800) );
na03f01  g3097 ( .o(n9827), .a(n9826), .b(n9825), .c(n9824_1) );
ao12f01  g3098 ( .o(n9828_1), .a(n9827), .b(n7306), .c(_net_5986) );
na04f01  g3099 ( .o(n4678), .a(n9828_1), .b(n9823), .c(n9822), .d(n9821) );
no02f01  g3100 ( .o(n4703), .a(n7232), .b(n7159) );
ao22f01  g3101 ( .o(n9831), .a(n6777), .b(net_6429), .c(n6776), .d(net_6493) );
ao22f01  g3102 ( .o(n9832), .a(n6780), .b(net_6461), .c(n6779_1), .d(net_6525) );
ao12f01  g3103 ( .o(n9833_1), .a(n6764), .b(n9832), .c(n9831) );
no02f01  g3104 ( .o(n9834), .a(n9181), .b(n6766) );
in01f01  g3105 ( .o(n9835), .a(_net_6073) );
oa22f01  g3106 ( .o(n9836), .a(n7964), .b(n6775), .c(n6784), .d(n9835) );
no03f01  g3107 ( .o(n9837_1), .a(n9836), .b(n9834), .c(n9833_1) );
in01f01  g3108 ( .o(n9838), .a(net_6477) );
in01f01  g3109 ( .o(n9839), .a(net_6445) );
oa22f01  g3110 ( .o(n9840_1), .a(n6790), .b(n9839), .c(n6789), .d(n9838) );
in01f01  g3111 ( .o(n9841), .a(net_6541) );
in01f01  g3112 ( .o(n9842), .a(net_6509) );
oa22f01  g3113 ( .o(n9843), .a(n6795), .b(n9841), .c(n6794), .d(n9842) );
no02f01  g3114 ( .o(n9844_1), .a(n9843), .b(n9840_1) );
na02f01  g3115 ( .o(n4708), .a(n9844_1), .b(n9837_1) );
in01f01  g3116 ( .o(n9846), .a(_net_7692) );
na02f01  g3117 ( .o(n9847), .a(n7207_1), .b(_net_7794) );
oa12f01  g3118 ( .o(n4727), .a(n9847), .b(n7207_1), .c(n9846) );
in01f01  g3119 ( .o(n9849_1), .a(_net_7286) );
na02f01  g3120 ( .o(n9850), .a(n8960), .b(n7180) );
oa12f01  g3121 ( .o(n4732), .a(n9850), .b(n7180), .c(n9849_1) );
no03f01  g3122 ( .o(n9852), .a(n6898), .b(n9592_1), .c(n8094) );
na02f01  g3123 ( .o(n9853_1), .a(n9852), .b(n7026) );
in01f01  g3124 ( .o(n9854), .a(_net_7381) );
no02f01  g3125 ( .o(n9855), .a(n9854), .b(_net_7382) );
no02f01  g3126 ( .o(n9856), .a(_net_7381), .b(n7026) );
na02f01  g3127 ( .o(n9857), .a(n6897), .b(_net_267) );
no02f01  g3128 ( .o(n9858_1), .a(n9857), .b(n6899_1) );
oa12f01  g3129 ( .o(n9859), .a(n9858_1), .b(n9856), .c(n9855) );
no02f01  g3130 ( .o(n9860), .a(n6897), .b(n8094) );
na02f01  g3131 ( .o(n9861), .a(n9860), .b(_net_7382) );
na03f01  g3132 ( .o(n4737), .a(n9861), .b(n9859), .c(n9853_1) );
in01f01  g3133 ( .o(n9863_1), .a(_net_7706) );
na02f01  g3134 ( .o(n9864), .a(n7207_1), .b(_net_7808) );
oa12f01  g3135 ( .o(n4760), .a(n9864), .b(n7207_1), .c(n9863_1) );
in01f01  g3136 ( .o(n9866), .a(_net_7559) );
na02f01  g3137 ( .o(n9867_1), .a(n9493), .b(n7519) );
oa12f01  g3138 ( .o(n4787), .a(n9867_1), .b(n7519), .c(n9866) );
in01f01  g3139 ( .o(n9869), .a(_net_7452) );
in01f01  g3140 ( .o(n9870), .a(net_365) );
in01f01  g3141 ( .o(n9871_1), .a(net_353) );
oa22f01  g3142 ( .o(n9872), .a(n6867_1), .b(n9871_1), .c(n8192_1), .d(n9870) );
na02f01  g3143 ( .o(n9873), .a(n9872), .b(n7197) );
oa12f01  g3144 ( .o(n4800), .a(n9873), .b(n7197), .c(n9869) );
in01f01  g3145 ( .o(n9875_1), .a(_net_7655) );
na02f01  g3146 ( .o(n9876), .a(n9493), .b(n7446_1) );
oa12f01  g3147 ( .o(n4809), .a(n9876), .b(n7446_1), .c(n9875_1) );
in01f01  g3148 ( .o(n9878), .a(_net_7624) );
na02f01  g3149 ( .o(n9879), .a(n6965), .b(net_7544) );
ao22f01  g3150 ( .o(n9880_1), .a(net_374), .b(_net_292), .c(_net_291), .d(net_376) );
na02f01  g3151 ( .o(n9881), .a(n9880_1), .b(n9879) );
na02f01  g3152 ( .o(n9882), .a(n9881), .b(n7400_1) );
oa12f01  g3153 ( .o(n4818), .a(n9882), .b(n7400_1), .c(n9878) );
na02f01  g3154 ( .o(n9884), .a(n7306), .b(_net_6019) );
na02f01  g3155 ( .o(n9885_1), .a(n7293), .b(net_219) );
ao22f01  g3156 ( .o(n9886), .a(n7297_1), .b(net_182), .c(n7296), .d(net_256) );
ao22f01  g3157 ( .o(n9887), .a(n7298), .b(_net_7746), .c(n7291), .d(_net_7717) );
na04f01  g3158 ( .o(n4831), .a(n9887), .b(n9886), .c(n9885_1), .d(n9884) );
in01f01  g3159 ( .o(n9889_1), .a(_net_6019) );
na02f01  g3160 ( .o(n9890), .a(n7348), .b(_net_7819) );
oa12f01  g3161 ( .o(n4843), .a(n9890), .b(n7348), .c(n9889_1) );
in01f01  g3162 ( .o(n9892), .a(n6802) );
na03f01  g3163 ( .o(n9893), .a(n8316_1), .b(n7281), .c(x1322) );
no02f01  g3164 ( .o(n4857), .a(n9893), .b(n9892) );
in01f01  g3165 ( .o(n9895), .a(_net_284) );
na02f01  g3166 ( .o(n9896), .a(n7440), .b(net_7807) );
oa12f01  g3167 ( .o(n4872), .a(n9896), .b(n7440), .c(n9895) );
ao12f01  g3168 ( .o(n9898), .a(x38), .b(n9259), .c(_net_6406) );
oa12f01  g3169 ( .o(n4877), .a(n9898), .b(n9259), .c(_net_6406) );
ao22f01  g3170 ( .o(n9900), .a(n7225), .b(_net_7410), .c(n7224), .d(_net_7442) );
ao22f01  g3171 ( .o(n9901), .a(n7229), .b(_net_7506), .c(n7228), .d(_net_7474) );
na02f01  g3172 ( .o(n4886), .a(n9901), .b(n9900) );
no02f01  g3173 ( .o(n4908), .a(n9893), .b(n8315) );
na02f01  g3174 ( .o(n9904), .a(n7348), .b(_net_7814) );
oa12f01  g3175 ( .o(n4917), .a(n9904), .b(n7348), .c(n7265_1) );
no02f01  g3176 ( .o(n9906), .a(n7125_1), .b(net_6826) );
no02f01  g3177 ( .o(n9907_1), .a(n9906), .b(n8323) );
no04f01  g3178 ( .o(n9908), .a(n8322), .b(n8321), .c(n7125_1), .d(net_6826) );
oa12f01  g3179 ( .o(n9909), .a(n8326), .b(n9908), .c(n9907_1) );
no02f01  g3180 ( .o(n9910), .a(n9908), .b(n9907_1) );
na02f01  g3181 ( .o(n9911_1), .a(n9910), .b(n2948) );
na02f01  g3182 ( .o(n4922), .a(n9911_1), .b(n9909) );
na02f01  g3183 ( .o(n9913), .a(n9311), .b(n9305) );
no02f01  g3184 ( .o(n9914_1), .a(n9308), .b(n9307_1) );
in01f01  g3185 ( .o(n9915), .a(n9914_1) );
na02f01  g3186 ( .o(n9916), .a(n9915), .b(n9309) );
oa22f01  g3187 ( .o(n4927), .a(n9916), .b(n9913), .c(n9313), .d(n9308) );
in01f01  g3188 ( .o(n9918_1), .a(_net_7659) );
na02f01  g3189 ( .o(n9919), .a(n7446_1), .b(n6971) );
oa12f01  g3190 ( .o(n4936), .a(n9919), .b(n7446_1), .c(n9918_1) );
in01f01  g3191 ( .o(n9921), .a(_net_295) );
na02f01  g3192 ( .o(n9922), .a(n7440), .b(_net_7815) );
oa12f01  g3193 ( .o(n4952), .a(n9922), .b(n7440), .c(n9921) );
in01f01  g3194 ( .o(n9924), .a(_net_7651) );
na02f01  g3195 ( .o(n9925), .a(n9154), .b(n7446_1) );
oa12f01  g3196 ( .o(n4961), .a(n9925), .b(n7446_1), .c(n9924) );
no02f01  g3197 ( .o(n9927), .a(n8060), .b(n7012) );
in01f01  g3198 ( .o(n9928), .a(net_6977) );
in01f01  g3199 ( .o(n9929), .a(net_7041) );
oa22f01  g3200 ( .o(n9930_1), .a(n6987), .b(n9928), .c(n6985), .d(n9929) );
in01f01  g3201 ( .o(n9931), .a(net_7073) );
in01f01  g3202 ( .o(n9932), .a(net_7009) );
oa22f01  g3203 ( .o(n9933), .a(n6992), .b(n9932), .c(n6991), .d(n9931) );
no02f01  g3204 ( .o(n9934), .a(n9933), .b(n9930_1) );
no02f01  g3205 ( .o(n9935_1), .a(n9934), .b(n6980) );
in01f01  g3206 ( .o(n9936), .a(_net_6157) );
oa22f01  g3207 ( .o(n9937), .a(n8069), .b(n6997), .c(n6995_1), .d(n9936) );
no03f01  g3208 ( .o(n9938), .a(n9937), .b(n9935_1), .c(n9927) );
in01f01  g3209 ( .o(n9939_1), .a(net_6989) );
in01f01  g3210 ( .o(n9940), .a(net_7021) );
oa22f01  g3211 ( .o(n9941), .a(n8075_1), .b(n9939_1), .c(n8074), .d(n9940) );
in01f01  g3212 ( .o(n9942), .a(net_7085) );
in01f01  g3213 ( .o(n9943), .a(net_7053) );
oa22f01  g3214 ( .o(n9944_1), .a(n8080_1), .b(n9942), .c(n8079), .d(n9943) );
no02f01  g3215 ( .o(n9945), .a(n9944_1), .b(n9941) );
na02f01  g3216 ( .o(n4974), .a(n9945), .b(n9938) );
in01f01  g3217 ( .o(n9947), .a(_net_7571) );
na02f01  g3218 ( .o(n9948), .a(n7519), .b(n7144) );
oa12f01  g3219 ( .o(n4987), .a(n9948), .b(n7519), .c(n9947) );
in01f01  g3220 ( .o(n9950), .a(_net_6029) );
no02f01  g3221 ( .o(n9951), .a(n7287), .b(n9950) );
in01f01  g3222 ( .o(n9952), .a(_net_7721) );
no04f01  g3223 ( .o(n9953_1), .a(n9705), .b(n7293), .c(n7292_1), .d(n9952) );
na02f01  g3224 ( .o(n9954), .a(x38), .b(n7300) );
no02f01  g3225 ( .o(n9955), .a(n9954), .b(n7301) );
no03f01  g3226 ( .o(n9956), .a(n9955), .b(n9953_1), .c(n9951) );
na02f01  g3227 ( .o(n9957_1), .a(n7302_1), .b(_net_115) );
in01f01  g3228 ( .o(n9958), .a(net_157) );
no04f01  g3229 ( .o(n9959), .a(n7307_1), .b(n7292_1), .c(n9958), .d(x1322) );
in01f01  g3230 ( .o(n9960), .a(net_231) );
no03f01  g3231 ( .o(n9961_1), .a(n7295), .b(n7294), .c(n9960) );
in01f01  g3232 ( .o(n9962), .a(net_194) );
no04f01  g3233 ( .o(n9963), .a(n7307_1), .b(n7292_1), .c(n9962), .d(n6800) );
no03f01  g3234 ( .o(n9964), .a(n9963), .b(n9961_1), .c(n9959) );
oa12f01  g3235 ( .o(n9965), .a(n9964), .b(n7305), .c(n7980_1) );
in01f01  g3236 ( .o(n9966_1), .a(_net_268) );
oa22f01  g3237 ( .o(n9967), .a(n7290), .b(n9846), .c(n7285), .d(n9966_1) );
no02f01  g3238 ( .o(n9968), .a(n9967), .b(n9965) );
na03f01  g3239 ( .o(n4992), .a(n9968), .b(n9957_1), .c(n9956) );
in01f01  g3240 ( .o(n9970), .a(_net_7727) );
in01f01  g3241 ( .o(n9971_1), .a(_net_6005) );
ao12f01  g3242 ( .o(n5013), .a(n7343), .b(n9971_1), .c(n9970) );
in01f01  g3243 ( .o(n9973), .a(_net_6693) );
in01f01  g3244 ( .o(n9974), .a(n513) );
ao12f01  g3245 ( .o(n9975), .a(n9973), .b(_net_6692), .c(net_6691) );
no03f01  g3246 ( .o(n9976_1), .a(n7663), .b(_net_6693), .c(n7153) );
no02f01  g3247 ( .o(n9977), .a(n9976_1), .b(n9975) );
na02f01  g3248 ( .o(n9978), .a(_net_5995), .b(n7067_1) );
oa22f01  g3249 ( .o(n5018), .a(n9978), .b(n9973), .c(n9977), .d(n9974) );
in01f01  g3250 ( .o(n9980), .a(net_355) );
no02f01  g3251 ( .o(n5027), .a(n6867_1), .b(n9980) );
in01f01  g3252 ( .o(n9982), .a(net_7799) );
na02f01  g3253 ( .o(n9983), .a(n6803), .b(_net_6034) );
oa12f01  g3254 ( .o(n5040), .a(n9983), .b(n6803), .c(n9982) );
in01f01  g3255 ( .o(n9985_1), .a(_net_7507) );
na02f01  g3256 ( .o(n9986), .a(n9786), .b(n7626_1) );
oa12f01  g3257 ( .o(n5061), .a(n9986), .b(n7626_1), .c(n9985_1) );
in01f01  g3258 ( .o(n9988_1), .a(_net_7508) );
na02f01  g3259 ( .o(n9989), .a(n7626_1), .b(n7553_1) );
oa12f01  g3260 ( .o(n5075), .a(n9989), .b(n7626_1), .c(n9988_1) );
in01f01  g3261 ( .o(n9991), .a(_net_7514) );
na02f01  g3262 ( .o(n9992_1), .a(n9487_1), .b(n7626_1) );
oa12f01  g3263 ( .o(n5080), .a(n9992_1), .b(n7626_1), .c(n9991) );
in01f01  g3264 ( .o(n9994), .a(net_7758) );
na04f01  g3265 ( .o(n9995), .a(_net_6028), .b(_net_7791), .c(net_303), .d(n9994) );
ao12f01  g3266 ( .o(n5085), .a(n9995), .b(net_305), .c(_net_6029) );
in01f01  g3267 ( .o(n9997_1), .a(_net_7433) );
na02f01  g3268 ( .o(n9998), .a(n7779_1), .b(n7197) );
oa12f01  g3269 ( .o(n5094), .a(n9998), .b(n7197), .c(n9997_1) );
na02f01  g3270 ( .o(n10000), .a(n7298), .b(net_7739) );
ao22f01  g3271 ( .o(n10001_1), .a(n7306), .b(_net_6009), .c(n7291), .d(net_7710) );
na02f01  g3272 ( .o(n10002), .a(n7302_1), .b(net_149) );
na02f01  g3273 ( .o(n10003), .a(n7296), .b(net_249) );
na03f01  g3274 ( .o(n10004), .a(n7308), .b(_net_175), .c(n6800) );
na03f01  g3275 ( .o(n10005), .a(n7308), .b(_net_212), .c(x1322) );
na03f01  g3276 ( .o(n10006_1), .a(n10005), .b(n10004), .c(n10003) );
ao12f01  g3277 ( .o(n10007), .a(n10006_1), .b(n7286), .c(_net_292) );
na04f01  g3278 ( .o(n5103), .a(n10007), .b(n10002), .c(n10001_1), .d(n10000) );
ao22f01  g3279 ( .o(n10009), .a(n7225), .b(_net_7416), .c(n7224), .d(_net_7448) );
ao22f01  g3280 ( .o(n10010_1), .a(n7229), .b(_net_7512), .c(n7228), .d(_net_7480) );
na02f01  g3281 ( .o(n5107), .a(n10010_1), .b(n10009) );
in01f01  g3282 ( .o(n10012), .a(_net_6415) );
na02f01  g3283 ( .o(n10013), .a(n7357), .b(net_6417) );
na02f01  g3284 ( .o(n10014_1), .a(n9305), .b(net_6417) );
in01f01  g3285 ( .o(n10015), .a(net_6412) );
in01f01  g3286 ( .o(n10016), .a(_net_6413) );
no02f01  g3287 ( .o(n10017), .a(n10016), .b(n10015) );
na03f01  g3288 ( .o(n10018), .a(n10017), .b(_net_6414), .c(_net_6415) );
in01f01  g3289 ( .o(n10019_1), .a(_net_6414) );
in01f01  g3290 ( .o(n10020), .a(n10017) );
oa12f01  g3291 ( .o(n10021), .a(n10012), .b(n10020), .c(n10019_1) );
na02f01  g3292 ( .o(n10022), .a(n10021), .b(n10018) );
oa22f01  g3293 ( .o(n5112), .a(n10022), .b(n10014_1), .c(n10013), .d(n10012) );
na02f01  g3294 ( .o(n10024), .a(n7339), .b(x1231) );
no04f01  g3295 ( .o(n5117), .a(n10024), .b(n7292_1), .c(x1215), .d(n6800) );
no02f01  g3296 ( .o(n10026), .a(n7339), .b(n7112) );
no03f01  g3297 ( .o(n5130), .a(n10026), .b(n7336), .c(x149) );
ao22f01  g3298 ( .o(n10028_1), .a(n7225), .b(_net_7426), .c(n7224), .d(net_7458) );
ao22f01  g3299 ( .o(n10029), .a(n7229), .b(net_7522), .c(n7228), .d(net_7490) );
na02f01  g3300 ( .o(n5134), .a(n10029), .b(n10028_1) );
in01f01  g3301 ( .o(n10031), .a(_net_7272) );
na02f01  g3302 ( .o(n10032_1), .a(n2913), .b(n6901) );
oa12f01  g3303 ( .o(n5143), .a(n10032_1), .b(n6901), .c(n10031) );
in01f01  g3304 ( .o(n10034), .a(_net_271) );
na02f01  g3305 ( .o(n10035), .a(n7440), .b(_net_7797) );
oa12f01  g3306 ( .o(n5164), .a(n10035), .b(n7440), .c(n10034) );
in01f01  g3307 ( .o(n10037_1), .a(_net_7435) );
na02f01  g3308 ( .o(n10038), .a(n9700_1), .b(n7197) );
oa12f01  g3309 ( .o(n5169), .a(n10038), .b(n7197), .c(n10037_1) );
na02f01  g3310 ( .o(n10040), .a(n6933), .b(_net_6084) );
na02f01  g3311 ( .o(n10041), .a(n6942), .b(n6917) );
na02f01  g3312 ( .o(n5198), .a(n10041), .b(n10040) );
no03f01  g3313 ( .o(n10043), .a(n6965), .b(n7654_1), .c(n8236) );
na02f01  g3314 ( .o(n10044), .a(n7444), .b(_net_7686) );
na02f01  g3315 ( .o(n10045), .a(n7445), .b(n8348) );
na03f01  g3316 ( .o(n10046), .a(n10045), .b(n10044), .c(n10043) );
no02f01  g3317 ( .o(n10047_1), .a(n8232_1), .b(n6966) );
na03f01  g3318 ( .o(n10048), .a(_net_7685), .b(_net_7684), .c(_net_7683) );
na02f01  g3319 ( .o(n10049), .a(n10048), .b(n8348) );
in01f01  g3320 ( .o(n10050), .a(n10048) );
na02f01  g3321 ( .o(n10051), .a(n10050), .b(_net_7686) );
na03f01  g3322 ( .o(n10052_1), .a(n10051), .b(n10049), .c(n10047_1) );
na02f01  g3323 ( .o(n10053), .a(n8237_1), .b(_net_7686) );
na03f01  g3324 ( .o(n5207), .a(n10053), .b(n10052_1), .c(n10046) );
no02f01  g3325 ( .o(n10055), .a(n9502_1), .b(n7468_1) );
no02f01  g3326 ( .o(n10056_1), .a(n9467_1), .b(n7470) );
in01f01  g3327 ( .o(n10057), .a(_net_6114) );
oa22f01  g3328 ( .o(n10058), .a(n8557_1), .b(n7123), .c(n7118), .d(n10057) );
no03f01  g3329 ( .o(n10059), .a(n10058), .b(n10056_1), .c(n10055) );
in01f01  g3330 ( .o(n10060), .a(net_6716) );
in01f01  g3331 ( .o(n10061_1), .a(net_6748) );
oa22f01  g3332 ( .o(n10062), .a(n7492_1), .b(n10060), .c(n7491), .d(n10061_1) );
in01f01  g3333 ( .o(n10063), .a(net_6812) );
in01f01  g3334 ( .o(n10064), .a(net_6780) );
oa22f01  g3335 ( .o(n10065), .a(n7497), .b(n10063), .c(n7496_1), .d(n10064) );
no02f01  g3336 ( .o(n10066_1), .a(n10065), .b(n10062) );
na02f01  g3337 ( .o(n5212), .a(n10066_1), .b(n10059) );
in01f01  g3338 ( .o(n10068), .a(_net_7593) );
na02f01  g3339 ( .o(n10069), .a(n6965), .b(net_7545) );
ao22f01  g3340 ( .o(n10070_1), .a(_net_292), .b(net_375), .c(_net_291), .d(net_377) );
na02f01  g3341 ( .o(n10071), .a(n10070_1), .b(n10069) );
na02f01  g3342 ( .o(n10072), .a(n10071), .b(n6968) );
oa12f01  g3343 ( .o(n5225), .a(n10072), .b(n6968), .c(n10068) );
in01f01  g3344 ( .o(n10074_1), .a(_net_7422) );
na02f01  g3345 ( .o(n10075), .a(n5027), .b(n7550) );
oa12f01  g3346 ( .o(n5230), .a(n10075), .b(n7550), .c(n10074_1) );
in01f01  g3347 ( .o(n10077), .a(_net_7297) );
na02f01  g3348 ( .o(n10078), .a(n9537_1), .b(n7180) );
oa12f01  g3349 ( .o(n5251), .a(n10078), .b(n7180), .c(n10077) );
in01f01  g3350 ( .o(n10080), .a(_net_7567) );
na02f01  g3351 ( .o(n10081), .a(n8639), .b(n7519) );
oa12f01  g3352 ( .o(n5256), .a(n10081), .b(n7519), .c(n10080) );
in01f01  g3353 ( .o(n10083), .a(_net_7416) );
na02f01  g3354 ( .o(n10084_1), .a(n7638), .b(n7550) );
oa12f01  g3355 ( .o(n5265), .a(n10084_1), .b(n7550), .c(n10083) );
in01f01  g3356 ( .o(n10086), .a(_net_7292) );
na02f01  g3357 ( .o(n10087), .a(n6898), .b(net_7244) );
ao22f01  g3358 ( .o(n10088), .a(net_338), .b(_net_269), .c(_net_270), .d(net_336) );
na02f01  g3359 ( .o(n10089_1), .a(n10088), .b(n10087) );
na02f01  g3360 ( .o(n10090), .a(n10089_1), .b(n7180) );
oa12f01  g3361 ( .o(n5274), .a(n10090), .b(n7180), .c(n10086) );
in01f01  g3362 ( .o(n10092), .a(net_6025) );
in01f01  g3363 ( .o(n10093), .a(_net_7731) );
ao12f01  g3364 ( .o(n5279), .a(n7343), .b(n10093), .c(n10092) );
in01f01  g3365 ( .o(n10095), .a(_net_6283) );
no02f01  g3366 ( .o(n5284), .a(_net_392), .b(n10095) );
in01f01  g3367 ( .o(n10097), .a(_net_7599) );
na02f01  g3368 ( .o(n10098), .a(n8639), .b(n6968) );
oa12f01  g3369 ( .o(n5293), .a(n10098), .b(n6968), .c(n10097) );
in01f01  g3370 ( .o(n10100), .a(_net_7411) );
na02f01  g3371 ( .o(n10101), .a(n9786), .b(n7550) );
oa12f01  g3372 ( .o(n5307), .a(n10101), .b(n7550), .c(n10100) );
in01f01  g3373 ( .o(n10103_1), .a(net_7750) );
na04f01  g3374 ( .o(n10104), .a(_net_7791), .b(net_303), .c(_net_5984), .d(n10103_1) );
ao12f01  g3375 ( .o(n5316), .a(n10104), .b(net_309), .c(_net_5985) );
na02f01  g3376 ( .o(n10106), .a(n10043), .b(n6959) );
no02f01  g3377 ( .o(n10107_1), .a(_net_7684), .b(n8231) );
no02f01  g3378 ( .o(n10108), .a(n6959), .b(_net_7683) );
oa12f01  g3379 ( .o(n10109), .a(n10047_1), .b(n10108), .c(n10107_1) );
na02f01  g3380 ( .o(n10110), .a(n8237_1), .b(_net_7684) );
na03f01  g3381 ( .o(n5321), .a(n10110), .b(n10109), .c(n10106) );
in01f01  g3382 ( .o(n10112_1), .a(_net_7662) );
na02f01  g3383 ( .o(n10113), .a(n9373_1), .b(n7446_1) );
oa12f01  g3384 ( .o(n5330), .a(n10113), .b(n7446_1), .c(n10112_1) );
in01f01  g3385 ( .o(n10115), .a(_net_6420) );
na02f01  g3386 ( .o(n10116_1), .a(n9412), .b(n10115) );
na02f01  g3387 ( .o(n10117), .a(n10116_1), .b(n9664_1) );
oa22f01  g3388 ( .o(n5344), .a(n10117), .b(n9411), .c(n9409), .d(n10115) );
in01f01  g3389 ( .o(n10119), .a(_net_7280) );
na02f01  g3390 ( .o(n10120_1), .a(n875), .b(n6901) );
oa12f01  g3391 ( .o(n5353), .a(n10120_1), .b(n6901), .c(n10119) );
in01f01  g3392 ( .o(n10122), .a(_net_7657) );
na02f01  g3393 ( .o(n10123), .a(n10071), .b(n7446_1) );
oa12f01  g3394 ( .o(n5370), .a(n10123), .b(n7446_1), .c(n10122) );
no02f01  g3395 ( .o(n10125), .a(n9292), .b(n6945) );
in01f01  g3396 ( .o(n10126), .a(net_6633) );
in01f01  g3397 ( .o(n10127), .a(net_6569) );
oa22f01  g3398 ( .o(n10128_1), .a(n6922), .b(n10127), .c(n6919_1), .d(n10126) );
in01f01  g3399 ( .o(n10129), .a(net_6665) );
in01f01  g3400 ( .o(n10130), .a(net_6601) );
oa22f01  g3401 ( .o(n10131), .a(n6927), .b(n10130), .c(n6925), .d(n10129) );
no02f01  g3402 ( .o(n10132_1), .a(n10131), .b(n10128_1) );
no02f01  g3403 ( .o(n10133), .a(n10132_1), .b(n6934_1) );
in01f01  g3404 ( .o(n10134), .a(_net_6096) );
oa22f01  g3405 ( .o(n10135), .a(n7042), .b(n6916), .c(n6932), .d(n10134) );
no03f01  g3406 ( .o(n10136), .a(n10135), .b(n10133), .c(n10125) );
in01f01  g3407 ( .o(n10137_1), .a(net_6583) );
in01f01  g3408 ( .o(n10138), .a(net_6615) );
oa22f01  g3409 ( .o(n10139), .a(n7058_1), .b(n10137_1), .c(n7057), .d(n10138) );
in01f01  g3410 ( .o(n10140), .a(net_6679) );
in01f01  g3411 ( .o(n10141_1), .a(net_6647) );
oa22f01  g3412 ( .o(n10142), .a(n7063), .b(n10140), .c(n7062_1), .d(n10141_1) );
no02f01  g3413 ( .o(n10143), .a(n10142), .b(n10139) );
na02f01  g3414 ( .o(n5388), .a(n10143), .b(n10136) );
ao22f01  g3415 ( .o(n10145_1), .a(n6877), .b(_net_7253), .c(n6876_1), .d(_net_7317) );
ao22f01  g3416 ( .o(n10146), .a(n6881_1), .b(_net_7285), .c(n6880), .d(_net_7349) );
na02f01  g3417 ( .o(n5397), .a(n10146), .b(n10145_1) );
in01f01  g3418 ( .o(n10148), .a(_net_7429) );
na02f01  g3419 ( .o(n10149), .a(n7550), .b(n420) );
oa12f01  g3420 ( .o(n5406), .a(n10149), .b(n7550), .c(n10148) );
in01f01  g3421 ( .o(n10151), .a(_net_7631) );
na02f01  g3422 ( .o(n10152), .a(n8639), .b(n7400_1) );
oa12f01  g3423 ( .o(n5411), .a(n10152), .b(n7400_1), .c(n10151) );
in01f01  g3424 ( .o(n10154_1), .a(_net_7295) );
na02f01  g3425 ( .o(n10155), .a(n7994_1), .b(n7180) );
oa12f01  g3426 ( .o(n5420), .a(n10155), .b(n7180), .c(n10154_1) );
in01f01  g3427 ( .o(n10157), .a(_net_7795) );
na02f01  g3428 ( .o(n10158_1), .a(n6803), .b(_net_6030) );
oa12f01  g3429 ( .o(n5429), .a(n10158_1), .b(n6803), .c(n10157) );
in01f01  g3430 ( .o(n10160), .a(_net_119) );
na02f01  g3431 ( .o(n10161), .a(net_315), .b(_net_154) );
oa12f01  g3432 ( .o(n5446), .a(n10161), .b(n10160), .c(_net_154) );
in01f01  g3433 ( .o(n10163), .a(_net_5987) );
na02f01  g3434 ( .o(n10164), .a(n7348), .b(_net_7796) );
oa12f01  g3435 ( .o(n5455), .a(n10164), .b(n7348), .c(n10163) );
in01f01  g3436 ( .o(n10166), .a(_net_7587) );
na02f01  g3437 ( .o(n10167), .a(n9154), .b(n6968) );
oa12f01  g3438 ( .o(n5477), .a(n10167), .b(n6968), .c(n10166) );
in01f01  g3439 ( .o(n10169), .a(_net_7513) );
na02f01  g3440 ( .o(n10170), .a(n7626_1), .b(n6872_1) );
oa12f01  g3441 ( .o(n5490), .a(n10170), .b(n7626_1), .c(n10169) );
na02f01  g3442 ( .o(n10172), .a(n7440), .b(_net_7796) );
oa12f01  g3443 ( .o(n5495), .a(n10172), .b(n7440), .c(n7253) );
in01f01  g3444 ( .o(n10174), .a(_net_7467) );
na02f01  g3445 ( .o(n10175), .a(n9700_1), .b(n6869) );
oa12f01  g3446 ( .o(n5508), .a(n10175), .b(n6869), .c(n10174) );
na02f01  g3447 ( .o(n10177), .a(n7298), .b(net_7738) );
ao22f01  g3448 ( .o(n10178), .a(n7306), .b(_net_6008), .c(n7291), .d(net_7709) );
na02f01  g3449 ( .o(n10179), .a(n7302_1), .b(net_148) );
na02f01  g3450 ( .o(n10180), .a(n7296), .b(net_248) );
na03f01  g3451 ( .o(n10181), .a(n7308), .b(_net_174), .c(n6800) );
na03f01  g3452 ( .o(n10182), .a(n7308), .b(_net_211), .c(x1322) );
na03f01  g3453 ( .o(n10183), .a(n10182), .b(n10181), .c(n10180) );
ao12f01  g3454 ( .o(n10184), .a(n10183), .b(n7286), .c(_net_291) );
na04f01  g3455 ( .o(n5517), .a(n10184), .b(n10179), .c(n10178), .d(n10177) );
na02f01  g3456 ( .o(n10186), .a(n7302_1), .b(net_153) );
na02f01  g3457 ( .o(n10187), .a(n7306), .b(net_6024) );
na02f01  g3458 ( .o(n10188), .a(n7296), .b(net_261) );
ao22f01  g3459 ( .o(n10189), .a(n7297_1), .b(net_187), .c(n7293), .d(net_224) );
na04f01  g3460 ( .o(n5525), .a(n10189), .b(n10188), .c(n10187), .d(n10186) );
in01f01  g3461 ( .o(n10191), .a(_net_293) );
no02f01  g3462 ( .o(n10192), .a(n10191), .b(_net_294) );
na02f01  g3463 ( .o(n10193), .a(_net_289), .b(_net_295) );
ao12f01  g3464 ( .o(n10194), .a(n10193), .b(_net_266), .c(n7653) );
na02f01  g3465 ( .o(n10195), .a(n10194), .b(n10192) );
in01f01  g3466 ( .o(n10196), .a(n10193) );
no02f01  g3467 ( .o(n10197), .a(n10191), .b(n9540) );
na03f01  g3468 ( .o(n10198), .a(n10197), .b(n10196), .c(_net_263) );
na03f01  g3469 ( .o(n10199), .a(_net_265), .b(_net_266), .c(n7653) );
na04f01  g3470 ( .o(n10200), .a(n10199), .b(n10196), .c(n10191), .d(n9540) );
oa12f01  g3471 ( .o(n10201), .a(n7653), .b(_net_265), .c(_net_266) );
na04f01  g3472 ( .o(n10202), .a(n10201), .b(n10196), .c(n10191), .d(_net_294) );
na04f01  g3473 ( .o(n10203), .a(n10202), .b(n10200), .c(n10198), .d(n10195) );
in01f01  g3474 ( .o(n10204), .a(n10203) );
no02f01  g3475 ( .o(n5529), .a(n10204), .b(x837) );
na02f01  g3476 ( .o(n10206), .a(n7232), .b(net_7771) );
no02f01  g3477 ( .o(n10207), .a(n10206), .b(n6885) );
no02f01  g3478 ( .o(n10208), .a(n10207), .b(_net_7721) );
no02f01  g3479 ( .o(n5534), .a(n10208), .b(n7343) );
in01f01  g3480 ( .o(n10210), .a(_net_7577) );
na02f01  g3481 ( .o(n10211), .a(n3015), .b(n7519) );
oa12f01  g3482 ( .o(n5543), .a(n10211), .b(n7519), .c(n10210) );
no02f01  g3483 ( .o(n5552), .a(n6867_1), .b(n9870) );
in01f01  g3484 ( .o(n10214), .a(_net_7430) );
in01f01  g3485 ( .o(n10215), .a(net_363) );
no02f01  g3486 ( .o(n6437), .a(n6867_1), .b(n10215) );
na02f01  g3487 ( .o(n10217), .a(n6437), .b(n7550) );
oa12f01  g3488 ( .o(n5565), .a(n10217), .b(n7550), .c(n10214) );
in01f01  g3489 ( .o(n10219), .a(_net_7502) );
na02f01  g3490 ( .o(n10220), .a(n7860), .b(n7626_1) );
oa12f01  g3491 ( .o(n5570), .a(n10220), .b(n7626_1), .c(n10219) );
in01f01  g3492 ( .o(n10222), .a(_net_7622) );
na02f01  g3493 ( .o(n10223), .a(n7644_1), .b(n7400_1) );
oa12f01  g3494 ( .o(n5579), .a(n10223), .b(n7400_1), .c(n10222) );
no02f01  g3495 ( .o(n10225), .a(n8610), .b(n7012) );
no02f01  g3496 ( .o(n10226), .a(n8619), .b(n6997) );
in01f01  g3497 ( .o(n10227), .a(_net_6162) );
no02f01  g3498 ( .o(n10228), .a(n7020), .b(n7017) );
oa22f01  g3499 ( .o(n10229), .a(n10228), .b(n6980), .c(n6995_1), .d(n10227) );
no03f01  g3500 ( .o(n10230), .a(n10229), .b(n10226), .c(n10225) );
in01f01  g3501 ( .o(n10231), .a(net_7026) );
in01f01  g3502 ( .o(n10232), .a(net_6994) );
oa22f01  g3503 ( .o(n10233), .a(n8075_1), .b(n10232), .c(n8074), .d(n10231) );
in01f01  g3504 ( .o(n10234), .a(net_7058) );
in01f01  g3505 ( .o(n10235), .a(net_7090) );
oa22f01  g3506 ( .o(n10236), .a(n8080_1), .b(n10235), .c(n8079), .d(n10234) );
no02f01  g3507 ( .o(n10237), .a(n10236), .b(n10233) );
na02f01  g3508 ( .o(n5596), .a(n10237), .b(n10230) );
in01f01  g3509 ( .o(n10239), .a(_net_7420) );
na02f01  g3510 ( .o(n10240), .a(n9872), .b(n7550) );
oa12f01  g3511 ( .o(n5601), .a(n10240), .b(n7550), .c(n10239) );
no02f01  g3512 ( .o(n10242), .a(n8452), .b(n6824) );
in01f01  g3513 ( .o(n10243), .a(net_6841) );
in01f01  g3514 ( .o(n10244), .a(net_6905) );
oa22f01  g3515 ( .o(n10245), .a(n6810), .b(n10243), .c(n6807), .d(n10244) );
in01f01  g3516 ( .o(n10246), .a(net_6873) );
in01f01  g3517 ( .o(n10247), .a(net_6937) );
oa22f01  g3518 ( .o(n10248), .a(n6815), .b(n10246), .c(n6813_1), .d(n10247) );
no02f01  g3519 ( .o(n10249), .a(n10248), .b(n10245) );
no02f01  g3520 ( .o(n10250), .a(n10249), .b(n6826_1) );
in01f01  g3521 ( .o(n10251), .a(_net_6138) );
oa22f01  g3522 ( .o(n10252), .a(n9127), .b(n6836_1), .c(n6844), .d(n10251) );
no03f01  g3523 ( .o(n10253), .a(n10252), .b(n10250), .c(n10242) );
in01f01  g3524 ( .o(n10254), .a(net_6855) );
in01f01  g3525 ( .o(n10255), .a(net_6887) );
oa22f01  g3526 ( .o(n10256), .a(n6850_1), .b(n10254), .c(n6849), .d(n10255) );
in01f01  g3527 ( .o(n10257), .a(net_6951) );
in01f01  g3528 ( .o(n10258), .a(net_6919) );
oa22f01  g3529 ( .o(n10259), .a(n6855_1), .b(n10257), .c(n6854), .d(n10258) );
no02f01  g3530 ( .o(n10260), .a(n10259), .b(n10256) );
na02f01  g3531 ( .o(n5623), .a(n10260), .b(n10253) );
in01f01  g3532 ( .o(n10262), .a(_net_7736) );
ao12f01  g3533 ( .o(n5633), .a(n7343), .b(n10262), .c(n8875) );
in01f01  g3534 ( .o(n10264), .a(_net_6204) );
no02f01  g3535 ( .o(n5638), .a(_net_392), .b(n10264) );
in01f01  g3536 ( .o(n10266), .a(_net_7634) );
na02f01  g3537 ( .o(n10267), .a(n7892), .b(n7400_1) );
oa12f01  g3538 ( .o(n5643), .a(n10267), .b(n7400_1), .c(n10266) );
no02f01  g3539 ( .o(n5660), .a(n7332), .b(n8803) );
no02f01  g3540 ( .o(n10270), .a(n6880), .b(n9440) );
no03f01  g3541 ( .o(n10271), .a(_net_7380), .b(n6879), .c(n6875) );
no02f01  g3542 ( .o(n10272), .a(n10271), .b(n10270) );
oa22f01  g3543 ( .o(n5669), .a(n10272), .b(n8096), .c(n8097_1), .d(n9440) );
in01f01  g3544 ( .o(n10274), .a(_net_7564) );
na02f01  g3545 ( .o(n10275), .a(n8043), .b(n7519) );
oa12f01  g3546 ( .o(n5674), .a(n10275), .b(n7519), .c(n10274) );
in01f01  g3547 ( .o(n10277), .a(_net_6282) );
no02f01  g3548 ( .o(n5691), .a(n10277), .b(_net_392) );
ao22f01  g3549 ( .o(n10279), .a(n6877), .b(_net_7263), .c(n6876_1), .d(_net_7327) );
ao22f01  g3550 ( .o(n10280), .a(n6881_1), .b(_net_7295), .c(n6880), .d(_net_7359) );
na02f01  g3551 ( .o(n5700), .a(n10280), .b(n10279) );
in01f01  g3552 ( .o(n5709), .a(n10014_1) );
in01f01  g3553 ( .o(n10283), .a(_net_269) );
na02f01  g3554 ( .o(n10284), .a(n7440), .b(_net_7795) );
oa12f01  g3555 ( .o(n5722), .a(n10284), .b(n7440), .c(n10283) );
in01f01  g3556 ( .o(n10286), .a(_net_5998) );
na02f01  g3557 ( .o(n10287), .a(n7348), .b(_net_7804) );
oa12f01  g3558 ( .o(n5739), .a(n10287), .b(n7348), .c(n10286) );
no02f01  g3559 ( .o(n10289), .a(n8711_1), .b(n8713) );
na02f01  g3560 ( .o(n10290), .a(n10289), .b(n9605) );
no03f01  g3561 ( .o(n10291), .a(n7467), .b(n7117), .c(n7121) );
no02f01  g3562 ( .o(n10292), .a(n7132), .b(n9600) );
no02f01  g3563 ( .o(n10293), .a(n7133_1), .b(_net_6825) );
no02f01  g3564 ( .o(n10294), .a(n10293), .b(n10292) );
ao22f01  g3565 ( .o(n10295), .a(n10294), .b(n10291), .c(n8716), .d(_net_6825) );
na02f01  g3566 ( .o(n5748), .a(n10295), .b(n10290) );
no02f01  g3567 ( .o(n10297), .a(n10017), .b(n10019_1) );
no02f01  g3568 ( .o(n10298), .a(n10020), .b(_net_6414) );
no02f01  g3569 ( .o(n10299), .a(n10298), .b(n10297) );
oa22f01  g3570 ( .o(n5753), .a(n10299), .b(n10014_1), .c(n10013), .d(n10019_1) );
no02f01  g3571 ( .o(n10301), .a(n7012), .b(n9626) );
no02f01  g3572 ( .o(n10302), .a(n8782), .b(n6997) );
in01f01  g3573 ( .o(n10303), .a(_net_6154) );
oa22f01  g3574 ( .o(n10304), .a(n8790), .b(n6980), .c(n6995_1), .d(n10303) );
no03f01  g3575 ( .o(n10305), .a(n10304), .b(n10302), .c(n10301) );
in01f01  g3576 ( .o(n10306), .a(net_6986) );
in01f01  g3577 ( .o(n10307), .a(net_7018) );
oa22f01  g3578 ( .o(n10308), .a(n8075_1), .b(n10306), .c(n8074), .d(n10307) );
in01f01  g3579 ( .o(n10309), .a(net_7082) );
in01f01  g3580 ( .o(n10310), .a(net_7050) );
oa22f01  g3581 ( .o(n10311), .a(n8080_1), .b(n10309), .c(n8079), .d(n10310) );
no02f01  g3582 ( .o(n10312), .a(n10311), .b(n10308) );
na02f01  g3583 ( .o(n5775), .a(n10312), .b(n10305) );
in01f01  g3584 ( .o(n10314), .a(_net_7561) );
na02f01  g3585 ( .o(n10315), .a(n10071), .b(n7519) );
oa12f01  g3586 ( .o(n5809), .a(n10315), .b(n7519), .c(n10314) );
in01f01  g3587 ( .o(n10317), .a(net_382) );
no02f01  g3588 ( .o(n5814), .a(n6966), .b(n10317) );
ao22f01  g3589 ( .o(n10319), .a(n6736_1), .b(_net_7633), .c(n6734), .d(_net_7601) );
ao22f01  g3590 ( .o(n10320), .a(n6739), .b(_net_7665), .c(n6738), .d(_net_7569) );
na02f01  g3591 ( .o(n5819), .a(n10320), .b(n10319) );
ao22f01  g3592 ( .o(n10322), .a(n6877), .b(_net_7258), .c(n6876_1), .d(_net_7322) );
ao22f01  g3593 ( .o(n10323), .a(n6881_1), .b(_net_7290), .c(n6880), .d(_net_7354) );
na02f01  g3594 ( .o(n5828), .a(n10323), .b(n10322) );
ao22f01  g3595 ( .o(n10325), .a(n6736_1), .b(net_7645), .c(n6734), .d(net_7613) );
ao22f01  g3596 ( .o(n10326), .a(n6739), .b(net_7677), .c(n6738), .d(_net_7581) );
na02f01  g3597 ( .o(n5845), .a(n10326), .b(n10325) );
in01f01  g3598 ( .o(n10328), .a(_net_7734) );
in01f01  g3599 ( .o(n10329), .a(net_6036) );
ao12f01  g3600 ( .o(n5850), .a(n7343), .b(n10329), .c(n10328) );
na02f01  g3601 ( .o(n10331), .a(n8177), .b(n8086) );
no03f01  g3602 ( .o(n10332), .a(_net_6407), .b(_net_6405), .c(_net_6406) );
na02f01  g3603 ( .o(n10333), .a(n10332), .b(n8088_1) );
no04f01  g3604 ( .o(n10334), .a(_net_6407), .b(_net_6405), .c(_net_6406), .d(_net_6404) );
ao12f01  g3605 ( .o(n5855), .a(n10331), .b(n10334), .c(n10333) );
no02f01  g3606 ( .o(n10336), .a(_net_7232), .b(n7579) );
no02f01  g3607 ( .o(n10337), .a(n9116), .b(_net_7229) );
no02f01  g3608 ( .o(n10338), .a(n10337), .b(n10336) );
no02f01  g3609 ( .o(n10339), .a(n7576), .b(net_7231) );
no02f01  g3610 ( .o(n10340), .a(n10339), .b(n10338) );
no04f01  g3611 ( .o(n10341), .a(n10337), .b(n10336), .c(n7576), .d(net_7231) );
oa12f01  g3612 ( .o(n10342), .a(n9641), .b(n10341), .c(n10340) );
no02f01  g3613 ( .o(n10343), .a(n10341), .b(n10340) );
na02f01  g3614 ( .o(n10344), .a(n10343), .b(n4276) );
na02f01  g3615 ( .o(n5885), .a(n10344), .b(n10342) );
na02f01  g3616 ( .o(n10346), .a(n7440), .b(_net_7806) );
oa12f01  g3617 ( .o(n5890), .a(n10346), .b(n7440), .c(n7415) );
in01f01  g3618 ( .o(n10348), .a(_net_7407) );
na02f01  g3619 ( .o(n10349), .a(n7550), .b(n7387) );
oa12f01  g3620 ( .o(n5899), .a(n10349), .b(n7550), .c(n10348) );
in01f01  g3621 ( .o(n10351), .a(net_7802) );
na02f01  g3622 ( .o(n10352), .a(n6803), .b(_net_6040) );
oa12f01  g3623 ( .o(n5925), .a(n10352), .b(n6803), .c(n10351) );
in01f01  g3624 ( .o(n10354), .a(_net_7553) );
na02f01  g3625 ( .o(n10355), .a(n8246), .b(n7519) );
oa12f01  g3626 ( .o(n5938), .a(n10355), .b(n7519), .c(n10354) );
na02f01  g3627 ( .o(n10357), .a(n7348), .b(_net_7809) );
oa12f01  g3628 ( .o(n5960), .a(n10357), .b(n7348), .c(n7121) );
in01f01  g3629 ( .o(n10359), .a(_net_7360) );
na02f01  g3630 ( .o(n10360), .a(n7437_1), .b(n7030) );
oa12f01  g3631 ( .o(n5973), .a(n10360), .b(n7030), .c(n10359) );
na02f01  g3632 ( .o(n10362), .a(n8120), .b(n6921) );
na02f01  g3633 ( .o(n10363), .a(n8122), .b(_net_6689) );
na02f01  g3634 ( .o(n10364), .a(n10363), .b(n10362) );
na02f01  g3635 ( .o(n10365), .a(n10364), .b(n8125_1) );
na02f01  g3636 ( .o(n10366), .a(n6927), .b(n6919_1) );
ao22f01  g3637 ( .o(n10367), .a(n10366), .b(n8127), .c(n8132), .d(_net_6689) );
na02f01  g3638 ( .o(n5982), .a(n10367), .b(n10365) );
ao12f01  g3639 ( .o(n10369), .a(x38), .b(n9546_1), .c(_net_6410) );
oa12f01  g3640 ( .o(n5987), .a(n10369), .b(n9546_1), .c(_net_6410) );
in01f01  g3641 ( .o(n10371), .a(_net_7357) );
na02f01  g3642 ( .o(n10372), .a(n8809_1), .b(n7030) );
oa12f01  g3643 ( .o(n5992), .a(n10372), .b(n7030), .c(n10371) );
na02f01  g3644 ( .o(n10374), .a(n8116_1), .b(n8028_1) );
ao22f01  g3645 ( .o(n10375), .a(n9810), .b(n8033_1), .c(n8034), .d(_net_6066) );
na02f01  g3646 ( .o(n5997), .a(n10375), .b(n10374) );
in01f01  g3647 ( .o(n10377), .a(_net_7596) );
na02f01  g3648 ( .o(n10378), .a(n8043), .b(n6968) );
oa12f01  g3649 ( .o(n6024), .a(n10378), .b(n6968), .c(n10377) );
no02f01  g3650 ( .o(n10380), .a(n7085_1), .b(n6764) );
no02f01  g3651 ( .o(n10381), .a(n7094), .b(n6766) );
in01f01  g3652 ( .o(n10382), .a(_net_6081) );
oa22f01  g3653 ( .o(n10383), .a(n9047_1), .b(n6775), .c(n6784), .d(n10382) );
no03f01  g3654 ( .o(n10384), .a(n10383), .b(n10381), .c(n10380) );
in01f01  g3655 ( .o(n10385), .a(net_6453) );
in01f01  g3656 ( .o(n10386), .a(net_6485) );
oa22f01  g3657 ( .o(n10387), .a(n6790), .b(n10385), .c(n6789), .d(n10386) );
in01f01  g3658 ( .o(n10388), .a(net_6517) );
in01f01  g3659 ( .o(n10389), .a(net_6549) );
oa22f01  g3660 ( .o(n10390), .a(n6795), .b(n10389), .c(n6794), .d(n10388) );
no02f01  g3661 ( .o(n10391), .a(n10390), .b(n10387) );
na02f01  g3662 ( .o(n6029), .a(n10391), .b(n10384) );
ao22f01  g3663 ( .o(n10393), .a(n6736_1), .b(net_7637), .c(n6734), .d(net_7605) );
ao22f01  g3664 ( .o(n10394), .a(n6739), .b(net_7669), .c(n6738), .d(_net_7573) );
na02f01  g3665 ( .o(n6038), .a(n10394), .b(n10393) );
ao12f01  g3666 ( .o(n10396), .a(n6824), .b(n9202), .c(n9201_1) );
no02f01  g3667 ( .o(n10397), .a(n8435_1), .b(n6826_1) );
in01f01  g3668 ( .o(n10398), .a(_net_6132) );
oa22f01  g3669 ( .o(n10399), .a(n8443_1), .b(n6836_1), .c(n6844), .d(n10398) );
no03f01  g3670 ( .o(n10400), .a(n10399), .b(n10397), .c(n10396) );
in01f01  g3671 ( .o(n10401), .a(net_6849) );
in01f01  g3672 ( .o(n10402), .a(net_6881) );
oa22f01  g3673 ( .o(n10403), .a(n6850_1), .b(n10401), .c(n6849), .d(n10402) );
in01f01  g3674 ( .o(n10404), .a(net_6913) );
in01f01  g3675 ( .o(n10405), .a(net_6945) );
oa22f01  g3676 ( .o(n10406), .a(n6855_1), .b(n10405), .c(n6854), .d(n10404) );
no02f01  g3677 ( .o(n10407), .a(n10406), .b(n10403) );
na02f01  g3678 ( .o(n6052), .a(n10407), .b(n10400) );
in01f01  g3679 ( .o(n10409), .a(_net_7482) );
na02f01  g3680 ( .o(n10410), .a(n9487_1), .b(n6869) );
oa12f01  g3681 ( .o(n6061), .a(n10410), .b(n6869), .c(n10409) );
in01f01  g3682 ( .o(n10412), .a(n2222) );
ao12f01  g3683 ( .o(n10413), .a(n7756_1), .b(_net_6557), .c(net_6556) );
no03f01  g3684 ( .o(n10414), .a(n7765), .b(_net_6558), .c(n7762) );
no02f01  g3685 ( .o(n10415), .a(n10414), .b(n10413) );
na02f01  g3686 ( .o(n10416), .a(_net_5984), .b(n8330) );
oa22f01  g3687 ( .o(n6074), .a(n10416), .b(n7756_1), .c(n10415), .d(n10412) );
ao22f01  g3688 ( .o(n10418), .a(n6736_1), .b(net_7647), .c(n6734), .d(net_7615) );
ao22f01  g3689 ( .o(n10419), .a(n6739), .b(net_7679), .c(n6738), .d(_net_7583) );
na02f01  g3690 ( .o(n6083), .a(n10419), .b(n10418) );
in01f01  g3691 ( .o(n10421), .a(_net_6407) );
na04f01  g3692 ( .o(n10422), .a(n10421), .b(_net_6410), .c(n9258_1), .d(n8084) );
in01f01  g3693 ( .o(n10423), .a(_net_6408) );
na02f01  g3694 ( .o(n10424), .a(_net_6409), .b(n10423) );
no03f01  g3695 ( .o(n6088), .a(n10424), .b(n10422), .c(n8090) );
in01f01  g3696 ( .o(n10426), .a(_net_7405) );
na02f01  g3697 ( .o(n10427), .a(n8817), .b(n7550) );
oa12f01  g3698 ( .o(n6093), .a(n10427), .b(n7550), .c(n10426) );
no02f01  g3699 ( .o(n10429), .a(n8291), .b(n7721) );
in01f01  g3700 ( .o(n10430), .a(net_7114) );
in01f01  g3701 ( .o(n10431), .a(net_7178) );
oa22f01  g3702 ( .o(n10432), .a(n7580), .b(n10430), .c(n7577_1), .d(n10431) );
in01f01  g3703 ( .o(n10433), .a(net_7146) );
in01f01  g3704 ( .o(n10434), .a(net_7210) );
oa22f01  g3705 ( .o(n10435), .a(n7585), .b(n10433), .c(n7583), .d(n10434) );
no02f01  g3706 ( .o(n10436), .a(n10435), .b(n10432) );
no02f01  g3707 ( .o(n10437), .a(n10436), .b(n7592) );
in01f01  g3708 ( .o(n10438), .a(_net_6181) );
no02f01  g3709 ( .o(n10439), .a(n8508_1), .b(n8505) );
oa22f01  g3710 ( .o(n10440), .a(n10439), .b(n7574), .c(n7590), .d(n10438) );
no03f01  g3711 ( .o(n10441), .a(n10440), .b(n10437), .c(n10429) );
in01f01  g3712 ( .o(n10442), .a(net_7128) );
in01f01  g3713 ( .o(n10443), .a(net_7160) );
oa22f01  g3714 ( .o(n10444), .a(n7740), .b(n10442), .c(n7739), .d(n10443) );
in01f01  g3715 ( .o(n10445), .a(net_7224) );
in01f01  g3716 ( .o(n10446), .a(net_7192) );
oa22f01  g3717 ( .o(n10447), .a(n7745), .b(n10445), .c(n7744), .d(n10446) );
no02f01  g3718 ( .o(n10448), .a(n10447), .b(n10444) );
na02f01  g3719 ( .o(n6119), .a(n10448), .b(n10441) );
in01f01  g3720 ( .o(n10450), .a(_net_7729) );
ao12f01  g3721 ( .o(n6124), .a(n7343), .b(n10450), .c(n8419) );
no02f01  g3722 ( .o(n10452), .a(n6736_1), .b(n6734) );
in01f01  g3723 ( .o(n10453), .a(_net_264) );
no02f01  g3724 ( .o(n8038), .a(n8236), .b(n10453) );
in01f01  g3725 ( .o(n10455), .a(n8038) );
na02f01  g3726 ( .o(n10456), .a(_net_289), .b(n10453) );
oa22f01  g3727 ( .o(n6140), .a(n10456), .b(n6735), .c(n10455), .d(n10452) );
in01f01  g3728 ( .o(n10458), .a(_net_6292) );
no02f01  g3729 ( .o(n6153), .a(_net_392), .b(n10458) );
in01f01  g3730 ( .o(n10460), .a(_net_6208) );
no02f01  g3731 ( .o(n6166), .a(_net_392), .b(n10460) );
oa12f01  g3732 ( .o(n10462), .a(n8028_1), .b(n9180), .c(n9177) );
na02f01  g3733 ( .o(n10463), .a(n9832), .b(n9831) );
ao22f01  g3734 ( .o(n10464), .a(n10463), .b(n8033_1), .c(n8034), .d(_net_6071) );
na02f01  g3735 ( .o(n10465), .a(n9050), .b(n9049) );
ao22f01  g3736 ( .o(n10466), .a(n10465), .b(n8113), .c(n8031), .d(n8110) );
na03f01  g3737 ( .o(n6171), .a(n10466), .b(n10464), .c(n10462) );
na02f01  g3738 ( .o(n10468), .a(n8211_1), .b(_net_6124) );
na02f01  g3739 ( .o(n10469), .a(n9658), .b(n8213) );
na02f01  g3740 ( .o(n6186), .a(n10469), .b(n10468) );
ao22f01  g3741 ( .o(n10471), .a(n7000_1), .b(net_6969), .c(n6999), .d(net_7033) );
ao22f01  g3742 ( .o(n10472), .a(n7003), .b(net_7001), .c(n7002), .d(net_7065) );
na02f01  g3743 ( .o(n10473), .a(n10472), .b(n10471) );
na02f01  g3744 ( .o(n10474), .a(n10473), .b(n6981) );
ao22f01  g3745 ( .o(n10475), .a(n7323), .b(n6998), .c(n6996), .d(_net_6149) );
na02f01  g3746 ( .o(n10476), .a(n7327), .b(n7013_1) );
oa12f01  g3747 ( .o(n10477), .a(n7022), .b(n8478), .c(n8475) );
na04f01  g3748 ( .o(n6191), .a(n10477), .b(n10476), .c(n10475), .d(n10474) );
in01f01  g3749 ( .o(n10479), .a(_net_7693) );
na02f01  g3750 ( .o(n10480), .a(n7207_1), .b(_net_7795) );
oa12f01  g3751 ( .o(n6200), .a(n10480), .b(n7207_1), .c(n10479) );
in01f01  g3752 ( .o(n10482), .a(_net_7254) );
na02f01  g3753 ( .o(n10483), .a(n8960), .b(n6901) );
oa12f01  g3754 ( .o(n6209), .a(n10483), .b(n6901), .c(n10482) );
no02f01  g3755 ( .o(n10485), .a(n7822_1), .b(n6945) );
no02f01  g3756 ( .o(n10486), .a(n8746), .b(n6934_1) );
in01f01  g3757 ( .o(n10487), .a(_net_6099) );
in01f01  g3758 ( .o(n10488), .a(net_6574) );
in01f01  g3759 ( .o(n10489), .a(net_6638) );
oa22f01  g3760 ( .o(n10490), .a(n6922), .b(n10488), .c(n6919_1), .d(n10489) );
in01f01  g3761 ( .o(n10491), .a(net_6606) );
in01f01  g3762 ( .o(n10492), .a(net_6670) );
oa22f01  g3763 ( .o(n10493), .a(n6927), .b(n10491), .c(n6925), .d(n10492) );
no02f01  g3764 ( .o(n10494), .a(n10493), .b(n10490) );
oa22f01  g3765 ( .o(n10495), .a(n10494), .b(n6916), .c(n6932), .d(n10487) );
no03f01  g3766 ( .o(n10496), .a(n10495), .b(n10486), .c(n10485) );
in01f01  g3767 ( .o(n10497), .a(net_6586) );
in01f01  g3768 ( .o(n10498), .a(net_6618) );
oa22f01  g3769 ( .o(n10499), .a(n7058_1), .b(n10497), .c(n7057), .d(n10498) );
in01f01  g3770 ( .o(n10500), .a(net_6650) );
in01f01  g3771 ( .o(n10501), .a(net_6682) );
oa22f01  g3772 ( .o(n10502), .a(n7063), .b(n10501), .c(n7062_1), .d(n10500) );
no02f01  g3773 ( .o(n10503), .a(n10502), .b(n10499) );
na02f01  g3774 ( .o(n6218), .a(n10503), .b(n10496) );
ao22f01  g3775 ( .o(n10505), .a(n6877), .b(_net_7280), .c(n6876_1), .d(net_7344) );
ao22f01  g3776 ( .o(n10506), .a(n6881_1), .b(net_7312), .c(n6880), .d(net_7376) );
na02f01  g3777 ( .o(n6227), .a(n10506), .b(n10505) );
ao22f01  g3778 ( .o(n10508), .a(n7225), .b(_net_7418), .c(n7224), .d(_net_7450) );
ao22f01  g3779 ( .o(n10509), .a(n7229), .b(_net_7514), .c(n7228), .d(_net_7482) );
na02f01  g3780 ( .o(n6244), .a(n10509), .b(n10508) );
ao22f01  g3781 ( .o(n10511), .a(n7225), .b(_net_7409), .c(n7224), .d(_net_7441) );
ao22f01  g3782 ( .o(n10512), .a(n7229), .b(_net_7505), .c(n7228), .d(_net_7473) );
na02f01  g3783 ( .o(n6249), .a(n10512), .b(n10511) );
in01f01  g3784 ( .o(n10514), .a(_net_7434) );
na02f01  g3785 ( .o(n10515), .a(n7883_1), .b(n7197) );
oa12f01  g3786 ( .o(n6266), .a(n10515), .b(n7197), .c(n10514) );
ao22f01  g3787 ( .o(n10517), .a(n6877), .b(_net_7261), .c(n6876_1), .d(_net_7325) );
ao22f01  g3788 ( .o(n10518), .a(n6881_1), .b(_net_7293), .c(n6880), .d(_net_7357) );
na02f01  g3789 ( .o(n6271), .a(n10518), .b(n10517) );
ao22f01  g3790 ( .o(n10520), .a(n6877), .b(_net_7268), .c(n6876_1), .d(_net_7332) );
ao22f01  g3791 ( .o(n10521), .a(n6881_1), .b(_net_7300), .c(n6880), .d(_net_7364) );
na02f01  g3792 ( .o(n6281), .a(n10521), .b(n10520) );
ao22f01  g3793 ( .o(n10523), .a(n7298), .b(_net_7723), .c(n7288_1), .d(_net_6031) );
ao22f01  g3794 ( .o(n10524), .a(n7306), .b(_net_5987), .c(n7286), .d(_net_270) );
na02f01  g3795 ( .o(n10525), .a(n7302_1), .b(_net_117) );
na03f01  g3796 ( .o(n10526), .a(n7308), .b(net_159), .c(n6800) );
na03f01  g3797 ( .o(n10527), .a(n7308), .b(net_196), .c(x1322) );
na02f01  g3798 ( .o(n10528), .a(n7296), .b(net_233) );
na03f01  g3799 ( .o(n10529), .a(n10528), .b(n10527), .c(n10526) );
ao12f01  g3800 ( .o(n10530), .a(n10529), .b(n7291), .c(_net_7694) );
na04f01  g3801 ( .o(n6290), .a(n10530), .b(n10525), .c(n10524), .d(n10523) );
in01f01  g3802 ( .o(n10532), .a(_net_7787) );
no04f01  g3803 ( .o(n10533), .a(n7360), .b(n7355), .c(n10532), .d(n7359_1) );
no02f01  g3804 ( .o(n10534), .a(n10533), .b(_net_7789) );
in01f01  g3805 ( .o(n10535), .a(_net_7789) );
in01f01  g3806 ( .o(n10536), .a(n10533) );
no02f01  g3807 ( .o(n10537), .a(n10536), .b(n10535) );
no03f01  g3808 ( .o(n6294), .a(n10537), .b(n10534), .c(n7358) );
ao12f01  g3809 ( .o(n10539), .a(n8330), .b(_net_6555), .c(_net_6558) );
oa12f01  g3810 ( .o(n10540), .a(n10539), .b(_net_6555), .c(_net_6558) );
na02f01  g3811 ( .o(n10541), .a(n8472), .b(n9269) );
oa12f01  g3812 ( .o(n6311), .a(n8366), .b(n10541), .c(n10540) );
in01f01  g3813 ( .o(n10543), .a(_net_6001) );
na02f01  g3814 ( .o(n10544), .a(n7348), .b(net_7807) );
oa12f01  g3815 ( .o(n6324), .a(n10544), .b(n7348), .c(n10543) );
no02f01  g3816 ( .o(n10546), .a(n8104), .b(n8101) );
no02f01  g3817 ( .o(n10547), .a(n10546), .b(n6764) );
in01f01  g3818 ( .o(n10548), .a(net_6432) );
in01f01  g3819 ( .o(n10549), .a(net_6496) );
oa22f01  g3820 ( .o(n10550), .a(n6750), .b(n10548), .c(n6748), .d(n10549) );
in01f01  g3821 ( .o(n10551), .a(net_6528) );
in01f01  g3822 ( .o(n10552), .a(net_6464) );
oa22f01  g3823 ( .o(n10553), .a(n6755), .b(n10552), .c(n6754), .d(n10551) );
no02f01  g3824 ( .o(n10554), .a(n10553), .b(n10550) );
no02f01  g3825 ( .o(n10555), .a(n10554), .b(n6766) );
in01f01  g3826 ( .o(n10556), .a(_net_6074) );
oa22f01  g3827 ( .o(n10557), .a(n9225_1), .b(n6775), .c(n6784), .d(n10556) );
no03f01  g3828 ( .o(n10558), .a(n10557), .b(n10555), .c(n10547) );
in01f01  g3829 ( .o(n10559), .a(net_6478) );
in01f01  g3830 ( .o(n10560), .a(net_6446) );
oa22f01  g3831 ( .o(n10561), .a(n6790), .b(n10560), .c(n6789), .d(n10559) );
in01f01  g3832 ( .o(n10562), .a(net_6510) );
in01f01  g3833 ( .o(n10563), .a(net_6542) );
oa22f01  g3834 ( .o(n10564), .a(n6795), .b(n10563), .c(n6794), .d(n10562) );
no02f01  g3835 ( .o(n10565), .a(n10564), .b(n10561) );
na02f01  g3836 ( .o(n6337), .a(n10565), .b(n10558) );
in01f01  g3837 ( .o(n10567), .a(_net_7353) );
na02f01  g3838 ( .o(n10568), .a(n9587), .b(n7030) );
oa12f01  g3839 ( .o(n6346), .a(n10568), .b(n7030), .c(n10567) );
in01f01  g3840 ( .o(n10570), .a(_net_7440) );
na02f01  g3841 ( .o(n10571), .a(n8141), .b(n7197) );
oa12f01  g3842 ( .o(n6362), .a(n10571), .b(n7197), .c(n10570) );
in01f01  g3843 ( .o(n10573), .a(_net_7098) );
in01f01  g3844 ( .o(n10574), .a(n2590) );
ao12f01  g3845 ( .o(n10575), .a(n10573), .b(_net_7097), .c(net_7096) );
no03f01  g3846 ( .o(n10576), .a(n8760), .b(_net_7098), .c(n8385) );
no02f01  g3847 ( .o(n10577), .a(n10576), .b(n10575) );
na02f01  g3848 ( .o(n10578), .a(_net_6028), .b(n8650_1) );
oa22f01  g3849 ( .o(n6371), .a(n10578), .b(n10573), .c(n10577), .d(n10574) );
in01f01  g3850 ( .o(n10580), .a(_net_7661) );
na02f01  g3851 ( .o(n10581), .a(n7446_1), .b(n7428) );
oa12f01  g3852 ( .o(n6381), .a(n10581), .b(n7446_1), .c(n10580) );
no02f01  g3853 ( .o(n10583), .a(n8746), .b(n6945) );
no02f01  g3854 ( .o(n10584), .a(n10494), .b(n6934_1) );
in01f01  g3855 ( .o(n10585), .a(_net_6101) );
in01f01  g3856 ( .o(n10586), .a(net_6576) );
in01f01  g3857 ( .o(n10587), .a(net_6640) );
oa22f01  g3858 ( .o(n10588), .a(n6922), .b(n10586), .c(n6919_1), .d(n10587) );
in01f01  g3859 ( .o(n10589), .a(net_6608) );
in01f01  g3860 ( .o(n10590), .a(net_6672) );
oa22f01  g3861 ( .o(n10591), .a(n6927), .b(n10589), .c(n6925), .d(n10590) );
no02f01  g3862 ( .o(n10592), .a(n10591), .b(n10588) );
oa22f01  g3863 ( .o(n10593), .a(n10592), .b(n6916), .c(n6932), .d(n10585) );
no03f01  g3864 ( .o(n10594), .a(n10593), .b(n10584), .c(n10583) );
in01f01  g3865 ( .o(n10595), .a(net_6588) );
in01f01  g3866 ( .o(n10596), .a(net_6620) );
oa22f01  g3867 ( .o(n10597), .a(n7058_1), .b(n10595), .c(n7057), .d(n10596) );
in01f01  g3868 ( .o(n10598), .a(net_6652) );
in01f01  g3869 ( .o(n10599), .a(net_6684) );
oa22f01  g3870 ( .o(n10600), .a(n7063), .b(n10599), .c(n7062_1), .d(n10598) );
no02f01  g3871 ( .o(n10601), .a(n10600), .b(n10597) );
na02f01  g3872 ( .o(n6395), .a(n10601), .b(n10594) );
in01f01  g3873 ( .o(n10603), .a(_net_7438) );
na02f01  g3874 ( .o(n10604), .a(n7860), .b(n7197) );
oa12f01  g3875 ( .o(n6411), .a(n10604), .b(n7197), .c(n10603) );
ao22f01  g3876 ( .o(n10606), .a(n6877), .b(_net_7250), .c(n6876_1), .d(_net_7314) );
ao22f01  g3877 ( .o(n10607), .a(n6881_1), .b(_net_7282), .c(n6880), .d(_net_7346) );
na02f01  g3878 ( .o(n6432), .a(n10607), .b(n10606) );
no02f01  g3879 ( .o(n10609), .a(_net_6692), .b(n7153) );
no02f01  g3880 ( .o(n10610), .a(n7663), .b(net_6691) );
no02f01  g3881 ( .o(n10611), .a(n10610), .b(n10609) );
oa22f01  g3882 ( .o(n6450), .a(n10611), .b(n9974), .c(n9978), .d(n7663) );
in01f01  g3883 ( .o(n10613), .a(_net_7257) );
na02f01  g3884 ( .o(n10614), .a(n9587), .b(n6901) );
oa12f01  g3885 ( .o(n6455), .a(n10614), .b(n6901), .c(n10613) );
ao22f01  g3886 ( .o(n10616), .a(n7225), .b(_net_7413), .c(n7224), .d(_net_7445) );
ao22f01  g3887 ( .o(n10617), .a(n7229), .b(_net_7509), .c(n7228), .d(_net_7477) );
na02f01  g3888 ( .o(n6493), .a(n10617), .b(n10616) );
in01f01  g3889 ( .o(n10619), .a(_net_5857) );
in01f01  g3890 ( .o(n10620), .a(x1034) );
in01f01  g3891 ( .o(n10621), .a(_net_5999) );
no02f01  g3892 ( .o(n10622), .a(n10621), .b(_net_6000) );
na02f01  g3893 ( .o(n10623), .a(_net_5995), .b(_net_6001) );
ao12f01  g3894 ( .o(n10624), .a(n10623), .b(n7191), .c(_net_5966) );
na02f01  g3895 ( .o(n10625), .a(n10624), .b(n10622) );
in01f01  g3896 ( .o(n10626), .a(n10623) );
na03f01  g3897 ( .o(n10627), .a(n7191), .b(_net_5966), .c(_net_5965) );
na04f01  g3898 ( .o(n10628), .a(n10627), .b(n10626), .c(n10621), .d(n7673) );
oa12f01  g3899 ( .o(n10629), .a(n7191), .b(_net_5966), .c(_net_5965) );
na04f01  g3900 ( .o(n10630), .a(n10629), .b(n10626), .c(n10621), .d(_net_6000) );
no02f01  g3901 ( .o(n10631), .a(n10621), .b(n7673) );
na03f01  g3902 ( .o(n10632), .a(n10631), .b(n10626), .c(_net_5964) );
na04f01  g3903 ( .o(n10633), .a(n10632), .b(n10630), .c(n10628), .d(n10625) );
na03f01  g3904 ( .o(n10634), .a(n10633), .b(net_7773), .c(n10620) );
oa12f01  g3905 ( .o(n6527), .a(n10634), .b(n10619), .c(x1034) );
na02f01  g3906 ( .o(n10636), .a(n9211_1), .b(n8213) );
ao22f01  g3907 ( .o(n10637), .a(n9658), .b(n9200), .c(n8211_1), .d(_net_6126) );
na02f01  g3908 ( .o(n6540), .a(n10637), .b(n10636) );
in01f01  g3909 ( .o(n10639), .a(_net_118) );
na02f01  g3910 ( .o(n10640), .a(net_314), .b(_net_154) );
oa12f01  g3911 ( .o(n6545), .a(n10640), .b(n10639), .c(_net_154) );
in01f01  g3912 ( .o(n10642), .a(_net_7654) );
na02f01  g3913 ( .o(n10643), .a(n7644_1), .b(n7446_1) );
oa12f01  g3914 ( .o(n6558), .a(n10643), .b(n7446_1), .c(n10642) );
na02f01  g3915 ( .o(n10645), .a(n7009_1), .b(n6981) );
ao22f01  g3916 ( .o(n10646), .a(n9719_1), .b(n6998), .c(n6996), .d(_net_6146) );
na02f01  g3917 ( .o(n6570), .a(n10646), .b(n10645) );
na03f01  g3918 ( .o(n10648), .a(_net_6407), .b(_net_6405), .c(_net_6406) );
no02f01  g3919 ( .o(n10649), .a(n8087), .b(_net_6411) );
ao12f01  g3920 ( .o(n6583), .a(n8177), .b(n10649), .c(n10648) );
ao22f01  g3921 ( .o(n10651), .a(n6877), .b(_net_7251), .c(n6876_1), .d(_net_7315) );
ao22f01  g3922 ( .o(n10652), .a(n6881_1), .b(_net_7283), .c(n6880), .d(_net_7347) );
na02f01  g3923 ( .o(n6591), .a(n10652), .b(n10651) );
in01f01  g3924 ( .o(n10654), .a(net_6769) );
in01f01  g3925 ( .o(n10655), .a(net_6705) );
oa22f01  g3926 ( .o(n10656), .a(n7129), .b(n10655), .c(n7126), .d(n10654) );
in01f01  g3927 ( .o(n10657), .a(net_6737) );
in01f01  g3928 ( .o(n10658), .a(net_6801) );
oa22f01  g3929 ( .o(n10659), .a(n7134), .b(n10657), .c(n7132), .d(n10658) );
no02f01  g3930 ( .o(n10660), .a(n10659), .b(n10656) );
no02f01  g3931 ( .o(n10661), .a(n10660), .b(n7468_1) );
no02f01  g3932 ( .o(n10662), .a(n8665), .b(n7470) );
in01f01  g3933 ( .o(n10663), .a(_net_6119) );
oa22f01  g3934 ( .o(n10664), .a(n8673), .b(n7123), .c(n7118), .d(n10663) );
no03f01  g3935 ( .o(n10665), .a(n10664), .b(n10662), .c(n10661) );
in01f01  g3936 ( .o(n10666), .a(net_6721) );
in01f01  g3937 ( .o(n10667), .a(net_6753) );
oa22f01  g3938 ( .o(n10668), .a(n7492_1), .b(n10666), .c(n7491), .d(n10667) );
in01f01  g3939 ( .o(n10669), .a(net_6817) );
in01f01  g3940 ( .o(n10670), .a(net_6785) );
oa22f01  g3941 ( .o(n10671), .a(n7497), .b(n10669), .c(n7496_1), .d(n10670) );
no02f01  g3942 ( .o(n10672), .a(n10671), .b(n10668) );
na02f01  g3943 ( .o(n6596), .a(n10672), .b(n10665) );
in01f01  g3944 ( .o(n10674), .a(_net_7448) );
na02f01  g3945 ( .o(n10675), .a(n7638), .b(n7197) );
oa12f01  g3946 ( .o(n6601), .a(n10675), .b(n7197), .c(n10674) );
na02f01  g3947 ( .o(n10677), .a(n9518), .b(_net_7098) );
na03f01  g3948 ( .o(n10678), .a(n9517_1), .b(n9516), .c(n10573) );
na02f01  g3949 ( .o(n10679), .a(n8199), .b(net_7096) );
na03f01  g3950 ( .o(n10680), .a(n8198), .b(n8197_1), .c(n8385) );
ao22f01  g3951 ( .o(n10681), .a(n10680), .b(n10679), .c(n7011), .d(_net_7092) );
na02f01  g3952 ( .o(n10682), .a(n7214), .b(n8760) );
na03f01  g3953 ( .o(n10683), .a(n7213), .b(n7211), .c(_net_7097) );
na03f01  g3954 ( .o(n10684), .a(n10683), .b(n10682), .c(n10681) );
ao12f01  g3955 ( .o(n6606), .a(n10684), .b(n10678), .c(n10677) );
ao22f01  g3956 ( .o(n10686), .a(n6877), .b(_net_7262), .c(n6876_1), .d(_net_7326) );
ao22f01  g3957 ( .o(n10687), .a(n6881_1), .b(_net_7294), .c(n6880), .d(_net_7358) );
na02f01  g3958 ( .o(n6624), .a(n10687), .b(n10686) );
oa12f01  g3959 ( .o(n10689), .a(n7575), .b(n9756), .c(n9753) );
ao22f01  g3960 ( .o(n10690), .a(n7908), .b(n7593), .c(n7591_1), .d(_net_6170) );
na02f01  g3961 ( .o(n10691), .a(n7732_1), .b(n7731) );
ao22f01  g3962 ( .o(n10692), .a(n7912), .b(n7914), .c(n7920_1), .d(n10691) );
na03f01  g3963 ( .o(n6634), .a(n10692), .b(n10690), .c(n10689) );
no03f01  g3964 ( .o(n10694), .a(n6912), .b(_net_5999), .c(n7673) );
no02f01  g3965 ( .o(n10695), .a(n7191), .b(n6912) );
ao22f01  g3966 ( .o(n10696), .a(n10695), .b(n10631), .c(n10694), .d(n10629) );
ao12f01  g3967 ( .o(n10697), .a(n6912), .b(n7191), .c(_net_5966) );
no03f01  g3968 ( .o(n10698), .a(n6912), .b(_net_5999), .c(_net_6000) );
ao22f01  g3969 ( .o(n10699), .a(n10698), .b(n10627), .c(n10697), .d(n10622) );
na02f01  g3970 ( .o(n6643), .a(n10699), .b(n10696) );
in01f01  g3971 ( .o(n10701), .a(_net_124) );
na02f01  g3972 ( .o(n10702), .a(net_320), .b(_net_154) );
oa12f01  g3973 ( .o(n6652), .a(n10702), .b(n10701), .c(_net_154) );
na02f01  g3974 ( .o(n10704), .a(n6817), .b(n6812) );
na02f01  g3975 ( .o(n10705), .a(n8213), .b(n10704) );
ao22f01  g3976 ( .o(n10706), .a(n6811), .b(net_6832), .c(n6808), .d(net_6896) );
ao22f01  g3977 ( .o(n10707), .a(n6816), .b(net_6864), .c(n6814), .d(net_6928) );
na02f01  g3978 ( .o(n10708), .a(n10707), .b(n10706) );
ao22f01  g3979 ( .o(n10709), .a(n10708), .b(n9200), .c(n8211_1), .d(_net_6129) );
na02f01  g3980 ( .o(n10710), .a(n8216_1), .b(n9205) );
in01f01  g3981 ( .o(n10711), .a(net_6846) );
in01f01  g3982 ( .o(n10712), .a(net_6910) );
oa22f01  g3983 ( .o(n10713), .a(n6810), .b(n10711), .c(n6807), .d(n10712) );
in01f01  g3984 ( .o(n10714), .a(net_6942) );
in01f01  g3985 ( .o(n10715), .a(net_6878) );
oa22f01  g3986 ( .o(n10716), .a(n6815), .b(n10715), .c(n6813_1), .d(n10714) );
oa12f01  g3987 ( .o(n10717), .a(n9207), .b(n10716), .c(n10713) );
na04f01  g3988 ( .o(n6665), .a(n10717), .b(n10710), .c(n10709), .d(n10705) );
na02f01  g3989 ( .o(n10719), .a(n7440), .b(_net_7801) );
oa12f01  g3990 ( .o(n6682), .a(n10719), .b(n7440), .c(n7850) );
ao22f01  g3991 ( .o(n10721), .a(n7288_1), .b(_net_6033), .c(n7286), .d(_net_272) );
ao22f01  g3992 ( .o(n10722), .a(n7298), .b(_net_7725), .c(n7291), .d(_net_7696) );
na02f01  g3993 ( .o(n10723), .a(n7302_1), .b(_net_119) );
na03f01  g3994 ( .o(n10724), .a(n7308), .b(net_198), .c(x1322) );
na02f01  g3995 ( .o(n10725), .a(n7296), .b(net_235) );
na03f01  g3996 ( .o(n10726), .a(n7308), .b(net_161), .c(n6800) );
na03f01  g3997 ( .o(n10727), .a(n10726), .b(n10725), .c(n10724) );
ao12f01  g3998 ( .o(n10728), .a(n10727), .b(n7306), .c(_net_5989) );
na04f01  g3999 ( .o(n6691), .a(n10728), .b(n10723), .c(n10722), .d(n10721) );
in01f01  g4000 ( .o(n10730), .a(_net_7623) );
na02f01  g4001 ( .o(n10731), .a(n9493), .b(n7400_1) );
oa12f01  g4002 ( .o(n6695), .a(n10731), .b(n7400_1), .c(n10730) );
in01f01  g4003 ( .o(n10733), .a(_net_7279) );
na02f01  g4004 ( .o(n10734), .a(n1034), .b(n6901) );
oa12f01  g4005 ( .o(n6709), .a(n10734), .b(n6901), .c(n10733) );
ao22f01  g4006 ( .o(n10736), .a(n7130), .b(net_6699), .c(n7127), .d(net_6763) );
ao22f01  g4007 ( .o(n10737), .a(n7135), .b(net_6731), .c(n7133_1), .d(net_6795) );
ao12f01  g4008 ( .o(n10738), .a(n7468_1), .b(n10737), .c(n10736) );
in01f01  g4009 ( .o(n10739), .a(net_6765) );
in01f01  g4010 ( .o(n10740), .a(net_6701) );
oa22f01  g4011 ( .o(n10741), .a(n7129), .b(n10740), .c(n7126), .d(n10739) );
in01f01  g4012 ( .o(n10742), .a(net_6733) );
in01f01  g4013 ( .o(n10743), .a(net_6797) );
oa22f01  g4014 ( .o(n10744), .a(n7134), .b(n10742), .c(n7132), .d(n10743) );
no02f01  g4015 ( .o(n10745), .a(n10744), .b(n10741) );
no02f01  g4016 ( .o(n10746), .a(n10745), .b(n7470) );
in01f01  g4017 ( .o(n10747), .a(_net_6113) );
in01f01  g4018 ( .o(n10748), .a(net_6767) );
in01f01  g4019 ( .o(n10749), .a(net_6703) );
oa22f01  g4020 ( .o(n10750), .a(n7129), .b(n10749), .c(n7126), .d(n10748) );
in01f01  g4021 ( .o(n10751), .a(net_6799) );
in01f01  g4022 ( .o(n10752), .a(net_6735) );
oa22f01  g4023 ( .o(n10753), .a(n7134), .b(n10752), .c(n7132), .d(n10751) );
no02f01  g4024 ( .o(n10754), .a(n10753), .b(n10750) );
oa22f01  g4025 ( .o(n10755), .a(n10754), .b(n7123), .c(n7118), .d(n10747) );
no03f01  g4026 ( .o(n10756), .a(n10755), .b(n10746), .c(n10738) );
in01f01  g4027 ( .o(n10757), .a(net_6747) );
in01f01  g4028 ( .o(n10758), .a(net_6715) );
oa22f01  g4029 ( .o(n10759), .a(n7492_1), .b(n10758), .c(n7491), .d(n10757) );
in01f01  g4030 ( .o(n10760), .a(net_6779) );
in01f01  g4031 ( .o(n10761), .a(net_6811) );
oa22f01  g4032 ( .o(n10762), .a(n7497), .b(n10761), .c(n7496_1), .d(n10760) );
no02f01  g4033 ( .o(n10763), .a(n10762), .b(n10759) );
na02f01  g4034 ( .o(n6727), .a(n10763), .b(n10756) );
in01f01  g4035 ( .o(n10765), .a(_net_7620) );
na02f01  g4036 ( .o(n10766), .a(n8426_1), .b(n7400_1) );
oa12f01  g4037 ( .o(n6741), .a(n10766), .b(n7400_1), .c(n10765) );
no02f01  g4038 ( .o(n10768), .a(n8443_1), .b(n6824) );
no02f01  g4039 ( .o(n10769), .a(n8452), .b(n6826_1) );
in01f01  g4040 ( .o(n10770), .a(_net_6136) );
oa22f01  g4041 ( .o(n10771), .a(n10249), .b(n6836_1), .c(n6844), .d(n10770) );
no03f01  g4042 ( .o(n10772), .a(n10771), .b(n10769), .c(n10768) );
in01f01  g4043 ( .o(n10773), .a(net_6885) );
in01f01  g4044 ( .o(n10774), .a(net_6853) );
oa22f01  g4045 ( .o(n10775), .a(n6850_1), .b(n10774), .c(n6849), .d(n10773) );
in01f01  g4046 ( .o(n10776), .a(net_6949) );
in01f01  g4047 ( .o(n10777), .a(net_6917) );
oa22f01  g4048 ( .o(n10778), .a(n6855_1), .b(n10776), .c(n6854), .d(n10777) );
no02f01  g4049 ( .o(n10779), .a(n10778), .b(n10775) );
na02f01  g4050 ( .o(n6765), .a(n10779), .b(n10772) );
no02f01  g4051 ( .o(n10781), .a(n10754), .b(n7468_1) );
no02f01  g4052 ( .o(n10782), .a(n10660), .b(n7470) );
in01f01  g4053 ( .o(n10783), .a(_net_6117) );
oa22f01  g4054 ( .o(n10784), .a(n8665), .b(n7123), .c(n7118), .d(n10783) );
no03f01  g4055 ( .o(n10785), .a(n10784), .b(n10782), .c(n10781) );
in01f01  g4056 ( .o(n10786), .a(net_6751) );
in01f01  g4057 ( .o(n10787), .a(net_6719) );
oa22f01  g4058 ( .o(n10788), .a(n7492_1), .b(n10787), .c(n7491), .d(n10786) );
in01f01  g4059 ( .o(n10789), .a(net_6783) );
in01f01  g4060 ( .o(n10790), .a(net_6815) );
oa22f01  g4061 ( .o(n10791), .a(n7497), .b(n10790), .c(n7496_1), .d(n10789) );
no02f01  g4062 ( .o(n10792), .a(n10791), .b(n10788) );
na02f01  g4063 ( .o(n6774), .a(n10792), .b(n10785) );
in01f01  g4064 ( .o(n10794), .a(_net_7723) );
in01f01  g4065 ( .o(n10795), .a(_net_5993) );
ao12f01  g4066 ( .o(n6779), .a(n7343), .b(n10795), .c(n10794) );
in01f01  g4067 ( .o(n10797), .a(_net_7446) );
na02f01  g4068 ( .o(n10798), .a(n8994), .b(n7197) );
oa12f01  g4069 ( .o(n6788), .a(n10798), .b(n7197), .c(n10797) );
in01f01  g4070 ( .o(n10800), .a(_net_7258) );
na02f01  g4071 ( .o(n10801), .a(n7393), .b(n6901) );
oa12f01  g4072 ( .o(n6801), .a(n10801), .b(n6901), .c(n10800) );
in01f01  g4073 ( .o(n10803), .a(_net_7700) );
na02f01  g4074 ( .o(n10804), .a(n7207_1), .b(net_7802) );
oa12f01  g4075 ( .o(n6818), .a(n10804), .b(n7207_1), .c(n10803) );
in01f01  g4076 ( .o(n10806), .a(_net_7584) );
na02f01  g4077 ( .o(n10807), .a(n8842), .b(n6968) );
oa12f01  g4078 ( .o(n6831), .a(n10807), .b(n6968), .c(n10806) );
oa12f01  g4079 ( .o(n6840), .a(n10795), .b(n6761_1), .c(n7533) );
in01f01  g4080 ( .o(n10810), .a(_net_7325) );
na02f01  g4081 ( .o(n10811), .a(n8809_1), .b(n7150) );
oa12f01  g4082 ( .o(n6845), .a(n10811), .b(n7150), .c(n10810) );
ao22f01  g4083 ( .o(n10813), .a(n6736_1), .b(_net_7626), .c(n6734), .d(_net_7594) );
ao22f01  g4084 ( .o(n10814), .a(n6739), .b(_net_7658), .c(n6738), .d(_net_7562) );
na02f01  g4085 ( .o(n6850), .a(n10814), .b(n10813) );
in01f01  g4086 ( .o(n10816), .a(_net_5990) );
na02f01  g4087 ( .o(n10817), .a(n7348), .b(net_7799) );
oa12f01  g4088 ( .o(n6855), .a(n10817), .b(n7348), .c(n10816) );
ao22f01  g4089 ( .o(n10819), .a(n7225), .b(_net_7424), .c(n7224), .d(net_7456) );
ao22f01  g4090 ( .o(n10820), .a(n7229), .b(net_7520), .c(n7228), .d(net_7488) );
na02f01  g4091 ( .o(n6872), .a(n10820), .b(n10819) );
no02f01  g4092 ( .o(n10822), .a(n9934), .b(n7012) );
no02f01  g4093 ( .o(n10823), .a(n8471), .b(n6997) );
in01f01  g4094 ( .o(n10824), .a(_net_6161) );
oa22f01  g4095 ( .o(n10825), .a(n8479), .b(n6980), .c(n6995_1), .d(n10824) );
no03f01  g4096 ( .o(n10826), .a(n10825), .b(n10823), .c(n10822) );
in01f01  g4097 ( .o(n10827), .a(net_6993) );
in01f01  g4098 ( .o(n10828), .a(net_7025) );
oa22f01  g4099 ( .o(n10829), .a(n8075_1), .b(n10827), .c(n8074), .d(n10828) );
in01f01  g4100 ( .o(n10830), .a(net_7089) );
in01f01  g4101 ( .o(n10831), .a(net_7057) );
oa22f01  g4102 ( .o(n10832), .a(n8080_1), .b(n10830), .c(n8079), .d(n10831) );
no02f01  g4103 ( .o(n10833), .a(n10832), .b(n10829) );
na02f01  g4104 ( .o(n6881), .a(n10833), .b(n10826) );
in01f01  g4105 ( .o(n10835), .a(_net_7427) );
na02f01  g4106 ( .o(n10836), .a(n1173), .b(n7550) );
oa12f01  g4107 ( .o(n6890), .a(n10836), .b(n7550), .c(n10835) );
ao22f01  g4108 ( .o(n10838), .a(n7225), .b(_net_7423), .c(n7224), .d(net_7455) );
ao22f01  g4109 ( .o(n10839), .a(n7229), .b(net_7519), .c(n7228), .d(net_7487) );
na02f01  g4110 ( .o(n6915), .a(n10839), .b(n10838) );
in01f01  g4111 ( .o(n10841), .a(_net_7443) );
na02f01  g4112 ( .o(n10842), .a(n9786), .b(n7197) );
oa12f01  g4113 ( .o(n6924), .a(n10842), .b(n7197), .c(n10841) );
ao22f01  g4114 ( .o(n10844), .a(n6736_1), .b(_net_7630), .c(n6734), .d(_net_7598) );
ao22f01  g4115 ( .o(n10845), .a(n6739), .b(_net_7662), .c(n6738), .d(_net_7566) );
na02f01  g4116 ( .o(n6929), .a(n10845), .b(n10844) );
in01f01  g4117 ( .o(n10847), .a(_net_114) );
na02f01  g4118 ( .o(n10848), .a(net_310), .b(_net_154) );
oa12f01  g4119 ( .o(n6938), .a(n10848), .b(n10847), .c(_net_154) );
in01f01  g4120 ( .o(n10850), .a(_net_7589) );
na02f01  g4121 ( .o(n10851), .a(n7449), .b(n6968) );
oa12f01  g4122 ( .o(n6943), .a(n10851), .b(n6968), .c(n10850) );
in01f01  g4123 ( .o(n10853), .a(_net_7500) );
na02f01  g4124 ( .o(n10854), .a(n7952), .b(n7626_1) );
oa12f01  g4125 ( .o(n6952), .a(n10854), .b(n7626_1), .c(n10853) );
no02f01  g4126 ( .o(n10856), .a(n10132_1), .b(n6945) );
no02f01  g4127 ( .o(n10857), .a(n7042), .b(n6934_1) );
in01f01  g4128 ( .o(n10858), .a(_net_6098) );
oa22f01  g4129 ( .o(n10859), .a(n7050), .b(n6916), .c(n6932), .d(n10858) );
no03f01  g4130 ( .o(n10860), .a(n10859), .b(n10857), .c(n10856) );
in01f01  g4131 ( .o(n10861), .a(net_6617) );
in01f01  g4132 ( .o(n10862), .a(net_6585) );
oa22f01  g4133 ( .o(n10863), .a(n7058_1), .b(n10862), .c(n7057), .d(n10861) );
in01f01  g4134 ( .o(n10864), .a(net_6681) );
in01f01  g4135 ( .o(n10865), .a(net_6649) );
oa22f01  g4136 ( .o(n10866), .a(n7063), .b(n10864), .c(n7062_1), .d(n10865) );
no02f01  g4137 ( .o(n10867), .a(n10866), .b(n10863) );
na02f01  g4138 ( .o(n6964), .a(n10867), .b(n10860) );
ao22f01  g4139 ( .o(n10869), .a(n7225), .b(_net_7402), .c(n7224), .d(_net_7434) );
ao22f01  g4140 ( .o(n10870), .a(n7229), .b(_net_7498), .c(n7228), .d(_net_7466) );
na02f01  g4141 ( .o(n6969), .a(n10870), .b(n10869) );
in01f01  g4142 ( .o(n10872), .a(_net_7256) );
na02f01  g4143 ( .o(n10873), .a(n8208), .b(n6901) );
oa12f01  g4144 ( .o(n6995), .a(n10873), .b(n6901), .c(n10872) );
na02f01  g4145 ( .o(n10875), .a(n7440), .b(_net_7804) );
oa12f01  g4146 ( .o(n7000), .a(n10875), .b(n7440), .c(n8192_1) );
in01f01  g4147 ( .o(n10877), .a(_net_7408) );
na02f01  g4148 ( .o(n10878), .a(n8141), .b(n7550) );
oa12f01  g4149 ( .o(n7013), .a(n10878), .b(n7550), .c(n10877) );
no02f01  g4150 ( .o(n10880), .a(n10249), .b(n6824) );
no02f01  g4151 ( .o(n10881), .a(n9127), .b(n6826_1) );
in01f01  g4152 ( .o(n10882), .a(_net_6140) );
oa22f01  g4153 ( .o(n10883), .a(n9135), .b(n6836_1), .c(n6844), .d(n10882) );
no03f01  g4154 ( .o(n10884), .a(n10883), .b(n10881), .c(n10880) );
in01f01  g4155 ( .o(n10885), .a(net_6857) );
in01f01  g4156 ( .o(n10886), .a(net_6889) );
oa22f01  g4157 ( .o(n10887), .a(n6850_1), .b(n10885), .c(n6849), .d(n10886) );
in01f01  g4158 ( .o(n10888), .a(net_6953) );
in01f01  g4159 ( .o(n10889), .a(net_6921) );
oa22f01  g4160 ( .o(n10890), .a(n6855_1), .b(n10888), .c(n6854), .d(n10889) );
no02f01  g4161 ( .o(n10891), .a(n10890), .b(n10887) );
na02f01  g4162 ( .o(n7018), .a(n10891), .b(n10884) );
ao22f01  g4163 ( .o(n10893), .a(n7225), .b(_net_7430), .c(n7224), .d(net_7462) );
ao22f01  g4164 ( .o(n10894), .a(n7229), .b(net_7526), .c(n7228), .d(net_7494) );
na02f01  g4165 ( .o(n7023), .a(n10894), .b(n10893) );
in01f01  g4166 ( .o(n10896), .a(_net_7298) );
na02f01  g4167 ( .o(n10897), .a(n7242), .b(n7180) );
oa12f01  g4168 ( .o(n7032), .a(n10897), .b(n7180), .c(n10896) );
in01f01  g4169 ( .o(n10899), .a(_net_7579) );
na02f01  g4170 ( .o(n10900), .a(n1163), .b(n7519) );
oa12f01  g4171 ( .o(n7053), .a(n10900), .b(n7519), .c(n10899) );
in01f01  g4172 ( .o(n10902), .a(_net_7268) );
na02f01  g4173 ( .o(n10903), .a(n7256_1), .b(n6901) );
oa12f01  g4174 ( .o(n7058), .a(n10903), .b(n6901), .c(n10902) );
no02f01  g4175 ( .o(n10905), .a(n7477), .b(n7468_1) );
no02f01  g4176 ( .o(n10906), .a(n7486), .b(n7470) );
in01f01  g4177 ( .o(n10907), .a(_net_6122) );
no02f01  g4178 ( .o(n10908), .a(n8988), .b(n8985) );
oa22f01  g4179 ( .o(n10909), .a(n10908), .b(n7123), .c(n7118), .d(n10907) );
no03f01  g4180 ( .o(n10910), .a(n10909), .b(n10906), .c(n10905) );
in01f01  g4181 ( .o(n10911), .a(net_6724) );
in01f01  g4182 ( .o(n10912), .a(net_6756) );
oa22f01  g4183 ( .o(n10913), .a(n7492_1), .b(n10911), .c(n7491), .d(n10912) );
in01f01  g4184 ( .o(n10914), .a(net_6788) );
in01f01  g4185 ( .o(n10915), .a(net_6820) );
oa22f01  g4186 ( .o(n10916), .a(n7497), .b(n10915), .c(n7496_1), .d(n10914) );
no02f01  g4187 ( .o(n10917), .a(n10916), .b(n10913) );
na02f01  g4188 ( .o(n7067), .a(n10917), .b(n10910) );
no02f01  g4189 ( .o(n7072), .a(n6896), .b(n6895_1) );
in01f01  g4190 ( .o(n10920), .a(_net_6284) );
no02f01  g4191 ( .o(n7077), .a(_net_392), .b(n10920) );
ao22f01  g4192 ( .o(n10922), .a(n7225), .b(_net_7401), .c(n7224), .d(_net_7433) );
ao22f01  g4193 ( .o(n10923), .a(n7229), .b(_net_7497), .c(n7228), .d(_net_7465) );
na02f01  g4194 ( .o(n7102), .a(n10923), .b(n10922) );
in01f01  g4195 ( .o(n10925), .a(net_7767) );
na02f01  g4196 ( .o(n10926), .a(net_7769), .b(n8997) );
oa12f01  g4197 ( .o(n7107), .a(n10926), .b(n10206), .c(n10925) );
in01f01  g4198 ( .o(n10928), .a(_net_7705) );
na02f01  g4199 ( .o(n10929), .a(n7207_1), .b(net_7807) );
oa12f01  g4200 ( .o(n7133), .a(n10929), .b(n7207_1), .c(n10928) );
in01f01  g4201 ( .o(n10931), .a(_net_5848) );
ao12f01  g4202 ( .o(n7138), .a(n10925), .b(n10206), .c(n10931) );
na02f01  g4203 ( .o(n10933), .a(n7291), .b(_net_7719) );
na02f01  g4204 ( .o(n10934), .a(n7293), .b(_net_221) );
ao22f01  g4205 ( .o(n10935), .a(n7297_1), .b(_net_184), .c(n7296), .d(net_258) );
ao22f01  g4206 ( .o(n10936), .a(n7306), .b(_net_6021), .c(n7298), .d(_net_7748) );
na04f01  g4207 ( .o(n7164), .a(n10936), .b(n10935), .c(n10934), .d(n10933) );
na02f01  g4208 ( .o(n10938), .a(n6801_1), .b(x1261) );
no02f01  g4209 ( .o(n7172), .a(n10938), .b(n8317) );
ao22f01  g4210 ( .o(n10940), .a(n6877), .b(_net_7255), .c(n6876_1), .d(_net_7319) );
ao22f01  g4211 ( .o(n10941), .a(n6881_1), .b(_net_7287), .c(n6880), .d(_net_7351) );
na02f01  g4212 ( .o(n7177), .a(n10941), .b(n10940) );
na02f01  g4213 ( .o(n10943), .a(n8861), .b(n7768_1) );
na02f01  g4214 ( .o(n10944), .a(n6755), .b(n6748) );
ao22f01  g4215 ( .o(n10945), .a(n10944), .b(n8859), .c(n8862), .d(_net_6554) );
na02f01  g4216 ( .o(n7194), .a(n10945), .b(n10943) );
no02f01  g4217 ( .o(n10947), .a(n9233_1), .b(n6764) );
no02f01  g4218 ( .o(n10948), .a(n6766), .b(n6757) );
in01f01  g4219 ( .o(n10949), .a(_net_6080) );
oa22f01  g4220 ( .o(n10950), .a(n6784), .b(n10949), .c(n6775), .d(n6773) );
no03f01  g4221 ( .o(n10951), .a(n10950), .b(n10948), .c(n10947) );
in01f01  g4222 ( .o(n10952), .a(net_6452) );
in01f01  g4223 ( .o(n10953), .a(net_6484) );
oa22f01  g4224 ( .o(n10954), .a(n6790), .b(n10952), .c(n6789), .d(n10953) );
in01f01  g4225 ( .o(n10955), .a(net_6548) );
in01f01  g4226 ( .o(n10956), .a(net_6516) );
oa22f01  g4227 ( .o(n10957), .a(n6795), .b(n10955), .c(n6794), .d(n10956) );
no02f01  g4228 ( .o(n10958), .a(n10957), .b(n10954) );
na02f01  g4229 ( .o(n7207), .a(n10958), .b(n10951) );
in01f01  g4230 ( .o(n10960), .a(_net_7361) );
na02f01  g4231 ( .o(n10961), .a(n9537_1), .b(n7030) );
oa12f01  g4232 ( .o(n7216), .a(n10961), .b(n7030), .c(n10960) );
in01f01  g4233 ( .o(n10963), .a(_net_6210) );
no02f01  g4234 ( .o(n7221), .a(_net_392), .b(n10963) );
in01f01  g4235 ( .o(n10965), .a(_net_6239) );
no02f01  g4236 ( .o(n7226), .a(_net_392), .b(n10965) );
in01f01  g4237 ( .o(n10967), .a(_net_6294) );
no02f01  g4238 ( .o(n7235), .a(_net_392), .b(n10967) );
na02f01  g4239 ( .o(n10969), .a(n6996), .b(_net_6145) );
na02f01  g4240 ( .o(n10970), .a(n7327), .b(n6981) );
na02f01  g4241 ( .o(n7240), .a(n10970), .b(n10969) );
na02f01  g4242 ( .o(n10972), .a(n9667), .b(n9404) );
na03f01  g4243 ( .o(n10973), .a(n9665), .b(_net_6423), .c(_net_6422) );
na03f01  g4244 ( .o(n10974), .a(n10973), .b(n10972), .c(n9410_1) );
oa12f01  g4245 ( .o(n7245), .a(n10974), .b(n9409), .c(n9404) );
oa12f01  g4246 ( .o(n10977), .a(n6981), .b(n8051_1), .c(n8048) );
ao22f01  g4247 ( .o(n10978), .a(n10473), .b(n6998), .c(n6996), .d(_net_6151) );
na02f01  g4248 ( .o(n10979), .a(n8482), .b(n8481_1) );
ao22f01  g4249 ( .o(n10980), .a(n10979), .b(n7022), .c(n7323), .d(n7013_1) );
na03f01  g4250 ( .o(n7270), .a(n10980), .b(n10978), .c(n10977) );
in01f01  g4251 ( .o(n10982), .a(_net_6290) );
no02f01  g4252 ( .o(n7275), .a(_net_392), .b(n10982) );
oa12f01  g4253 ( .o(n7280), .a(n7335_1), .b(n6821), .c(n7687) );
na02f01  g4254 ( .o(n10985), .a(n6803), .b(_net_6028) );
oa12f01  g4255 ( .o(n7297), .a(n10985), .b(n6803), .c(n7330_1) );
in01f01  g4256 ( .o(n10987), .a(_net_6287) );
no02f01  g4257 ( .o(n7302), .a(n10987), .b(_net_392) );
in01f01  g4258 ( .o(n10989), .a(_net_7697) );
na02f01  g4259 ( .o(n10990), .a(n7207_1), .b(net_7799) );
oa12f01  g4260 ( .o(n7307), .a(n10990), .b(n7207_1), .c(n10989) );
in01f01  g4261 ( .o(n10992), .a(_net_7365) );
na02f01  g4262 ( .o(n10993), .a(n9685), .b(n7030) );
oa12f01  g4263 ( .o(n7321), .a(n10993), .b(n7030), .c(n10992) );
no02f01  g4264 ( .o(n10995), .a(n8282), .b(n7721) );
no02f01  g4265 ( .o(n10996), .a(n8291), .b(n7592) );
in01f01  g4266 ( .o(n10997), .a(_net_6179) );
oa22f01  g4267 ( .o(n10998), .a(n10436), .b(n7574), .c(n7590), .d(n10997) );
no03f01  g4268 ( .o(n10999), .a(n10998), .b(n10996), .c(n10995) );
in01f01  g4269 ( .o(n11000), .a(net_7126) );
in01f01  g4270 ( .o(n11001), .a(net_7158) );
oa22f01  g4271 ( .o(n11002), .a(n7740), .b(n11000), .c(n7739), .d(n11001) );
in01f01  g4272 ( .o(n11003), .a(net_7222) );
in01f01  g4273 ( .o(n11004), .a(net_7190) );
oa22f01  g4274 ( .o(n11005), .a(n7745), .b(n11003), .c(n7744), .d(n11004) );
no02f01  g4275 ( .o(n11006), .a(n11005), .b(n11002) );
na02f01  g4276 ( .o(n7340), .a(n11006), .b(n10999) );
ao22f01  g4277 ( .o(n11008), .a(n6736_1), .b(net_7636), .c(n6734), .d(net_7604) );
ao22f01  g4278 ( .o(n11009), .a(n6739), .b(net_7668), .c(n6738), .d(_net_7572) );
na02f01  g4279 ( .o(n7354), .a(n11009), .b(n11008) );
ao22f01  g4280 ( .o(n11011), .a(n6877), .b(_net_7279), .c(n6876_1), .d(net_7343) );
ao22f01  g4281 ( .o(n11012), .a(n6881_1), .b(net_7311), .c(n6880), .d(net_7375) );
na02f01  g4282 ( .o(n7363), .a(n11012), .b(n11011) );
in01f01  g4283 ( .o(n11014), .a(_net_7666) );
na02f01  g4284 ( .o(n11015), .a(n7892), .b(n7446_1) );
oa12f01  g4285 ( .o(n7381), .a(n11015), .b(n7446_1), .c(n11014) );
na02f01  g4286 ( .o(n11017), .a(n7119), .b(_net_6105) );
na02f01  g4287 ( .o(n11018), .a(n8187), .b(n7124) );
na02f01  g4288 ( .o(n7386), .a(n11018), .b(n11017) );
in01f01  g4289 ( .o(n11020), .a(_net_117) );
na02f01  g4290 ( .o(n11021), .a(net_313), .b(_net_154) );
oa12f01  g4291 ( .o(n7395), .a(n11021), .b(n11020), .c(_net_154) );
in01f01  g4292 ( .o(n11023), .a(_net_7473) );
na02f01  g4293 ( .o(n11024), .a(n7200), .b(n6869) );
oa12f01  g4294 ( .o(n7400), .a(n11024), .b(n6869), .c(n11023) );
no02f01  g4295 ( .o(n11026), .a(n6821), .b(n6819) );
na03f01  g4296 ( .o(n11027), .a(n6823), .b(n8344), .c(_net_6957) );
na02f01  g4297 ( .o(n11028), .a(n6823), .b(n8344) );
na02f01  g4298 ( .o(n11029), .a(n11028), .b(n6818_1) );
na03f01  g4299 ( .o(n11030), .a(n11029), .b(n11027), .c(n11026) );
na02f01  g4300 ( .o(n11031), .a(n8345_1), .b(_net_6957) );
na02f01  g4301 ( .o(n7422), .a(n11031), .b(n11030) );
no02f01  g4302 ( .o(n7432), .a(n7232), .b(n7158) );
na02f01  g4303 ( .o(n11034), .a(n10463), .b(n8028_1) );
ao22f01  g4304 ( .o(n11035), .a(n8031), .b(n8033_1), .c(n8034), .d(_net_6069) );
na02f01  g4305 ( .o(n11036), .a(n8037), .b(n8110) );
oa12f01  g4306 ( .o(n11037), .a(n8113), .b(n9046), .c(n9043) );
na04f01  g4307 ( .o(n7437), .a(n11037), .b(n11036), .c(n11035), .d(n11034) );
in01f01  g4308 ( .o(n11039), .a(_net_6007) );
na02f01  g4309 ( .o(n11040), .a(n7348), .b(_net_7810) );
oa12f01  g4310 ( .o(n7454), .a(n11040), .b(n7348), .c(n11039) );
in01f01  g4311 ( .o(n11042), .a(_net_7263) );
na02f01  g4312 ( .o(n11043), .a(n7994_1), .b(n6901) );
oa12f01  g4313 ( .o(n7459), .a(n11043), .b(n6901), .c(n11042) );
in01f01  g4314 ( .o(n11045), .a(_net_6221) );
no02f01  g4315 ( .o(n7473), .a(_net_392), .b(n11045) );
in01f01  g4316 ( .o(n11047), .a(_net_7351) );
na02f01  g4317 ( .o(n11048), .a(n8022), .b(n7030) );
oa12f01  g4318 ( .o(n7478), .a(n11048), .b(n7030), .c(n11047) );
no02f01  g4319 ( .o(n11050), .a(_net_6962), .b(n8252) );
no02f01  g4320 ( .o(n11051), .a(n8253_1), .b(net_6961) );
no02f01  g4321 ( .o(n11052), .a(n11051), .b(n11050) );
oa22f01  g4322 ( .o(n7487), .a(n11052), .b(n8250), .c(n8256), .d(n8253_1) );
na02f01  g4323 ( .o(n11054), .a(n8108), .b(n8028_1) );
ao22f01  g4324 ( .o(n11055), .a(n8116_1), .b(n8033_1), .c(n8034), .d(_net_6068) );
na02f01  g4325 ( .o(n11056), .a(n9810), .b(n8110) );
oa12f01  g4326 ( .o(n11057), .a(n8113), .b(n6772), .c(n6769) );
na04f01  g4327 ( .o(n7496), .a(n11057), .b(n11056), .c(n11055), .d(n11054) );
no04f01  g4328 ( .o(n7501), .a(n7340_1), .b(n7782), .c(n7294), .d(n7281) );
in01f01  g4329 ( .o(n11060), .a(_net_7471) );
na02f01  g4330 ( .o(n11061), .a(n7387), .b(n6869) );
oa12f01  g4331 ( .o(n7518), .a(n11061), .b(n6869), .c(n11060) );
ao22f01  g4332 ( .o(n11063), .a(n7288_1), .b(_net_6045), .c(n7286), .d(_net_284) );
ao22f01  g4333 ( .o(n11064), .a(n7298), .b(_net_7734), .c(n7291), .d(_net_7705) );
na02f01  g4334 ( .o(n11065), .a(n7302_1), .b(_net_128) );
na03f01  g4335 ( .o(n11066), .a(n7308), .b(net_207), .c(x1322) );
na02f01  g4336 ( .o(n11067), .a(n7296), .b(net_244) );
na03f01  g4337 ( .o(n11068), .a(n7308), .b(net_170), .c(n6800) );
na03f01  g4338 ( .o(n11069), .a(n11068), .b(n11067), .c(n11066) );
ao12f01  g4339 ( .o(n11070), .a(n11069), .b(n7306), .c(_net_6001) );
na04f01  g4340 ( .o(n7539), .a(n11070), .b(n11065), .c(n11064), .d(n11063) );
ao22f01  g4341 ( .o(n11072), .a(n6877), .b(_net_7271), .c(n6876_1), .d(net_7335) );
ao22f01  g4342 ( .o(n11073), .a(n6881_1), .b(net_7303), .c(n6880), .d(net_7367) );
na02f01  g4343 ( .o(n7543), .a(n11073), .b(n11072) );
ao22f01  g4344 ( .o(n11075), .a(n6736_1), .b(_net_7629), .c(n6734), .d(_net_7597) );
ao22f01  g4345 ( .o(n11076), .a(n6739), .b(_net_7661), .c(n6738), .d(_net_7565) );
na02f01  g4346 ( .o(n7548), .a(n11076), .b(n11075) );
in01f01  g4347 ( .o(n11078), .a(n9860) );
na02f01  g4348 ( .o(n11079), .a(n6899_1), .b(n9854) );
na02f01  g4349 ( .o(n11080), .a(n6898), .b(_net_7381) );
na02f01  g4350 ( .o(n11081), .a(n11080), .b(n11079) );
oa22f01  g4351 ( .o(n7558), .a(n11081), .b(n9857), .c(n11078), .d(n9854) );
in01f01  g4352 ( .o(n11083), .a(_net_7293) );
na02f01  g4353 ( .o(n11084), .a(n8809_1), .b(n7180) );
oa12f01  g4354 ( .o(n7563), .a(n11084), .b(n7180), .c(n11083) );
na02f01  g4355 ( .o(n11086), .a(n10708), .b(n8213) );
ao22f01  g4356 ( .o(n11087), .a(n8216_1), .b(n9200), .c(n8211_1), .d(_net_6127) );
na02f01  g4357 ( .o(n7572), .a(n11087), .b(n11086) );
in01f01  g4358 ( .o(n11089), .a(_net_7798) );
na02f01  g4359 ( .o(n11090), .a(n6803), .b(_net_6033) );
oa12f01  g4360 ( .o(n7586), .a(n11090), .b(n6803), .c(n11089) );
in01f01  g4361 ( .o(n11092), .a(_net_127) );
na02f01  g4362 ( .o(n11093), .a(_net_154), .b(net_323) );
oa12f01  g4363 ( .o(n7591), .a(n11093), .b(n11092), .c(_net_154) );
na03f01  g4364 ( .o(n11095), .a(n9707), .b(n9706), .c(_net_6022) );
na02f01  g4365 ( .o(n11096), .a(n7293), .b(net_222) );
ao22f01  g4366 ( .o(n11097), .a(n7297_1), .b(net_185), .c(n7296), .d(net_259) );
na03f01  g4367 ( .o(n7596), .a(n11097), .b(n11096), .c(n11095) );
na02f01  g4368 ( .o(n11099), .a(n8544_1), .b(n8338) );
na02f01  g4369 ( .o(n11100), .a(n6815), .b(n6807) );
ao22f01  g4370 ( .o(n11101), .a(n11100), .b(n8340_1), .c(n8345_1), .d(_net_6959) );
na02f01  g4371 ( .o(n7608), .a(n11101), .b(n11099) );
ao22f01  g4372 ( .o(n11103), .a(n7225), .b(_net_7407), .c(n7224), .d(_net_7439) );
ao22f01  g4373 ( .o(n11104), .a(n7229), .b(_net_7503), .c(n7228), .d(_net_7471) );
na02f01  g4374 ( .o(n7613), .a(n11104), .b(n11103) );
in01f01  g4375 ( .o(n11106), .a(_net_6206) );
no02f01  g4376 ( .o(n7622), .a(_net_392), .b(n11106) );
in01f01  g4377 ( .o(n11108), .a(_net_7331) );
na02f01  g4378 ( .o(n11109), .a(n7567_1), .b(n7150) );
oa12f01  g4379 ( .o(n7631), .a(n11109), .b(n7150), .c(n11108) );
na02f01  g4380 ( .o(n11111), .a(n7348), .b(_net_7805) );
oa12f01  g4381 ( .o(n7640), .a(n11111), .b(n7348), .c(n10621) );
in01f01  g4382 ( .o(n11113), .a(_net_6298) );
no02f01  g4383 ( .o(n7649), .a(n11113), .b(_net_392) );
na02f01  g4384 ( .o(n11115), .a(n8310), .b(n7576) );
ao22f01  g4385 ( .o(n11116), .a(n9111), .b(n8307_1), .c(n8312), .d(_net_7228) );
na02f01  g4386 ( .o(n7666), .a(n11116), .b(n11115) );
oa12f01  g4387 ( .o(n11118), .a(n6917), .b(n7804), .c(n7801) );
ao22f01  g4388 ( .o(n11119), .a(n6923), .b(net_6564), .c(n6920), .d(net_6628) );
ao22f01  g4389 ( .o(n11120), .a(n6928), .b(net_6596), .c(n6926), .d(net_6660) );
na02f01  g4390 ( .o(n11121), .a(n11120), .b(n11119) );
ao22f01  g4391 ( .o(n11122), .a(n11121), .b(n6935), .c(n6933), .d(_net_6091) );
in01f01  g4392 ( .o(n11123), .a(net_6578) );
in01f01  g4393 ( .o(n11124), .a(net_6642) );
oa22f01  g4394 ( .o(n11125), .a(n6922), .b(n11123), .c(n6919_1), .d(n11124) );
in01f01  g4395 ( .o(n11126), .a(net_6674) );
in01f01  g4396 ( .o(n11127), .a(net_6610) );
oa22f01  g4397 ( .o(n11128), .a(n6927), .b(n11127), .c(n6925), .d(n11126) );
no02f01  g4398 ( .o(n11129), .a(n11128), .b(n11125) );
no03f01  g4399 ( .o(n11130), .a(n11129), .b(n6947_1), .c(n6943_1) );
ao12f01  g4400 ( .o(n11131), .a(n11130), .b(n8005_1), .c(n6946) );
na03f01  g4401 ( .o(n7671), .a(n11131), .b(n11122), .c(n11118) );
no02f01  g4402 ( .o(n11133), .a(n10494), .b(n6945) );
no02f01  g4403 ( .o(n11134), .a(n10592), .b(n6934_1) );
in01f01  g4404 ( .o(n11135), .a(_net_6103) );
oa22f01  g4405 ( .o(n11136), .a(n11129), .b(n6916), .c(n6932), .d(n11135) );
no03f01  g4406 ( .o(n11137), .a(n11136), .b(n11134), .c(n11133) );
in01f01  g4407 ( .o(n11138), .a(net_6590) );
in01f01  g4408 ( .o(n11139), .a(net_6622) );
oa22f01  g4409 ( .o(n11140), .a(n7058_1), .b(n11138), .c(n7057), .d(n11139) );
in01f01  g4410 ( .o(n11141), .a(net_6654) );
in01f01  g4411 ( .o(n11142), .a(net_6686) );
oa22f01  g4412 ( .o(n11143), .a(n7063), .b(n11142), .c(n7062_1), .d(n11141) );
no02f01  g4413 ( .o(n11144), .a(n11143), .b(n11140) );
na02f01  g4414 ( .o(n7676), .a(n11144), .b(n11137) );
in01f01  g4415 ( .o(n11146), .a(_net_125) );
na02f01  g4416 ( .o(n11147), .a(net_321), .b(_net_154) );
oa12f01  g4417 ( .o(n7681), .a(n11147), .b(n11146), .c(_net_154) );
ao22f01  g4418 ( .o(n11149), .a(n6738), .b(_net_7553), .c(n6736_1), .d(_net_7617) );
ao22f01  g4419 ( .o(n11150), .a(n6739), .b(_net_7649), .c(n6734), .d(_net_7585) );
na02f01  g4420 ( .o(n7686), .a(n11150), .b(n11149) );
na02f01  g4421 ( .o(n11152), .a(n7348), .b(_net_7801) );
oa12f01  g4422 ( .o(n7695), .a(n11152), .b(n7348), .c(n6912) );
no03f01  g4423 ( .o(n11154), .a(_net_6043), .b(n7570), .c(n8699) );
no02f01  g4424 ( .o(n11155), .a(n7570), .b(n8695) );
ao22f01  g4425 ( .o(n11156), .a(n11155), .b(n8705), .c(n11154), .d(n8703_1) );
ao12f01  g4426 ( .o(n11157), .a(n7570), .b(_net_5982), .c(n8695) );
no03f01  g4427 ( .o(n11158), .a(_net_6043), .b(n7570), .c(_net_6044) );
ao22f01  g4428 ( .o(n11159), .a(n11158), .b(n8701), .c(n11157), .d(n8694_1) );
na02f01  g4429 ( .o(n7709), .a(n11159), .b(n11156) );
in01f01  g4430 ( .o(n11161), .a(_net_7273) );
na02f01  g4431 ( .o(n11162), .a(n518), .b(n6901) );
oa12f01  g4432 ( .o(n7723), .a(n11162), .b(n6901), .c(n11161) );
in01f01  g4433 ( .o(n11164), .a(_net_7289) );
na02f01  g4434 ( .o(n11165), .a(n9587), .b(n7180) );
oa12f01  g4435 ( .o(n7728), .a(n11165), .b(n7180), .c(n11164) );
ao22f01  g4436 ( .o(n11167), .a(n7288_1), .b(_net_6043), .c(n7286), .d(_net_282) );
ao22f01  g4437 ( .o(n11168), .a(n7298), .b(_net_7732), .c(n7291), .d(_net_7703) );
na02f01  g4438 ( .o(n11169), .a(n7302_1), .b(_net_126) );
na03f01  g4439 ( .o(n11170), .a(n7308), .b(net_205), .c(x1322) );
na02f01  g4440 ( .o(n11171), .a(n7296), .b(net_242) );
na03f01  g4441 ( .o(n11172), .a(n7308), .b(net_168), .c(n6800) );
na03f01  g4442 ( .o(n11173), .a(n11172), .b(n11171), .c(n11170) );
ao12f01  g4443 ( .o(n11174), .a(n11173), .b(n7306), .c(_net_5999) );
na04f01  g4444 ( .o(n7737), .a(n11174), .b(n11169), .c(n11168), .d(n11167) );
no02f01  g4445 ( .o(n7741), .a(n10333), .b(n10331) );
ao12f01  g4446 ( .o(n11177), .a(n9607), .b(net_6826), .c(_net_6827) );
no03f01  g4447 ( .o(n11178), .a(_net_6828), .b(n8220_1), .c(n8219) );
no02f01  g4448 ( .o(n11179), .a(n11178), .b(n11177) );
oa22f01  g4449 ( .o(n7746), .a(n11179), .b(n8226), .c(n8227), .d(n9607) );
in01f01  g4450 ( .o(n11181), .a(_net_7555) );
na02f01  g4451 ( .o(n11182), .a(n9154), .b(n7519) );
oa12f01  g4452 ( .o(n7751), .a(n11182), .b(n7519), .c(n11181) );
in01f01  g4453 ( .o(n11184), .a(_net_7699) );
na02f01  g4454 ( .o(n11185), .a(n7207_1), .b(_net_7801) );
oa12f01  g4455 ( .o(n7768), .a(n11185), .b(n7207_1), .c(n11184) );
na02f01  g4456 ( .o(n11187), .a(n7298), .b(_net_7736) );
ao22f01  g4457 ( .o(n11188), .a(n7306), .b(_net_6006), .c(n7291), .d(_net_7707) );
na02f01  g4458 ( .o(n11189), .a(n7302_1), .b(net_146) );
na02f01  g4459 ( .o(n11190), .a(n7296), .b(net_246) );
na03f01  g4460 ( .o(n11191), .a(n7308), .b(_net_172), .c(n6800) );
na03f01  g4461 ( .o(n11192), .a(n7308), .b(_net_209), .c(x1322) );
na03f01  g4462 ( .o(n11193), .a(n11192), .b(n11191), .c(n11190) );
ao12f01  g4463 ( .o(n11194), .a(n11193), .b(n7286), .c(_net_289) );
na04f01  g4464 ( .o(n7773), .a(n11194), .b(n11189), .c(n11188), .d(n11187) );
ao12f01  g4465 ( .o(n11196), .a(n6945), .b(n11120), .c(n11119) );
no02f01  g4466 ( .o(n11197), .a(n7805), .b(n6934_1) );
in01f01  g4467 ( .o(n11198), .a(_net_6093) );
oa22f01  g4468 ( .o(n11199), .a(n7813), .b(n6916), .c(n6932), .d(n11198) );
no03f01  g4469 ( .o(n11200), .a(n11199), .b(n11197), .c(n11196) );
in01f01  g4470 ( .o(n11201), .a(net_6612) );
in01f01  g4471 ( .o(n11202), .a(net_6580) );
oa22f01  g4472 ( .o(n11203), .a(n7058_1), .b(n11202), .c(n7057), .d(n11201) );
in01f01  g4473 ( .o(n11204), .a(net_6676) );
in01f01  g4474 ( .o(n11205), .a(net_6644) );
oa22f01  g4475 ( .o(n11206), .a(n7063), .b(n11204), .c(n7062_1), .d(n11205) );
no02f01  g4476 ( .o(n11207), .a(n11206), .b(n11203) );
na02f01  g4477 ( .o(n7788), .a(n11207), .b(n11200) );
in01f01  g4478 ( .o(n11209), .a(_net_6049) );
ao12f01  g4479 ( .o(n11210), .a(n9253), .b(_net_7230), .c(_net_7233) );
oa12f01  g4480 ( .o(n11211), .a(n11210), .b(_net_7230), .c(_net_7233) );
na02f01  g4481 ( .o(n11212), .a(n10338), .b(n4276) );
oa12f01  g4482 ( .o(n7793), .a(n11209), .b(n11212), .c(n11211) );
in01f01  g4483 ( .o(n11214), .a(_net_7442) );
na02f01  g4484 ( .o(n11215), .a(n7197), .b(n6891) );
oa12f01  g4485 ( .o(n7798), .a(n11215), .b(n7197), .c(n11214) );
no02f01  g4486 ( .o(n11217), .a(n6809_1), .b(_net_6962) );
no02f01  g4487 ( .o(n11218), .a(_net_6959), .b(n8253_1) );
no02f01  g4488 ( .o(n11219), .a(n11218), .b(n11217) );
no02f01  g4489 ( .o(n11220), .a(n6806_1), .b(net_6961) );
no02f01  g4490 ( .o(n11221), .a(n11220), .b(n11219) );
no04f01  g4491 ( .o(n11222), .a(n11218), .b(n11217), .c(n6806_1), .d(net_6961) );
no02f01  g4492 ( .o(n11223), .a(n6806_1), .b(n8252) );
no02f01  g4493 ( .o(n11224), .a(_net_6958), .b(net_6961) );
no02f01  g4494 ( .o(n11225), .a(n11224), .b(n11223) );
oa12f01  g4495 ( .o(n11226), .a(n11225), .b(n11222), .c(n11221) );
no02f01  g4496 ( .o(n11227), .a(n11222), .b(n11221) );
in01f01  g4497 ( .o(n9778), .a(n11225) );
na02f01  g4498 ( .o(n11229), .a(n9778), .b(n11227) );
na02f01  g4499 ( .o(n7822), .a(n11229), .b(n11226) );
in01f01  g4500 ( .o(n11231), .a(_net_7276) );
na02f01  g4501 ( .o(n11232), .a(n1639), .b(n6901) );
oa12f01  g4502 ( .o(n7835), .a(n11232), .b(n6901), .c(n11231) );
na02f01  g4503 ( .o(n11234), .a(n7291), .b(net_7715) );
na02f01  g4504 ( .o(n11235), .a(n7293), .b(_net_217) );
ao22f01  g4505 ( .o(n11236), .a(n7297_1), .b(_net_180), .c(n7296), .d(net_254) );
ao22f01  g4506 ( .o(n11237), .a(n7306), .b(_net_6017), .c(n7298), .d(net_7744) );
na04f01  g4507 ( .o(n7845), .a(n11237), .b(n11236), .c(n11235), .d(n11234) );
ao22f01  g4508 ( .o(n11239), .a(n7225), .b(_net_7408), .c(n7224), .d(_net_7440) );
ao22f01  g4509 ( .o(n11240), .a(n7229), .b(_net_7504), .c(n7228), .d(_net_7472) );
na02f01  g4510 ( .o(n7853), .a(n11240), .b(n11239) );
no02f01  g4511 ( .o(n7858), .a(n8317), .b(n9892) );
na03f01  g4512 ( .o(n11243), .a(n9260), .b(_net_6407), .c(_net_6408) );
ao12f01  g4513 ( .o(n11244), .a(x38), .b(n11243), .c(_net_6409) );
oa12f01  g4514 ( .o(n7863), .a(n11244), .b(n11243), .c(_net_6409) );
in01f01  g4515 ( .o(n11246), .a(_net_7484) );
na02f01  g4516 ( .o(n11247), .a(n9872), .b(n6869) );
oa12f01  g4517 ( .o(n7888), .a(n11247), .b(n6869), .c(n11246) );
in01f01  g4518 ( .o(n11249), .a(_net_5850) );
in01f01  g4519 ( .o(n11250), .a(x837) );
na03f01  g4520 ( .o(n11251), .a(n10203), .b(net_7780), .c(n11250) );
oa12f01  g4521 ( .o(n7897), .a(n11251), .b(n11249), .c(x837) );
in01f01  g4522 ( .o(n11253), .a(_net_7796) );
na02f01  g4523 ( .o(n11254), .a(n6803), .b(_net_6031) );
oa12f01  g4524 ( .o(n7902), .a(n11254), .b(n6803), .c(n11253) );
na02f01  g4525 ( .o(n11256), .a(n8857), .b(_net_6552) );
na02f01  g4526 ( .o(n11257), .a(n8856), .b(n6758) );
na02f01  g4527 ( .o(n11258), .a(n11257), .b(n11256) );
na02f01  g4528 ( .o(n11259), .a(n8862), .b(_net_6552) );
oa12f01  g4529 ( .o(n7911), .a(n11259), .b(n11258), .c(n8858) );
ao22f01  g4530 ( .o(n11261), .a(n6736_1), .b(_net_7623), .c(n6734), .d(_net_7591) );
ao22f01  g4531 ( .o(n11262), .a(n6739), .b(_net_7655), .c(n6738), .d(_net_7559) );
na02f01  g4532 ( .o(n7933), .a(n11262), .b(n11261) );
in01f01  g4533 ( .o(n11264), .a(net_7760) );
na04f01  g4534 ( .o(n11265), .a(_net_6039), .b(_net_7791), .c(net_303), .d(n11264) );
ao12f01  g4535 ( .o(n7950), .a(n11265), .b(net_304), .c(_net_6040) );
in01f01  g4536 ( .o(n11267), .a(_net_5855) );
in01f01  g4537 ( .o(n11268), .a(x977) );
na03f01  g4538 ( .o(n11269), .a(n9364), .b(net_7775), .c(n11268) );
oa12f01  g4539 ( .o(n7975), .a(n11269), .b(n11267), .c(x977) );
ao22f01  g4540 ( .o(n11271), .a(n6877), .b(_net_7252), .c(n6876_1), .d(_net_7316) );
ao22f01  g4541 ( .o(n11272), .a(n6881_1), .b(_net_7284), .c(n6880), .d(_net_7348) );
na02f01  g4542 ( .o(n7980), .a(n11272), .b(n11271) );
in01f01  g4543 ( .o(n11274), .a(_net_7425) );
na02f01  g4544 ( .o(n11275), .a(n2958), .b(n7550) );
oa12f01  g4545 ( .o(n7985), .a(n11275), .b(n7550), .c(n11274) );
in01f01  g4546 ( .o(n11277), .a(_net_5852) );
in01f01  g4547 ( .o(n11278), .a(x889) );
no02f01  g4548 ( .o(n11279), .a(n10034), .b(_net_272) );
na02f01  g4549 ( .o(n11280), .a(_net_267), .b(_net_273) );
ao12f01  g4550 ( .o(n11281), .a(n11280), .b(_net_192), .c(n9591) );
na02f01  g4551 ( .o(n11282), .a(n11281), .b(n11279) );
in01f01  g4552 ( .o(n11283), .a(n11280) );
no02f01  g4553 ( .o(n11284), .a(n10034), .b(n9019) );
na03f01  g4554 ( .o(n11285), .a(n11284), .b(n11283), .c(_net_189) );
na03f01  g4555 ( .o(n11286), .a(_net_192), .b(n9591), .c(_net_191) );
na04f01  g4556 ( .o(n11287), .a(n11286), .b(n11283), .c(n10034), .d(n9019) );
oa12f01  g4557 ( .o(n11288), .a(n9591), .b(_net_192), .c(_net_191) );
na04f01  g4558 ( .o(n11289), .a(n11288), .b(n11283), .c(n10034), .d(_net_272) );
na04f01  g4559 ( .o(n11290), .a(n11289), .b(n11287), .c(n11285), .d(n11282) );
na03f01  g4560 ( .o(n11291), .a(n11290), .b(net_7778), .c(n11278) );
oa12f01  g4561 ( .o(n8010), .a(n11291), .b(n11277), .c(x889) );
in01f01  g4562 ( .o(n11293), .a(_net_291) );
na02f01  g4563 ( .o(n11294), .a(n7440), .b(_net_7811) );
oa12f01  g4564 ( .o(n8019), .a(n11294), .b(n7440), .c(n11293) );
in01f01  g4565 ( .o(n11296), .a(_net_6286) );
no02f01  g4566 ( .o(n8024), .a(_net_392), .b(n11296) );
ao12f01  g4567 ( .o(n11298), .a(n6764), .b(n8107_1), .c(n8106) );
no02f01  g4568 ( .o(n11299), .a(n10546), .b(n6766) );
in01f01  g4569 ( .o(n11300), .a(_net_6072) );
oa22f01  g4570 ( .o(n11301), .a(n10554), .b(n6775), .c(n6784), .d(n11300) );
no03f01  g4571 ( .o(n11302), .a(n11301), .b(n11299), .c(n11298) );
in01f01  g4572 ( .o(n11303), .a(net_6476) );
in01f01  g4573 ( .o(n11304), .a(net_6444) );
oa22f01  g4574 ( .o(n11305), .a(n6790), .b(n11304), .c(n6789), .d(n11303) );
in01f01  g4575 ( .o(n11306), .a(net_6540) );
in01f01  g4576 ( .o(n11307), .a(net_6508) );
oa22f01  g4577 ( .o(n11308), .a(n6795), .b(n11306), .c(n6794), .d(n11307) );
no02f01  g4578 ( .o(n11309), .a(n11308), .b(n11305) );
na02f01  g4579 ( .o(n8033), .a(n11309), .b(n11302) );
in01f01  g4580 ( .o(n11311), .a(_net_7262) );
na02f01  g4581 ( .o(n11312), .a(n7926), .b(n6901) );
oa12f01  g4582 ( .o(n8080), .a(n11312), .b(n6901), .c(n11311) );
in01f01  g4583 ( .o(n11314), .a(_net_7573) );
na02f01  g4584 ( .o(n11315), .a(n7519), .b(n718) );
oa12f01  g4585 ( .o(n8097), .a(n11315), .b(n7519), .c(n11314) );
in01f01  g4586 ( .o(n11317), .a(_net_7499) );
na02f01  g4587 ( .o(n11318), .a(n9700_1), .b(n7626_1) );
oa12f01  g4588 ( .o(n8102), .a(n11318), .b(n7626_1), .c(n11317) );
in01f01  g4589 ( .o(n11320), .a(_net_7417) );
na02f01  g4590 ( .o(n11321), .a(n7550), .b(n6872_1) );
oa12f01  g4591 ( .o(n8107), .a(n11321), .b(n7550), .c(n11320) );
no02f01  g4592 ( .o(n11323), .a(n10745), .b(n7468_1) );
no02f01  g4593 ( .o(n11324), .a(n10754), .b(n7470) );
in01f01  g4594 ( .o(n11325), .a(_net_6115) );
oa22f01  g4595 ( .o(n11326), .a(n10660), .b(n7123), .c(n7118), .d(n11325) );
no03f01  g4596 ( .o(n11327), .a(n11326), .b(n11324), .c(n11323) );
in01f01  g4597 ( .o(n11328), .a(net_6717) );
in01f01  g4598 ( .o(n11329), .a(net_6749) );
oa22f01  g4599 ( .o(n11330), .a(n7492_1), .b(n11328), .c(n7491), .d(n11329) );
in01f01  g4600 ( .o(n11331), .a(net_6813) );
in01f01  g4601 ( .o(n11332), .a(net_6781) );
oa22f01  g4602 ( .o(n11333), .a(n7497), .b(n11331), .c(n7496_1), .d(n11332) );
no02f01  g4603 ( .o(n11334), .a(n11333), .b(n11330) );
na02f01  g4604 ( .o(n8112), .a(n11334), .b(n11327) );
in01f01  g4605 ( .o(n11336), .a(_net_7562) );
na02f01  g4606 ( .o(n11337), .a(n7707), .b(n7519) );
oa12f01  g4607 ( .o(n8121), .a(n11337), .b(n7519), .c(n11336) );
in01f01  g4608 ( .o(n11339), .a(_net_7291) );
na02f01  g4609 ( .o(n11340), .a(n7180), .b(n7033) );
oa12f01  g4610 ( .o(n8130), .a(n11340), .b(n7180), .c(n11339) );
in01f01  g4611 ( .o(n11342), .a(_net_7592) );
na02f01  g4612 ( .o(n11343), .a(n9881), .b(n6968) );
oa12f01  g4613 ( .o(n8135), .a(n11343), .b(n6968), .c(n11342) );
no04f01  g4614 ( .o(n8152), .a(n8362_1), .b(n8352), .c(n6966), .d(_net_7683) );
ao22f01  g4615 ( .o(n11346), .a(n6736_1), .b(_net_7628), .c(n6734), .d(_net_7596) );
ao22f01  g4616 ( .o(n11347), .a(n6739), .b(_net_7660), .c(n6738), .d(_net_7564) );
na02f01  g4617 ( .o(n8161), .a(n11347), .b(n11346) );
ao22f01  g4618 ( .o(n11349), .a(n7225), .b(_net_7429), .c(n7224), .d(net_7461) );
ao22f01  g4619 ( .o(n11350), .a(n7229), .b(net_7525), .c(n7228), .d(net_7493) );
na02f01  g4620 ( .o(n8170), .a(n11350), .b(n11349) );
ao22f01  g4621 ( .o(n11352), .a(n6877), .b(_net_7274), .c(n6876_1), .d(net_7338) );
ao22f01  g4622 ( .o(n11353), .a(n6881_1), .b(net_7306), .c(n6880), .d(net_7370) );
na02f01  g4623 ( .o(n8179), .a(n11353), .b(n11352) );
in01f01  g4624 ( .o(n11355), .a(_net_7275) );
na02f01  g4625 ( .o(n11356), .a(n2084), .b(n6901) );
oa12f01  g4626 ( .o(n8192), .a(n11356), .b(n6901), .c(n11355) );
no03f01  g4627 ( .o(n11358), .a(n8094), .b(_net_271), .c(n9019) );
no02f01  g4628 ( .o(n11359), .a(n8094), .b(n9591) );
ao22f01  g4629 ( .o(n11360), .a(n11359), .b(n11284), .c(n11358), .d(n11288) );
ao12f01  g4630 ( .o(n11361), .a(n8094), .b(_net_192), .c(n9591) );
no03f01  g4631 ( .o(n11362), .a(n8094), .b(_net_271), .c(_net_272) );
ao22f01  g4632 ( .o(n11363), .a(n11362), .b(n11286), .c(n11361), .d(n11279) );
na02f01  g4633 ( .o(n8197), .a(n11363), .b(n11360) );
no02f01  g4634 ( .o(n11365), .a(n8069), .b(n7012) );
no02f01  g4635 ( .o(n11366), .a(n9934), .b(n6997) );
in01f01  g4636 ( .o(n11367), .a(_net_6159) );
oa22f01  g4637 ( .o(n11368), .a(n8471), .b(n6980), .c(n6995_1), .d(n11367) );
no03f01  g4638 ( .o(n11369), .a(n11368), .b(n11366), .c(n11365) );
in01f01  g4639 ( .o(n11370), .a(net_6991) );
in01f01  g4640 ( .o(n11371), .a(net_7023) );
oa22f01  g4641 ( .o(n11372), .a(n8075_1), .b(n11370), .c(n8074), .d(n11371) );
in01f01  g4642 ( .o(n11373), .a(net_7055) );
in01f01  g4643 ( .o(n11374), .a(net_7087) );
oa22f01  g4644 ( .o(n11375), .a(n8080_1), .b(n11374), .c(n8079), .d(n11373) );
no02f01  g4645 ( .o(n11376), .a(n11375), .b(n11372) );
na02f01  g4646 ( .o(n8202), .a(n11376), .b(n11369) );
na02f01  g4647 ( .o(n11378), .a(_net_5990), .b(_net_5984) );
ao12f01  g4648 ( .o(n11379), .a(n11378), .b(_net_5962), .c(n7533) );
na02f01  g4649 ( .o(n11380), .a(n11379), .b(n7541) );
in01f01  g4650 ( .o(n11381), .a(n11378) );
na04f01  g4651 ( .o(n11382), .a(n11381), .b(n7543_1), .c(n7535_1), .d(n7538) );
na04f01  g4652 ( .o(n11383), .a(n11381), .b(n7534), .c(_net_5989), .d(n7538) );
na03f01  g4653 ( .o(n11384), .a(n11381), .b(n7539_1), .c(_net_5960) );
na04f01  g4654 ( .o(n11385), .a(n11384), .b(n11383), .c(n11382), .d(n11380) );
in01f01  g4655 ( .o(n11386), .a(n11385) );
no02f01  g4656 ( .o(n8211), .a(n11386), .b(x1062) );
in01f01  g4657 ( .o(n11388), .a(_net_7702) );
na02f01  g4658 ( .o(n11389), .a(n7207_1), .b(_net_7804) );
oa12f01  g4659 ( .o(n8216), .a(n11389), .b(n7207_1), .c(n11388) );
no02f01  g4660 ( .o(n8224), .a(n7161), .b(n7232) );
in01f01  g4661 ( .o(n11392), .a(_net_7580) );
na02f01  g4662 ( .o(n11393), .a(n5814), .b(n7519) );
oa12f01  g4663 ( .o(n8237), .a(n11393), .b(n7519), .c(n11392) );
in01f01  g4664 ( .o(n11395), .a(_net_7432) );
na02f01  g4665 ( .o(n11396), .a(n5552), .b(n7550) );
oa12f01  g4666 ( .o(n8253), .a(n11396), .b(n7550), .c(n11395) );
ao22f01  g4667 ( .o(n11398), .a(n7225), .b(_net_7404), .c(n7224), .d(_net_7436) );
ao22f01  g4668 ( .o(n11399), .a(n7229), .b(_net_7500), .c(n7228), .d(_net_7468) );
na02f01  g4669 ( .o(n8258), .a(n11399), .b(n11398) );
na02f01  g4670 ( .o(n11401), .a(n10016), .b(n10015) );
na02f01  g4671 ( .o(n11402), .a(n11401), .b(n10020) );
oa22f01  g4672 ( .o(n8284), .a(n11402), .b(n10014_1), .c(n10013), .d(n10016) );
in01f01  g4673 ( .o(n11404), .a(_net_7648) );
na02f01  g4674 ( .o(n11405), .a(n8842), .b(n7446_1) );
oa12f01  g4675 ( .o(n8294), .a(n11405), .b(n7446_1), .c(n11404) );
in01f01  g4676 ( .o(n11407), .a(_net_6020) );
na02f01  g4677 ( .o(n11408), .a(n7348), .b(_net_7820) );
oa12f01  g4678 ( .o(n8299), .a(n11408), .b(n7348), .c(n11407) );
in01f01  g4679 ( .o(n11410), .a(_net_6200) );
no02f01  g4680 ( .o(n8324), .a(_net_392), .b(n11410) );
no02f01  g4681 ( .o(n11412), .a(n8673), .b(n7468_1) );
no02f01  g4682 ( .o(n11413), .a(n8682), .b(n7470) );
ao22f01  g4683 ( .o(n11414), .a(n7130), .b(net_6713), .c(n7127), .d(net_6777) );
ao22f01  g4684 ( .o(n11415), .a(n7135), .b(net_6745), .c(n7133_1), .d(net_6809) );
ao12f01  g4685 ( .o(n11416), .a(n7123), .b(n11415), .c(n11414) );
in01f01  g4686 ( .o(n11417), .a(_net_6123) );
no02f01  g4687 ( .o(n11418), .a(n7118), .b(n11417) );
no04f01  g4688 ( .o(n11419), .a(n11418), .b(n11416), .c(n11413), .d(n11412) );
in01f01  g4689 ( .o(n11420), .a(net_6725) );
in01f01  g4690 ( .o(n11421), .a(net_6757) );
oa22f01  g4691 ( .o(n11422), .a(n7492_1), .b(n11420), .c(n7491), .d(n11421) );
in01f01  g4692 ( .o(n11423), .a(net_6821) );
in01f01  g4693 ( .o(n11424), .a(net_6789) );
oa22f01  g4694 ( .o(n11425), .a(n7497), .b(n11423), .c(n7496_1), .d(n11424) );
no02f01  g4695 ( .o(n11426), .a(n11425), .b(n11422) );
na02f01  g4696 ( .o(n8345), .a(n11426), .b(n11419) );
na02f01  g4697 ( .o(n11428), .a(n10291), .b(n7125_1) );
ao22f01  g4698 ( .o(n11429), .a(n10289), .b(n9611_1), .c(n8716), .d(_net_6823) );
na02f01  g4699 ( .o(n8354), .a(n11429), .b(n11428) );
in01f01  g4700 ( .o(n11431), .a(n9444) );
no02f01  g4701 ( .o(n8367), .a(n11431), .b(n9439) );
oa12f01  g4702 ( .o(n11433), .a(n7397), .b(n6959), .c(n8231) );
na03f01  g4703 ( .o(n11434), .a(n11433), .b(n10048), .c(n10047_1) );
na02f01  g4704 ( .o(n11435), .a(n7399), .b(n6961) );
ao22f01  g4705 ( .o(n11436), .a(n11435), .b(n10043), .c(n8237_1), .d(_net_7685) );
na02f01  g4706 ( .o(n8372), .a(n11436), .b(n11434) );
in01f01  g4707 ( .o(n11438), .a(_net_7735) );
ao12f01  g4708 ( .o(n8377), .a(n7343), .b(n11438), .c(n7315) );
in01f01  g4709 ( .o(n11440), .a(_net_7602) );
na02f01  g4710 ( .o(n11441), .a(n7892), .b(n6968) );
oa12f01  g4711 ( .o(n8382), .a(n11441), .b(n6968), .c(n11440) );
ao12f01  g4712 ( .o(n11443), .a(n7682), .b(_net_6960), .c(_net_6963) );
oa12f01  g4713 ( .o(n11444), .a(n11443), .b(_net_6960), .c(_net_6963) );
na02f01  g4714 ( .o(n11445), .a(n9778), .b(n11219) );
oa12f01  g4715 ( .o(n8387), .a(n9526), .b(n11445), .c(n11444) );
in01f01  g4716 ( .o(n11447), .a(_net_7568) );
na02f01  g4717 ( .o(n11448), .a(n7519), .b(n7403) );
oa12f01  g4718 ( .o(n8396), .a(n11448), .b(n7519), .c(n11447) );
na02f01  g4719 ( .o(n11450), .a(n8340_1), .b(n6806_1) );
ao22f01  g4720 ( .o(n11451), .a(n8538), .b(n8338), .c(n8345_1), .d(_net_6958) );
na02f01  g4721 ( .o(n8405), .a(n11451), .b(n11450) );
in01f01  g4722 ( .o(n11453), .a(_net_7333) );
na02f01  g4723 ( .o(n11454), .a(n9685), .b(n7150) );
oa12f01  g4724 ( .o(n8410), .a(n11454), .b(n7150), .c(n11453) );
na02f01  g4725 ( .o(n11456), .a(n11121), .b(n6917) );
ao22f01  g4726 ( .o(n11457), .a(n8005_1), .b(n6935), .c(n6933), .d(_net_6089) );
no03f01  g4727 ( .o(n11458), .a(n10592), .b(n6947_1), .c(n6943_1) );
ao12f01  g4728 ( .o(n11459), .a(n11458), .b(n8009), .c(n6946) );
na03f01  g4729 ( .o(n8426), .a(n11459), .b(n11457), .c(n11456) );
na02f01  g4730 ( .o(n11461), .a(n7298), .b(net_7741) );
ao22f01  g4731 ( .o(n11462), .a(n7306), .b(_net_6011), .c(n7291), .d(net_7712) );
na02f01  g4732 ( .o(n11463), .a(n7302_1), .b(net_151) );
na02f01  g4733 ( .o(n11464), .a(n7296), .b(net_251) );
na03f01  g4734 ( .o(n11465), .a(n7308), .b(_net_177), .c(n6800) );
na03f01  g4735 ( .o(n11466), .a(n7308), .b(_net_214), .c(x1322) );
na03f01  g4736 ( .o(n11467), .a(n11466), .b(n11465), .c(n11464) );
ao12f01  g4737 ( .o(n11468), .a(n11467), .b(n7286), .c(_net_294) );
na04f01  g4738 ( .o(n8435), .a(n11468), .b(n11463), .c(n11462), .d(n11461) );
no03f01  g4739 ( .o(n8443), .a(n7114), .b(_net_7688), .c(x1155) );
in01f01  g4740 ( .o(n11471), .a(_net_7450) );
na02f01  g4741 ( .o(n11472), .a(n9487_1), .b(n7197) );
oa12f01  g4742 ( .o(n8481), .a(n11472), .b(n7197), .c(n11471) );
in01f01  g4743 ( .o(n11474), .a(net_7173) );
in01f01  g4744 ( .o(n11475), .a(net_7109) );
oa22f01  g4745 ( .o(n11476), .a(n7580), .b(n11475), .c(n7577_1), .d(n11474) );
in01f01  g4746 ( .o(n11477), .a(net_7141) );
in01f01  g4747 ( .o(n11478), .a(net_7205) );
oa22f01  g4748 ( .o(n11479), .a(n7585), .b(n11477), .c(n7583), .d(n11478) );
no02f01  g4749 ( .o(n11480), .a(n11479), .b(n11476) );
no02f01  g4750 ( .o(n11481), .a(n11480), .b(n7721) );
no02f01  g4751 ( .o(n11482), .a(n7935), .b(n7592) );
in01f01  g4752 ( .o(n11483), .a(_net_6178) );
oa22f01  g4753 ( .o(n11484), .a(n7718), .b(n7574), .c(n7590), .d(n11483) );
no03f01  g4754 ( .o(n11485), .a(n11484), .b(n11482), .c(n11481) );
in01f01  g4755 ( .o(n11486), .a(net_7157) );
in01f01  g4756 ( .o(n11487), .a(net_7125) );
oa22f01  g4757 ( .o(n11488), .a(n7740), .b(n11487), .c(n7739), .d(n11486) );
in01f01  g4758 ( .o(n11489), .a(net_7189) );
in01f01  g4759 ( .o(n11490), .a(net_7221) );
oa22f01  g4760 ( .o(n11491), .a(n7745), .b(n11490), .c(n7744), .d(n11489) );
no02f01  g4761 ( .o(n11492), .a(n11491), .b(n11488) );
na02f01  g4762 ( .o(n8486), .a(n11492), .b(n11485) );
in01f01  g4763 ( .o(n11494), .a(_net_7801) );
na02f01  g4764 ( .o(n11495), .a(n6803), .b(_net_6039) );
oa12f01  g4765 ( .o(n8499), .a(n11495), .b(n6803), .c(n11494) );
no02f01  g4766 ( .o(n11497), .a(_net_6557), .b(n7762) );
no02f01  g4767 ( .o(n11498), .a(n7765), .b(net_6556) );
no02f01  g4768 ( .o(n11499), .a(n11498), .b(n11497) );
oa22f01  g4769 ( .o(n8508), .a(n11499), .b(n10412), .c(n10416), .d(n7765) );
in01f01  g4770 ( .o(n11501), .a(_net_7575) );
na02f01  g4771 ( .o(n11502), .a(n7519), .b(n793) );
oa12f01  g4772 ( .o(n8517), .a(n11502), .b(n7519), .c(n11501) );
in01f01  g4773 ( .o(n11504), .a(_net_7349) );
na02f01  g4774 ( .o(n11505), .a(n7183), .b(n7030) );
oa12f01  g4775 ( .o(n8526), .a(n11505), .b(n7030), .c(n11504) );
in01f01  g4776 ( .o(n11507), .a(_net_7284) );
na02f01  g4777 ( .o(n11508), .a(n7180), .b(n6904) );
oa12f01  g4778 ( .o(n8531), .a(n11508), .b(n7180), .c(n11507) );
ao22f01  g4779 ( .o(n11510), .a(n6736_1), .b(_net_7625), .c(n6734), .d(_net_7593) );
ao22f01  g4780 ( .o(n11511), .a(n6739), .b(_net_7657), .c(n6738), .d(_net_7561) );
na02f01  g4781 ( .o(n8540), .a(n11511), .b(n11510) );
ao22f01  g4782 ( .o(n11513), .a(n6877), .b(_net_7260), .c(n6876_1), .d(_net_7324) );
ao22f01  g4783 ( .o(n11514), .a(n6881_1), .b(_net_7292), .c(n6880), .d(_net_7356) );
na02f01  g4784 ( .o(n8557), .a(n11514), .b(n11513) );
in01f01  g4785 ( .o(n11516), .a(_net_122) );
na02f01  g4786 ( .o(n11517), .a(net_318), .b(_net_154) );
oa12f01  g4787 ( .o(n8570), .a(n11517), .b(n11516), .c(_net_154) );
in01f01  g4788 ( .o(n11519), .a(_net_6281) );
no02f01  g4789 ( .o(n8583), .a(_net_392), .b(n11519) );
in01f01  g4790 ( .o(n11521), .a(n11290) );
no02f01  g4791 ( .o(n8588), .a(n11521), .b(x889) );
in01f01  g4792 ( .o(n11523), .a(_net_7695) );
na02f01  g4793 ( .o(n11524), .a(n7207_1), .b(_net_7797) );
oa12f01  g4794 ( .o(n8593), .a(n11524), .b(n7207_1), .c(n11523) );
in01f01  g4795 ( .o(n11526), .a(_net_7319) );
na02f01  g4796 ( .o(n11527), .a(n8022), .b(n7150) );
oa12f01  g4797 ( .o(n8602), .a(n11527), .b(n7150), .c(n11526) );
ao22f01  g4798 ( .o(n11529), .a(n6877), .b(_net_7275), .c(n6876_1), .d(net_7339) );
ao22f01  g4799 ( .o(n11530), .a(n6881_1), .b(net_7307), .c(n6880), .d(net_7371) );
na02f01  g4800 ( .o(n8607), .a(n11530), .b(n11529) );
in01f01  g4801 ( .o(n11532), .a(_net_6164) );
no02f01  g4802 ( .o(n8616), .a(n11532), .b(n7168) );
no02f01  g4803 ( .o(n11534), .a(n8087), .b(_net_6410) );
ao12f01  g4804 ( .o(n8625), .a(n8084), .b(n11534), .c(n8179_1) );
no02f01  g4805 ( .o(n11536), .a(n8397), .b(n6824) );
no02f01  g4806 ( .o(n11537), .a(n8406), .b(n6826_1) );
in01f01  g4807 ( .o(n11538), .a(_net_6141) );
no02f01  g4808 ( .o(n11539), .a(n10716), .b(n10713) );
oa22f01  g4809 ( .o(n11540), .a(n11539), .b(n6836_1), .c(n6844), .d(n11538) );
no03f01  g4810 ( .o(n11541), .a(n11540), .b(n11537), .c(n11536) );
in01f01  g4811 ( .o(n11542), .a(net_6890) );
in01f01  g4812 ( .o(n11543), .a(net_6858) );
oa22f01  g4813 ( .o(n11544), .a(n6850_1), .b(n11543), .c(n6849), .d(n11542) );
in01f01  g4814 ( .o(n11545), .a(net_6922) );
in01f01  g4815 ( .o(n11546), .a(net_6954) );
oa22f01  g4816 ( .o(n11547), .a(n6855_1), .b(n11546), .c(n6854), .d(n11545) );
no02f01  g4817 ( .o(n11548), .a(n11547), .b(n11544) );
na02f01  g4818 ( .o(n8645), .a(n11548), .b(n11541) );
ao22f01  g4819 ( .o(n11550), .a(n7225), .b(_net_7406), .c(n7224), .d(_net_7438) );
ao22f01  g4820 ( .o(n11551), .a(n7229), .b(_net_7502), .c(n7228), .d(_net_7470) );
na02f01  g4821 ( .o(n8662), .a(n11551), .b(n11550) );
in01f01  g4822 ( .o(n11553), .a(_net_7267) );
na02f01  g4823 ( .o(n11554), .a(n7567_1), .b(n6901) );
oa12f01  g4824 ( .o(n8671), .a(n11554), .b(n6901), .c(n11553) );
na02f01  g4825 ( .o(n11556), .a(n9410_1), .b(n9405_1) );
oa12f01  g4826 ( .o(n8676), .a(n11556), .b(n9409), .c(n9405_1) );
in01f01  g4827 ( .o(n11558), .a(_net_7627) );
na02f01  g4828 ( .o(n11559), .a(n7400_1), .b(n6971) );
oa12f01  g4829 ( .o(n8689), .a(n11559), .b(n7400_1), .c(n11558) );
na02f01  g4830 ( .o(n11561), .a(n6996), .b(_net_6144) );
na02f01  g4831 ( .o(n11562), .a(n9719_1), .b(n6981) );
na02f01  g4832 ( .o(n8694), .a(n11562), .b(n11561) );
na02f01  g4833 ( .o(n11564), .a(n7348), .b(_net_7813) );
oa12f01  g4834 ( .o(n8703), .a(n11564), .b(n7348), .c(n7259) );
ao22f01  g4835 ( .o(n11566), .a(n7298), .b(_net_7731), .c(n7288_1), .d(_net_6042) );
ao22f01  g4836 ( .o(n11567), .a(n7306), .b(_net_5998), .c(n7286), .d(_net_281) );
na02f01  g4837 ( .o(n11568), .a(n7302_1), .b(_net_125) );
na03f01  g4838 ( .o(n11569), .a(n7308), .b(net_167), .c(n6800) );
na03f01  g4839 ( .o(n11570), .a(n7308), .b(net_204), .c(x1322) );
na02f01  g4840 ( .o(n11571), .a(n7296), .b(net_241) );
na03f01  g4841 ( .o(n11572), .a(n11571), .b(n11570), .c(n11569) );
ao12f01  g4842 ( .o(n11573), .a(n11572), .b(n7291), .c(_net_7702) );
na04f01  g4843 ( .o(n8708), .a(n11573), .b(n11568), .c(n11567), .d(n11566) );
in01f01  g4844 ( .o(n11575), .a(_net_7477) );
na02f01  g4845 ( .o(n11576), .a(n8633), .b(n6869) );
oa12f01  g4846 ( .o(n8720), .a(n11576), .b(n6869), .c(n11575) );
na02f01  g4847 ( .o(n11578), .a(n10289), .b(n9617) );
na02f01  g4848 ( .o(n11579), .a(n7134), .b(n7126) );
ao22f01  g4849 ( .o(n11580), .a(n11579), .b(n10291), .c(n8716), .d(_net_6824) );
na02f01  g4850 ( .o(n8725), .a(n11580), .b(n11578) );
na02f01  g4851 ( .o(n11582), .a(n10737), .b(n10736) );
na02f01  g4852 ( .o(n11583), .a(n11582), .b(n7124) );
ao22f01  g4853 ( .o(n11584), .a(n8183_1), .b(n8159), .c(n7119), .d(_net_6109) );
na02f01  g4854 ( .o(n11585), .a(n8187), .b(n8164) );
oa12f01  g4855 ( .o(n11586), .a(n8167), .b(n8681_1), .c(n8678) );
na04f01  g4856 ( .o(n8730), .a(n11586), .b(n11585), .c(n11584), .d(n11583) );
in01f01  g4857 ( .o(n11588), .a(_net_7805) );
na02f01  g4858 ( .o(n11589), .a(n6803), .b(_net_6043) );
oa12f01  g4859 ( .o(n8743), .a(n11589), .b(n6803), .c(n11588) );
in01f01  g4860 ( .o(n11591), .a(_net_7476) );
na02f01  g4861 ( .o(n11592), .a(n7553_1), .b(n6869) );
oa12f01  g4862 ( .o(n8748), .a(n11592), .b(n6869), .c(n11591) );
in01f01  g4863 ( .o(n11594), .a(_net_7585) );
na02f01  g4864 ( .o(n11595), .a(n8246), .b(n6968) );
oa12f01  g4865 ( .o(n8753), .a(n11595), .b(n6968), .c(n11594) );
in01f01  g4866 ( .o(n11597), .a(_net_6288) );
no02f01  g4867 ( .o(n8762), .a(_net_392), .b(n11597) );
ao12f01  g4868 ( .o(n11599), .a(n9671), .b(n10332), .c(n10423) );
no02f01  g4869 ( .o(n11600), .a(n11599), .b(_net_6411) );
no02f01  g4870 ( .o(n8771), .a(n11600), .b(n8177) );
na02f01  g4871 ( .o(n11602), .a(n9105), .b(n8307_1) );
no02f01  g4872 ( .o(n11603), .a(n7583), .b(n9102) );
no02f01  g4873 ( .o(n11604), .a(n7584), .b(_net_7230) );
no02f01  g4874 ( .o(n11605), .a(n11604), .b(n11603) );
ao22f01  g4875 ( .o(n11606), .a(n11605), .b(n8310), .c(n8312), .d(_net_7230) );
na02f01  g4876 ( .o(n8775), .a(n11606), .b(n11602) );
in01f01  g4877 ( .o(n11608), .a(_net_7265) );
na02f01  g4878 ( .o(n11609), .a(n9537_1), .b(n6901) );
oa12f01  g4879 ( .o(n8780), .a(n11609), .b(n6901), .c(n11608) );
na04f01  g4880 ( .o(n8809), .a(n10016), .b(_net_6414), .c(net_6412), .d(n10012) );
in01f01  g4881 ( .o(n11612), .a(_net_7409) );
na02f01  g4882 ( .o(n11613), .a(n7550), .b(n7200) );
oa12f01  g4883 ( .o(n8818), .a(n11613), .b(n7550), .c(n11612) );
ao22f01  g4884 ( .o(n11615), .a(n7225), .b(_net_7403), .c(n7224), .d(_net_7435) );
ao22f01  g4885 ( .o(n11616), .a(n7229), .b(_net_7499), .c(n7228), .d(_net_7467) );
na02f01  g4886 ( .o(n8831), .a(n11616), .b(n11615) );
in01f01  g4887 ( .o(n11618), .a(_net_7664) );
na02f01  g4888 ( .o(n11619), .a(n7446_1), .b(n7403) );
oa12f01  g4889 ( .o(n8840), .a(n11619), .b(n7446_1), .c(n11618) );
in01f01  g4890 ( .o(n11621), .a(_net_6048) );
oa12f01  g4891 ( .o(n8845), .a(n11621), .b(n7572_1), .c(n8695) );
in01f01  g4892 ( .o(n11623), .a(_net_7363) );
na02f01  g4893 ( .o(n11624), .a(n7567_1), .b(n7030) );
oa12f01  g4894 ( .o(n8855), .a(n11624), .b(n7030), .c(n11623) );
in01f01  g4895 ( .o(n11626), .a(_net_7625) );
na02f01  g4896 ( .o(n11627), .a(n10071), .b(n7400_1) );
oa12f01  g4897 ( .o(n8860), .a(n11627), .b(n7400_1), .c(n11626) );
in01f01  g4898 ( .o(n11629), .a(_net_6185) );
no02f01  g4899 ( .o(n8869), .a(_net_392), .b(n11629) );
in01f01  g4900 ( .o(n11631), .a(_net_6297) );
no02f01  g4901 ( .o(n8895), .a(_net_392), .b(n11631) );
na02f01  g4902 ( .o(n11633), .a(n7912), .b(n7575) );
ao22f01  g4903 ( .o(n11634), .a(n7917), .b(n7593), .c(n7591_1), .d(_net_6166) );
na02f01  g4904 ( .o(n8917), .a(n11634), .b(n11633) );
no03f01  g4905 ( .o(n11636), .a(n7360), .b(n10532), .c(n7359_1) );
no02f01  g4906 ( .o(n11637), .a(n7361), .b(_net_7787) );
no03f01  g4907 ( .o(n8922), .a(n11637), .b(n11636), .c(n7358) );
in01f01  g4908 ( .o(n11639), .a(_net_7322) );
na02f01  g4909 ( .o(n11640), .a(n7393), .b(n7150) );
oa12f01  g4910 ( .o(n8948), .a(n11640), .b(n7150), .c(n11639) );
in01f01  g4911 ( .o(n11642), .a(_net_7451) );
na02f01  g4912 ( .o(n11643), .a(n8193), .b(n7197) );
oa12f01  g4913 ( .o(n8953), .a(n11643), .b(n7197), .c(n11642) );
ao22f01  g4914 ( .o(n11645), .a(n7225), .b(_net_7417), .c(n7224), .d(_net_7449) );
ao22f01  g4915 ( .o(n11646), .a(n7229), .b(_net_7513), .c(n7228), .d(_net_7481) );
na02f01  g4916 ( .o(n8967), .a(n11646), .b(n11645) );
in01f01  g4917 ( .o(n11648), .a(_net_7466) );
na02f01  g4918 ( .o(n11649), .a(n7883_1), .b(n6869) );
oa12f01  g4919 ( .o(n8976), .a(n11649), .b(n6869), .c(n11648) );
in01f01  g4920 ( .o(n11651), .a(_net_7581) );
na02f01  g4921 ( .o(n11652), .a(n7519), .b(n698) );
oa12f01  g4922 ( .o(n8986), .a(n11652), .b(n7519), .c(n11651) );
na02f01  g4923 ( .o(n11654), .a(n7440), .b(_net_7813) );
oa12f01  g4924 ( .o(n8995), .a(n11654), .b(n7440), .c(n10191) );
na02f01  g4925 ( .o(n11656), .a(n7440), .b(_net_7794) );
oa12f01  g4926 ( .o(n9000), .a(n11656), .b(n7440), .c(n9966_1) );
na02f01  g4927 ( .o(n11658), .a(n9915), .b(n9306) );
na02f01  g4928 ( .o(n11659), .a(n9914_1), .b(_net_7783) );
na02f01  g4929 ( .o(n11660), .a(n11659), .b(n11658) );
oa22f01  g4930 ( .o(n9005), .a(n11660), .b(n9913), .c(n9313), .d(n9306) );
na02f01  g4931 ( .o(n11662), .a(n7306), .b(_net_6018) );
na02f01  g4932 ( .o(n11663), .a(n7293), .b(net_218) );
ao22f01  g4933 ( .o(n11664), .a(n7297_1), .b(net_181), .c(n7296), .d(net_255) );
ao22f01  g4934 ( .o(n11665), .a(n7298), .b(_net_7745), .c(n7291), .d(_net_7716) );
na04f01  g4935 ( .o(n9030), .a(n11665), .b(n11664), .c(n11663), .d(n11662) );
ao22f01  g4936 ( .o(n11667), .a(n6738), .b(_net_7552), .c(n6736_1), .d(_net_7616) );
ao22f01  g4937 ( .o(n11668), .a(n6739), .b(_net_7648), .c(n6734), .d(_net_7584) );
na02f01  g4938 ( .o(n9042), .a(n11668), .b(n11667) );
in01f01  g4939 ( .o(n11670), .a(_net_7423) );
na02f01  g4940 ( .o(n11671), .a(n7550), .b(n634) );
oa12f01  g4941 ( .o(n9052), .a(n11671), .b(n7550), .c(n11670) );
in01f01  g4942 ( .o(n11673), .a(_net_115) );
na02f01  g4943 ( .o(n11674), .a(net_311), .b(_net_154) );
oa12f01  g4944 ( .o(n9074), .a(n11674), .b(n11673), .c(_net_154) );
ao22f01  g4945 ( .o(n11676), .a(n6736_1), .b(net_7642), .c(n6734), .d(net_7610) );
ao22f01  g4946 ( .o(n11677), .a(n6739), .b(net_7674), .c(n6738), .d(_net_7578) );
na02f01  g4947 ( .o(n9096), .a(n11677), .b(n11676) );
na02f01  g4948 ( .o(n11679), .a(n7440), .b(_net_7809) );
oa12f01  g4949 ( .o(n9101), .a(n11679), .b(n7440), .c(n8236) );
in01f01  g4950 ( .o(n11681), .a(_net_7716) );
na02f01  g4951 ( .o(n11682), .a(n7207_1), .b(_net_7818) );
oa12f01  g4952 ( .o(n9106), .a(n11682), .b(n7207_1), .c(n11681) );
na02f01  g4953 ( .o(n11684), .a(n7440), .b(_net_7812) );
oa12f01  g4954 ( .o(n9115), .a(n11684), .b(n7440), .c(n7143) );
in01f01  g4955 ( .o(n11686), .a(_net_7558) );
na02f01  g4956 ( .o(n11687), .a(n7644_1), .b(n7519) );
oa12f01  g4957 ( .o(n9124), .a(n11687), .b(n7519), .c(n11686) );
in01f01  g4958 ( .o(n11689), .a(_net_7660) );
na02f01  g4959 ( .o(n11690), .a(n8043), .b(n7446_1) );
oa12f01  g4960 ( .o(n9129), .a(n11690), .b(n7446_1), .c(n11689) );
ao22f01  g4961 ( .o(n11692), .a(n6877), .b(_net_7256), .c(n6876_1), .d(_net_7320) );
ao22f01  g4962 ( .o(n11693), .a(n6881_1), .b(_net_7288), .c(n6880), .d(_net_7352) );
na02f01  g4963 ( .o(n9151), .a(n11693), .b(n11692) );
in01f01  g4964 ( .o(n11695), .a(_net_7259) );
na02f01  g4965 ( .o(n11696), .a(n7033), .b(n6901) );
oa12f01  g4966 ( .o(n9156), .a(n11696), .b(n6901), .c(n11695) );
in01f01  g4967 ( .o(n11698), .a(_net_6187) );
no02f01  g4968 ( .o(n9173), .a(_net_392), .b(n11698) );
in01f01  g4969 ( .o(n11700), .a(_net_7260) );
na02f01  g4970 ( .o(n11701), .a(n10089_1), .b(n6901) );
oa12f01  g4971 ( .o(n9187), .a(n11701), .b(n6901), .c(n11700) );
ao22f01  g4972 ( .o(n11703), .a(n6877), .b(_net_7266), .c(n6876_1), .d(_net_7330) );
ao22f01  g4973 ( .o(n11704), .a(n6881_1), .b(_net_7298), .c(n6880), .d(_net_7362) );
na02f01  g4974 ( .o(n9192), .a(n11704), .b(n11703) );
no02f01  g4975 ( .o(n11706), .a(n6739), .b(n8349) );
no03f01  g4976 ( .o(n11707), .a(_net_7682), .b(n6733), .c(n6735) );
no02f01  g4977 ( .o(n11708), .a(n11707), .b(n11706) );
oa22f01  g4978 ( .o(n9201), .a(n11708), .b(n10455), .c(n10456), .d(n8349) );
in01f01  g4979 ( .o(n11710), .a(_net_5986) );
na02f01  g4980 ( .o(n11711), .a(n7348), .b(_net_7795) );
oa12f01  g4981 ( .o(n9206), .a(n11711), .b(n7348), .c(n11710) );
in01f01  g4982 ( .o(n11713), .a(n9347) );
no02f01  g4983 ( .o(n9211), .a(n11713), .b(x940) );
no02f01  g4984 ( .o(n11715), .a(n9283), .b(n6945) );
no02f01  g4985 ( .o(n11716), .a(n9292), .b(n6934_1) );
in01f01  g4986 ( .o(n11717), .a(_net_6094) );
oa22f01  g4987 ( .o(n11718), .a(n10132_1), .b(n6916), .c(n6932), .d(n11717) );
no03f01  g4988 ( .o(n11719), .a(n11718), .b(n11716), .c(n11715) );
in01f01  g4989 ( .o(n11720), .a(net_6613) );
in01f01  g4990 ( .o(n11721), .a(net_6581) );
oa22f01  g4991 ( .o(n11722), .a(n7058_1), .b(n11721), .c(n7057), .d(n11720) );
in01f01  g4992 ( .o(n11723), .a(net_6677) );
in01f01  g4993 ( .o(n11724), .a(net_6645) );
oa22f01  g4994 ( .o(n11725), .a(n7063), .b(n11723), .c(n7062_1), .d(n11724) );
no02f01  g4995 ( .o(n11726), .a(n11725), .b(n11722) );
na02f01  g4996 ( .o(n9220), .a(n11726), .b(n11719) );
in01f01  g4997 ( .o(n11728), .a(_net_7701) );
na02f01  g4998 ( .o(n11729), .a(n7207_1), .b(_net_7803) );
oa12f01  g4999 ( .o(n9233), .a(n11729), .b(n7207_1), .c(n11728) );
na02f01  g5000 ( .o(n11731), .a(_net_6405), .b(n8088_1) );
na03f01  g5001 ( .o(n9258), .a(n11731), .b(n8090), .c(n6910_1) );
in01f01  g5002 ( .o(n11733), .a(_net_7515) );
na02f01  g5003 ( .o(n11734), .a(n8193), .b(n7626_1) );
oa12f01  g5004 ( .o(n9263), .a(n11734), .b(n7626_1), .c(n11733) );
no02f01  g5005 ( .o(n11736), .a(n7228), .b(n7224) );
oa22f01  g5006 ( .o(n9272), .a(n11736), .b(n8872), .c(n8873_1), .d(n7227) );
na02f01  g5007 ( .o(n11738), .a(n8162), .b(n7124) );
ao22f01  g5008 ( .o(n11739), .a(n8159), .b(n7137), .c(n7119), .d(_net_6106) );
na02f01  g5009 ( .o(n9277), .a(n11739), .b(n11738) );
no02f01  g5010 ( .o(n11741), .a(n6843), .b(n6824) );
no02f01  g5011 ( .o(n11742), .a(n7612), .b(n6826_1) );
in01f01  g5012 ( .o(n11743), .a(_net_6137) );
oa22f01  g5013 ( .o(n11744), .a(n8397), .b(n6836_1), .c(n6844), .d(n11743) );
no03f01  g5014 ( .o(n11745), .a(n11744), .b(n11742), .c(n11741) );
in01f01  g5015 ( .o(n11746), .a(net_6886) );
in01f01  g5016 ( .o(n11747), .a(net_6854) );
oa22f01  g5017 ( .o(n11748), .a(n6850_1), .b(n11747), .c(n6849), .d(n11746) );
in01f01  g5018 ( .o(n11749), .a(net_6918) );
in01f01  g5019 ( .o(n11750), .a(net_6950) );
oa22f01  g5020 ( .o(n11751), .a(n6855_1), .b(n11750), .c(n6854), .d(n11749) );
no02f01  g5021 ( .o(n11752), .a(n11751), .b(n11748) );
na02f01  g5022 ( .o(n9282), .a(n11752), .b(n11745) );
in01f01  g5023 ( .o(n11754), .a(_net_7516) );
na02f01  g5024 ( .o(n11755), .a(n9872), .b(n7626_1) );
oa12f01  g5025 ( .o(n9307), .a(n11755), .b(n7626_1), .c(n11754) );
in01f01  g5026 ( .o(n11757), .a(_net_7726) );
ao12f01  g5027 ( .o(n9312), .a(n7343), .b(n11757), .c(n7190_1) );
ao22f01  g5028 ( .o(n11759), .a(n7225), .b(_net_7427), .c(n7224), .d(net_7459) );
ao22f01  g5029 ( .o(n11760), .a(n7229), .b(net_7523), .c(n7228), .d(net_7491) );
na02f01  g5030 ( .o(n9321), .a(n11760), .b(n11759) );
no02f01  g5031 ( .o(n9330), .a(n10938), .b(n9893) );
in01f01  g5032 ( .o(n11763), .a(net_6003) );
in01f01  g5033 ( .o(n11764), .a(_net_7725) );
ao12f01  g5034 ( .o(n9335), .a(n7343), .b(n11764), .c(n11763) );
in01f01  g5035 ( .o(n11766), .a(_net_7504) );
na02f01  g5036 ( .o(n11767), .a(n8141), .b(n7626_1) );
oa12f01  g5037 ( .o(n9352), .a(n11767), .b(n7626_1), .c(n11766) );
in01f01  g5038 ( .o(n11769), .a(_net_7569) );
na02f01  g5039 ( .o(n11770), .a(n9318), .b(n7519) );
oa12f01  g5040 ( .o(n9410), .a(n11770), .b(n7519), .c(n11769) );
na02f01  g5041 ( .o(n11772), .a(n6933), .b(_net_6085) );
na02f01  g5042 ( .o(n11773), .a(n8009), .b(n6917) );
na02f01  g5043 ( .o(n9415), .a(n11773), .b(n11772) );
in01f01  g5044 ( .o(n11775), .a(_net_7317) );
na02f01  g5045 ( .o(n11776), .a(n7183), .b(n7150) );
oa12f01  g5046 ( .o(n9420), .a(n11776), .b(n7150), .c(n11775) );
in01f01  g5047 ( .o(n11778), .a(_net_7745) );
in01f01  g5048 ( .o(n11779), .a(_net_288) );
ao12f01  g5049 ( .o(n9436), .a(n7343), .b(n11779), .c(n11778) );
ao22f01  g5050 ( .o(n11781), .a(n7288_1), .b(net_6035), .c(n7286), .d(net_274) );
ao22f01  g5051 ( .o(n11782), .a(n7298), .b(_net_7727), .c(n7291), .d(_net_7698) );
na02f01  g5052 ( .o(n11783), .a(n7302_1), .b(_net_121) );
na03f01  g5053 ( .o(n11784), .a(n7308), .b(net_200), .c(x1322) );
na02f01  g5054 ( .o(n11785), .a(n7296), .b(net_237) );
na03f01  g5055 ( .o(n11786), .a(n7308), .b(net_163), .c(n6800) );
na03f01  g5056 ( .o(n11787), .a(n11786), .b(n11785), .c(n11784) );
ao12f01  g5057 ( .o(n11788), .a(n11787), .b(n7306), .c(_net_5991) );
na04f01  g5058 ( .o(n9441), .a(n11788), .b(n11783), .c(n11782), .d(n11781) );
in01f01  g5059 ( .o(n11790), .a(_net_6319) );
no02f01  g5060 ( .o(n9449), .a(_net_392), .b(n11790) );
ao12f01  g5061 ( .o(n11792), .a(n7067_1), .b(_net_6693), .c(_net_6690) );
oa12f01  g5062 ( .o(n11793), .a(n11792), .b(_net_6693), .c(_net_6690) );
na02f01  g5063 ( .o(n11794), .a(n7665), .b(n548) );
oa12f01  g5064 ( .o(n9454), .a(n9971_1), .b(n11794), .c(n11793) );
in01f01  g5065 ( .o(n11796), .a(_net_7415) );
na02f01  g5066 ( .o(n11797), .a(n7550), .b(n7504) );
oa12f01  g5067 ( .o(n9487), .a(n11797), .b(n7550), .c(n11796) );
in01f01  g5068 ( .o(n11799), .a(_net_7282) );
na02f01  g5069 ( .o(n11800), .a(n8731), .b(n7180) );
oa12f01  g5070 ( .o(n9492), .a(n11800), .b(n7180), .c(n11799) );
in01f01  g5071 ( .o(n11802), .a(_net_7597) );
na02f01  g5072 ( .o(n11803), .a(n7428), .b(n6968) );
oa12f01  g5073 ( .o(n9497), .a(n11803), .b(n6968), .c(n11802) );
in01f01  g5074 ( .o(n11805), .a(_net_7617) );
na02f01  g5075 ( .o(n11806), .a(n8246), .b(n7400_1) );
oa12f01  g5076 ( .o(n9507), .a(n11806), .b(n7400_1), .c(n11805) );
in01f01  g5077 ( .o(n11808), .a(_net_7616) );
na02f01  g5078 ( .o(n11809), .a(n8842), .b(n7400_1) );
oa12f01  g5079 ( .o(n9512), .a(n11809), .b(n7400_1), .c(n11808) );
ao22f01  g5080 ( .o(n11811), .a(n7225), .b(_net_7425), .c(n7224), .d(net_7457) );
ao22f01  g5081 ( .o(n11812), .a(n7229), .b(net_7521), .c(n7228), .d(net_7489) );
na02f01  g5082 ( .o(n9533), .a(n11812), .b(n11811) );
ao22f01  g5083 ( .o(n11814), .a(net_7739), .b(net_7710), .c(net_7737), .d(net_7708) );
ao22f01  g5084 ( .o(n11815), .a(net_7740), .b(net_7711), .c(net_7742), .d(net_7713) );
ao22f01  g5085 ( .o(n11816), .a(_net_7705), .b(_net_7734), .c(_net_7736), .d(_net_7707) );
ao22f01  g5086 ( .o(n11817), .a(net_7709), .b(net_7738), .c(_net_7733), .d(_net_7704) );
na04f01  g5087 ( .o(n11818), .a(n11817), .b(n11816), .c(n11815), .d(n11814) );
na02f01  g5088 ( .o(n11819), .a(_net_7745), .b(_net_7716) );
ao22f01  g5089 ( .o(n11820), .a(_net_7717), .b(_net_7746), .c(_net_7719), .d(_net_7748) );
ao22f01  g5090 ( .o(n11821), .a(net_7715), .b(net_7744), .c(net_7714), .d(net_7743) );
ao22f01  g5091 ( .o(n11822), .a(net_7712), .b(net_7741), .c(_net_7718), .d(_net_7747) );
na04f01  g5092 ( .o(n11823), .a(n11822), .b(n11821), .c(n11820), .d(n11819) );
no02f01  g5093 ( .o(n11824), .a(n11823), .b(n11818) );
ao22f01  g5094 ( .o(n11825), .a(_net_7723), .b(_net_7694), .c(net_7691), .d(_net_7720) );
ao22f01  g5095 ( .o(n11826), .a(_net_7693), .b(_net_7722), .c(_net_7721), .d(_net_7692) );
ao22f01  g5096 ( .o(n11827), .a(_net_7695), .b(_net_7724), .c(_net_7727), .d(_net_7698) );
na03f01  g5097 ( .o(n11828), .a(n11827), .b(n11826), .c(n11825) );
ao22f01  g5098 ( .o(n11829), .a(_net_7702), .b(_net_7731), .c(_net_7700), .d(_net_7729) );
ao22f01  g5099 ( .o(n11830), .a(_net_7735), .b(_net_7706), .c(_net_7703), .d(_net_7732) );
ao22f01  g5100 ( .o(n11831), .a(_net_7726), .b(_net_7697), .c(_net_7699), .d(_net_7728) );
ao22f01  g5101 ( .o(n11832), .a(_net_7725), .b(_net_7696), .c(_net_7701), .d(_net_7730) );
na04f01  g5102 ( .o(n11833), .a(n11832), .b(n11831), .c(n11830), .d(n11829) );
no02f01  g5103 ( .o(n11834), .a(n11833), .b(n11828) );
na02f01  g5104 ( .o(n9546), .a(n11834), .b(n11824) );
in01f01  g5105 ( .o(n11836), .a(net_7756) );
na04f01  g5106 ( .o(n11837), .a(_net_6017), .b(_net_7791), .c(net_303), .d(n11836) );
ao12f01  g5107 ( .o(n9554), .a(n11837), .b(net_306), .c(_net_6018) );
no04f01  g5108 ( .o(n9559), .a(n10024), .b(n7292_1), .c(x1215), .d(x1322) );
na02f01  g5109 ( .o(n11840), .a(n7348), .b(_net_7821) );
oa12f01  g5110 ( .o(n9564), .a(n11840), .b(n7348), .c(n7692) );
in01f01  g5111 ( .o(n11842), .a(_net_7509) );
na02f01  g5112 ( .o(n11843), .a(n8633), .b(n7626_1) );
oa12f01  g5113 ( .o(n9569), .a(n11843), .b(n7626_1), .c(n11842) );
no03f01  g5114 ( .o(n11845), .a(n8236), .b(_net_293), .c(n9540) );
no02f01  g5115 ( .o(n11846), .a(n8236), .b(n7653) );
ao22f01  g5116 ( .o(n11847), .a(n11846), .b(n10197), .c(n11845), .d(n10201) );
ao12f01  g5117 ( .o(n11848), .a(n8236), .b(_net_266), .c(n7653) );
no03f01  g5118 ( .o(n11849), .a(n8236), .b(_net_293), .c(_net_294) );
ao22f01  g5119 ( .o(n11850), .a(n11849), .b(n10199), .c(n11848), .d(n10192) );
na02f01  g5120 ( .o(n9574), .a(n11850), .b(n11847) );
in01f01  g5121 ( .o(n11852), .a(_net_7506) );
na02f01  g5122 ( .o(n11853), .a(n7626_1), .b(n6891) );
oa12f01  g5123 ( .o(n9583), .a(n11853), .b(n7626_1), .c(n11852) );
no03f01  g5124 ( .o(n11855), .a(n9339_1), .b(n6976), .c(_net_6032) );
no02f01  g5125 ( .o(n11856), .a(n6976), .b(n7316_1) );
ao22f01  g5126 ( .o(n11857), .a(n11856), .b(n9345), .c(n11855), .d(n9343_1) );
ao12f01  g5127 ( .o(n11858), .a(n6976), .b(n7316_1), .c(_net_5978) );
no03f01  g5128 ( .o(n11859), .a(_net_6033), .b(n6976), .c(_net_6032) );
ao22f01  g5129 ( .o(n11860), .a(n11859), .b(n9341), .c(n11858), .d(n9335_1) );
na02f01  g5130 ( .o(n9592), .a(n11860), .b(n11857) );
ao12f01  g5131 ( .o(n11862), .a(n7012), .b(n10472), .c(n10471) );
no02f01  g5132 ( .o(n11863), .a(n8052), .b(n6997) );
in01f01  g5133 ( .o(n11864), .a(_net_6153) );
oa22f01  g5134 ( .o(n11865), .a(n8060), .b(n6980), .c(n6995_1), .d(n11864) );
no03f01  g5135 ( .o(n11866), .a(n11865), .b(n11863), .c(n11862) );
in01f01  g5136 ( .o(n11867), .a(net_6985) );
in01f01  g5137 ( .o(n11868), .a(net_7017) );
oa22f01  g5138 ( .o(n11869), .a(n8075_1), .b(n11867), .c(n8074), .d(n11868) );
in01f01  g5139 ( .o(n11870), .a(net_7081) );
in01f01  g5140 ( .o(n11871), .a(net_7049) );
oa22f01  g5141 ( .o(n11872), .a(n8080_1), .b(n11870), .c(n8079), .d(n11871) );
no02f01  g5142 ( .o(n11873), .a(n11872), .b(n11869) );
na02f01  g5143 ( .o(n9597), .a(n11873), .b(n11866) );
in01f01  g5144 ( .o(n11875), .a(_net_7324) );
na02f01  g5145 ( .o(n11876), .a(n10089_1), .b(n7150) );
oa12f01  g5146 ( .o(n9602), .a(n11876), .b(n7150), .c(n11875) );
in01f01  g5147 ( .o(n11878), .a(n8177) );
no03f01  g5148 ( .o(n9616), .a(n9819_1), .b(n8178), .c(n11878) );
in01f01  g5149 ( .o(n11880), .a(_net_7436) );
na02f01  g5150 ( .o(n11881), .a(n7952), .b(n7197) );
oa12f01  g5151 ( .o(n9633), .a(n11881), .b(n7197), .c(n11880) );
in01f01  g5152 ( .o(n11883), .a(_net_7414) );
na02f01  g5153 ( .o(n11884), .a(n8994), .b(n7550) );
oa12f01  g5154 ( .o(n9638), .a(n11884), .b(n7550), .c(n11883) );
in01f01  g5155 ( .o(n11886), .a(_net_7327) );
na02f01  g5156 ( .o(n11887), .a(n7994_1), .b(n7150) );
oa12f01  g5157 ( .o(n9655), .a(n11887), .b(n7150), .c(n11886) );
in01f01  g5158 ( .o(n11889), .a(_net_7656) );
na02f01  g5159 ( .o(n11890), .a(n9881), .b(n7446_1) );
oa12f01  g5160 ( .o(n9664), .a(n11890), .b(n7446_1), .c(n11889) );
in01f01  g5161 ( .o(n11892), .a(_net_7588) );
na02f01  g5162 ( .o(n11893), .a(n8426_1), .b(n6968) );
oa12f01  g5163 ( .o(n9673), .a(n11893), .b(n6968), .c(n11892) );
no04f01  g5164 ( .o(n9678), .a(n8925), .b(n8915), .c(n6867_1), .d(_net_7532) );
in01f01  g5165 ( .o(n11896), .a(_net_7560) );
na02f01  g5166 ( .o(n11897), .a(n9881), .b(n7519) );
oa12f01  g5167 ( .o(n9683), .a(n11897), .b(n7519), .c(n11896) );
na02f01  g5168 ( .o(n11899), .a(n8124), .b(_net_6693) );
na03f01  g5169 ( .o(n11900), .a(n8123), .b(n8121_1), .c(n9973) );
na02f01  g5170 ( .o(n11901), .a(n8936), .b(net_6691) );
na03f01  g5171 ( .o(n11902), .a(n8935), .b(n8934_1), .c(n7153) );
ao22f01  g5172 ( .o(n11903), .a(n11902), .b(n11901), .c(n6944), .d(_net_6687) );
na02f01  g5173 ( .o(n11904), .a(n10364), .b(n7663) );
na03f01  g5174 ( .o(n11905), .a(n10363), .b(n10362), .c(_net_6692) );
na03f01  g5175 ( .o(n11906), .a(n11905), .b(n11904), .c(n11903) );
ao12f01  g5176 ( .o(n9700), .a(n11906), .b(n11900), .c(n11899) );
na02f01  g5177 ( .o(n11908), .a(n10421), .b(_net_6406) );
no04f01  g5178 ( .o(n9709), .a(n11908), .b(n10424), .c(n11878), .d(n8090) );
no02f01  g5179 ( .o(n11910), .a(n8406), .b(n6824) );
no02f01  g5180 ( .o(n11911), .a(n11539), .b(n6826_1) );
ao22f01  g5181 ( .o(n11912), .a(n6811), .b(net_6848), .c(n6808), .d(net_6912) );
ao22f01  g5182 ( .o(n11913), .a(n6816), .b(net_6880), .c(n6814), .d(net_6944) );
ao12f01  g5183 ( .o(n11914), .a(n6836_1), .b(n11913), .c(n11912) );
in01f01  g5184 ( .o(n11915), .a(_net_6143) );
no02f01  g5185 ( .o(n11916), .a(n6844), .b(n11915) );
no04f01  g5186 ( .o(n11917), .a(n11916), .b(n11914), .c(n11911), .d(n11910) );
in01f01  g5187 ( .o(n11918), .a(net_6860) );
in01f01  g5188 ( .o(n11919), .a(net_6892) );
oa22f01  g5189 ( .o(n11920), .a(n6850_1), .b(n11918), .c(n6849), .d(n11919) );
in01f01  g5190 ( .o(n11921), .a(net_6924) );
in01f01  g5191 ( .o(n11922), .a(net_6956) );
oa22f01  g5192 ( .o(n11923), .a(n6855_1), .b(n11922), .c(n6854), .d(n11921) );
no02f01  g5193 ( .o(n11924), .a(n11923), .b(n11920) );
na02f01  g5194 ( .o(n9714), .a(n11924), .b(n11917) );
no02f01  g5195 ( .o(n11926), .a(n9757), .b(n7721) );
no02f01  g5196 ( .o(n11927), .a(n9766), .b(n7592) );
in01f01  g5197 ( .o(n11928), .a(_net_6174) );
oa22f01  g5198 ( .o(n11929), .a(n11480), .b(n7574), .c(n7590), .d(n11928) );
no03f01  g5199 ( .o(n11930), .a(n11929), .b(n11927), .c(n11926) );
in01f01  g5200 ( .o(n11931), .a(net_7153) );
in01f01  g5201 ( .o(n11932), .a(net_7121) );
oa22f01  g5202 ( .o(n11933), .a(n7740), .b(n11932), .c(n7739), .d(n11931) );
in01f01  g5203 ( .o(n11934), .a(net_7217) );
in01f01  g5204 ( .o(n11935), .a(net_7185) );
oa22f01  g5205 ( .o(n11936), .a(n7745), .b(n11934), .c(n7744), .d(n11935) );
no02f01  g5206 ( .o(n11937), .a(n11936), .b(n11933) );
na02f01  g5207 ( .o(n9719), .a(n11937), .b(n11930) );
no02f01  g5208 ( .o(n11939), .a(n7026), .b(net_7378) );
in01f01  g5209 ( .o(n11940), .a(n11939) );
no02f01  g5210 ( .o(n11941), .a(n11940), .b(n9437) );
no02f01  g5211 ( .o(n11942), .a(n11939), .b(n9438) );
oa12f01  g5212 ( .o(n11943), .a(n9197), .b(n11942), .c(n11941) );
no02f01  g5213 ( .o(n11944), .a(n11942), .b(n11941) );
na02f01  g5214 ( .o(n11945), .a(n11944), .b(n3464) );
na02f01  g5215 ( .o(n9733), .a(n11945), .b(n11943) );
ao22f01  g5216 ( .o(n11947), .a(n6877), .b(_net_7264), .c(n6876_1), .d(_net_7328) );
ao22f01  g5217 ( .o(n11948), .a(n6881_1), .b(_net_7296), .c(n6880), .d(_net_7360) );
na02f01  g5218 ( .o(n9742), .a(n11948), .b(n11947) );
in01f01  g5219 ( .o(n11950), .a(_net_7576) );
na02f01  g5220 ( .o(n11951), .a(n2404), .b(n7519) );
oa12f01  g5221 ( .o(n9763), .a(n11951), .b(n7519), .c(n11950) );
in01f01  g5222 ( .o(n11953), .a(_net_7283) );
na02f01  g5223 ( .o(n11954), .a(n7659), .b(n7180) );
oa12f01  g5224 ( .o(n9768), .a(n11954), .b(n7180), .c(n11953) );
in01f01  g5225 ( .o(n11956), .a(_net_6002) );
na02f01  g5226 ( .o(n11957), .a(n7348), .b(_net_7808) );
oa12f01  g5227 ( .o(n9773), .a(n11957), .b(n7348), .c(n11956) );
in01f01  g5228 ( .o(n11959), .a(_net_7566) );
na02f01  g5229 ( .o(n11960), .a(n9373_1), .b(n7519) );
oa12f01  g5230 ( .o(n9787), .a(n11960), .b(n7519), .c(n11959) );
na02f01  g5231 ( .o(n11962), .a(n7348), .b(_net_7798) );
oa12f01  g5232 ( .o(n9792), .a(n11962), .b(n7348), .c(n7535_1) );
na02f01  g5233 ( .o(n11964), .a(n7028), .b(_net_7384) );
na02f01  g5234 ( .o(n11965), .a(n7029), .b(n9441_1) );
na03f01  g5235 ( .o(n11966), .a(n11965), .b(n11964), .c(n9852) );
na03f01  g5236 ( .o(n11967), .a(_net_7383), .b(_net_7381), .c(_net_7382) );
na02f01  g5237 ( .o(n11968), .a(n11967), .b(n9441_1) );
in01f01  g5238 ( .o(n11969), .a(n11967) );
na02f01  g5239 ( .o(n11970), .a(n11969), .b(_net_7384) );
na03f01  g5240 ( .o(n11971), .a(n11970), .b(n11968), .c(n9858_1) );
na02f01  g5241 ( .o(n11972), .a(n9860), .b(_net_7384) );
na03f01  g5242 ( .o(n9801), .a(n11972), .b(n11971), .c(n11966) );
in01f01  g5243 ( .o(n11974), .a(_net_5859) );
in01f01  g5244 ( .o(n11975), .a(x1062) );
na03f01  g5245 ( .o(n11976), .a(n11385), .b(net_7772), .c(n11975) );
oa12f01  g5246 ( .o(n9814), .a(n11976), .b(n11974), .c(x1062) );
na02f01  g5247 ( .o(n11978), .a(n7852), .b(n7194_1) );
no02f01  g5248 ( .o(n11979), .a(_net_7533), .b(n7846) );
no02f01  g5249 ( .o(n11980), .a(n7194_1), .b(_net_7532) );
oa12f01  g5250 ( .o(n11981), .a(n7845_1), .b(n11980), .c(n11979) );
na02f01  g5251 ( .o(n11982), .a(n7854), .b(_net_7533) );
na03f01  g5252 ( .o(n9819), .a(n11982), .b(n11981), .c(n11978) );
oa12f01  g5253 ( .o(n11984), .a(n7027_1), .b(n9854), .c(n7026) );
na03f01  g5254 ( .o(n11985), .a(n11984), .b(n11967), .c(n9858_1) );
na02f01  g5255 ( .o(n11986), .a(n7179), .b(n7149) );
ao22f01  g5256 ( .o(n11987), .a(n11986), .b(n9852), .c(n9860), .d(_net_7383) );
na02f01  g5257 ( .o(n9824), .a(n11987), .b(n11985) );
in01f01  g5258 ( .o(n11989), .a(_net_7421) );
na02f01  g5259 ( .o(n11990), .a(n1277), .b(n7550) );
oa12f01  g5260 ( .o(n9849), .a(n11990), .b(n7550), .c(n11989) );
na02f01  g5261 ( .o(n11992), .a(n9260), .b(n10421) );
oa12f01  g5262 ( .o(n11993), .a(_net_6407), .b(n9259), .c(n9258_1) );
na03f01  g5263 ( .o(n9858), .a(n11993), .b(n11992), .c(n6910_1) );
no02f01  g5264 ( .o(n11995), .a(_net_7097), .b(n8385) );
no02f01  g5265 ( .o(n11996), .a(n8760), .b(net_7096) );
no02f01  g5266 ( .o(n11997), .a(n11996), .b(n11995) );
oa22f01  g5267 ( .o(n9863), .a(n11997), .b(n10574), .c(n10578), .d(n8760) );
in01f01  g5268 ( .o(n11999), .a(n9665) );
na02f01  g5269 ( .o(n12000), .a(n9664_1), .b(n9663) );
na02f01  g5270 ( .o(n12001), .a(n12000), .b(n11999) );
oa22f01  g5271 ( .o(n9880), .a(n12001), .b(n9411), .c(n9409), .d(n9663) );
oa12f01  g5272 ( .o(n12003), .a(n7124), .b(n10744), .c(n10741) );
ao22f01  g5273 ( .o(n12004), .a(n11582), .b(n8159), .c(n7119), .d(_net_6111) );
na02f01  g5274 ( .o(n12005), .a(n11415), .b(n11414) );
ao22f01  g5275 ( .o(n12006), .a(n12005), .b(n8167), .c(n8183_1), .d(n8164) );
na03f01  g5276 ( .o(n9889), .a(n12006), .b(n12004), .c(n12003) );
in01f01  g5277 ( .o(n12008), .a(_net_287) );
na02f01  g5278 ( .o(n12009), .a(_net_225), .b(_net_227) );
na02f01  g5279 ( .o(n9894), .a(n12009), .b(n12008) );
na02f01  g5280 ( .o(n12011), .a(n7298), .b(net_7740) );
ao22f01  g5281 ( .o(n12012), .a(n7306), .b(_net_6010), .c(n7291), .d(net_7711) );
na02f01  g5282 ( .o(n12013), .a(n7302_1), .b(net_150) );
na02f01  g5283 ( .o(n12014), .a(n7296), .b(net_250) );
na03f01  g5284 ( .o(n12015), .a(n7308), .b(_net_176), .c(n6800) );
na03f01  g5285 ( .o(n12016), .a(n7308), .b(_net_213), .c(x1322) );
na03f01  g5286 ( .o(n12017), .a(n12016), .b(n12015), .c(n12014) );
ao12f01  g5287 ( .o(n12018), .a(n12017), .b(n7286), .c(_net_293) );
na04f01  g5288 ( .o(n9907), .a(n12018), .b(n12013), .c(n12012), .d(n12011) );
oa12f01  g5289 ( .o(n9939), .a(n11779), .b(n7851), .c(n7410) );
in01f01  g5290 ( .o(n12021), .a(_net_7348) );
na02f01  g5291 ( .o(n12022), .a(n7030), .b(n6904) );
oa12f01  g5292 ( .o(n9949), .a(n12022), .b(n7030), .c(n12021) );
in01f01  g5293 ( .o(n12024), .a(_net_7402) );
na02f01  g5294 ( .o(n12025), .a(n7883_1), .b(n7550) );
oa12f01  g5295 ( .o(n9966), .a(n12025), .b(n7550), .c(n12024) );
no02f01  g5296 ( .o(n12027), .a(n10554), .b(n6764) );
no02f01  g5297 ( .o(n12028), .a(n9225_1), .b(n6766) );
in01f01  g5298 ( .o(n12029), .a(_net_6076) );
oa22f01  g5299 ( .o(n12030), .a(n9233_1), .b(n6775), .c(n6784), .d(n12029) );
no03f01  g5300 ( .o(n12031), .a(n12030), .b(n12028), .c(n12027) );
in01f01  g5301 ( .o(n12032), .a(net_6448) );
in01f01  g5302 ( .o(n12033), .a(net_6480) );
oa22f01  g5303 ( .o(n12034), .a(n6790), .b(n12032), .c(n6789), .d(n12033) );
in01f01  g5304 ( .o(n12035), .a(net_6512) );
in01f01  g5305 ( .o(n12036), .a(net_6544) );
oa22f01  g5306 ( .o(n12037), .a(n6795), .b(n12036), .c(n6794), .d(n12035) );
no02f01  g5307 ( .o(n12038), .a(n12037), .b(n12034) );
na02f01  g5308 ( .o(n9971), .a(n12038), .b(n12031) );
no02f01  g5309 ( .o(n12040), .a(n11636), .b(_net_7788) );
no03f01  g5310 ( .o(n9981), .a(n12040), .b(n10533), .c(n7358) );
in01f01  g5311 ( .o(n12042), .a(_net_7717) );
na02f01  g5312 ( .o(n12043), .a(n7207_1), .b(_net_7819) );
oa12f01  g5313 ( .o(n9997), .a(n12043), .b(n7207_1), .c(n12042) );
na02f01  g5314 ( .o(n12045), .a(n7440), .b(_net_7793) );
oa12f01  g5315 ( .o(n10019), .a(n12045), .b(n7440), .c(n8094) );
in01f01  g5316 ( .o(n12047), .a(_net_7582) );
na02f01  g5317 ( .o(n12048), .a(n3604), .b(n7519) );
oa12f01  g5318 ( .o(n10032), .a(n12048), .b(n7519), .c(n12047) );
na02f01  g5319 ( .o(n12050), .a(n7348), .b(_net_7817) );
oa12f01  g5320 ( .o(n10037), .a(n12050), .b(n7348), .c(n6819) );
in01f01  g5321 ( .o(n12052), .a(_net_6202) );
no02f01  g5322 ( .o(n10042), .a(_net_392), .b(n12052) );
in01f01  g5323 ( .o(n12054), .a(_net_7287) );
na02f01  g5324 ( .o(n12055), .a(n8022), .b(n7180) );
oa12f01  g5325 ( .o(n10052), .a(n12055), .b(n7180), .c(n12054) );
in01f01  g5326 ( .o(n12057), .a(n10633) );
no02f01  g5327 ( .o(n10061), .a(n12057), .b(x1034) );
ao22f01  g5328 ( .o(n12059), .a(n7306), .b(_net_5995), .c(n7291), .d(_net_7699) );
ao22f01  g5329 ( .o(n12060), .a(n7288_1), .b(_net_6039), .c(n7286), .d(_net_278) );
na02f01  g5330 ( .o(n12061), .a(n7302_1), .b(_net_122) );
na03f01  g5331 ( .o(n12062), .a(n7308), .b(_net_201), .c(x1322) );
na02f01  g5332 ( .o(n12063), .a(n7296), .b(net_238) );
na03f01  g5333 ( .o(n12064), .a(n7308), .b(net_164), .c(n6800) );
na03f01  g5334 ( .o(n12065), .a(n12064), .b(n12063), .c(n12062) );
ao12f01  g5335 ( .o(n12066), .a(n12065), .b(n7298), .c(_net_7728) );
na04f01  g5336 ( .o(n10066), .a(n12066), .b(n12061), .c(n12060), .d(n12059) );
in01f01  g5337 ( .o(n12068), .a(_net_7251) );
na02f01  g5338 ( .o(n12069), .a(n7659), .b(n6901) );
oa12f01  g5339 ( .o(n10074), .a(n12069), .b(n6901), .c(n12068) );
na02f01  g5340 ( .o(n12071), .a(n8861), .b(n7754) );
no02f01  g5341 ( .o(n12072), .a(n6754), .b(n7749) );
no02f01  g5342 ( .o(n12073), .a(n6779_1), .b(_net_6555) );
no02f01  g5343 ( .o(n12074), .a(n12073), .b(n12072) );
ao22f01  g5344 ( .o(n12075), .a(n12074), .b(n8859), .c(n8862), .d(_net_6555) );
na02f01  g5345 ( .o(n10079), .a(n12075), .b(n12071) );
oa12f01  g5346 ( .o(n12077), .a(n8213), .b(n6832), .c(n6829) );
ao22f01  g5347 ( .o(n12078), .a(n8211_1), .b(_net_6131), .c(n9200), .d(n10704) );
na02f01  g5348 ( .o(n12079), .a(n11913), .b(n11912) );
ao22f01  g5349 ( .o(n12080), .a(n12079), .b(n9207), .c(n10708), .d(n9205) );
na03f01  g5350 ( .o(n10084), .a(n12080), .b(n12078), .c(n12077) );
no02f01  g5351 ( .o(n12082), .a(n10436), .b(n7721) );
no02f01  g5352 ( .o(n12083), .a(n10439), .b(n7592) );
in01f01  g5353 ( .o(n12084), .a(_net_6183) );
no02f01  g5354 ( .o(n12085), .a(n9074_1), .b(n9071) );
oa22f01  g5355 ( .o(n12086), .a(n12085), .b(n7574), .c(n7590), .d(n12084) );
no03f01  g5356 ( .o(n12087), .a(n12086), .b(n12083), .c(n12082) );
in01f01  g5357 ( .o(n12088), .a(net_7162) );
in01f01  g5358 ( .o(n12089), .a(net_7130) );
oa22f01  g5359 ( .o(n12090), .a(n7740), .b(n12089), .c(n7739), .d(n12088) );
in01f01  g5360 ( .o(n12091), .a(net_7194) );
in01f01  g5361 ( .o(n12092), .a(net_7226) );
oa22f01  g5362 ( .o(n12093), .a(n7745), .b(n12092), .c(n7744), .d(n12091) );
no02f01  g5363 ( .o(n12094), .a(n12093), .b(n12090) );
na02f01  g5364 ( .o(n10089), .a(n12094), .b(n12087) );
in01f01  g5365 ( .o(n12096), .a(_net_7264) );
na02f01  g5366 ( .o(n12097), .a(n7437_1), .b(n6901) );
oa12f01  g5367 ( .o(n10094), .a(n12097), .b(n6901), .c(n12096) );
in01f01  g5368 ( .o(n12099), .a(_net_7479) );
na02f01  g5369 ( .o(n12100), .a(n7504), .b(n6869) );
oa12f01  g5370 ( .o(n10099), .a(n12100), .b(n6869), .c(n12099) );
ao22f01  g5371 ( .o(n12102), .a(n6736_1), .b(_net_7634), .c(n6734), .d(_net_7602) );
ao22f01  g5372 ( .o(n12103), .a(n6739), .b(_net_7666), .c(n6738), .d(_net_7570) );
na02f01  g5373 ( .o(n10116), .a(n12103), .b(n12102) );
in01f01  g5374 ( .o(n12105), .a(_net_7356) );
na02f01  g5375 ( .o(n12106), .a(n10089_1), .b(n7030) );
oa12f01  g5376 ( .o(n10128), .a(n12106), .b(n7030), .c(n12105) );
no02f01  g5377 ( .o(n12108), .a(n9766), .b(n7721) );
no02f01  g5378 ( .o(n12109), .a(n11480), .b(n7592) );
in01f01  g5379 ( .o(n12110), .a(_net_6176) );
oa22f01  g5380 ( .o(n12111), .a(n7935), .b(n7574), .c(n7590), .d(n12110) );
no03f01  g5381 ( .o(n12112), .a(n12111), .b(n12109), .c(n12108) );
in01f01  g5382 ( .o(n12113), .a(net_7123) );
in01f01  g5383 ( .o(n12114), .a(net_7155) );
oa22f01  g5384 ( .o(n12115), .a(n7740), .b(n12113), .c(n7739), .d(n12114) );
in01f01  g5385 ( .o(n12116), .a(net_7219) );
in01f01  g5386 ( .o(n12117), .a(net_7187) );
oa22f01  g5387 ( .o(n12118), .a(n7745), .b(n12116), .c(n7744), .d(n12117) );
no02f01  g5388 ( .o(n12119), .a(n12118), .b(n12115) );
na02f01  g5389 ( .o(n10137), .a(n12119), .b(n12112) );
na02f01  g5390 ( .o(n12121), .a(n7917), .b(n7575) );
oa12f01  g5391 ( .o(n10150), .a(n12121), .b(n7590), .c(n11532) );
bf01f01  g5392 ( .o(x124), .a(_net_5857) );
bf01f01  g5393 ( .o(x84), .a(_net_5852) );
bf01f01  g5394 ( .o(x131), .a(_net_5859) );
bf01f01  g5395 ( .o(x145), .a(x130657) );
bf01f01  g5396 ( .o(x63), .a(_net_5850) );
bf01f01  g5397 ( .o(x96), .a(_net_5853) );
bf01f01  g5398 ( .o(x106), .a(_net_5855) );
bf01f01  g5399 ( .o(x101), .a(_net_5854) );
bf01f01  g5400 ( .o(x114), .a(_net_5856) );
bf01f01  g5401 ( .o(x77), .a(_net_5851) );
bf01f01  g5402 ( .o(n276), .a(net_7807) );
bf01f01  g5403 ( .o(n286), .a(_net_6104) );
bf01f01  g5404 ( .o(n291), .a(net_6453) );
bf01f01  g5405 ( .o(n305), .a(_net_7820) );
bf01f01  g5406 ( .o(n310), .a(net_6704) );
bf01f01  g5407 ( .o(n324), .a(net_7802) );
bf01f01  g5408 ( .o(n334), .a(net_133) );
bf01f01  g5409 ( .o(n339), .a(_net_6168) );
bf01f01  g5410 ( .o(n344), .a(_net_6080) );
bf01f01  g5411 ( .o(n349), .a(net_6474) );
bf01f01  g5412 ( .o(n352), .a(x1542) );
bf01f01  g5413 ( .o(n357), .a(net_7114) );
bf01f01  g5414 ( .o(n361), .a(_net_7819) );
bf01f01  g5415 ( .o(n366), .a(net_6996) );
bf01f01  g5416 ( .o(n395), .a(_net_7820) );
bf01f01  g5417 ( .o(n405), .a(net_6395) );
bf01f01  g5418 ( .o(n410), .a(_net_6117) );
bf01f01  g5419 ( .o(n415), .a(_net_7795) );
bf01f01  g5420 ( .o(n424), .a(_net_7819) );
bf01f01  g5421 ( .o(n429), .a(_net_7806) );
bf01f01  g5422 ( .o(n434), .a(net_7713) );
bf01f01  g5423 ( .o(n438), .a(_net_7815) );
bf01f01  g5424 ( .o(n443), .a(net_7000) );
bf01f01  g5425 ( .o(n451), .a(x1527) );
bf01f01  g5426 ( .o(n455), .a(_net_7798) );
bf01f01  g5427 ( .o(n470), .a(net_7388) );
bf01f01  g5428 ( .o(n474), .a(net_6397) );
bf01f01  g5429 ( .o(n479), .a(_net_7818) );
bf01f01  g5430 ( .o(n484), .a(net_6870) );
bf01f01  g5431 ( .o(n488), .a(_net_7794) );
bf01f01  g5432 ( .o(n493), .a(_net_7822) );
bf01f01  g5433 ( .o(n498), .a(net_6059) );
bf01f01  g5434 ( .o(n503), .a(_net_6091) );
bf01f01  g5435 ( .o(n508), .a(_net_6112) );
bf01f01  g5436 ( .o(n556), .a(_net_7794) );
bf01f01  g5437 ( .o(n566), .a(_net_7808) );
bf01f01  g5438 ( .o(n571), .a(net_152) );
bf01f01  g5439 ( .o(n580), .a(x1587) );
bf01f01  g5440 ( .o(n585), .a(_net_6177) );
bf01f01  g5441 ( .o(n590), .a(net_6400) );
bf01f01  g5442 ( .o(n610), .a(_net_7800) );
bf01f01  g5443 ( .o(n625), .a(net_7246) );
bf01f01  g5444 ( .o(n664), .a(net_6383) );
bf01f01  g5445 ( .o(n669), .a(net_6440) );
bf01f01  g5446 ( .o(n678), .a(_net_7823) );
bf01f01  g5447 ( .o(n683), .a(_net_7796) );
bf01f01  g5448 ( .o(n703), .a(_net_6127) );
bf01f01  g5449 ( .o(n722), .a(net_6396) );
bf01f01  g5450 ( .o(n741), .a(net_147) );
bf01f01  g5451 ( .o(n751), .a(_net_5976) );
bf01f01  g5452 ( .o(n761), .a(net_6468) );
bf01f01  g5453 ( .o(n774), .a(x806) );
bf01f01  g5454 ( .o(n779), .a(net_6385) );
bf01f01  g5455 ( .o(n783), .a(net_7802) );
bf01f01  g5456 ( .o(n798), .a(net_7134) );
bf01f01  g5457 ( .o(n802), .a(net_7133) );
bf01f01  g5458 ( .o(n811), .a(net_6399) );
bf01f01  g5459 ( .o(n815), .a(_net_6084) );
bf01f01  g5460 ( .o(n830), .a(net_7396) );
bf01f01  g5461 ( .o(n839), .a(_net_7818) );
bf01f01  g5462 ( .o(n844), .a(net_6381) );
bf01f01  g5463 ( .o(n854), .a(net_7390) );
bf01f01  g5464 ( .o(n857), .a(_net_7794) );
bf01f01  g5465 ( .o(n867), .a(net_6711) );
bf01f01  g5466 ( .o(n870), .a(_net_7818) );
bf01f01  g5467 ( .o(n880), .a(_net_7816) );
bf01f01  g5468 ( .o(n890), .a(net_6616) );
bf01f01  g5469 ( .o(n894), .a(net_6382) );
bf01f01  g5470 ( .o(n899), .a(net_6739) );
bf01f01  g5471 ( .o(n907), .a(_net_7800) );
bf01f01  g5472 ( .o(n911), .a(_net_7806) );
bf01f01  g5473 ( .o(n916), .a(net_6746) );
bf01f01  g5474 ( .o(n920), .a(_net_6160) );
bf01f01  g5475 ( .o(n935), .a(net_7799) );
bf01f01  g5476 ( .o(n940), .a(net_6979) );
bf01f01  g5477 ( .o(n948), .a(x1467) );
bf01f01  g5478 ( .o(n953), .a(net_6989) );
bf01f01  g5479 ( .o(n956), .a(_net_7823) );
bf01f01  g5480 ( .o(n976), .a(_net_7813) );
bf01f01  g5481 ( .o(n981), .a(net_6999) );
bf01f01  g5482 ( .o(n1000), .a(net_388) );
bf01f01  g5483 ( .o(n1005), .a(net_6391) );
bf01f01  g5484 ( .o(n1020), .a(net_6998) );
bf01f01  g5485 ( .o(n1053), .a(net_6386) );
bf01f01  g5486 ( .o(n1062), .a(_net_7812) );
bf01f01  g5487 ( .o(n1077), .a(net_7004) );
bf01f01  g5488 ( .o(n1081), .a(net_7010) );
bf01f01  g5489 ( .o(n1085), .a(net_6461) );
bf01f01  g5490 ( .o(n1089), .a(net_6832) );
bf01f01  g5491 ( .o(n1093), .a(net_6977) );
bf01f01  g5492 ( .o(n1097), .a(_net_7801) );
bf01f01  g5493 ( .o(n1102), .a(net_6856) );
bf01f01  g5494 ( .o(n1111), .a(_net_6183) );
bf01f01  g5495 ( .o(n1121), .a(net_6847) );
bf01f01  g5496 ( .o(n1130), .a(_net_7809) );
bf01f01  g5497 ( .o(n1140), .a(net_6986) );
bf01f01  g5498 ( .o(n1144), .a(_net_6099) );
bf01f01  g5499 ( .o(n1148), .a(_net_7815) );
bf01f01  g5500 ( .o(n1158), .a(_net_6066) );
bf01f01  g5501 ( .o(n1168), .a(net_6398) );
bf01f01  g5502 ( .o(n1183), .a(net_144) );
bf01f01  g5503 ( .o(n1187), .a(net_6400) );
bf01f01  g5504 ( .o(n1191), .a(_net_7823) );
bf01f01  g5505 ( .o(n1195), .a(_net_7822) );
bf01f01  g5506 ( .o(n1200), .a(_net_6064) );
bf01f01  g5507 ( .o(n1205), .a(_net_7814) );
bf01f01  g5508 ( .o(n1210), .a(net_6845) );
bf01f01  g5509 ( .o(n1224), .a(net_6608) );
bf01f01  g5510 ( .o(n1232), .a(_net_7795) );
no02f01  g5511 ( .o(n1236), .a(n6966), .b(n7599_1) );
bf01f01  g5512 ( .o(n1240), .a(_net_7820) );
bf01f01  g5513 ( .o(n1244), .a(net_6395) );
bf01f01  g5514 ( .o(n1248), .a(_net_7794) );
bf01f01  g5515 ( .o(n1258), .a(net_7019) );
bf01f01  g5516 ( .o(n1262), .a(_net_6158) );
bf01f01  g5517 ( .o(n1287), .a(net_7119) );
bf01f01  g5518 ( .o(n1291), .a(net_6574) );
bf01f01  g5519 ( .o(n1300), .a(_net_7803) );
bf01f01  g5520 ( .o(n1305), .a(net_7395) );
bf01f01  g5521 ( .o(n1318), .a(_net_7812) );
bf01f01  g5522 ( .o(n1322), .a(_net_7798) );
bf01f01  g5523 ( .o(n1326), .a(_net_7820) );
bf01f01  g5524 ( .o(n1331), .a(net_6859) );
bf01f01  g5525 ( .o(n1355), .a(net_6877) );
bf01f01  g5526 ( .o(n1359), .a(net_7234) );
bf01f01  g5527 ( .o(n1378), .a(_net_5960) );
bf01f01  g5528 ( .o(n1383), .a(net_6694) );
bf01f01  g5529 ( .o(n1386), .a(net_6400) );
bf01f01  g5530 ( .o(n1400), .a(_net_7794) );
bf01f01  g5531 ( .o(n1414), .a(_net_7815) );
bf01f01  g5532 ( .o(n1423), .a(_net_7809) );
bf01f01  g5533 ( .o(n1438), .a(net_6745) );
bf01f01  g5534 ( .o(n1446), .a(_net_7813) );
bf01f01  g5535 ( .o(n1455), .a(_net_7803) );
bf01f01  g5536 ( .o(n1460), .a(_net_6132) );
bf01f01  g5537 ( .o(n1465), .a(_net_7821) );
bf01f01  g5538 ( .o(n1469), .a(net_6392) );
bf01f01  g5539 ( .o(n1474), .a(net_6612) );
bf01f01  g5540 ( .o(n1478), .a(_net_6106) );
bf01f01  g5541 ( .o(n1482), .a(x1417) );
bf01f01  g5542 ( .o(n1491), .a(_net_7803) );
bf01f01  g5543 ( .o(n1506), .a(net_7550) );
bf01f01  g5544 ( .o(n1510), .a(_net_7824) );
bf01f01  g5545 ( .o(n1515), .a(net_6619) );
bf01f01  g5546 ( .o(n1524), .a(net_7106) );
bf01f01  g5547 ( .o(n1528), .a(_net_6179) );
bf01f01  g5548 ( .o(n1538), .a(net_7247) );
bf01f01  g5549 ( .o(n1551), .a(net_7146) );
bf01f01  g5550 ( .o(n1560), .a(net_7126) );
bf01f01  g5551 ( .o(n1564), .a(net_6482) );
bf01f01  g5552 ( .o(n1568), .a(net_6888) );
bf01f01  g5553 ( .o(n1577), .a(net_6388) );
bf01f01  g5554 ( .o(n1587), .a(net_6584) );
bf01f01  g5555 ( .o(n1591), .a(net_6387) );
bf01f01  g5556 ( .o(n1596), .a(net_6732) );
bf01f01  g5557 ( .o(n1615), .a(_net_7814) );
bf01f01  g5558 ( .o(n1619), .a(_net_7796) );
bf01f01  g5559 ( .o(n1629), .a(_net_7810) );
bf01f01  g5560 ( .o(n1649), .a(net_7124) );
bf01f01  g5561 ( .o(n1653), .a(net_135) );
bf01f01  g5562 ( .o(n1663), .a(net_6061) );
bf01f01  g5563 ( .o(n1668), .a(_net_5980) );
bf01f01  g5564 ( .o(n1673), .a(net_6723) );
bf01f01  g5565 ( .o(n1681), .a(_net_7824) );
bf01f01  g5566 ( .o(n1686), .a(_net_7817) );
bf01f01  g5567 ( .o(n1691), .a(_net_7805) );
bf01f01  g5568 ( .o(n1701), .a(net_6432) );
bf01f01  g5569 ( .o(n1704), .a(_net_7805) );
bf01f01  g5570 ( .o(n1709), .a(_net_7800) );
bf01f01  g5571 ( .o(n1718), .a(_net_7803) );
bf01f01  g5572 ( .o(n1722), .a(_net_7818) );
bf01f01  g5573 ( .o(n1732), .a(_net_7809) );
bf01f01  g5574 ( .o(n1756), .a(_net_7796) );
bf01f01  g5575 ( .o(n1761), .a(net_6570) );
bf01f01  g5576 ( .o(n1765), .a(_net_7821) );
bf01f01  g5577 ( .o(n1775), .a(net_6602) );
bf01f01  g5578 ( .o(n1779), .a(net_7551) );
bf01f01  g5579 ( .o(n1782), .a(_net_7800) );
bf01f01  g5580 ( .o(n1797), .a(_net_6120) );
bf01f01  g5581 ( .o(n1817), .a(_net_6175) );
bf01f01  g5582 ( .o(n1822), .a(_net_6093) );
bf01f01  g5583 ( .o(n1827), .a(_net_6072) );
bf01f01  g5584 ( .o(n1836), .a(x1432) );
bf01f01  g5585 ( .o(n1855), .a(x1382) );
bf01f01  g5586 ( .o(n1865), .a(net_6699) );
bf01f01  g5587 ( .o(n1874), .a(net_6599) );
bf01f01  g5588 ( .o(n1903), .a(_net_6082) );
bf01f01  g5589 ( .o(n1913), .a(_net_7816) );
bf01f01  g5590 ( .o(n1918), .a(net_7116) );
bf01f01  g5591 ( .o(n1932), .a(net_6995) );
bf01f01  g5592 ( .o(n1941), .a(net_6433) );
bf01f01  g5593 ( .o(n1954), .a(_net_7817) );
bf01f01  g5594 ( .o(n1964), .a(_net_6150) );
bf01f01  g5595 ( .o(n1973), .a(_net_7803) );
bf01f01  g5596 ( .o(n1978), .a(_net_7804) );
bf01f01  g5597 ( .o(n1983), .a(_net_6098) );
bf01f01  g5598 ( .o(n1998), .a(net_6737) );
bf01f01  g5599 ( .o(n2002), .a(_net_6107) );
bf01f01  g5600 ( .o(n2007), .a(_net_7815) );
bf01f01  g5601 ( .o(n2011), .a(_net_7818) );
bf01f01  g5602 ( .o(n2031), .a(_net_6122) );
bf01f01  g5603 ( .o(n2036), .a(net_6394) );
bf01f01  g5604 ( .o(n2051), .a(net_7391) );
bf01f01  g5605 ( .o(n2074), .a(net_7799) );
bf01f01  g5606 ( .o(n2079), .a(_net_5968) );
bf01f01  g5607 ( .o(n2088), .a(_net_7796) );
bf01f01  g5608 ( .o(n2093), .a(_net_7793) );
bf01f01  g5609 ( .o(n2098), .a(net_6709) );
bf01f01  g5610 ( .o(n2102), .a(net_6741) );
bf01f01  g5611 ( .o(n2106), .a(net_6056) );
bf01f01  g5612 ( .o(n2111), .a(net_7003) );
bf01f01  g5613 ( .o(n2115), .a(net_6452) );
bf01f01  g5614 ( .o(n2119), .a(net_6603) );
bf01f01  g5615 ( .o(n2122), .a(_net_7809) );
bf01f01  g5616 ( .o(n2127), .a(_net_6114) );
bf01f01  g5617 ( .o(n2132), .a(net_7147) );
bf01f01  g5618 ( .o(n2136), .a(net_6730) );
bf01f01  g5619 ( .o(n2144), .a(_net_7809) );
bf01f01  g5620 ( .o(n2149), .a(net_7144) );
no02f01  g5621 ( .o(n2152), .a(n6966), .b(n7250) );
bf01f01  g5622 ( .o(n2157), .a(_net_6140) );
bf01f01  g5623 ( .o(n2186), .a(net_6443) );
bf01f01  g5624 ( .o(n2189), .a(_net_7813) );
bf01f01  g5625 ( .o(n2203), .a(_net_7796) );
bf01f01  g5626 ( .o(n2218), .a(net_6456) );
no02f01  g5627 ( .o(n2260), .a(n6966), .b(n7351) );
bf01f01  g5628 ( .o(n2284), .a(net_6397) );
bf01f01  g5629 ( .o(n2288), .a(_net_7805) );
bf01f01  g5630 ( .o(n2293), .a(_net_6170) );
bf01f01  g5631 ( .o(n2307), .a(_net_7824) );
bf01f01  g5632 ( .o(n2316), .a(_net_7800) );
bf01f01  g5633 ( .o(n2321), .a(net_7159) );
bf01f01  g5634 ( .o(n2324), .a(net_6398) );
bf01f01  g5635 ( .o(n2338), .a(_net_7820) );
bf01f01  g5636 ( .o(n2342), .a(_net_7806) );
bf01f01  g5637 ( .o(n2347), .a(net_6849) );
bf01f01  g5638 ( .o(n2350), .a(net_142) );
bf01f01  g5639 ( .o(n2355), .a(_net_6101) );
bf01f01  g5640 ( .o(n2360), .a(_net_7812) );
bf01f01  g5641 ( .o(n2370), .a(net_6593) );
bf01f01  g5642 ( .o(n2373), .a(net_6397) );
no02f01  g5643 ( .o(n2381), .a(n6867_1), .b(n7978) );
bf01f01  g5644 ( .o(n2391), .a(net_6576) );
bf01f01  g5645 ( .o(n2399), .a(_net_7793) );
bf01f01  g5646 ( .o(n2417), .a(_net_7818) );
bf01f01  g5647 ( .o(n2422), .a(net_7016) );
bf01f01  g5648 ( .o(n2426), .a(net_6833) );
bf01f01  g5649 ( .o(n2440), .a(net_7240) );
bf01f01  g5650 ( .o(n2448), .a(net_6392) );
bf01f01  g5651 ( .o(n2452), .a(_net_7824) );
bf01f01  g5652 ( .o(n2462), .a(net_6426) );
bf01f01  g5653 ( .o(n2465), .a(_net_7818) );
bf01f01  g5654 ( .o(n2474), .a(_net_7810) );
bf01f01  g5655 ( .o(n2488), .a(net_7799) );
bf01f01  g5656 ( .o(n2493), .a(net_6435) );
bf01f01  g5657 ( .o(n2496), .a(_net_7805) );
no02f01  g5658 ( .o(n2500), .a(n6966), .b(n7351) );
bf01f01  g5659 ( .o(n2519), .a(_net_7795) );
bf01f01  g5660 ( .o(n2539), .a(_net_7797) );
bf01f01  g5661 ( .o(n2543), .a(net_7807) );
no02f01  g5662 ( .o(n2547), .a(n6899_1), .b(n7069) );
bf01f01  g5663 ( .o(n2556), .a(_net_7819) );
bf01f01  g5664 ( .o(n2561), .a(net_6390) );
bf01f01  g5665 ( .o(n2570), .a(_net_7798) );
bf01f01  g5666 ( .o(n2594), .a(net_6390) );
bf01f01  g5667 ( .o(n2597), .a(_net_7797) );
bf01f01  g5668 ( .o(n2601), .a(_net_7822) );
bf01f01  g5669 ( .o(n2605), .a(_net_7818) );
bf01f01  g5670 ( .o(n2610), .a(_net_6181) );
bf01f01  g5671 ( .o(n2615), .a(net_6967) );
bf01f01  g5672 ( .o(n2618), .a(_net_7793) );
bf01f01  g5673 ( .o(n2622), .a(_net_7822) );
bf01f01  g5674 ( .o(n2627), .a(_net_6126) );
bf01f01  g5675 ( .o(n2642), .a(_net_6145) );
bf01f01  g5676 ( .o(n2647), .a(net_6588) );
bf01f01  g5677 ( .o(n2656), .a(net_6606) );
bf01f01  g5678 ( .o(n2660), .a(net_149) );
bf01f01  g5679 ( .o(n2670), .a(_net_6134) );
bf01f01  g5680 ( .o(n2675), .a(net_6890) );
bf01f01  g5681 ( .o(n2679), .a(net_6964) );
bf01f01  g5682 ( .o(n2682), .a(_net_7822) );
bf01f01  g5683 ( .o(n2692), .a(net_7393) );
bf01f01  g5684 ( .o(n2701), .a(net_6981) );
bf01f01  g5685 ( .o(n2705), .a(net_6434) );
bf01f01  g5686 ( .o(n2709), .a(net_6969) );
bf01f01  g5687 ( .o(n2727), .a(net_6381) );
bf01f01  g5688 ( .o(n2737), .a(net_7708) );
bf01f01  g5689 ( .o(n2741), .a(net_6586) );
bf01f01  g5690 ( .o(n2745), .a(net_6725) );
bf01f01  g5691 ( .o(n2748), .a(_net_7823) );
bf01f01  g5692 ( .o(n2762), .a(_net_7823) );
bf01f01  g5693 ( .o(n2767), .a(net_7108) );
bf01f01  g5694 ( .o(n2781), .a(net_6880) );
no02f01  g5695 ( .o(n2784), .a(n6899_1), .b(n7509_1) );
bf01f01  g5696 ( .o(n2788), .a(_net_7801) );
bf01f01  g5697 ( .o(n2792), .a(net_7802) );
bf01f01  g5698 ( .o(n2801), .a(_net_7797) );
bf01f01  g5699 ( .o(n2805), .a(x1374) );
bf01f01  g5700 ( .o(n2814), .a(_net_7812) );
bf01f01  g5701 ( .o(n2819), .a(net_6579) );
bf01f01  g5702 ( .o(n2823), .a(net_7024) );
bf01f01  g5703 ( .o(n2827), .a(net_7153) );
bf01f01  g5704 ( .o(n2840), .a(_net_7801) );
bf01f01  g5705 ( .o(n2860), .a(net_7236) );
bf01f01  g5706 ( .o(n2864), .a(_net_6070) );
bf01f01  g5707 ( .o(n2869), .a(net_6478) );
bf01f01  g5708 ( .o(n2873), .a(net_6578) );
bf01f01  g5709 ( .o(n2877), .a(_net_6068) );
bf01f01  g5710 ( .o(n2882), .a(net_7547) );
bf01f01  g5711 ( .o(n2885), .a(_net_7816) );
bf01f01  g5712 ( .o(n2895), .a(_net_5972) );
no02f01  g5713 ( .o(n2904), .a(n6867_1), .b(n6974_1) );
bf01f01  g5714 ( .o(n2908), .a(_net_7814) );
bf01f01  g5715 ( .o(n2922), .a(net_7022) );
bf01f01  g5716 ( .o(n2926), .a(net_6755) );
bf01f01  g5717 ( .o(n2935), .a(net_390) );
bf01f01  g5718 ( .o(n2939), .a(_net_7816) );
bf01f01  g5719 ( .o(n2944), .a(net_7158) );
bf01f01  g5720 ( .o(n2963), .a(_net_6142) );
bf01f01  g5721 ( .o(n2967), .a(net_6392) );
bf01f01  g5722 ( .o(n2972), .a(net_7007) );
bf01f01  g5723 ( .o(n2996), .a(net_6438) );
bf01f01  g5724 ( .o(n3030), .a(net_7105) );
bf01f01  g5725 ( .o(n3033), .a(_net_7806) );
bf01f01  g5726 ( .o(n3037), .a(_net_7809) );
bf01f01  g5727 ( .o(n3052), .a(net_7136) );
bf01f01  g5728 ( .o(n3061), .a(net_7121) );
bf01f01  g5729 ( .o(n3069), .a(_net_7806) );
bf01f01  g5730 ( .o(n3074), .a(net_6717) );
bf01f01  g5731 ( .o(n3082), .a(net_7799) );
bf01f01  g5732 ( .o(n3102), .a(net_6706) );
bf01f01  g5733 ( .o(n3105), .a(net_6396) );
bf01f01  g5734 ( .o(n3110), .a(net_6473) );
bf01f01  g5735 ( .o(n3114), .a(net_6743) );
bf01f01  g5736 ( .o(n3117), .a(_net_7824) );
no02f01  g5737 ( .o(n3121), .a(n6966), .b(n7599_1) );
bf01f01  g5738 ( .o(n3126), .a(net_7387) );
bf01f01  g5739 ( .o(n3134), .a(_net_7809) );
bf01f01  g5740 ( .o(n3143), .a(_net_7819) );
bf01f01  g5741 ( .o(n3152), .a(_net_7805) );
bf01f01  g5742 ( .o(n3162), .a(net_6751) );
in01f01  g5743 ( .o(n3165), .a(n7343) );
bf01f01  g5744 ( .o(n3174), .a(_net_7815) );
bf01f01  g5745 ( .o(n3178), .a(net_6450) );
bf01f01  g5746 ( .o(n3186), .a(_net_7798) );
bf01f01  g5747 ( .o(n3190), .a(net_6861) );
bf01f01  g5748 ( .o(n3199), .a(net_7536) );
bf01f01  g5749 ( .o(n3207), .a(_net_7793) );
bf01f01  g5750 ( .o(n3226), .a(net_139) );
bf01f01  g5751 ( .o(n3235), .a(x1443) );
bf01f01  g5752 ( .o(n3244), .a(_net_7822) );
bf01f01  g5753 ( .o(n3249), .a(_net_6083) );
bf01f01  g5754 ( .o(n3258), .a(x1366) );
bf01f01  g5755 ( .o(n3272), .a(net_7799) );
no02f01  g5756 ( .o(n3276), .a(n6867_1), .b(n8170_1) );
bf01f01  g5757 ( .o(n3280), .a(_net_7795) );
bf01f01  g5758 ( .o(n3290), .a(net_7710) );
bf01f01  g5759 ( .o(n3299), .a(_net_7793) );
bf01f01  g5760 ( .o(n3303), .a(_net_7809) );
bf01f01  g5761 ( .o(n3318), .a(net_6883) );
no02f01  g5762 ( .o(n3325), .a(n6899_1), .b(n7173) );
bf01f01  g5763 ( .o(n3330), .a(net_6868) );
no02f01  g5764 ( .o(n3333), .a(n6899_1), .b(n7254) );
bf01f01  g5765 ( .o(n3343), .a(_net_6063) );
bf01f01  g5766 ( .o(n3348), .a(net_7140) );
bf01f01  g5767 ( .o(n3361), .a(_net_6071) );
bf01f01  g5768 ( .o(n3365), .a(_net_7821) );
no02f01  g5769 ( .o(n3374), .a(n6867_1), .b(n7650) );
bf01f01  g5770 ( .o(n3379), .a(net_6698) );
bf01f01  g5771 ( .o(n3383), .a(net_6485) );
bf01f01  g5772 ( .o(n3386), .a(net_7807) );
bf01f01  g5773 ( .o(n3390), .a(x1424) );
bf01f01  g5774 ( .o(n3404), .a(net_6386) );
bf01f01  g5775 ( .o(n3408), .a(_net_7820) );
bf01f01  g5776 ( .o(n3413), .a(net_148) );
bf01f01  g5777 ( .o(n3418), .a(net_7248) );
in01f01  g5778 ( .o(n3431), .a(n7343) );
bf01f01  g5779 ( .o(n3436), .a(net_7120) );
bf01f01  g5780 ( .o(n3445), .a(net_6389) );
bf01f01  g5781 ( .o(n3450), .a(_net_6173) );
bf01f01  g5782 ( .o(n3469), .a(_net_7811) );
bf01f01  g5783 ( .o(n3479), .a(_net_6136) );
bf01f01  g5784 ( .o(n3494), .a(net_7241) );
bf01f01  g5785 ( .o(n3497), .a(_net_7803) );
bf01f01  g5786 ( .o(n3502), .a(_net_263) );
bf01f01  g5787 ( .o(n3511), .a(_net_7793) );
bf01f01  g5788 ( .o(n3520), .a(_net_7800) );
bf01f01  g5789 ( .o(n3524), .a(net_150) );
bf01f01  g5790 ( .o(n3528), .a(_net_7815) );
bf01f01  g5791 ( .o(n3532), .a(net_6384) );
bf01f01  g5792 ( .o(n3537), .a(_net_6078) );
bf01f01  g5793 ( .o(n3542), .a(net_6885) );
bf01f01  g5794 ( .o(n3555), .a(net_6385) );
bf01f01  g5795 ( .o(n3559), .a(_net_7810) );
bf01f01  g5796 ( .o(n3564), .a(net_6873) );
no02f01  g5797 ( .o(n3567), .a(n6966), .b(n8514) );
bf01f01  g5798 ( .o(n3587), .a(net_6476) );
bf01f01  g5799 ( .o(n3590), .a(_net_7803) );
bf01f01  g5800 ( .o(n3600), .a(net_6583) );
bf01f01  g5801 ( .o(n3618), .a(_net_7812) );
bf01f01  g5802 ( .o(n3623), .a(_net_6124) );
in01f01  g5803 ( .o(n3642), .a(n7343) );
bf01f01  g5804 ( .o(n3651), .a(net_7157) );
bf01f01  g5805 ( .o(n3655), .a(net_6591) );
bf01f01  g5806 ( .o(n3658), .a(net_6394) );
no02f01  g5807 ( .o(n3661), .a(n6867_1), .b(n8173) );
bf01f01  g5808 ( .o(n3670), .a(_net_7794) );
bf01f01  g5809 ( .o(n3679), .a(_net_7801) );
bf01f01  g5810 ( .o(n3689), .a(net_6605) );
bf01f01  g5811 ( .o(n3703), .a(net_6976) );
bf01f01  g5812 ( .o(n3707), .a(net_6721) );
bf01f01  g5813 ( .o(n3716), .a(net_6486) );
bf01f01  g5814 ( .o(n3720), .a(_net_6092) );
bf01f01  g5815 ( .o(n3725), .a(net_6881) );
bf01f01  g5816 ( .o(n3729), .a(_net_7813) );
bf01f01  g5817 ( .o(n3733), .a(x1550) );
bf01f01  g5818 ( .o(n3747), .a(_net_6129) );
bf01f01  g5819 ( .o(n3752), .a(_net_6069) );
bf01f01  g5820 ( .o(n3756), .a(net_6391) );
bf01f01  g5821 ( .o(n3761), .a(net_6442) );
bf01f01  g5822 ( .o(n3770), .a(net_6991) );
bf01f01  g5823 ( .o(n3773), .a(_net_7796) );
bf01f01  g5824 ( .o(n3777), .a(_net_7798) );
bf01f01  g5825 ( .o(n3791), .a(_net_7804) );
bf01f01  g5826 ( .o(n3801), .a(net_7149) );
bf01f01  g5827 ( .o(n3805), .a(net_7714) );
bf01f01  g5828 ( .o(n3809), .a(net_6429) );
bf01f01  g5829 ( .o(n3817), .a(net_6394) );
bf01f01  g5830 ( .o(n3822), .a(_net_6076) );
bf01f01  g5831 ( .o(n3831), .a(net_7802) );
bf01f01  g5832 ( .o(n3851), .a(net_6829) );
bf01f01  g5833 ( .o(n3855), .a(net_6595) );
bf01f01  g5834 ( .o(n3864), .a(net_6850) );
bf01f01  g5835 ( .o(n3867), .a(_net_7806) );
bf01f01  g5836 ( .o(n3881), .a(net_7799) );
bf01f01  g5837 ( .o(n3896), .a(net_6855) );
bf01f01  g5838 ( .o(n3899), .a(net_7799) );
bf01f01  g5839 ( .o(n3904), .a(net_7239) );
bf01f01  g5840 ( .o(n3917), .a(_net_7814) );
bf01f01  g5841 ( .o(n3936), .a(_net_7823) );
bf01f01  g5842 ( .o(n3945), .a(net_6384) );
bf01f01  g5843 ( .o(n3949), .a(_net_7822) );
bf01f01  g5844 ( .o(n3953), .a(_net_7815) );
bf01f01  g5845 ( .o(n3957), .a(net_6387) );
bf01f01  g5846 ( .o(n3962), .a(_net_6176) );
bf01f01  g5847 ( .o(n3972), .a(net_7537) );
bf01f01  g5848 ( .o(n3985), .a(_net_7815) );
bf01f01  g5849 ( .o(n3989), .a(net_6392) );
bf01f01  g5850 ( .o(n3993), .a(_net_7795) );
bf01f01  g5851 ( .o(n4002), .a(_net_7817) );
bf01f01  g5852 ( .o(n4007), .a(net_6852) );
bf01f01  g5853 ( .o(n4011), .a(_net_6103) );
bf01f01  g5854 ( .o(n4020), .a(_net_7813) );
bf01f01  g5855 ( .o(n4024), .a(_net_7804) );
bf01f01  g5856 ( .o(n4033), .a(_net_7821) );
bf01f01  g5857 ( .o(n4037), .a(_net_7793) );
bf01f01  g5858 ( .o(n4046), .a(net_6390) );
bf01f01  g5859 ( .o(n4051), .a(net_6613) );
bf01f01  g5860 ( .o(n4055), .a(net_7711) );
bf01f01  g5861 ( .o(n4059), .a(net_7013) );
bf01f01  g5862 ( .o(n4068), .a(net_6444) );
bf01f01  g5863 ( .o(n4071), .a(_net_7814) );
bf01f01  g5864 ( .o(n4075), .a(net_6399) );
no02f01  g5865 ( .o(n4079), .a(n6966), .b(n7188) );
bf01f01  g5866 ( .o(n4098), .a(_net_7798) );
bf01f01  g5867 ( .o(n4102), .a(_net_7813) );
bf01f01  g5868 ( .o(n4112), .a(net_6867) );
bf01f01  g5869 ( .o(n4131), .a(net_7400) );
bf01f01  g5870 ( .o(n4145), .a(net_6592) );
bf01f01  g5871 ( .o(n4148), .a(_net_7793) );
bf01f01  g5872 ( .o(n4153), .a(net_145) );
bf01f01  g5873 ( .o(n4158), .a(net_6714) );
bf01f01  g5874 ( .o(n4161), .a(net_6382) );
bf01f01  g5875 ( .o(n4176), .a(_net_6087) );
bf01f01  g5876 ( .o(n4191), .a(net_7123) );
bf01f01  g5877 ( .o(n4194), .a(_net_7822) );
bf01f01  g5878 ( .o(n4199), .a(net_6447) );
bf01f01  g5879 ( .o(n4207), .a(_net_7808) );
bf01f01  g5880 ( .o(n4221), .a(_net_7814) );
bf01f01  g5881 ( .o(n4231), .a(net_5858) );
bf01f01  g5882 ( .o(n4235), .a(_net_7813) );
bf01f01  g5883 ( .o(n4245), .a(net_7398) );
bf01f01  g5884 ( .o(n4253), .a(net_6391) );
bf01f01  g5885 ( .o(n4258), .a(_net_7816) );
bf01f01  g5886 ( .o(n4267), .a(_net_7796) );
bf01f01  g5887 ( .o(n4271), .a(net_6387) );
bf01f01  g5888 ( .o(n4280), .a(_net_7794) );
bf01f01  g5889 ( .o(n4284), .a(x1459) );
bf01f01  g5890 ( .o(n4309), .a(net_6753) );
bf01f01  g5891 ( .o(n4318), .a(net_6471) );
bf01f01  g5892 ( .o(n4326), .a(net_6387) );
bf01f01  g5893 ( .o(n4330), .a(net_6978) );
no02f01  g5894 ( .o(n4333), .a(n6966), .b(n8899_1) );
bf01f01  g5895 ( .o(n4338), .a(_net_7808) );
bf01f01  g5896 ( .o(n4343), .a(_net_7791) );
no02f01  g5897 ( .o(n4352), .a(n6966), .b(n7891) );
bf01f01  g5898 ( .o(n4362), .a(net_6863) );
bf01f01  g5899 ( .o(n4365), .a(_net_7797) );
bf01f01  g5900 ( .o(n4370), .a(_net_7811) );
bf01f01  g5901 ( .o(n4374), .a(_net_7818) );
bf01f01  g5902 ( .o(n4384), .a(net_6974) );
bf01f01  g5903 ( .o(n4388), .a(net_6431) );
bf01f01  g5904 ( .o(n4397), .a(net_6564) );
bf01f01  g5905 ( .o(n4401), .a(net_7162) );
bf01f01  g5906 ( .o(n4410), .a(net_7111) );
bf01f01  g5907 ( .o(n4419), .a(_net_6151) );
no02f01  g5908 ( .o(n4428), .a(n6899_1), .b(n7507) );
bf01f01  g5909 ( .o(n4448), .a(net_6886) );
no02f01  g5910 ( .o(n4451), .a(n6899_1), .b(n7173) );
in01f01  g5911 ( .o(n4459), .a(n7343) );
bf01f01  g5912 ( .o(n4469), .a(_net_6147) );
bf01f01  g5913 ( .o(n4473), .a(_net_7797) );
bf01f01  g5914 ( .o(n4478), .a(net_6448) );
bf01f01  g5915 ( .o(n4487), .a(net_7129) );
bf01f01  g5916 ( .o(n4496), .a(net_386) );
bf01f01  g5917 ( .o(n4505), .a(_net_7808) );
bf01f01  g5918 ( .o(n4524), .a(_net_7801) );
bf01f01  g5919 ( .o(n4548), .a(_net_7794) );
bf01f01  g5920 ( .o(n4558), .a(_net_7809) );
bf01f01  g5921 ( .o(n4562), .a(_net_7796) );
bf01f01  g5922 ( .o(n4567), .a(net_131) );
bf01f01  g5923 ( .o(n4577), .a(_net_6109) );
bf01f01  g5924 ( .o(n4581), .a(_net_7812) );
bf01f01  g5925 ( .o(n4600), .a(_net_7801) );
bf01f01  g5926 ( .o(n4604), .a(_net_7805) );
bf01f01  g5927 ( .o(n4613), .a(_net_7811) );
bf01f01  g5928 ( .o(n4617), .a(net_7807) );
bf01f01  g5929 ( .o(n4622), .a(_net_6097) );
bf01f01  g5930 ( .o(n4631), .a(_net_7821) );
bf01f01  g5931 ( .o(n4651), .a(_net_6171) );
bf01f01  g5932 ( .o(n4660), .a(_net_7795) );
bf01f01  g5933 ( .o(n4665), .a(net_6736) );
bf01f01  g5934 ( .o(n4669), .a(net_6581) );
bf01f01  g5935 ( .o(n4681), .a(x1564) );
bf01f01  g5936 ( .o(n4686), .a(net_6393) );
no02f01  g5937 ( .o(n4690), .a(n6899_1), .b(n7560) );
no02f01  g5938 ( .o(n4694), .a(n6867_1), .b(n6974_1) );
bf01f01  g5939 ( .o(n4699), .a(net_6993) );
bf01f01  g5940 ( .o(n4713), .a(net_7142) );
bf01f01  g5941 ( .o(n4717), .a(_net_7817) );
bf01f01  g5942 ( .o(n4722), .a(_net_6095) );
bf01f01  g5943 ( .o(n4742), .a(net_6735) );
bf01f01  g5944 ( .o(n4745), .a(net_7807) );
bf01f01  g5945 ( .o(n4750), .a(_net_6138) );
bf01f01  g5946 ( .o(n4755), .a(_net_6153) );
bf01f01  g5947 ( .o(n4765), .a(net_137) );
no02f01  g5948 ( .o(n4769), .a(n6867_1), .b(n7203_1) );
bf01f01  g5949 ( .o(n4774), .a(net_7545) );
bf01f01  g5950 ( .o(n4778), .a(net_6449) );
bf01f01  g5951 ( .o(n4782), .a(_net_6156) );
bf01f01  g5952 ( .o(n4791), .a(net_7799) );
bf01f01  g5953 ( .o(n4795), .a(_net_7803) );
bf01f01  g5954 ( .o(n4805), .a(net_7014) );
bf01f01  g5955 ( .o(n4814), .a(net_7128) );
no02f01  g5956 ( .o(n4822), .a(n6899_1), .b(n8826_1) );
bf01f01  g5957 ( .o(n4827), .a(net_6567) );
bf01f01  g5958 ( .o(n4834), .a(_net_7820) );
bf01f01  g5959 ( .o(n4838), .a(_net_7814) );
bf01f01  g5960 ( .o(n4848), .a(_net_6074) );
bf01f01  g5961 ( .o(n4853), .a(net_6875) );
bf01f01  g5962 ( .o(n4862), .a(_net_6402) );
bf01f01  g5963 ( .o(n4867), .a(_net_7819) );
bf01f01  g5964 ( .o(n4881), .a(net_6384) );
bf01f01  g5965 ( .o(n4890), .a(_net_7801) );
bf01f01  g5966 ( .o(n4895), .a(net_7154) );
bf01f01  g5967 ( .o(n4899), .a(_net_6143) );
bf01f01  g5968 ( .o(n4904), .a(net_7001) );
bf01f01  g5969 ( .o(n4913), .a(net_6573) );
bf01f01  g5970 ( .o(n4931), .a(_net_7823) );
bf01f01  g5971 ( .o(n4940), .a(_net_7812) );
bf01f01  g5972 ( .o(n4944), .a(net_7807) );
bf01f01  g5973 ( .o(n4947), .a(_net_7818) );
bf01f01  g5974 ( .o(n4957), .a(net_6718) );
bf01f01  g5975 ( .o(n4965), .a(_net_7823) );
bf01f01  g5976 ( .o(n4969), .a(_net_7811) );
bf01f01  g5977 ( .o(n4979), .a(net_6484) );
bf01f01  g5978 ( .o(n4983), .a(net_6858) );
bf01f01  g5979 ( .o(n4996), .a(_net_6065) );
bf01f01  g5980 ( .o(n5001), .a(net_6617) );
bf01f01  g5981 ( .o(n5005), .a(net_6854) );
bf01f01  g5982 ( .o(n5008), .a(net_6386) );
bf01f01  g5983 ( .o(n5023), .a(net_7539) );
bf01f01  g5984 ( .o(n5031), .a(_net_7819) );
bf01f01  g5985 ( .o(n5035), .a(_net_7817) );
bf01f01  g5986 ( .o(n5045), .a(net_7399) );
no02f01  g5987 ( .o(n5048), .a(n6966), .b(n7891) );
bf01f01  g5988 ( .o(n5053), .a(net_6970) );
no02f01  g5989 ( .o(n5056), .a(n6899_1), .b(n7254) );
bf01f01  g5990 ( .o(n5066), .a(_net_6115) );
bf01f01  g5991 ( .o(n5070), .a(_net_7801) );
bf01f01  g5992 ( .o(n5090), .a(net_7011) );
bf01f01  g5993 ( .o(n5098), .a(net_6399) );
bf01f01  g5994 ( .o(n5121), .a(net_6391) );
bf01f01  g5995 ( .o(n5126), .a(net_6589) );
bf01f01  g5996 ( .o(n5139), .a(net_6985) );
bf01f01  g5997 ( .o(n5148), .a(net_6572) );
bf01f01  g5998 ( .o(n5151), .a(_net_7821) );
bf01f01  g5999 ( .o(n5156), .a(net_6428) );
bf01f01  g6000 ( .o(n5159), .a(_net_7793) );
bf01f01  g6001 ( .o(n5173), .a(_net_7808) );
bf01f01  g6002 ( .o(n5178), .a(net_6841) );
bf01f01  g6003 ( .o(n5181), .a(x1519) );
bf01f01  g6004 ( .o(n5186), .a(net_7691) );
bf01f01  g6005 ( .o(n5189), .a(_net_7794) );
bf01f01  g6006 ( .o(n5193), .a(net_7802) );
bf01f01  g6007 ( .o(n5202), .a(_net_7811) );
bf01f01  g6008 ( .o(n5217), .a(net_6569) );
bf01f01  g6009 ( .o(n5221), .a(net_6857) );
bf01f01  g6010 ( .o(n5234), .a(_net_7806) );
bf01f01  g6011 ( .o(n5239), .a(net_6487) );
bf01f01  g6012 ( .o(n5242), .a(_net_7814) );
bf01f01  g6013 ( .o(n5246), .a(_net_7797) );
bf01f01  g6014 ( .o(n5261), .a(net_6843) );
bf01f01  g6015 ( .o(n5269), .a(_net_7798) );
bf01f01  g6016 ( .o(n5288), .a(net_6395) );
bf01f01  g6017 ( .o(n5298), .a(net_6965) );
bf01f01  g6018 ( .o(n5302), .a(_net_6128) );
bf01f01  g6019 ( .o(n5312), .a(net_7006) );
bf01f01  g6020 ( .o(n5326), .a(net_6844) );
bf01f01  g6021 ( .o(n5335), .a(net_7002) );
bf01f01  g6022 ( .o(n5339), .a(_net_6161) );
bf01f01  g6023 ( .o(n5349), .a(net_6987) );
bf01f01  g6024 ( .o(n5358), .a(net_6454) );
bf01f01  g6025 ( .o(n5362), .a(net_6460) );
bf01f01  g6026 ( .o(n5366), .a(net_6860) );
bf01f01  g6027 ( .o(n5375), .a(net_143) );
bf01f01  g6028 ( .o(n5380), .a(net_6729) );
bf01f01  g6029 ( .o(n5383), .a(_net_7819) );
bf01f01  g6030 ( .o(n5393), .a(net_7021) );
bf01f01  g6031 ( .o(n5402), .a(net_7151) );
bf01f01  g6032 ( .o(n5415), .a(_net_7804) );
bf01f01  g6033 ( .o(n5424), .a(_net_7797) );
bf01f01  g6034 ( .o(n5433), .a(_net_7801) );
bf01f01  g6035 ( .o(n5437), .a(net_6395) );
bf01f01  g6036 ( .o(n5441), .a(_net_7824) );
bf01f01  g6037 ( .o(n5451), .a(net_6436) );
bf01f01  g6038 ( .o(n5460), .a(_net_6075) );
no02f01  g6039 ( .o(n5464), .a(n6899_1), .b(n7246) );
bf01f01  g6040 ( .o(n5469), .a(net_6610) );
no02f01  g6041 ( .o(n5472), .a(n6966), .b(n7520) );
bf01f01  g6042 ( .o(n5481), .a(_net_7815) );
bf01f01  g6043 ( .o(n5486), .a(net_387) );
bf01f01  g6044 ( .o(n5500), .a(net_6575) );
bf01f01  g6045 ( .o(n5504), .a(net_7100) );
bf01f01  g6046 ( .o(n5513), .a(net_6024) );
bf01f01  g6047 ( .o(n5521), .a(net_7018) );
bf01f01  g6048 ( .o(n5539), .a(net_6839) );
bf01f01  g6049 ( .o(n5547), .a(_net_7808) );
bf01f01  g6050 ( .o(n5556), .a(net_6398) );
bf01f01  g6051 ( .o(n5560), .a(_net_7824) );
bf01f01  g6052 ( .o(n5575), .a(net_6620) );
bf01f01  g6053 ( .o(n5584), .a(net_7546) );
bf01f01  g6054 ( .o(n5588), .a(net_7235) );
no02f01  g6055 ( .o(n5591), .a(n6966), .b(n8514) );
bf01f01  g6056 ( .o(n5606), .a(_net_6172) );
bf01f01  g6057 ( .o(n5610), .a(_net_7796) );
bf01f01  g6058 ( .o(n5613), .a(_net_7813) );
bf01f01  g6059 ( .o(n5618), .a(_net_6067) );
bf01f01  g6060 ( .o(n5648), .a(net_6983) );
bf01f01  g6061 ( .o(n5651), .a(_net_7800) );
bf01f01  g6062 ( .o(n5655), .a(_net_7795) );
bf01f01  g6063 ( .o(n5664), .a(_net_7813) );
bf01f01  g6064 ( .o(n5679), .a(net_6727) );
bf01f01  g6065 ( .o(n5682), .a(_net_7795) );
bf01f01  g6066 ( .o(n5686), .a(x1358) );
bf01f01  g6067 ( .o(n5696), .a(net_6609) );
bf01f01  g6068 ( .o(n5704), .a(_net_7810) );
bf01f01  g6069 ( .o(n5713), .a(_net_7806) );
bf01f01  g6070 ( .o(n5717), .a(_net_7796) );
bf01f01  g6071 ( .o(n5727), .a(net_6598) );
bf01f01  g6072 ( .o(n5731), .a(net_7107) );
bf01f01  g6073 ( .o(n5735), .a(net_7026) );
bf01f01  g6074 ( .o(n5744), .a(net_7244) );
bf01f01  g6075 ( .o(n5758), .a(_net_6131) );
bf01f01  g6076 ( .o(n5763), .a(net_6560) );
bf01f01  g6077 ( .o(n5767), .a(net_6590) );
bf01f01  g6078 ( .o(n5771), .a(net_6480) );
bf01f01  g6079 ( .o(n5779), .a(_net_7812) );
bf01f01  g6080 ( .o(n5783), .a(net_6388) );
bf01f01  g6081 ( .o(n5787), .a(_net_7814) );
bf01f01  g6082 ( .o(n5796), .a(net_7802) );
bf01f01  g6083 ( .o(n5801), .a(net_7012) );
bf01f01  g6084 ( .o(n5805), .a(net_6437) );
bf01f01  g6085 ( .o(n5824), .a(net_7113) );
bf01f01  g6086 ( .o(n5833), .a(net_6878) );
bf01f01  g6087 ( .o(n5836), .a(net_7802) );
bf01f01  g6088 ( .o(n5840), .a(_net_7793) );
bf01f01  g6089 ( .o(n5860), .a(net_6479) );
bf01f01  g6090 ( .o(n5864), .a(net_7102) );
no02f01  g6091 ( .o(n5867), .a(n6899_1), .b(n7560) );
bf01f01  g6092 ( .o(n5872), .a(_net_6144) );
bf01f01  g6093 ( .o(n5876), .a(_net_7822) );
bf01f01  g6094 ( .o(n5881), .a(net_6720) );
bf01f01  g6095 ( .o(n5894), .a(net_6391) );
bf01f01  g6096 ( .o(n5903), .a(net_7790) );
bf01f01  g6097 ( .o(n5908), .a(_net_6180) );
bf01f01  g6098 ( .o(n5912), .a(_net_7811) );
bf01f01  g6099 ( .o(n5917), .a(net_6971) );
bf01f01  g6100 ( .o(n5920), .a(_net_7795) );
bf01f01  g6101 ( .o(n5930), .a(net_6580) );
bf01f01  g6102 ( .o(n5934), .a(net_7127) );
bf01f01  g6103 ( .o(n5943), .a(net_6887) );
bf01f01  g6104 ( .o(n5947), .a(net_6562) );
bf01f01  g6105 ( .o(n5951), .a(net_6973) );
bf01f01  g6106 ( .o(n5955), .a(_net_6079) );
bf01f01  g6107 ( .o(n5964), .a(x1557) );
bf01f01  g6108 ( .o(n5968), .a(_net_7821) );
bf01f01  g6109 ( .o(n5978), .a(net_6618) );
bf01f01  g6110 ( .o(n6002), .a(net_7712) );
bf01f01  g6111 ( .o(n6006), .a(net_7115) );
bf01f01  g6112 ( .o(n6009), .a(net_7802) );
bf01f01  g6113 ( .o(n6014), .a(net_5861) );
bf01f01  g6114 ( .o(n6019), .a(_net_6118) );
bf01f01  g6115 ( .o(n6034), .a(net_7125) );
bf01f01  g6116 ( .o(n6043), .a(net_6733) );
bf01f01  g6117 ( .o(n6047), .a(_net_6166) );
bf01f01  g6118 ( .o(n6056), .a(_net_7805) );
bf01f01  g6119 ( .o(n6066), .a(net_6466) );
bf01f01  g6120 ( .o(n6069), .a(_net_7800) );
bf01f01  g6121 ( .o(n6078), .a(x1572) );
bf01f01  g6122 ( .o(n6098), .a(_net_6139) );
bf01f01  g6123 ( .o(n6102), .a(_net_7798) );
bf01f01  g6124 ( .o(n6106), .a(_net_7824) );
no02f01  g6125 ( .o(n6110), .a(n6899_1), .b(n7895) );
bf01f01  g6126 ( .o(n6114), .a(net_7807) );
bf01f01  g6127 ( .o(n6128), .a(_net_7803) );
bf01f01  g6128 ( .o(n6132), .a(x1479) );
bf01f01  g6129 ( .o(n6136), .a(net_6384) );
bf01f01  g6130 ( .o(n6145), .a(net_6594) );
bf01f01  g6131 ( .o(n6148), .a(_net_7800) );
bf01f01  g6132 ( .o(n6158), .a(net_6892) );
bf01f01  g6133 ( .o(n6161), .a(_net_7816) );
bf01f01  g6134 ( .o(n6176), .a(_net_6105) );
bf01f01  g6135 ( .o(n6181), .a(_net_6113) );
bf01f01  g6136 ( .o(n6195), .a(_net_7813) );
bf01f01  g6137 ( .o(n6204), .a(net_6397) );
bf01f01  g6138 ( .o(n6214), .a(net_7385) );
no02f01  g6139 ( .o(n6222), .a(n6966), .b(n7142_1) );
in01f01  g6140 ( .o(n6231), .a(n7343) );
bf01f01  g6141 ( .o(n6235), .a(net_7799) );
bf01f01  g6142 ( .o(n6239), .a(net_6400) );
bf01f01  g6143 ( .o(n6254), .a(net_6697) );
bf01f01  g6144 ( .o(n6258), .a(net_6750) );
bf01f01  g6145 ( .o(n6261), .a(x1534) );
bf01f01  g6146 ( .o(n6276), .a(_net_5964) );
bf01f01  g6147 ( .o(n6285), .a(net_146) );
bf01f01  g6148 ( .o(n6299), .a(net_7130) );
no02f01  g6149 ( .o(n6302), .a(n6867_1), .b(n9980) );
bf01f01  g6150 ( .o(n6306), .a(net_6393) );
bf01f01  g6151 ( .o(n6316), .a(net_7770) );
bf01f01  g6152 ( .o(n6319), .a(net_389) );
bf01f01  g6153 ( .o(n6329), .a(net_7161) );
bf01f01  g6154 ( .o(n6332), .a(net_6396) );
bf01f01  g6155 ( .o(n6342), .a(net_6469) );
bf01f01  g6156 ( .o(n6350), .a(_net_7794) );
bf01f01  g6157 ( .o(n6354), .a(net_6747) );
bf01f01  g6158 ( .o(n6357), .a(_net_7817) );
bf01f01  g6159 ( .o(n6367), .a(net_6439) );
bf01f01  g6160 ( .o(n6386), .a(net_7117) );
bf01f01  g6161 ( .o(n6390), .a(_net_6165) );
bf01f01  g6162 ( .o(n6399), .a(net_6398) );
bf01f01  g6163 ( .o(n6403), .a(net_6738) );
bf01f01  g6164 ( .o(n6407), .a(net_6481) );
bf01f01  g6165 ( .o(n6415), .a(_net_7806) );
bf01f01  g6166 ( .o(n6419), .a(_net_7795) );
bf01f01  g6167 ( .o(n6423), .a(net_6382) );
bf01f01  g6168 ( .o(n6441), .a(net_7802) );
bf01f01  g6169 ( .o(n6446), .a(net_6702) );
bf01f01  g6170 ( .o(n6460), .a(_net_6152) );
bf01f01  g6171 ( .o(n6464), .a(_net_7817) );
bf01f01  g6172 ( .o(n6469), .a(net_6980) );
bf01f01  g6173 ( .o(n6472), .a(_net_7812) );
bf01f01  g6174 ( .o(n6477), .a(net_7148) );
bf01f01  g6175 ( .o(n6480), .a(_net_7796) );
bf01f01  g6176 ( .o(n6485), .a(net_6462) );
bf01f01  g6177 ( .o(n6489), .a(net_7242) );
bf01f01  g6178 ( .o(n6498), .a(_net_6159) );
bf01f01  g6179 ( .o(n6502), .a(net_7807) );
bf01f01  g6180 ( .o(n6507), .a(net_6563) );
bf01f01  g6181 ( .o(n6511), .a(net_6604) );
bf01f01  g6182 ( .o(n6515), .a(net_6836) );
bf01f01  g6183 ( .o(n6519), .a(net_6866) );
bf01f01  g6184 ( .o(n6522), .a(x1501) );
bf01f01  g6185 ( .o(n6531), .a(net_6385) );
no02f01  g6186 ( .o(n6535), .a(n6966), .b(n8812) );
bf01f01  g6187 ( .o(n6550), .a(net_7397) );
bf01f01  g6188 ( .o(n6554), .a(net_6713) );
bf01f01  g6189 ( .o(n6563), .a(net_6846) );
bf01f01  g6190 ( .o(n6566), .a(net_6381) );
no02f01  g6191 ( .o(n6574), .a(n6867_1), .b(n7650) );
bf01f01  g6192 ( .o(n6578), .a(net_132) );
bf01f01  g6193 ( .o(n6586), .a(_net_7817) );
bf01f01  g6194 ( .o(n6611), .a(_net_6096) );
bf01f01  g6195 ( .o(n6615), .a(_net_7817) );
bf01f01  g6196 ( .o(n6619), .a(_net_7793) );
bf01f01  g6197 ( .o(n6629), .a(_net_6085) );
bf01f01  g6198 ( .o(n6638), .a(_net_7817) );
bf01f01  g6199 ( .o(n6648), .a(net_7145) );
no02f01  g6200 ( .o(n6656), .a(n6966), .b(n8812) );
bf01f01  g6201 ( .o(n6661), .a(net_6424) );
bf01f01  g6202 ( .o(n6669), .a(net_6390) );
bf01f01  g6203 ( .o(n6674), .a(net_6834) );
bf01f01  g6204 ( .o(n6678), .a(net_6708) );
bf01f01  g6205 ( .o(n6687), .a(net_6997) );
bf01f01  g6206 ( .o(n6700), .a(_net_6157) );
bf01f01  g6207 ( .o(n6704), .a(_net_7794) );
bf01f01  g6208 ( .o(n6713), .a(_net_7793) );
bf01f01  g6209 ( .o(n6717), .a(_net_7796) );
bf01f01  g6210 ( .o(n6732), .a(_net_7810) );
bf01f01  g6211 ( .o(n6736), .a(net_7799) );
bf01f01  g6212 ( .o(n6746), .a(net_7549) );
bf01f01  g6213 ( .o(n6749), .a(_net_7810) );
bf01f01  g6214 ( .o(n6752), .a(_net_7794) );
bf01f01  g6215 ( .o(n6756), .a(net_6389) );
bf01f01  g6216 ( .o(n6761), .a(net_6728) );
bf01f01  g6217 ( .o(n6770), .a(net_6830) );
bf01f01  g6218 ( .o(n6783), .a(_net_7824) );
bf01f01  g6219 ( .o(n6793), .a(net_7394) );
bf01f01  g6220 ( .o(n6796), .a(_net_7801) );
bf01f01  g6221 ( .o(n6806), .a(net_6990) );
bf01f01  g6222 ( .o(n6809), .a(net_7799) );
bf01f01  g6223 ( .o(n6813), .a(_net_7798) );
bf01f01  g6224 ( .o(n6822), .a(net_6392) );
bf01f01  g6225 ( .o(n6826), .a(_net_7809) );
bf01f01  g6226 ( .o(n6836), .a(net_7025) );
bf01f01  g6227 ( .o(n6860), .a(net_6470) );
bf01f01  g6228 ( .o(n6863), .a(_net_7796) );
bf01f01  g6229 ( .o(n6867), .a(_net_7823) );
bf01f01  g6230 ( .o(n6876), .a(net_7807) );
bf01f01  g6231 ( .o(n6886), .a(net_6712) );
bf01f01  g6232 ( .o(n6895), .a(net_7009) );
bf01f01  g6233 ( .o(n6899), .a(net_6607) );
bf01f01  g6234 ( .o(n6902), .a(net_6395) );
bf01f01  g6235 ( .o(n6906), .a(_net_7804) );
bf01f01  g6236 ( .o(n6910), .a(_net_7818) );
no02f01  g6237 ( .o(n6919), .a(n6899_1), .b(n8964) );
bf01f01  g6238 ( .o(n6934), .a(net_7150) );
bf01f01  g6239 ( .o(n6947), .a(net_6390) );
bf01f01  g6240 ( .o(n6957), .a(net_6587) );
bf01f01  g6241 ( .o(n6960), .a(_net_7812) );
bf01f01  g6242 ( .o(n6974), .a(net_7245) );
bf01f01  g6243 ( .o(n6977), .a(_net_7816) );
bf01f01  g6244 ( .o(n6982), .a(_net_6146) );
bf01f01  g6245 ( .o(n6986), .a(net_7802) );
bf01f01  g6246 ( .o(n6990), .a(_net_7800) );
bf01f01  g6247 ( .o(n7005), .a(net_6621) );
bf01f01  g6248 ( .o(n7009), .a(net_6597) );
bf01f01  g6249 ( .o(n7027), .a(net_7802) );
bf01f01  g6250 ( .o(n7036), .a(net_6388) );
bf01f01  g6251 ( .o(n7041), .a(net_6889) );
bf01f01  g6252 ( .o(n7045), .a(_net_6182) );
bf01f01  g6253 ( .o(n7049), .a(net_6393) );
bf01f01  g6254 ( .o(n7062), .a(_net_7804) );
bf01f01  g6255 ( .o(n7082), .a(net_6872) );
no02f01  g6256 ( .o(n7085), .a(n6867_1), .b(n7175) );
bf01f01  g6257 ( .o(n7089), .a(_net_7811) );
bf01f01  g6258 ( .o(n7093), .a(net_6398) );
bf01f01  g6259 ( .o(n7098), .a(net_7152) );
bf01f01  g6260 ( .o(n7111), .a(_net_7821) );
bf01f01  g6261 ( .o(n7116), .a(_net_6133) );
bf01f01  g6262 ( .o(n7120), .a(_net_7803) );
bf01f01  g6263 ( .o(n7125), .a(net_6561) );
bf01f01  g6264 ( .o(n7128), .a(_net_7798) );
no02f01  g6265 ( .o(n7142), .a(n6867_1), .b(n9870) );
bf01f01  g6266 ( .o(n7147), .a(_net_6073) );
bf01f01  g6267 ( .o(n7151), .a(_net_7816) );
bf01f01  g6268 ( .o(n7155), .a(_net_7824) );
bf01f01  g6269 ( .o(n7160), .a(net_6862) );
bf01f01  g6270 ( .o(n7167), .a(net_141) );
bf01f01  g6271 ( .o(n7182), .a(net_7543) );
no02f01  g6272 ( .o(n7185), .a(n6899_1), .b(n8229) );
bf01f01  g6273 ( .o(n7190), .a(net_6430) );
bf01f01  g6274 ( .o(n7199), .a(net_7238) );
bf01f01  g6275 ( .o(n7203), .a(net_6477) );
bf01f01  g6276 ( .o(n7212), .a(net_6559) );
bf01f01  g6277 ( .o(n7230), .a(_net_7823) );
bf01f01  g6278 ( .o(n7249), .a(x1486) );
bf01f01  g6279 ( .o(n7252), .a(_net_7804) );
bf01f01  g6280 ( .o(n7256), .a(net_7792) );
bf01f01  g6281 ( .o(n7260), .a(_net_7797) );
bf01f01  g6282 ( .o(n7284), .a(_net_7816) );
bf01f01  g6283 ( .o(n7288), .a(net_6397) );
bf01f01  g6284 ( .o(n7292), .a(x1406) );
bf01f01  g6285 ( .o(n7312), .a(net_6869) );
bf01f01  g6286 ( .o(n7316), .a(_net_6178) );
bf01f01  g6287 ( .o(n7326), .a(net_6715) );
bf01f01  g6288 ( .o(n7330), .a(_net_6088) );
bf01f01  g6289 ( .o(n7335), .a(net_5860) );
bf01f01  g6290 ( .o(n7344), .a(_net_7803) );
bf01f01  g6291 ( .o(n7349), .a(net_6058) );
bf01f01  g6292 ( .o(n7359), .a(net_7008) );
bf01f01  g6293 ( .o(n7368), .a(_net_6121) );
bf01f01  g6294 ( .o(n7372), .a(_net_7798) );
bf01f01  g6295 ( .o(n7376), .a(net_134) );
bf01f01  g6296 ( .o(n7391), .a(net_7118) );
bf01f01  g6297 ( .o(n7404), .a(_net_7808) );
bf01f01  g6298 ( .o(n7408), .a(_net_7819) );
bf01f01  g6299 ( .o(n7413), .a(net_6994) );
bf01f01  g6300 ( .o(n7417), .a(_net_6081) );
bf01f01  g6301 ( .o(n7427), .a(_net_6149) );
bf01f01  g6302 ( .o(n7442), .a(net_6700) );
bf01f01  g6303 ( .o(n7446), .a(net_6696) );
bf01f01  g6304 ( .o(n7450), .a(net_6740) );
bf01f01  g6305 ( .o(n7463), .a(_net_7814) );
bf01f01  g6306 ( .o(n7468), .a(_net_6141) );
bf01f01  g6307 ( .o(n7482), .a(_net_7810) );
bf01f01  g6308 ( .o(n7492), .a(net_6726) );
bf01f01  g6309 ( .o(n7505), .a(net_6383) );
bf01f01  g6310 ( .o(n7509), .a(_net_7809) );
bf01f01  g6311 ( .o(n7513), .a(_net_7823) );
bf01f01  g6312 ( .o(n7522), .a(_net_7809) );
bf01f01  g6313 ( .o(n7527), .a(net_6451) );
bf01f01  g6314 ( .o(n7530), .a(_net_7808) );
bf01f01  g6315 ( .o(n7535), .a(net_6757) );
bf01f01  g6316 ( .o(n7553), .a(_net_6090) );
bf01f01  g6317 ( .o(n7567), .a(x1345) );
bf01f01  g6318 ( .o(n7577), .a(_net_6123) );
bf01f01  g6319 ( .o(n7581), .a(_net_7814) );
no02f01  g6320 ( .o(n7599), .a(n6867_1), .b(n10215) );
bf01f01  g6321 ( .o(n7604), .a(net_6716) );
bf01f01  g6322 ( .o(n7618), .a(net_7392) );
no02f01  g6323 ( .o(n7626), .a(n6867_1), .b(n8845_1) );
no02f01  g6324 ( .o(n7635), .a(n6966), .b(n7188) );
bf01f01  g6325 ( .o(n7644), .a(net_6396) );
bf01f01  g6326 ( .o(n7654), .a(net_7139) );
bf01f01  g6327 ( .o(n7658), .a(net_6467) );
no02f01  g6328 ( .o(n7661), .a(n6867_1), .b(n9980) );
bf01f01  g6329 ( .o(n7700), .a(net_6748) );
bf01f01  g6330 ( .o(n7704), .a(_net_6108) );
bf01f01  g6331 ( .o(n7714), .a(_net_226) );
bf01f01  g6332 ( .o(n7719), .a(net_6837) );
no02f01  g6333 ( .o(n7732), .a(n6867_1), .b(n10215) );
bf01f01  g6334 ( .o(n7756), .a(net_6441) );
bf01f01  g6335 ( .o(n7760), .a(net_7143) );
bf01f01  g6336 ( .o(n7764), .a(net_7160) );
bf01f01  g6337 ( .o(n7776), .a(net_6396) );
bf01f01  g6338 ( .o(n7779), .a(_net_7824) );
bf01f01  g6339 ( .o(n7784), .a(net_6710) );
bf01f01  g6340 ( .o(n7802), .a(_net_7800) );
bf01f01  g6341 ( .o(n7806), .a(_net_7815) );
bf01f01  g6342 ( .o(n7810), .a(_net_7797) );
bf01f01  g6343 ( .o(n7815), .a(net_6734) );
bf01f01  g6344 ( .o(n7818), .a(net_6386) );
bf01f01  g6345 ( .o(n7826), .a(_net_7801) );
bf01f01  g6346 ( .o(n7831), .a(net_6566) );
bf01f01  g6347 ( .o(n7840), .a(_net_6135) );
bf01f01  g6348 ( .o(n7848), .a(net_6382) );
bf01f01  g6349 ( .o(n7867), .a(net_6393) );
bf01f01  g6350 ( .o(n7871), .a(_net_7800) );
bf01f01  g6351 ( .o(n7875), .a(net_6874) );
no02f01  g6352 ( .o(n7878), .a(n6966), .b(n8899_1) );
bf01f01  g6353 ( .o(n7883), .a(_net_6148) );
bf01f01  g6354 ( .o(n7893), .a(net_7249) );
bf01f01  g6355 ( .o(n7906), .a(_net_7822) );
bf01f01  g6356 ( .o(n7916), .a(_net_6167) );
bf01f01  g6357 ( .o(n7920), .a(net_6386) );
no02f01  g6358 ( .o(n7924), .a(n6867_1), .b(n8170_1) );
bf01f01  g6359 ( .o(n7929), .a(net_6568) );
bf01f01  g6360 ( .o(n7937), .a(_net_7798) );
bf01f01  g6361 ( .o(n7942), .a(net_7540) );
bf01f01  g6362 ( .o(n7945), .a(net_6390) );
bf01f01  g6363 ( .o(n7955), .a(net_6724) );
bf01f01  g6364 ( .o(n7958), .a(net_138) );
bf01f01  g6365 ( .o(n7962), .a(_net_7811) );
bf01f01  g6366 ( .o(n7967), .a(net_6992) );
no02f01  g6367 ( .o(n7970), .a(n6867_1), .b(n7601) );
bf01f01  g6368 ( .o(n7989), .a(_net_7821) );
bf01f01  g6369 ( .o(n7994), .a(net_6585) );
bf01f01  g6370 ( .o(n7997), .a(_net_7820) );
bf01f01  g6371 ( .o(n8002), .a(net_6975) );
bf01f01  g6372 ( .o(n8005), .a(net_6394) );
bf01f01  g6373 ( .o(n8015), .a(net_7131) );
bf01f01  g6374 ( .o(n8028), .a(_net_7815) );
in01f01  g6375 ( .o(n8042), .a(n7343) );
bf01f01  g6376 ( .o(n8047), .a(_net_6169) );
bf01f01  g6377 ( .o(n8051), .a(net_6399) );
bf01f01  g6378 ( .o(n8056), .a(net_6988) );
bf01f01  g6379 ( .o(n8059), .a(_net_7819) );
bf01f01  g6380 ( .o(n8064), .a(net_6968) );
bf01f01  g6381 ( .o(n8067), .a(_net_7813) );
bf01f01  g6382 ( .o(n8072), .a(net_6614) );
bf01f01  g6383 ( .o(n8075), .a(_net_7824) );
bf01f01  g6384 ( .o(n8085), .a(net_6596) );
bf01f01  g6385 ( .o(n8088), .a(_net_7808) );
bf01f01  g6386 ( .o(n8092), .a(_net_7801) );
bf01f01  g6387 ( .o(n8116), .a(_net_7801) );
bf01f01  g6388 ( .o(n8125), .a(_net_7795) );
bf01f01  g6389 ( .o(n8140), .a(net_7141) );
bf01f01  g6390 ( .o(n8144), .a(net_6571) );
bf01f01  g6391 ( .o(n8147), .a(_net_7808) );
no02f01  g6392 ( .o(n8156), .a(n6899_1), .b(n8229) );
bf01f01  g6393 ( .o(n8166), .a(net_7715) );
bf01f01  g6394 ( .o(n8174), .a(_net_7820) );
bf01f01  g6395 ( .o(n8183), .a(net_7802) );
bf01f01  g6396 ( .o(n8188), .a(net_6835) );
bf01f01  g6397 ( .o(n8206), .a(_net_7816) );
bf01f01  g6398 ( .o(n8220), .a(net_6389) );
bf01f01  g6399 ( .o(n8228), .a(_net_7810) );
bf01f01  g6400 ( .o(n8232), .a(net_7807) );
bf01f01  g6401 ( .o(n8241), .a(net_6385) );
bf01f01  g6402 ( .o(n8245), .a(net_7799) );
bf01f01  g6403 ( .o(n8249), .a(net_6388) );
no02f01  g6404 ( .o(n8262), .a(n6966), .b(n7142_1) );
bf01f01  g6405 ( .o(n8266), .a(net_7799) );
bf01f01  g6406 ( .o(n8271), .a(_net_6116) );
bf01f01  g6407 ( .o(n8276), .a(net_6615) );
bf01f01  g6408 ( .o(n8280), .a(net_7538) );
bf01f01  g6409 ( .o(n8289), .a(_net_6125) );
bf01f01  g6410 ( .o(n8303), .a(_net_7810) );
bf01f01  g6411 ( .o(n8307), .a(_net_7811) );
bf01f01  g6412 ( .o(n8311), .a(_net_7816) );
bf01f01  g6413 ( .o(n8316), .a(net_6853) );
bf01f01  g6414 ( .o(n8320), .a(net_7138) );
bf01f01  g6415 ( .o(n8329), .a(_net_6100) );
bf01f01  g6416 ( .o(n8334), .a(net_6851) );
bf01f01  g6417 ( .o(n8337), .a(_net_7806) );
bf01f01  g6418 ( .o(n8340), .a(_net_7812) );
bf01f01  g6419 ( .o(n8350), .a(net_7023) );
bf01f01  g6420 ( .o(n8359), .a(net_6427) );
no02f01  g6421 ( .o(n8362), .a(n6966), .b(n7276) );
bf01f01  g6422 ( .o(n8392), .a(net_6425) );
bf01f01  g6423 ( .o(n8401), .a(net_7104) );
bf01f01  g6424 ( .o(n8415), .a(net_7137) );
bf01f01  g6425 ( .o(n8418), .a(net_6392) );
bf01f01  g6426 ( .o(n8422), .a(net_7237) );
bf01f01  g6427 ( .o(n8430), .a(net_6387) );
bf01f01  g6428 ( .o(n8438), .a(net_391) );
no02f01  g6429 ( .o(n8447), .a(n6899_1), .b(n7509_1) );
no02f01  g6430 ( .o(n8451), .a(n6867_1), .b(n7601) );
bf01f01  g6431 ( .o(n8455), .a(_net_7813) );
bf01f01  g6432 ( .o(n8459), .a(_net_7823) );
bf01f01  g6433 ( .o(n8464), .a(net_6742) );
bf01f01  g6434 ( .o(n8467), .a(_net_7804) );
bf01f01  g6435 ( .o(n8477), .a(net_6754) );
bf01f01  g6436 ( .o(n8491), .a(net_7020) );
bf01f01  g6437 ( .o(n8494), .a(_net_7810) );
bf01f01  g6438 ( .o(n8504), .a(net_6622) );
bf01f01  g6439 ( .o(n8513), .a(net_6744) );
bf01f01  g6440 ( .o(n8522), .a(net_6838) );
bf01f01  g6441 ( .o(n8535), .a(_net_7806) );
bf01f01  g6442 ( .o(n8544), .a(_net_7804) );
bf01f01  g6443 ( .o(n8549), .a(net_6707) );
bf01f01  g6444 ( .o(n8552), .a(_net_7795) );
bf01f01  g6445 ( .o(n8561), .a(_net_7824) );
bf01f01  g6446 ( .o(n8565), .a(_net_7797) );
bf01f01  g6447 ( .o(n8575), .a(net_6475) );
bf01f01  g6448 ( .o(n8578), .a(net_6385) );
bf01f01  g6449 ( .o(n8598), .a(net_6695) );
bf01f01  g6450 ( .o(n8612), .a(net_6463) );
bf01f01  g6451 ( .o(n8621), .a(net_6831) );
bf01f01  g6452 ( .o(n8628), .a(_net_7814) );
bf01f01  g6453 ( .o(n8632), .a(_net_7821) );
bf01f01  g6454 ( .o(n8637), .a(net_6013) );
bf01f01  g6455 ( .o(n8641), .a(net_6756) );
bf01f01  g6456 ( .o(n8650), .a(net_6865) );
bf01f01  g6457 ( .o(n8654), .a(net_6577) );
bf01f01  g6458 ( .o(n8658), .a(net_6600) );
no02f01  g6459 ( .o(n8666), .a(n6899_1), .b(n8964) );
bf01f01  g6460 ( .o(n8681), .a(net_6891) );
bf01f01  g6461 ( .o(n8685), .a(net_6722) );
bf01f01  g6462 ( .o(n8698), .a(x1451) );
no02f01  g6463 ( .o(n8711), .a(n6867_1), .b(n8845_1) );
bf01f01  g6464 ( .o(n8715), .a(net_6388) );
no02f01  g6465 ( .o(n8734), .a(n6899_1), .b(n7895) );
bf01f01  g6466 ( .o(n8739), .a(net_7389) );
bf01f01  g6467 ( .o(n8757), .a(net_140) );
bf01f01  g6468 ( .o(n8767), .a(net_7110) );
bf01f01  g6469 ( .o(n8784), .a(x1390) );
bf01f01  g6470 ( .o(n8788), .a(_net_7808) );
bf01f01  g6471 ( .o(n8793), .a(net_6882) );
bf01f01  g6472 ( .o(n8797), .a(net_6457) );
bf01f01  g6473 ( .o(n8800), .a(_net_7808) );
bf01f01  g6474 ( .o(n8805), .a(net_6982) );
bf01f01  g6475 ( .o(n8813), .a(_net_7797) );
bf01f01  g6476 ( .o(n8823), .a(net_7542) );
bf01f01  g6477 ( .o(n8826), .a(_net_7822) );
bf01f01  g6478 ( .o(n8835), .a(_net_7811) );
bf01f01  g6479 ( .o(n8864), .a(x1494) );
bf01f01  g6480 ( .o(n8873), .a(net_151) );
bf01f01  g6481 ( .o(n8877), .a(net_6389) );
bf01f01  g6482 ( .o(n8882), .a(net_6060) );
bf01f01  g6483 ( .o(n8886), .a(_net_7819) );
bf01f01  g6484 ( .o(n8891), .a(net_7132) );
no02f01  g6485 ( .o(n8899), .a(n6899_1), .b(n7507) );
bf01f01  g6486 ( .o(n8903), .a(_net_7822) );
bf01f01  g6487 ( .o(n8908), .a(_net_6119) );
bf01f01  g6488 ( .o(n8912), .a(_net_7804) );
bf01f01  g6489 ( .o(n8926), .a(_net_7809) );
bf01f01  g6490 ( .o(n8931), .a(net_7243) );
no02f01  g6491 ( .o(n8934), .a(n6899_1), .b(n8826_1) );
bf01f01  g6492 ( .o(n8939), .a(net_6458) );
bf01f01  g6493 ( .o(n8943), .a(_net_6086) );
bf01f01  g6494 ( .o(n8958), .a(_net_6130) );
bf01f01  g6495 ( .o(n8963), .a(net_7544) );
bf01f01  g6496 ( .o(n8971), .a(net_7807) );
bf01f01  g6497 ( .o(n8981), .a(_net_6154) );
bf01f01  g6498 ( .o(n8990), .a(net_6386) );
bf01f01  g6499 ( .o(n9010), .a(net_6582) );
bf01f01  g6500 ( .o(n9014), .a(net_7017) );
bf01f01  g6501 ( .o(n9017), .a(net_136) );
bf01f01  g6502 ( .o(n9022), .a(net_6445) );
bf01f01  g6503 ( .o(n9025), .a(_net_7800) );
bf01f01  g6504 ( .o(n9034), .a(net_6864) );
bf01f01  g6505 ( .o(n9037), .a(_net_7805) );
bf01f01  g6506 ( .o(n9047), .a(_net_189) );
bf01f01  g6507 ( .o(n9057), .a(net_6966) );
no02f01  g6508 ( .o(n9060), .a(n6899_1), .b(n7069) );
bf01f01  g6509 ( .o(n9065), .a(net_6984) );
bf01f01  g6510 ( .o(n9069), .a(_net_6110) );
bf01f01  g6511 ( .o(n9079), .a(net_7101) );
bf01f01  g6512 ( .o(n9082), .a(_net_7817) );
bf01f01  g6513 ( .o(n9086), .a(_net_7819) );
bf01f01  g6514 ( .o(n9091), .a(_net_6094) );
bf01f01  g6515 ( .o(n9110), .a(x1511) );
bf01f01  g6516 ( .o(n9120), .a(net_7155) );
bf01f01  g6517 ( .o(n9134), .a(_net_6137) );
bf01f01  g6518 ( .o(n9138), .a(_net_7793) );
bf01f01  g6519 ( .o(n9143), .a(net_6876) );
bf01f01  g6520 ( .o(n9146), .a(_net_7803) );
bf01f01  g6521 ( .o(n9160), .a(net_6393) );
bf01f01  g6522 ( .o(n9164), .a(_net_7811) );
bf01f01  g6523 ( .o(n9169), .a(net_6565) );
bf01f01  g6524 ( .o(n9178), .a(_net_6077) );
bf01f01  g6525 ( .o(n9182), .a(_net_7797) );
bf01f01  g6526 ( .o(n9196), .a(net_6383) );
no02f01  g6527 ( .o(n9215), .a(n6899_1), .b(n7246) );
bf01f01  g6528 ( .o(n9225), .a(net_7156) );
no02f01  g6529 ( .o(n9228), .a(n6867_1), .b(n7978) );
bf01f01  g6530 ( .o(n9238), .a(net_6705) );
bf01f01  g6531 ( .o(n9242), .a(net_6483) );
bf01f01  g6532 ( .o(n9245), .a(_net_7800) );
bf01f01  g6533 ( .o(n9250), .a(net_6701) );
bf01f01  g6534 ( .o(n9254), .a(net_7103) );
bf01f01  g6535 ( .o(n9267), .a(net_7807) );
bf01f01  g6536 ( .o(n9287), .a(net_6848) );
bf01f01  g6537 ( .o(n9290), .a(_net_7820) );
bf01f01  g6538 ( .o(n9294), .a(_net_7816) );
no02f01  g6539 ( .o(n9298), .a(n6966), .b(n10317) );
no02f01  g6540 ( .o(n9302), .a(n6867_1), .b(n7203_1) );
no02f01  g6541 ( .o(n9316), .a(n6899_1), .b(n7514) );
bf01f01  g6542 ( .o(n9326), .a(net_6749) );
bf01f01  g6543 ( .o(n9339), .a(_net_7800) );
bf01f01  g6544 ( .o(n9343), .a(_net_7808) );
bf01f01  g6545 ( .o(n9348), .a(net_7541) );
bf01f01  g6546 ( .o(n9356), .a(_net_7794) );
bf01f01  g6547 ( .o(n9361), .a(net_6464) );
bf01f01  g6548 ( .o(n9365), .a(_net_6089) );
bf01f01  g6549 ( .o(n9370), .a(net_7099) );
bf01f01  g6550 ( .o(n9373), .a(_net_7810) );
bf01f01  g6551 ( .o(n9377), .a(_net_7820) );
bf01f01  g6552 ( .o(n9381), .a(_net_7821) );
bf01f01  g6553 ( .o(n9385), .a(_net_7805) );
bf01f01  g6554 ( .o(n9390), .a(net_6601) );
bf01f01  g6555 ( .o(n9393), .a(_net_7804) );
bf01f01  g6556 ( .o(n9398), .a(_net_6102) );
bf01f01  g6557 ( .o(n9402), .a(x0) );
bf01f01  g6558 ( .o(n9405), .a(_net_7808) );
bf01f01  g6559 ( .o(n9425), .a(net_6459) );
bf01f01  g6560 ( .o(n9428), .a(_net_7808) );
bf01f01  g6561 ( .o(n9431), .a(_net_7810) );
bf01f01  g6562 ( .o(n9445), .a(net_6731) );
bf01f01  g6563 ( .o(n9459), .a(net_7709) );
bf01f01  g6564 ( .o(n9462), .a(_net_7816) );
bf01f01  g6565 ( .o(n9467), .a(net_6972) );
bf01f01  g6566 ( .o(n9470), .a(net_6394) );
bf01f01  g6567 ( .o(n9475), .a(net_6842) );
no02f01  g6568 ( .o(n9478), .a(n6867_1), .b(n9870) );
bf01f01  g6569 ( .o(n9483), .a(net_6611) );
bf01f01  g6570 ( .o(n9502), .a(_net_6163) );
bf01f01  g6571 ( .o(n9517), .a(net_6871) );
bf01f01  g6572 ( .o(n9520), .a(net_6391) );
bf01f01  g6573 ( .o(n9525), .a(net_7015) );
bf01f01  g6574 ( .o(n9528), .a(_net_7805) );
bf01f01  g6575 ( .o(n9537), .a(_net_7817) );
bf01f01  g6576 ( .o(n9541), .a(_net_7813) );
no02f01  g6577 ( .o(n9549), .a(n6867_1), .b(n7175) );
bf01f01  g6578 ( .o(n9579), .a(net_6840) );
bf01f01  g6579 ( .o(n9588), .a(net_6455) );
bf01f01  g6580 ( .o(n9606), .a(_net_7821) );
bf01f01  g6581 ( .o(n9611), .a(_net_6111) );
bf01f01  g6582 ( .o(n9620), .a(_net_7820) );
bf01f01  g6583 ( .o(n9624), .a(_net_7803) );
bf01f01  g6584 ( .o(n9628), .a(net_153) );
bf01f01  g6585 ( .o(n9642), .a(_net_7814) );
bf01f01  g6586 ( .o(n9647), .a(net_7386) );
bf01f01  g6587 ( .o(n9651), .a(net_7548) );
bf01f01  g6588 ( .o(n9660), .a(net_7005) );
bf01f01  g6589 ( .o(n9668), .a(net_6383) );
bf01f01  g6590 ( .o(n9687), .a(net_6392) );
bf01f01  g6591 ( .o(n9692), .a(net_6703) );
bf01f01  g6592 ( .o(n9695), .a(net_6381) );
bf01f01  g6593 ( .o(n9704), .a(_net_7804) );
bf01f01  g6594 ( .o(n9724), .a(_net_6162) );
bf01f01  g6595 ( .o(n9729), .a(net_6472) );
bf01f01  g6596 ( .o(n9737), .a(x1398) );
bf01f01  g6597 ( .o(n9746), .a(_net_7812) );
bf01f01  g6598 ( .o(n9750), .a(_net_7795) );
no02f01  g6599 ( .o(n9754), .a(n6867_1), .b(n8173) );
no02f01  g6600 ( .o(n9758), .a(n6966), .b(n7276) );
bf01f01  g6601 ( .o(n9783), .a(net_7027) );
bf01f01  g6602 ( .o(n9796), .a(_net_7810) );
bf01f01  g6603 ( .o(n9805), .a(net_6399) );
bf01f01  g6604 ( .o(n9809), .a(net_6388) );
no02f01  g6605 ( .o(n9828), .a(n6966), .b(n7520) );
bf01f01  g6606 ( .o(n9833), .a(net_7135) );
bf01f01  g6607 ( .o(n9837), .a(net_7122) );
bf01f01  g6608 ( .o(n9840), .a(net_6396) );
bf01f01  g6609 ( .o(n9844), .a(net_6387) );
no02f01  g6610 ( .o(n9853), .a(n6966), .b(n10317) );
bf01f01  g6611 ( .o(n9867), .a(_net_7811) );
bf01f01  g6612 ( .o(n9871), .a(_net_7797) );
bf01f01  g6613 ( .o(n9875), .a(_net_7806) );
bf01f01  g6614 ( .o(n9885), .a(net_7109) );
bf01f01  g6615 ( .o(n9899), .a(net_6752) );
bf01f01  g6616 ( .o(n9902), .a(_net_7798) );
bf01f01  g6617 ( .o(n9911), .a(net_6446) );
bf01f01  g6618 ( .o(n9914), .a(_net_7819) );
bf01f01  g6619 ( .o(n9918), .a(x1580) );
bf01f01  g6620 ( .o(n9923), .a(net_6719) );
bf01f01  g6621 ( .o(n9926), .a(net_6389) );
bf01f01  g6622 ( .o(n9930), .a(net_6393) );
bf01f01  g6623 ( .o(n9935), .a(net_6465) );
bf01f01  g6624 ( .o(n9944), .a(_net_6174) );
in01f01  g6625 ( .o(n9953), .a(n7343) );
bf01f01  g6626 ( .o(n9957), .a(net_6389) );
bf01f01  g6627 ( .o(n9961), .a(_net_7804) );
bf01f01  g6628 ( .o(n9976), .a(net_6057) );
bf01f01  g6629 ( .o(n9985), .a(net_6380) );
bf01f01  g6630 ( .o(n9988), .a(_net_7805) );
bf01f01  g6631 ( .o(n9992), .a(_net_7805) );
bf01f01  g6632 ( .o(n10001), .a(_net_7812) );
bf01f01  g6633 ( .o(n10006), .a(_net_6062) );
bf01f01  g6634 ( .o(n10010), .a(net_7802) );
bf01f01  g6635 ( .o(n10014), .a(x1351) );
bf01f01  g6636 ( .o(n10023), .a(net_130) );
bf01f01  g6637 ( .o(n10028), .a(net_6879) );
bf01f01  g6638 ( .o(n10047), .a(_net_6155) );
no02f01  g6639 ( .o(n10056), .a(n6966), .b(n7250) );
bf01f01  g6640 ( .o(n10070), .a(net_6884) );
bf01f01  g6641 ( .o(n10103), .a(_net_7815) );
bf01f01  g6642 ( .o(n10107), .a(_net_7818) );
bf01f01  g6643 ( .o(n10112), .a(net_7112) );
bf01f01  g6644 ( .o(n10120), .a(_net_7815) );
bf01f01  g6645 ( .o(n10124), .a(_net_7811) );
bf01f01  g6646 ( .o(n10132), .a(_net_7805) );
bf01f01  g6647 ( .o(n10141), .a(x1595) );
no02f01  g6648 ( .o(n10145), .a(n6899_1), .b(n7514) );
bf01f01  g6649 ( .o(n10154), .a(net_7807) );
bf01f01  g6650 ( .o(n10158), .a(_net_7806) );
ms00f80  l0001 ( .o(net_249), .ck(clk), .d(n266) );
ms00f80  l0002 ( .o(net_254), .ck(clk), .d(n271) );
ms00f80  l0003 ( .o(net_6907), .ck(clk), .d(n276) );
ms00f80  l0004 ( .o(_net_6082), .ck(clk), .d(n281) );
ms00f80  l0005 ( .o(net_6300), .ck(clk), .d(n286) );
ms00f80  l0006 ( .o(net_6453), .ck(clk), .d(n291) );
ms00f80  l0007 ( .o(_net_6032), .ck(clk), .d(n295) );
ms00f80  l0008 ( .o(_net_6133), .ck(clk), .d(n300) );
ms00f80  l0009 ( .o(net_7222), .ck(clk), .d(n305) );
ms00f80  l0010 ( .o(net_6704), .ck(clk), .d(n310) );
ms00f80  l0011 ( .o(_net_7481), .ck(clk), .d(n314) );
ms00f80  l0012 ( .o(_net_175), .ck(clk), .d(n319) );
ms00f80  l0013 ( .o(net_7204), .ck(clk), .d(n324) );
ms00f80  l0014 ( .o(_net_6062), .ck(clk), .d(n329) );
ms00f80  l0015 ( .o(net_6227), .ck(clk), .d(n334) );
ms00f80  l0016 ( .o(net_6364), .ck(clk), .d(n339) );
ms00f80  l0017 ( .o(net_6256), .ck(clk), .d(n344) );
ms00f80  l0018 ( .o(net_6474), .ck(clk), .d(n349) );
ms00f80  l0019 ( .o(_net_7800), .ck(clk), .d(n352) );
ms00f80  l0020 ( .o(net_7114), .ck(clk), .d(n357) );
ms00f80  l0021 ( .o(net_6784), .ck(clk), .d(n361) );
ms00f80  l0022 ( .o(net_6996), .ck(clk), .d(n366) );
ms00f80  l0023 ( .o(_net_7474), .ck(clk), .d(n370) );
ms00f80  l0024 ( .o(_net_7252), .ck(clk), .d(n375) );
ms00f80  l0025 ( .o(_net_298), .ck(clk), .d(n380) );
ms00f80  l0026 ( .o(_net_6404), .ck(clk), .d(n385) );
ms00f80  l0027 ( .o(_net_6088), .ck(clk), .d(n390) );
ms00f80  l0028 ( .o(net_7055), .ck(clk), .d(n395) );
ms00f80  l0029 ( .o(_net_7595), .ck(clk), .d(n400) );
ms00f80  l0030 ( .o(net_6396), .ck(clk), .d(n405) );
ms00f80  l0031 ( .o(net_6313), .ck(clk), .d(n410) );
ms00f80  l0032 ( .o(net_7062), .ck(clk), .d(n415) );
ms00f80  l0033 ( .o(net_7525), .ck(clk), .d(n420) );
ms00f80  l0034 ( .o(net_6514), .ck(clk), .d(n424) );
ms00f80  l0035 ( .o(net_6803), .ck(clk), .d(n429) );
ms00f80  l0036 ( .o(net_7713), .ck(clk), .d(n434) );
ms00f80  l0037 ( .o(net_6510), .ck(clk), .d(n438) );
ms00f80  l0038 ( .o(net_7000), .ck(clk), .d(n443) );
ms00f80  l0039 ( .o(_net_6150), .ck(clk), .d(n447) );
ms00f80  l0040 ( .o(net_7802), .ck(clk), .d(n451) );
ms00f80  l0041 ( .o(net_6628), .ck(clk), .d(n455) );
ms00f80  l0042 ( .o(_net_7355), .ck(clk), .d(n460) );
ms00f80  l0043 ( .o(_net_6100), .ck(clk), .d(n465) );
ms00f80  l0044 ( .o(net_7388), .ck(clk), .d(n470) );
ms00f80  l0045 ( .o(net_362), .ck(clk), .d(n474) );
ms00f80  l0046 ( .o(net_6783), .ck(clk), .d(n479) );
ms00f80  l0047 ( .o(net_6870), .ck(clk), .d(n484) );
ms00f80  l0048 ( .o(net_7196), .ck(clk), .d(n488) );
ms00f80  l0049 ( .o(net_7224), .ck(clk), .d(n493) );
ms00f80  l0050 ( .o(_net_6194), .ck(clk), .d(n498) );
ms00f80  l0051 ( .o(net_6267), .ck(clk), .d(n503) );
ms00f80  l0052 ( .o(net_6308), .ck(clk), .d(n508) );
ms00f80  l0053 ( .o(net_6691), .ck(clk), .d(n513) );
ms00f80  l0054 ( .o(net_7369), .ck(clk), .d(n518) );
ms00f80  l0055 ( .o(_net_6079), .ck(clk), .d(n523) );
ms00f80  l0056 ( .o(_net_7689), .ck(clk), .d(n528) );
ms00f80  l0057 ( .o(_net_6104), .ck(clk), .d(n533) );
ms00f80  l0058 ( .o(_net_7603), .ck(clk), .d(n538) );
ms00f80  l0059 ( .o(_net_7316), .ck(clk), .d(n543) );
ms00f80  l0060 ( .o(_net_5965), .ck(clk), .d(n548) );
ms00f80  l0061 ( .o(x14), .ck(clk), .d(n553) );
ms00f80  l0062 ( .o(net_6791), .ck(clk), .d(n556) );
ms00f80  l0063 ( .o(_net_6294), .ck(clk), .d(n561) );
ms00f80  l0064 ( .o(net_6773), .ck(clk), .d(n566) );
ms00f80  l0065 ( .o(net_6218), .ck(clk), .d(n571) );
ms00f80  l0066 ( .o(net_7342), .ck(clk), .d(n576) );
ms00f80  l0067 ( .o(_net_7794), .ck(clk), .d(n580) );
ms00f80  l0068 ( .o(net_6373), .ck(clk), .d(n585) );
ms00f80  l0069 ( .o(net_365), .ck(clk), .d(n590) );
ms00f80  l0070 ( .o(net_7492), .ck(clk), .d(n595) );
ms00f80  l0071 ( .o(_net_7285), .ck(clk), .d(n600) );
ms00f80  l0072 ( .o(_net_6210), .ck(clk), .d(n605) );
ms00f80  l0073 ( .o(net_6900), .ck(clk), .d(n610) );
ms00f80  l0074 ( .o(net_7604), .ck(clk), .d(n615) );
ms00f80  l0075 ( .o(_net_6004), .ck(clk), .d(n620) );
ms00f80  l0076 ( .o(net_7246), .ck(clk), .d(n625) );
ms00f80  l0077 ( .o(_net_7441), .ck(clk), .d(n629) );
ms00f80  l0078 ( .o(net_7487), .ck(clk), .d(n634) );
ms00f80  l0079 ( .o(_net_7694), .ck(clk), .d(n639) );
ms00f80  l0080 ( .o(_net_7094), .ck(clk), .d(n644) );
ms00f80  l0081 ( .o(_net_212), .ck(clk), .d(n649) );
ms00f80  l0082 ( .o(_net_7753), .ck(clk), .d(n654) );
ms00f80  l0083 ( .o(net_160), .ck(clk), .d(n659) );
ms00f80  l0084 ( .o(net_6384), .ck(clk), .d(n664) );
ms00f80  l0085 ( .o(net_6440), .ck(clk), .d(n669) );
ms00f80  l0086 ( .o(_net_6208), .ck(clk), .d(n673) );
ms00f80  l0087 ( .o(net_6653), .ck(clk), .d(n678) );
ms00f80  l0088 ( .o(net_6491), .ck(clk), .d(n683) );
ms00f80  l0089 ( .o(_net_7330), .ck(clk), .d(n688) );
ms00f80  l0090 ( .o(_net_7271), .ck(clk), .d(n693) );
ms00f80  l0091 ( .o(net_7645), .ck(clk), .d(n698) );
ms00f80  l0092 ( .o(net_6323), .ck(clk), .d(n703) );
ms00f80  l0093 ( .o(_net_7300), .ck(clk), .d(n708) );
ms00f80  l0094 ( .o(net_7774), .ck(clk), .d(n713) );
ms00f80  l0095 ( .o(net_7637), .ck(clk), .d(n718) );
ms00f80  l0096 ( .o(net_361), .ck(clk), .d(n722) );
ms00f80  l0097 ( .o(net_236), .ck(clk), .d(n727) );
ms00f80  l0098 ( .o(x561), .ck(clk), .d(n732) );
ms00f80  l0099 ( .o(_net_6037), .ck(clk), .d(n736) );
ms00f80  l0100 ( .o(net_6213), .ck(clk), .d(n741) );
ms00f80  l0101 ( .o(net_235), .ck(clk), .d(n746) );
ms00f80  l0102 ( .o(net_7758), .ck(clk), .d(n751) );
ms00f80  l0103 ( .o(_net_6147), .ck(clk), .d(n756) );
ms00f80  l0104 ( .o(net_6468), .ck(clk), .d(n761) );
ms00f80  l0105 ( .o(_net_113), .ck(clk), .d(n765) );
ms00f80  l0106 ( .o(_net_7732), .ck(clk), .d(n770) );
ms00f80  l0107 ( .o(net_6380), .ck(clk), .d(n774) );
ms00f80  l0108 ( .o(net_6386), .ck(clk), .d(n779) );
ms00f80  l0109 ( .o(net_139), .ck(clk), .d(n783) );
ms00f80  l0110 ( .o(_net_6012), .ck(clk), .d(n788) );
ms00f80  l0111 ( .o(net_7607), .ck(clk), .d(n793) );
ms00f80  l0112 ( .o(net_7134), .ck(clk), .d(n798) );
ms00f80  l0113 ( .o(net_7133), .ck(clk), .d(n802) );
ms00f80  l0114 ( .o(_net_7786), .ck(clk), .d(n806) );
ms00f80  l0115 ( .o(net_6400), .ck(clk), .d(n811) );
ms00f80  l0116 ( .o(net_6260), .ck(clk), .d(n815) );
ms00f80  l0117 ( .o(_net_121), .ck(clk), .d(n820) );
ms00f80  l0118 ( .o(_net_120), .ck(clk), .d(n825) );
ms00f80  l0119 ( .o(net_7396), .ck(clk), .d(n830) );
ms00f80  l0120 ( .o(net_220), .ck(clk), .d(n834) );
ms00f80  l0121 ( .o(net_6545), .ck(clk), .d(n839) );
ms00f80  l0122 ( .o(net_326), .ck(clk), .d(n844) );
ms00f80  l0123 ( .o(net_171), .ck(clk), .d(n849) );
ms00f80  l0124 ( .o(net_7390), .ck(clk), .d(n854) );
ms00f80  l0125 ( .o(net_6521), .ck(clk), .d(n857) );
ms00f80  l0126 ( .o(_net_6086), .ck(clk), .d(n862) );
ms00f80  l0127 ( .o(net_6711), .ck(clk), .d(n867) );
ms00f80  l0128 ( .o(net_6815), .ck(clk), .d(n870) );
ms00f80  l0129 ( .o(net_7312), .ck(clk), .d(n875) );
ms00f80  l0130 ( .o(net_6646), .ck(clk), .d(n880) );
ms00f80  l0131 ( .o(_net_6008), .ck(clk), .d(n885) );
ms00f80  l0132 ( .o(net_6616), .ck(clk), .d(n890) );
ms00f80  l0133 ( .o(net_347), .ck(clk), .d(n894) );
ms00f80  l0134 ( .o(net_6739), .ck(clk), .d(n899) );
ms00f80  l0135 ( .o(_net_7439), .ck(clk), .d(n903) );
ms00f80  l0136 ( .o(net_7067), .ck(clk), .d(n907) );
ms00f80  l0137 ( .o(net_7073), .ck(clk), .d(n911) );
ms00f80  l0138 ( .o(net_6746), .ck(clk), .d(n916) );
ms00f80  l0139 ( .o(net_6356), .ck(clk), .d(n920) );
ms00f80  l0140 ( .o(_net_7354), .ck(clk), .d(n925) );
ms00f80  l0141 ( .o(_net_7632), .ck(clk), .d(n930) );
ms00f80  l0142 ( .o(net_7066), .ck(clk), .d(n935) );
ms00f80  l0143 ( .o(net_6979), .ck(clk), .d(n940) );
ms00f80  l0144 ( .o(_net_5851), .ck(clk), .d(n944) );
ms00f80  l0145 ( .o(_net_7809), .ck(clk), .d(n948) );
ms00f80  l0146 ( .o(net_6989), .ck(clk), .d(n953) );
ms00f80  l0147 ( .o(net_7058), .ck(clk), .d(n956) );
ms00f80  l0148 ( .o(_net_7629), .ck(clk), .d(n961) );
ms00f80  l0149 ( .o(net_204), .ck(clk), .d(n966) );
ms00f80  l0150 ( .o(_net_7296), .ck(clk), .d(n971) );
ms00f80  l0151 ( .o(net_150), .ck(clk), .d(n976) );
ms00f80  l0152 ( .o(net_6999), .ck(clk), .d(n981) );
ms00f80  l0153 ( .o(_net_282), .ck(clk), .d(n985) );
ms00f80  l0154 ( .o(_net_7653), .ck(clk), .d(n990) );
ms00f80  l0155 ( .o(_net_5856), .ck(clk), .d(n995) );
ms00f80  l0156 ( .o(net_391), .ck(clk), .d(n1000) );
ms00f80  l0157 ( .o(net_6392), .ck(clk), .d(n1005) );
ms00f80  l0158 ( .o(_net_7621), .ck(clk), .d(n1010) );
ms00f80  l0159 ( .o(_net_6120), .ck(clk), .d(n1015) );
ms00f80  l0160 ( .o(net_6998), .ck(clk), .d(n1020) );
ms00f80  l0161 ( .o(_net_7447), .ck(clk), .d(n1024) );
ms00f80  l0162 ( .o(net_7334), .ck(clk), .d(n1029) );
ms00f80  l0163 ( .o(net_7311), .ck(clk), .d(n1034) );
ms00f80  l0164 ( .o(_net_6220), .ck(clk), .d(n1039) );
ms00f80  l0165 ( .o(_net_7281), .ck(clk), .d(n1044) );
ms00f80  l0166 ( .o(_net_7578), .ck(clk), .d(n1049) );
ms00f80  l0167 ( .o(net_351), .ck(clk), .d(n1053) );
ms00f80  l0168 ( .o(x657), .ck(clk), .d(n1058) );
ms00f80  l0169 ( .o(net_6944), .ck(clk), .d(n1062) );
ms00f80  l0170 ( .o(net_5992), .ck(clk), .d(n1067) );
ms00f80  l0171 ( .o(_net_6286), .ck(clk), .d(n1072) );
ms00f80  l0172 ( .o(net_7004), .ck(clk), .d(n1077) );
ms00f80  l0173 ( .o(net_7010), .ck(clk), .d(n1081) );
ms00f80  l0174 ( .o(net_6461), .ck(clk), .d(n1085) );
ms00f80  l0175 ( .o(net_6832), .ck(clk), .d(n1089) );
ms00f80  l0176 ( .o(net_6977), .ck(clk), .d(n1093) );
ms00f80  l0177 ( .o(net_6901), .ck(clk), .d(n1097) );
ms00f80  l0178 ( .o(net_6856), .ck(clk), .d(n1102) );
ms00f80  l0179 ( .o(_net_7412), .ck(clk), .d(n1106) );
ms00f80  l0180 ( .o(net_6379), .ck(clk), .d(n1111) );
ms00f80  l0181 ( .o(net_6060), .ck(clk), .d(n1116) );
ms00f80  l0182 ( .o(net_6847), .ck(clk), .d(n1121) );
ms00f80  l0183 ( .o(_net_7274), .ck(clk), .d(n1125) );
ms00f80  l0184 ( .o(net_6671), .ck(clk), .d(n1130) );
ms00f80  l0185 ( .o(_net_7299), .ck(clk), .d(n1135) );
ms00f80  l0186 ( .o(net_6986), .ck(clk), .d(n1140) );
ms00f80  l0187 ( .o(net_6275), .ck(clk), .d(n1144) );
ms00f80  l0188 ( .o(net_6677), .ck(clk), .d(n1148) );
ms00f80  l0189 ( .o(_net_6167), .ck(clk), .d(n1153) );
ms00f80  l0190 ( .o(net_6242), .ck(clk), .d(n1158) );
ms00f80  l0191 ( .o(net_7611), .ck(clk), .d(n1163) );
ms00f80  l0192 ( .o(net_363), .ck(clk), .d(n1168) );
ms00f80  l0193 ( .o(net_7523), .ck(clk), .d(n1173) );
ms00f80  l0194 ( .o(_net_6135), .ck(clk), .d(n1178) );
ms00f80  l0195 ( .o(net_6238), .ck(clk), .d(n1183) );
ms00f80  l0196 ( .o(net_345), .ck(clk), .d(n1187) );
ms00f80  l0197 ( .o(net_6788), .ck(clk), .d(n1191) );
ms00f80  l0198 ( .o(net_6922), .ck(clk), .d(n1195) );
ms00f80  l0199 ( .o(net_6240), .ck(clk), .d(n1200) );
ms00f80  l0200 ( .o(net_7081), .ck(clk), .d(n1205) );
ms00f80  l0201 ( .o(net_6845), .ck(clk), .d(n1210) );
ms00f80  l0202 ( .o(_net_7503), .ck(clk), .d(n1214) );
ms00f80  l0203 ( .o(_net_7428), .ck(clk), .d(n1219) );
ms00f80  l0204 ( .o(net_6608), .ck(clk), .d(n1224) );
ms00f80  l0205 ( .o(_net_7730), .ck(clk), .d(n1228) );
ms00f80  l0206 ( .o(net_132), .ck(clk), .d(n1232) );
ms00f80  l0207 ( .o(net_7675), .ck(clk), .d(n1236) );
ms00f80  l0208 ( .o(net_6952), .ck(clk), .d(n1240) );
ms00f80  l0209 ( .o(net_360), .ck(clk), .d(n1244) );
ms00f80  l0210 ( .o(net_6759), .ck(clk), .d(n1248) );
ms00f80  l0211 ( .o(_net_7512), .ck(clk), .d(n1253) );
ms00f80  l0212 ( .o(net_7019), .ck(clk), .d(n1258) );
ms00f80  l0213 ( .o(net_6354), .ck(clk), .d(n1262) );
ms00f80  l0214 ( .o(_net_7590), .ck(clk), .d(n1267) );
ms00f80  l0215 ( .o(_net_273), .ck(clk), .d(n1272) );
ms00f80  l0216 ( .o(net_7453), .ck(clk), .d(n1277) );
ms00f80  l0217 ( .o(_net_299), .ck(clk), .d(n1282) );
ms00f80  l0218 ( .o(net_7119), .ck(clk), .d(n1287) );
ms00f80  l0219 ( .o(net_6574), .ck(clk), .d(n1291) );
ms00f80  l0220 ( .o(_net_7315), .ck(clk), .d(n1295) );
ms00f80  l0221 ( .o(net_7070), .ck(clk), .d(n1300) );
ms00f80  l0222 ( .o(net_7395), .ck(clk), .d(n1305) );
ms00f80  l0223 ( .o(_net_5966), .ck(clk), .d(n1309) );
ms00f80  l0224 ( .o(_net_6000), .ck(clk), .d(n1314) );
ms00f80  l0225 ( .o(net_7182), .ck(clk), .d(n1318) );
ms00f80  l0226 ( .o(net_7200), .ck(clk), .d(n1322) );
ms00f80  l0227 ( .o(net_6515), .ck(clk), .d(n1326) );
ms00f80  l0228 ( .o(net_6859), .ck(clk), .d(n1331) );
ms00f80  l0229 ( .o(_net_5991), .ck(clk), .d(n1335) );
ms00f80  l0230 ( .o(_net_7707), .ck(clk), .d(n1340) );
ms00f80  l0231 ( .o(net_6961), .ck(clk), .d(n1345) );
ms00f80  l0232 ( .o(net_7303), .ck(clk), .d(n1350) );
ms00f80  l0233 ( .o(net_6877), .ck(clk), .d(n1355) );
ms00f80  l0234 ( .o(net_7234), .ck(clk), .d(n1359) );
ms00f80  l0235 ( .o(_net_213), .ck(clk), .d(n1363) );
ms00f80  l0236 ( .o(net_6025), .ck(clk), .d(n1368) );
ms00f80  l0237 ( .o(_net_5997), .ck(clk), .d(n1373) );
ms00f80  l0238 ( .o(net_7750), .ck(clk), .d(n1378) );
ms00f80  l0239 ( .o(net_6694), .ck(clk), .d(n1383) );
ms00f80  l0240 ( .o(net_325), .ck(clk), .d(n1386) );
ms00f80  l0241 ( .o(_net_7658), .ck(clk), .d(n1391) );
ms00f80  l0242 ( .o(net_6190), .ck(clk), .d(n1396) );
ms00f80  l0243 ( .o(net_6624), .ck(clk), .d(n1400) );
ms00f80  l0244 ( .o(_net_6182), .ck(clk), .d(n1405) );
ms00f80  l0245 ( .o(_net_5960), .ck(clk), .d(n1410) );
ms00f80  l0246 ( .o(net_7217), .ck(clk), .d(n1414) );
ms00f80  l0247 ( .o(_net_7253), .ck(clk), .d(n1419) );
ms00f80  l0248 ( .o(net_6941), .ck(clk), .d(n1423) );
ms00f80  l0249 ( .o(_net_7497), .ck(clk), .d(n1428) );
ms00f80  l0250 ( .o(_net_7768), .ck(clk), .d(n1433) );
ms00f80  l0251 ( .o(net_6745), .ck(clk), .d(n1438) );
ms00f80  l0252 ( .o(_net_7565), .ck(clk), .d(n1442) );
ms00f80  l0253 ( .o(net_6913), .ck(clk), .d(n1446) );
ms00f80  l0254 ( .o(_net_6044), .ck(clk), .d(n1451) );
ms00f80  l0255 ( .o(net_6633), .ck(clk), .d(n1455) );
ms00f80  l0256 ( .o(net_6328), .ck(clk), .d(n1460) );
ms00f80  l0257 ( .o(net_6953), .ck(clk), .d(n1465) );
ms00f80  l0258 ( .o(net_357), .ck(clk), .d(n1469) );
ms00f80  l0259 ( .o(net_6612), .ck(clk), .d(n1474) );
ms00f80  l0260 ( .o(net_6302), .ck(clk), .d(n1478) );
ms00f80  l0261 ( .o(_net_7815), .ck(clk), .d(n1482) );
ms00f80  l0262 ( .o(_net_7746), .ck(clk), .d(n1487) );
ms00f80  l0263 ( .o(net_6768), .ck(clk), .d(n1491) );
ms00f80  l0264 ( .o(net_6059), .ck(clk), .d(n1496) );
ms00f80  l0265 ( .o(_net_7698), .ck(clk), .d(n1501) );
ms00f80  l0266 ( .o(net_7550), .ck(clk), .d(n1506) );
ms00f80  l0267 ( .o(net_7091), .ck(clk), .d(n1510) );
ms00f80  l0268 ( .o(net_6619), .ck(clk), .d(n1515) );
ms00f80  l0269 ( .o(_net_6095), .ck(clk), .d(n1519) );
ms00f80  l0270 ( .o(net_7106), .ck(clk), .d(n1524) );
ms00f80  l0271 ( .o(net_6375), .ck(clk), .d(n1528) );
ms00f80  l0272 ( .o(net_203), .ck(clk), .d(n1533) );
ms00f80  l0273 ( .o(net_7247), .ck(clk), .d(n1538) );
ms00f80  l0274 ( .o(x287), .ck(clk), .d(n1542) );
ms00f80  l0275 ( .o(_net_7534), .ck(clk), .d(n1546) );
ms00f80  l0276 ( .o(net_7146), .ck(clk), .d(n1551) );
ms00f80  l0277 ( .o(_net_7406), .ck(clk), .d(n1555) );
ms00f80  l0278 ( .o(net_7126), .ck(clk), .d(n1560) );
ms00f80  l0279 ( .o(net_6482), .ck(clk), .d(n1564) );
ms00f80  l0280 ( .o(net_6888), .ck(clk), .d(n1568) );
ms00f80  l0281 ( .o(net_258), .ck(clk), .d(n1572) );
ms00f80  l0282 ( .o(net_353), .ck(clk), .d(n1577) );
ms00f80  l0283 ( .o(_net_7535), .ck(clk), .d(n1582) );
ms00f80  l0284 ( .o(net_6584), .ck(clk), .d(n1587) );
ms00f80  l0285 ( .o(net_352), .ck(clk), .d(n1591) );
ms00f80  l0286 ( .o(net_6732), .ck(clk), .d(n1596) );
ms00f80  l0287 ( .o(_net_7759), .ck(clk), .d(n1600) );
ms00f80  l0288 ( .o(net_165), .ck(clk), .d(n1605) );
ms00f80  l0289 ( .o(_net_7498), .ck(clk), .d(n1610) );
ms00f80  l0290 ( .o(net_6914), .ck(clk), .d(n1615) );
ms00f80  l0291 ( .o(net_7198), .ck(clk), .d(n1619) );
ms00f80  l0292 ( .o(_net_7696), .ck(clk), .d(n1624) );
ms00f80  l0293 ( .o(net_6537), .ck(clk), .d(n1629) );
ms00f80  l0294 ( .o(_net_7570), .ck(clk), .d(n1634) );
ms00f80  l0295 ( .o(net_7308), .ck(clk), .d(n1639) );
ms00f80  l0296 ( .o(net_260), .ck(clk), .d(n1644) );
ms00f80  l0297 ( .o(net_7124), .ck(clk), .d(n1649) );
ms00f80  l0298 ( .o(net_6229), .ck(clk), .d(n1653) );
ms00f80  l0299 ( .o(net_245), .ck(clk), .d(n1658) );
ms00f80  l0300 ( .o(net_6197), .ck(clk), .d(n1663) );
ms00f80  l0301 ( .o(net_7760), .ck(clk), .d(n1668) );
ms00f80  l0302 ( .o(net_6723), .ck(clk), .d(n1673) );
ms00f80  l0303 ( .o(_net_6042), .ck(clk), .d(n1677) );
ms00f80  l0304 ( .o(net_6654), .ck(clk), .d(n1681) );
ms00f80  l0305 ( .o(net_6512), .ck(clk), .d(n1686) );
ms00f80  l0306 ( .o(net_6770), .ck(clk), .d(n1691) );
ms00f80  l0307 ( .o(_net_6168), .ck(clk), .d(n1696) );
ms00f80  l0308 ( .o(net_6432), .ck(clk), .d(n1701) );
ms00f80  l0309 ( .o(net_6500), .ck(clk), .d(n1704) );
ms00f80  l0310 ( .o(net_7170), .ck(clk), .d(n1709) );
ms00f80  l0311 ( .o(_net_7358), .ck(clk), .d(n1714) );
ms00f80  l0312 ( .o(net_6903), .ck(clk), .d(n1718) );
ms00f80  l0313 ( .o(net_7220), .ck(clk), .d(n1722) );
ms00f80  l0314 ( .o(_net_6180), .ck(clk), .d(n1727) );
ms00f80  l0315 ( .o(net_6806), .ck(clk), .d(n1732) );
ms00f80  l0316 ( .o(_net_7468), .ck(clk), .d(n1737) );
ms00f80  l0317 ( .o(_net_5996), .ck(clk), .d(n1742) );
ms00f80  l0318 ( .o(_net_6077), .ck(clk), .d(n1747) );
ms00f80  l0319 ( .o(net_7495), .ck(clk), .d(n1752) );
ms00f80  l0320 ( .o(net_6896), .ck(clk), .d(n1756) );
ms00f80  l0321 ( .o(net_6570), .ck(clk), .d(n1761) );
ms00f80  l0322 ( .o(net_7223), .ck(clk), .d(n1765) );
ms00f80  l0323 ( .o(_net_5985), .ck(clk), .d(n1770) );
ms00f80  l0324 ( .o(net_6602), .ck(clk), .d(n1775) );
ms00f80  l0325 ( .o(net_7551), .ck(clk), .d(n1779) );
ms00f80  l0326 ( .o(net_7035), .ck(clk), .d(n1782) );
ms00f80  l0327 ( .o(_net_6296), .ck(clk), .d(n1787) );
ms00f80  l0328 ( .o(net_7742), .ck(clk), .d(n1792) );
ms00f80  l0329 ( .o(net_6316), .ck(clk), .d(n1797) );
ms00f80  l0330 ( .o(_net_6185), .ck(clk), .d(n1802) );
ms00f80  l0331 ( .o(_net_7328), .ck(clk), .d(n1807) );
ms00f80  l0332 ( .o(_net_7359), .ck(clk), .d(n1812) );
ms00f80  l0333 ( .o(net_6371), .ck(clk), .d(n1817) );
ms00f80  l0334 ( .o(net_6269), .ck(clk), .d(n1822) );
ms00f80  l0335 ( .o(net_6248), .ck(clk), .d(n1827) );
ms00f80  l0336 ( .o(_net_7650), .ck(clk), .d(n1832) );
ms00f80  l0337 ( .o(_net_7813), .ck(clk), .d(n1836) );
ms00f80  l0338 ( .o(_net_6087), .ck(clk), .d(n1841) );
ms00f80  l0339 ( .o(_net_6292), .ck(clk), .d(n1846) );
ms00f80  l0340 ( .o(net_6223), .ck(clk), .d(n1851) );
ms00f80  l0341 ( .o(_net_7819), .ck(clk), .d(n1855) );
ms00f80  l0342 ( .o(net_7767), .ck(clk), .d(n1860) );
ms00f80  l0343 ( .o(net_6699), .ck(clk), .d(n1865) );
ms00f80  l0344 ( .o(_net_7255), .ck(clk), .d(n1869) );
ms00f80  l0345 ( .o(net_6599), .ck(clk), .d(n1874) );
ms00f80  l0346 ( .o(_net_7600), .ck(clk), .d(n1878) );
ms00f80  l0347 ( .o(_net_6067), .ck(clk), .d(n1883) );
ms00f80  l0348 ( .o(_net_7628), .ck(clk), .d(n1888) );
ms00f80  l0349 ( .o(_net_6155), .ck(clk), .d(n1893) );
ms00f80  l0350 ( .o(net_6053), .ck(clk), .d(n1898) );
ms00f80  l0351 ( .o(net_6258), .ck(clk), .d(n1903) );
ms00f80  l0352 ( .o(_net_7379), .ck(clk), .d(n1908) );
ms00f80  l0353 ( .o(net_6543), .ck(clk), .d(n1913) );
ms00f80  l0354 ( .o(net_7116), .ck(clk), .d(n1918) );
ms00f80  l0355 ( .o(_net_6070), .ck(clk), .d(n1922) );
ms00f80  l0356 ( .o(_net_6690), .ck(clk), .d(n1927) );
ms00f80  l0357 ( .o(net_6995), .ck(clk), .d(n1932) );
ms00f80  l0358 ( .o(net_241), .ck(clk), .d(n1936) );
ms00f80  l0359 ( .o(net_6433), .ck(clk), .d(n1941) );
ms00f80  l0360 ( .o(_net_7472), .ck(clk), .d(n1945) );
ms00f80  l0361 ( .o(_net_7532), .ck(clk), .d(n1950) );
ms00f80  l0362 ( .o(net_7052), .ck(clk), .d(n1954) );
ms00f80  l0363 ( .o(_net_129), .ck(clk), .d(n1959) );
ms00f80  l0364 ( .o(net_6346), .ck(clk), .d(n1964) );
ms00f80  l0365 ( .o(_net_7594), .ck(clk), .d(n1969) );
ms00f80  l0366 ( .o(net_6800), .ck(clk), .d(n1973) );
ms00f80  l0367 ( .o(net_7174), .ck(clk), .d(n1978) );
ms00f80  l0368 ( .o(net_6274), .ck(clk), .d(n1983) );
ms00f80  l0369 ( .o(_net_6108), .ck(clk), .d(n1988) );
ms00f80  l0370 ( .o(net_7520), .ck(clk), .d(n1993) );
ms00f80  l0371 ( .o(net_6737), .ck(clk), .d(n1998) );
ms00f80  l0372 ( .o(net_6303), .ck(clk), .d(n2002) );
ms00f80  l0373 ( .o(net_6812), .ck(clk), .d(n2007) );
ms00f80  l0374 ( .o(net_7188), .ck(clk), .d(n2011) );
ms00f80  l0375 ( .o(_net_7426), .ck(clk), .d(n2016) );
ms00f80  l0376 ( .o(net_7790), .ck(clk), .d(n2021) );
ms00f80  l0377 ( .o(_net_6107), .ck(clk), .d(n2026) );
ms00f80  l0378 ( .o(net_6318), .ck(clk), .d(n2031) );
ms00f80  l0379 ( .o(net_319), .ck(clk), .d(n2036) );
ms00f80  l0380 ( .o(_net_7483), .ck(clk), .d(n2041) );
ms00f80  l0381 ( .o(_net_7093), .ck(clk), .d(n2046) );
ms00f80  l0382 ( .o(net_7391), .ck(clk), .d(n2051) );
ms00f80  l0383 ( .o(_net_7465), .ck(clk), .d(n2055) );
ms00f80  l0384 ( .o(_net_7352), .ck(clk), .d(n2060) );
ms00f80  l0385 ( .o(_net_6125), .ck(clk), .d(n2065) );
ms00f80  l0386 ( .o(_net_6827), .ck(clk), .d(n2070) );
ms00f80  l0387 ( .o(net_7201), .ck(clk), .d(n2074) );
ms00f80  l0388 ( .o(net_7754), .ck(clk), .d(n2079) );
ms00f80  l0389 ( .o(net_7371), .ck(clk), .d(n2084) );
ms00f80  l0390 ( .o(net_7063), .ck(clk), .d(n2088) );
ms00f80  l0391 ( .o(net_6893), .ck(clk), .d(n2093) );
ms00f80  l0392 ( .o(net_6709), .ck(clk), .d(n2098) );
ms00f80  l0393 ( .o(net_6741), .ck(clk), .d(n2102) );
ms00f80  l0394 ( .o(net_6191), .ck(clk), .d(n2106) );
ms00f80  l0395 ( .o(net_7003), .ck(clk), .d(n2111) );
ms00f80  l0396 ( .o(net_6452), .ck(clk), .d(n2115) );
ms00f80  l0397 ( .o(net_6603), .ck(clk), .d(n2119) );
ms00f80  l0398 ( .o(net_7076), .ck(clk), .d(n2122) );
ms00f80  l0399 ( .o(net_6310), .ck(clk), .d(n2127) );
ms00f80  l0400 ( .o(net_7147), .ck(clk), .d(n2132) );
ms00f80  l0401 ( .o(net_6730), .ck(clk), .d(n2136) );
ms00f80  l0402 ( .o(_net_7683), .ck(clk), .d(n2140) );
ms00f80  l0403 ( .o(net_7179), .ck(clk), .d(n2144) );
ms00f80  l0404 ( .o(net_7144), .ck(clk), .d(n2149) );
ms00f80  l0405 ( .o(net_7613), .ck(clk), .d(n2152) );
ms00f80  l0406 ( .o(net_6336), .ck(clk), .d(n2157) );
ms00f80  l0407 ( .o(_net_7554), .ck(clk), .d(n2162) );
ms00f80  l0408 ( .o(_net_7649), .ck(clk), .d(n2167) );
ms00f80  l0409 ( .o(_net_6963), .ck(clk), .d(n2172) );
ms00f80  l0410 ( .o(x397), .ck(clk), .d(n2177) );
ms00f80  l0411 ( .o(_net_7763), .ck(clk), .d(n2181) );
ms00f80  l0412 ( .o(net_6443), .ck(clk), .d(n2186) );
ms00f80  l0413 ( .o(net_6540), .ck(clk), .d(n2189) );
ms00f80  l0414 ( .o(_net_6177), .ck(clk), .d(n2194) );
ms00f80  l0415 ( .o(_net_7229), .ck(clk), .d(n2199) );
ms00f80  l0416 ( .o(net_6658), .ck(clk), .d(n2203) );
ms00f80  l0417 ( .o(_net_5963), .ck(clk), .d(n2208) );
ms00f80  l0418 ( .o(_net_6016), .ck(clk), .d(n2213) );
ms00f80  l0419 ( .o(net_6456), .ck(clk), .d(n2218) );
ms00f80  l0420 ( .o(net_6556), .ck(clk), .d(n2222) );
ms00f80  l0421 ( .o(_net_6960), .ck(clk), .d(n2227) );
ms00f80  l0422 ( .o(_net_263), .ck(clk), .d(n2232) );
ms00f80  l0423 ( .o(_net_6184), .ck(clk), .d(n2237) );
ms00f80  l0424 ( .o(_net_7724), .ck(clk), .d(n2242) );
ms00f80  l0425 ( .o(x494), .ck(clk), .d(n2247) );
ms00f80  l0426 ( .o(_net_6401), .ck(clk), .d(n2251) );
ms00f80  l0427 ( .o(net_7458), .ck(clk), .d(n2256) );
ms00f80  l0428 ( .o(net_7671), .ck(clk), .d(n2260) );
ms00f80  l0429 ( .o(_net_7401), .ck(clk), .d(n2265) );
ms00f80  l0430 ( .o(_net_5977), .ck(clk), .d(n2270) );
ms00f80  l0431 ( .o(_net_6139), .ck(clk), .d(n2275) );
ms00f80  l0432 ( .o(_net_7748), .ck(clk), .d(n2280) );
ms00f80  l0433 ( .o(net_322), .ck(clk), .d(n2284) );
ms00f80  l0434 ( .o(net_142), .ck(clk), .d(n2288) );
ms00f80  l0435 ( .o(net_6366), .ck(clk), .d(n2293) );
ms00f80  l0436 ( .o(_net_6015), .ck(clk), .d(n2298) );
ms00f80  l0437 ( .o(_net_6187), .ck(clk), .d(n2303) );
ms00f80  l0438 ( .o(net_7194), .ck(clk), .d(n2307) );
ms00f80  l0439 ( .o(_net_7556), .ck(clk), .d(n2312) );
ms00f80  l0440 ( .o(net_6035), .ck(clk), .d(n2316) );
ms00f80  l0441 ( .o(net_7159), .ck(clk), .d(n2321) );
ms00f80  l0442 ( .o(net_323), .ck(clk), .d(n2324) );
ms00f80  l0443 ( .o(_net_6134), .ck(clk), .d(n2329) );
ms00f80  l0444 ( .o(_net_7747), .ck(clk), .d(n2334) );
ms00f80  l0445 ( .o(net_6920), .ck(clk), .d(n2338) );
ms00f80  l0446 ( .o(net_6501), .ck(clk), .d(n2342) );
ms00f80  l0447 ( .o(net_6849), .ck(clk), .d(n2347) );
ms00f80  l0448 ( .o(net_6236), .ck(clk), .d(n2350) );
ms00f80  l0449 ( .o(net_6277), .ck(clk), .d(n2355) );
ms00f80  l0450 ( .o(net_6912), .ck(clk), .d(n2360) );
ms00f80  l0451 ( .o(_net_6163), .ck(clk), .d(n2365) );
ms00f80  l0452 ( .o(net_6593), .ck(clk), .d(n2370) );
ms00f80  l0453 ( .o(net_6398), .ck(clk), .d(n2373) );
ms00f80  l0454 ( .o(_net_7720), .ck(clk), .d(n2377) );
ms00f80  l0455 ( .o(net_7527), .ck(clk), .d(n2381) );
ms00f80  l0456 ( .o(_net_6169), .ck(clk), .d(n2386) );
ms00f80  l0457 ( .o(net_6576), .ck(clk), .d(n2391) );
ms00f80  l0458 ( .o(net_183), .ck(clk), .d(n2395) );
ms00f80  l0459 ( .o(net_6758), .ck(clk), .d(n2399) );
ms00f80  l0460 ( .o(net_7608), .ck(clk), .d(n2404) );
ms00f80  l0461 ( .o(_net_7511), .ck(clk), .d(n2409) );
ms00f80  l0462 ( .o(x699), .ck(clk), .d(n2414) );
ms00f80  l0463 ( .o(net_6680), .ck(clk), .d(n2417) );
ms00f80  l0464 ( .o(net_7016), .ck(clk), .d(n2422) );
ms00f80  l0465 ( .o(net_6833), .ck(clk), .d(n2426) );
ms00f80  l0466 ( .o(_net_7431), .ck(clk), .d(n2430) );
ms00f80  l0467 ( .o(_net_279), .ck(clk), .d(n2435) );
ms00f80  l0468 ( .o(net_7240), .ck(clk), .d(n2440) );
ms00f80  l0469 ( .o(_net_5972), .ck(clk), .d(n2444) );
ms00f80  l0470 ( .o(net_377), .ck(clk), .d(n2448) );
ms00f80  l0471 ( .o(net_6821), .ck(clk), .d(n2452) );
ms00f80  l0472 ( .o(_net_5984), .ck(clk), .d(n2457) );
ms00f80  l0473 ( .o(net_6426), .ck(clk), .d(n2462) );
ms00f80  l0474 ( .o(net_6918), .ck(clk), .d(n2465) );
ms00f80  l0475 ( .o(_net_6118), .ck(clk), .d(n2470) );
ms00f80  l0476 ( .o(net_6672), .ck(clk), .d(n2474) );
ms00f80  l0477 ( .o(_net_7294), .ck(clk), .d(n2479) );
ms00f80  l0478 ( .o(net_224), .ck(clk), .d(n2484) );
ms00f80  l0479 ( .o(net_6764), .ck(clk), .d(n2488) );
ms00f80  l0480 ( .o(net_6435), .ck(clk), .d(n2493) );
ms00f80  l0481 ( .o(net_7207), .ck(clk), .d(n2496) );
ms00f80  l0482 ( .o(net_7639), .ck(clk), .d(n2500) );
ms00f80  l0483 ( .o(_net_7704), .ck(clk), .d(n2505) );
ms00f80  l0484 ( .o(net_252), .ck(clk), .d(n2510) );
ms00f80  l0485 ( .o(net_6014), .ck(clk), .d(n2515) );
ms00f80  l0486 ( .o(net_6522), .ck(clk), .d(n2519) );
ms00f80  l0487 ( .o(net_179), .ck(clk), .d(n2524) );
ms00f80  l0488 ( .o(_net_7419), .ck(clk), .d(n2529) );
ms00f80  l0489 ( .o(_net_6160), .ck(clk), .d(n2534) );
ms00f80  l0490 ( .o(net_134), .ck(clk), .d(n2539) );
ms00f80  l0491 ( .o(net_6939), .ck(clk), .d(n2543) );
ms00f80  l0492 ( .o(net_7337), .ck(clk), .d(n2547) );
ms00f80  l0493 ( .o(_net_7445), .ck(clk), .d(n2552) );
ms00f80  l0494 ( .o(net_6951), .ck(clk), .d(n2556) );
ms00f80  l0495 ( .o(net_300), .ck(clk), .d(n2561) );
ms00f80  l0496 ( .o(_net_7663), .ck(clk), .d(n2566) );
ms00f80  l0497 ( .o(net_6898), .ck(clk), .d(n2570) );
ms00f80  l0498 ( .o(_net_176), .ck(clk), .d(n2575) );
ms00f80  l0499 ( .o(net_207), .ck(clk), .d(n2580) );
ms00f80  l0500 ( .o(net_7779), .ck(clk), .d(n2585) );
ms00f80  l0501 ( .o(net_7096), .ck(clk), .d(n2590) );
ms00f80  l0502 ( .o(net_6391), .ck(clk), .d(n2594) );
ms00f80  l0503 ( .o(net_7032), .ck(clk), .d(n2597) );
ms00f80  l0504 ( .o(net_6517), .ck(clk), .d(n2601) );
ms00f80  l0505 ( .o(net_6513), .ck(clk), .d(n2605) );
ms00f80  l0506 ( .o(net_6377), .ck(clk), .d(n2610) );
ms00f80  l0507 ( .o(net_6967), .ck(clk), .d(n2615) );
ms00f80  l0508 ( .o(net_7060), .ck(clk), .d(n2618) );
ms00f80  l0509 ( .o(net_7089), .ck(clk), .d(n2622) );
ms00f80  l0510 ( .o(net_6322), .ck(clk), .d(n2627) );
ms00f80  l0511 ( .o(_net_7765), .ck(clk), .d(n2632) );
ms00f80  l0512 ( .o(net_257), .ck(clk), .d(n2637) );
ms00f80  l0513 ( .o(net_6341), .ck(clk), .d(n2642) );
ms00f80  l0514 ( .o(net_6588), .ck(clk), .d(n2647) );
ms00f80  l0515 ( .o(net_187), .ck(clk), .d(n2651) );
ms00f80  l0516 ( .o(net_6606), .ck(clk), .d(n2656) );
ms00f80  l0517 ( .o(net_6215), .ck(clk), .d(n2660) );
ms00f80  l0518 ( .o(_net_6121), .ck(clk), .d(n2665) );
ms00f80  l0519 ( .o(net_6330), .ck(clk), .d(n2670) );
ms00f80  l0520 ( .o(net_6890), .ck(clk), .d(n2675) );
ms00f80  l0521 ( .o(net_6964), .ck(clk), .d(n2679) );
ms00f80  l0522 ( .o(net_7057), .ck(clk), .d(n2682) );
ms00f80  l0523 ( .o(net_7777), .ck(clk), .d(n2687) );
ms00f80  l0524 ( .o(net_7393), .ck(clk), .d(n2692) );
ms00f80  l0525 ( .o(_net_6822), .ck(clk), .d(n2696) );
ms00f80  l0526 ( .o(net_6981), .ck(clk), .d(n2701) );
ms00f80  l0527 ( .o(net_6434), .ck(clk), .d(n2705) );
ms00f80  l0528 ( .o(net_6969), .ck(clk), .d(n2709) );
ms00f80  l0529 ( .o(_net_126), .ck(clk), .d(n2713) );
ms00f80  l0530 ( .o(net_238), .ck(clk), .d(n2718) );
ms00f80  l0531 ( .o(_net_280), .ck(clk), .d(n2723) );
ms00f80  l0532 ( .o(net_346), .ck(clk), .d(n2727) );
ms00f80  l0533 ( .o(_net_7314), .ck(clk), .d(n2732) );
ms00f80  l0534 ( .o(net_7708), .ck(clk), .d(n2737) );
ms00f80  l0535 ( .o(net_6586), .ck(clk), .d(n2741) );
ms00f80  l0536 ( .o(net_6725), .ck(clk), .d(n2745) );
ms00f80  l0537 ( .o(net_6955), .ck(clk), .d(n2748) );
ms00f80  l0538 ( .o(net_163), .ck(clk), .d(n2753) );
ms00f80  l0539 ( .o(_net_6097), .ck(clk), .d(n2758) );
ms00f80  l0540 ( .o(net_7225), .ck(clk), .d(n2762) );
ms00f80  l0541 ( .o(net_7108), .ck(clk), .d(n2767) );
ms00f80  l0542 ( .o(_net_6022), .ck(clk), .d(n2771) );
ms00f80  l0543 ( .o(_net_5978), .ck(clk), .d(n2776) );
ms00f80  l0544 ( .o(net_6880), .ck(clk), .d(n2781) );
ms00f80  l0545 ( .o(net_7343), .ck(clk), .d(n2784) );
ms00f80  l0546 ( .o(net_6496), .ck(clk), .d(n2788) );
ms00f80  l0547 ( .o(net_6664), .ck(clk), .d(n2792) );
ms00f80  l0548 ( .o(net_232), .ck(clk), .d(n2797) );
ms00f80  l0549 ( .o(net_6524), .ck(clk), .d(n2801) );
ms00f80  l0550 ( .o(_net_7820), .ck(clk), .d(n2805) );
ms00f80  l0551 ( .o(_net_214), .ck(clk), .d(n2810) );
ms00f80  l0552 ( .o(net_6539), .ck(clk), .d(n2814) );
ms00f80  l0553 ( .o(net_6579), .ck(clk), .d(n2819) );
ms00f80  l0554 ( .o(net_7024), .ck(clk), .d(n2823) );
ms00f80  l0555 ( .o(net_7153), .ck(clk), .d(n2827) );
ms00f80  l0556 ( .o(_net_6156), .ck(clk), .d(n2831) );
ms00f80  l0557 ( .o(_net_6029), .ck(clk), .d(n2836) );
ms00f80  l0558 ( .o(net_6631), .ck(clk), .d(n2840) );
ms00f80  l0559 ( .o(_net_7261), .ck(clk), .d(n2845) );
ms00f80  l0560 ( .o(net_7670), .ck(clk), .d(n2850) );
ms00f80  l0561 ( .o(_net_7501), .ck(clk), .d(n2855) );
ms00f80  l0562 ( .o(net_7236), .ck(clk), .d(n2860) );
ms00f80  l0563 ( .o(net_6246), .ck(clk), .d(n2864) );
ms00f80  l0564 ( .o(net_6478), .ck(clk), .d(n2869) );
ms00f80  l0565 ( .o(net_6578), .ck(clk), .d(n2873) );
ms00f80  l0566 ( .o(net_6244), .ck(clk), .d(n2877) );
ms00f80  l0567 ( .o(net_7547), .ck(clk), .d(n2882) );
ms00f80  l0568 ( .o(net_6813), .ck(clk), .d(n2885) );
ms00f80  l0569 ( .o(_net_7572), .ck(clk), .d(n2890) );
ms00f80  l0570 ( .o(net_7756), .ck(clk), .d(n2895) );
ms00f80  l0571 ( .o(_net_7722), .ck(clk), .d(n2900) );
ms00f80  l0572 ( .o(net_7461), .ck(clk), .d(n2904) );
ms00f80  l0573 ( .o(net_6946), .ck(clk), .d(n2908) );
ms00f80  l0574 ( .o(net_7336), .ck(clk), .d(n2913) );
ms00f80  l0575 ( .o(x315), .ck(clk), .d(n2918) );
ms00f80  l0576 ( .o(net_7022), .ck(clk), .d(n2922) );
ms00f80  l0577 ( .o(net_6755), .ck(clk), .d(n2926) );
ms00f80  l0578 ( .o(_net_6221), .ck(clk), .d(n2930) );
ms00f80  l0579 ( .o(_net_5920), .ck(clk), .d(n2935) );
ms00f80  l0580 ( .o(net_6781), .ck(clk), .d(n2939) );
ms00f80  l0581 ( .o(net_7158), .ck(clk), .d(n2944) );
ms00f80  l0582 ( .o(_net_5969), .ck(clk), .d(n2948) );
ms00f80  l0583 ( .o(_net_7552), .ck(clk), .d(n2953) );
ms00f80  l0584 ( .o(net_7457), .ck(clk), .d(n2958) );
ms00f80  l0585 ( .o(net_6338), .ck(clk), .d(n2963) );
ms00f80  l0586 ( .o(net_337), .ck(clk), .d(n2967) );
ms00f80  l0587 ( .o(net_7007), .ck(clk), .d(n2972) );
ms00f80  l0588 ( .o(_net_266), .ck(clk), .d(n2976) );
ms00f80  l0589 ( .o(_net_6553), .ck(clk), .d(n2981) );
ms00f80  l0590 ( .o(_net_6063), .ck(clk), .d(n2986) );
ms00f80  l0591 ( .o(_net_7531), .ck(clk), .d(n2991) );
ms00f80  l0592 ( .o(net_6438), .ck(clk), .d(n2996) );
ms00f80  l0593 ( .o(_net_6038), .ck(clk), .d(n3000) );
ms00f80  l0594 ( .o(_net_6090), .ck(clk), .d(n3005) );
ms00f80  l0595 ( .o(_net_7751), .ck(clk), .d(n3010) );
ms00f80  l0596 ( .o(net_7609), .ck(clk), .d(n3015) );
ms00f80  l0597 ( .o(_net_7320), .ck(clk), .d(n3020) );
ms00f80  l0598 ( .o(_net_173), .ck(clk), .d(n3025) );
ms00f80  l0599 ( .o(net_7105), .ck(clk), .d(n3030) );
ms00f80  l0600 ( .o(net_6906), .ck(clk), .d(n3033) );
ms00f80  l0601 ( .o(net_6909), .ck(clk), .d(n3037) );
ms00f80  l0602 ( .o(_net_6023), .ck(clk), .d(n3042) );
ms00f80  l0603 ( .o(_net_7667), .ck(clk), .d(n3047) );
ms00f80  l0604 ( .o(net_7136), .ck(clk), .d(n3052) );
ms00f80  l0605 ( .o(_net_226), .ck(clk), .d(n3056) );
ms00f80  l0606 ( .o(net_7121), .ck(clk), .d(n3061) );
ms00f80  l0607 ( .o(_net_184), .ck(clk), .d(n3065) );
ms00f80  l0608 ( .o(net_6938), .ck(clk), .d(n3069) );
ms00f80  l0609 ( .o(net_6717), .ck(clk), .d(n3074) );
ms00f80  l0610 ( .o(net_233), .ck(clk), .d(n3078) );
ms00f80  l0611 ( .o(net_6796), .ck(clk), .d(n3082) );
ms00f80  l0612 ( .o(_net_6688), .ck(clk), .d(n3087) );
ms00f80  l0613 ( .o(_net_6281), .ck(clk), .d(n3092) );
ms00f80  l0614 ( .o(_net_128), .ck(clk), .d(n3097) );
ms00f80  l0615 ( .o(net_6706), .ck(clk), .d(n3102) );
ms00f80  l0616 ( .o(net_303), .ck(clk), .d(n3105) );
ms00f80  l0617 ( .o(net_6473), .ck(clk), .d(n3110) );
ms00f80  l0618 ( .o(net_6743), .ck(clk), .d(n3114) );
ms00f80  l0619 ( .o(net_153), .ck(clk), .d(n3117) );
ms00f80  l0620 ( .o(net_7643), .ck(clk), .d(n3121) );
ms00f80  l0621 ( .o(net_7387), .ck(clk), .d(n3126) );
ms00f80  l0622 ( .o(_net_7410), .ck(clk), .d(n3130) );
ms00f80  l0623 ( .o(net_6639), .ck(clk), .d(n3134) );
ms00f80  l0624 ( .o(_net_7557), .ck(clk), .d(n3139) );
ms00f80  l0625 ( .o(net_6681), .ck(clk), .d(n3143) );
ms00f80  l0626 ( .o(_net_7449), .ck(clk), .d(n3148) );
ms00f80  l0627 ( .o(net_7040), .ck(clk), .d(n3152) );
ms00f80  l0628 ( .o(_net_7690), .ck(clk), .d(n3157) );
ms00f80  l0629 ( .o(net_6751), .ck(clk), .d(n3162) );
ms00f80  l0630 ( .o(net_7738), .ck(clk), .d(n3165) );
ms00f80  l0631 ( .o(_net_7470), .ck(clk), .d(n3170) );
ms00f80  l0632 ( .o(net_152), .ck(clk), .d(n3174) );
ms00f80  l0633 ( .o(net_6450), .ck(clk), .d(n3178) );
ms00f80  l0634 ( .o(_net_7350), .ck(clk), .d(n3182) );
ms00f80  l0635 ( .o(net_135), .ck(clk), .d(n3186) );
ms00f80  l0636 ( .o(net_6861), .ck(clk), .d(n3190) );
ms00f80  l0637 ( .o(_net_7277), .ck(clk), .d(n3194) );
ms00f80  l0638 ( .o(net_7536), .ck(clk), .d(n3199) );
ms00f80  l0639 ( .o(_net_178), .ck(clk), .d(n3203) );
ms00f80  l0640 ( .o(net_6488), .ck(clk), .d(n3207) );
ms00f80  l0641 ( .o(_net_7326), .ck(clk), .d(n3212) );
ms00f80  l0642 ( .o(_net_6110), .ck(clk), .d(n3217) );
ms00f80  l0643 ( .o(_net_7478), .ck(clk), .d(n3222) );
ms00f80  l0644 ( .o(net_6233), .ck(clk), .d(n3226) );
ms00f80  l0645 ( .o(_net_154), .ck(clk), .d(n3231) );
ms00f80  l0646 ( .o(_net_7812), .ck(clk), .d(n3235) );
ms00f80  l0647 ( .o(_net_6175), .ck(clk), .d(n3240) );
ms00f80  l0648 ( .o(net_6652), .ck(clk), .d(n3244) );
ms00f80  l0649 ( .o(_net_6259), .ck(clk), .d(n3249) );
ms00f80  l0650 ( .o(_net_272), .ck(clk), .d(n3254) );
ms00f80  l0651 ( .o(_net_7821), .ck(clk), .d(n3258) );
ms00f80  l0652 ( .o(_net_116), .ck(clk), .d(n3263) );
ms00f80  l0653 ( .o(_net_6102), .ck(clk), .d(n3268) );
ms00f80  l0654 ( .o(net_6661), .ck(clk), .d(n3272) );
ms00f80  l0655 ( .o(net_7488), .ck(clk), .d(n3276) );
ms00f80  l0656 ( .o(net_6760), .ck(clk), .d(n3280) );
ms00f80  l0657 ( .o(_net_6204), .ck(clk), .d(n3285) );
ms00f80  l0658 ( .o(net_7710), .ck(clk), .d(n3290) );
ms00f80  l0659 ( .o(_net_6083), .ck(clk), .d(n3294) );
ms00f80  l0660 ( .o(net_6623), .ck(clk), .d(n3299) );
ms00f80  l0661 ( .o(net_6536), .ck(clk), .d(n3303) );
ms00f80  l0662 ( .o(_net_7266), .ck(clk), .d(n3308) );
ms00f80  l0663 ( .o(_net_6171), .ck(clk), .d(n3313) );
ms00f80  l0664 ( .o(net_6883), .ck(clk), .d(n3318) );
ms00f80  l0665 ( .o(x447), .ck(clk), .d(n3322) );
ms00f80  l0666 ( .o(net_7310), .ck(clk), .d(n3325) );
ms00f80  l0667 ( .o(net_6868), .ck(clk), .d(n3330) );
ms00f80  l0668 ( .o(net_7344), .ck(clk), .d(n3333) );
ms00f80  l0669 ( .o(_net_6041), .ck(clk), .d(n3338) );
ms00f80  l0670 ( .o(_net_6199), .ck(clk), .d(n3343) );
ms00f80  l0671 ( .o(net_7140), .ck(clk), .d(n3348) );
ms00f80  l0672 ( .o(x589), .ck(clk), .d(n3352) );
ms00f80  l0673 ( .o(_net_7583), .ck(clk), .d(n3356) );
ms00f80  l0674 ( .o(net_6247), .ck(clk), .d(n3361) );
ms00f80  l0675 ( .o(net_6548), .ck(clk), .d(n3365) );
ms00f80  l0676 ( .o(_net_5980), .ck(clk), .d(n3370) );
ms00f80  l0677 ( .o(net_7517), .ck(clk), .d(n3374) );
ms00f80  l0678 ( .o(net_6698), .ck(clk), .d(n3379) );
ms00f80  l0679 ( .o(net_6485), .ck(clk), .d(n3383) );
ms00f80  l0680 ( .o(net_7042), .ck(clk), .d(n3386) );
ms00f80  l0681 ( .o(_net_7814), .ck(clk), .d(n3390) );
ms00f80  l0682 ( .o(_net_6142), .ck(clk), .d(n3395) );
ms00f80  l0683 ( .o(_net_7619), .ck(clk), .d(n3400) );
ms00f80  l0684 ( .o(net_371), .ck(clk), .d(n3404) );
ms00f80  l0685 ( .o(net_6547), .ck(clk), .d(n3408) );
ms00f80  l0686 ( .o(net_6214), .ck(clk), .d(n3413) );
ms00f80  l0687 ( .o(net_7248), .ck(clk), .d(n3418) );
ms00f80  l0688 ( .o(net_197), .ck(clk), .d(n3422) );
ms00f80  l0689 ( .o(_net_7618), .ck(clk), .d(n3427) );
ms00f80  l0690 ( .o(net_7743), .ck(clk), .d(n3431) );
ms00f80  l0691 ( .o(net_7120), .ck(clk), .d(n3436) );
ms00f80  l0692 ( .o(_net_211), .ck(clk), .d(n3440) );
ms00f80  l0693 ( .o(net_334), .ck(clk), .d(n3445) );
ms00f80  l0694 ( .o(net_6369), .ck(clk), .d(n3450) );
ms00f80  l0695 ( .o(x786), .ck(clk), .d(n3455) );
ms00f80  l0696 ( .o(_net_6075), .ck(clk), .d(n3459) );
ms00f80  l0697 ( .o(_net_191), .ck(clk), .d(n3464) );
ms00f80  l0698 ( .o(net_7213), .ck(clk), .d(n3469) );
ms00f80  l0699 ( .o(_net_6130), .ck(clk), .d(n3474) );
ms00f80  l0700 ( .o(net_6332), .ck(clk), .d(n3479) );
ms00f80  l0701 ( .o(_net_6290), .ck(clk), .d(n3484) );
ms00f80  l0702 ( .o(_net_7362), .ck(clk), .d(n3489) );
ms00f80  l0703 ( .o(net_7241), .ck(clk), .d(n3494) );
ms00f80  l0704 ( .o(net_140), .ck(clk), .d(n3497) );
ms00f80  l0705 ( .o(net_7766), .ck(clk), .d(n3502) );
ms00f80  l0706 ( .o(_net_6078), .ck(clk), .d(n3507) );
ms00f80  l0707 ( .o(net_7195), .ck(clk), .d(n3511) );
ms00f80  l0708 ( .o(_net_6687), .ck(clk), .d(n3516) );
ms00f80  l0709 ( .o(net_6765), .ck(clk), .d(n3520) );
ms00f80  l0710 ( .o(net_6216), .ck(clk), .d(n3524) );
ms00f80  l0711 ( .o(net_7082), .ck(clk), .d(n3528) );
ms00f80  l0712 ( .o(net_329), .ck(clk), .d(n3532) );
ms00f80  l0713 ( .o(net_6254), .ck(clk), .d(n3537) );
ms00f80  l0714 ( .o(net_6885), .ck(clk), .d(n3542) );
ms00f80  l0715 ( .o(net_7642), .ck(clk), .d(n3546) );
ms00f80  l0716 ( .o(net_7231), .ck(clk), .d(n3551) );
ms00f80  l0717 ( .o(net_310), .ck(clk), .d(n3555) );
ms00f80  l0718 ( .o(net_6505), .ck(clk), .d(n3559) );
ms00f80  l0719 ( .o(net_6873), .ck(clk), .d(n3564) );
ms00f80  l0720 ( .o(net_7672), .ck(clk), .d(n3567) );
ms00f80  l0721 ( .o(_net_7703), .ck(clk), .d(n3572) );
ms00f80  l0722 ( .o(_net_6408), .ck(clk), .d(n3577) );
ms00f80  l0723 ( .o(net_255), .ck(clk), .d(n3582) );
ms00f80  l0724 ( .o(net_6476), .ck(clk), .d(n3587) );
ms00f80  l0725 ( .o(net_6530), .ck(clk), .d(n3590) );
ms00f80  l0726 ( .o(_net_5962), .ck(clk), .d(n3595) );
ms00f80  l0727 ( .o(net_6583), .ck(clk), .d(n3600) );
ms00f80  l0728 ( .o(net_7678), .ck(clk), .d(n3604) );
ms00f80  l0729 ( .o(_net_6092), .ck(clk), .d(n3609) );
ms00f80  l0730 ( .o(_net_5988), .ck(clk), .d(n3614) );
ms00f80  l0731 ( .o(net_6674), .ck(clk), .d(n3618) );
ms00f80  l0732 ( .o(net_6320), .ck(clk), .d(n3623) );
ms00f80  l0733 ( .o(_net_7781), .ck(clk), .d(n3628) );
ms00f80  l0734 ( .o(_net_7665), .ck(clk), .d(n3633) );
ms00f80  l0735 ( .o(net_7378), .ck(clk), .d(n3638) );
ms00f80  l0736 ( .o(net_7737), .ck(clk), .d(n3642) );
ms00f80  l0737 ( .o(x217), .ck(clk), .d(n3647) );
ms00f80  l0738 ( .o(net_7157), .ck(clk), .d(n3651) );
ms00f80  l0739 ( .o(net_6591), .ck(clk), .d(n3655) );
ms00f80  l0740 ( .o(net_6395), .ck(clk), .d(n3658) );
ms00f80  l0741 ( .o(net_7490), .ck(clk), .d(n3661) );
ms00f80  l0742 ( .o(_net_7424), .ck(clk), .d(n3666) );
ms00f80  l0743 ( .o(net_7061), .ck(clk), .d(n3670) );
ms00f80  l0744 ( .o(_net_7728), .ck(clk), .d(n3675) );
ms00f80  l0745 ( .o(net_7171), .ck(clk), .d(n3679) );
ms00f80  l0746 ( .o(_net_5854), .ck(clk), .d(n3684) );
ms00f80  l0747 ( .o(net_6605), .ck(clk), .d(n3689) );
ms00f80  l0748 ( .o(_net_7250), .ck(clk), .d(n3693) );
ms00f80  l0749 ( .o(_net_5853), .ck(clk), .d(n3698) );
ms00f80  l0750 ( .o(net_6976), .ck(clk), .d(n3703) );
ms00f80  l0751 ( .o(net_6721), .ck(clk), .d(n3707) );
ms00f80  l0752 ( .o(net_7775), .ck(clk), .d(n3711) );
ms00f80  l0753 ( .o(net_6486), .ck(clk), .d(n3716) );
ms00f80  l0754 ( .o(net_6268), .ck(clk), .d(n3720) );
ms00f80  l0755 ( .o(net_6881), .ck(clk), .d(n3725) );
ms00f80  l0756 ( .o(net_7048), .ck(clk), .d(n3729) );
ms00f80  l0757 ( .o(net_7799), .ck(clk), .d(n3733) );
ms00f80  l0758 ( .o(_net_7444), .ck(clk), .d(n3737) );
ms00f80  l0759 ( .o(_net_7598), .ck(clk), .d(n3742) );
ms00f80  l0760 ( .o(net_6325), .ck(clk), .d(n3747) );
ms00f80  l0761 ( .o(net_6245), .ck(clk), .d(n3752) );
ms00f80  l0762 ( .o(net_336), .ck(clk), .d(n3756) );
ms00f80  l0763 ( .o(net_6442), .ck(clk), .d(n3761) );
ms00f80  l0764 ( .o(_net_290), .ck(clk), .d(n3765) );
ms00f80  l0765 ( .o(net_6991), .ck(clk), .d(n3770) );
ms00f80  l0766 ( .o(net_6928), .ck(clk), .d(n3773) );
ms00f80  l0767 ( .o(net_6525), .ck(clk), .d(n3777) );
ms00f80  l0768 ( .o(_net_7626), .ck(clk), .d(n3782) );
ms00f80  l0769 ( .o(_net_7092), .ck(clk), .d(n3787) );
ms00f80  l0770 ( .o(net_6666), .ck(clk), .d(n3791) );
ms00f80  l0771 ( .o(_net_7785), .ck(clk), .d(n3796) );
ms00f80  l0772 ( .o(net_7149), .ck(clk), .d(n3801) );
ms00f80  l0773 ( .o(net_7714), .ck(clk), .d(n3805) );
ms00f80  l0774 ( .o(net_6429), .ck(clk), .d(n3809) );
ms00f80  l0775 ( .o(net_182), .ck(clk), .d(n3813) );
ms00f80  l0776 ( .o(net_339), .ck(clk), .d(n3817) );
ms00f80  l0777 ( .o(net_6252), .ck(clk), .d(n3822) );
ms00f80  l0778 ( .o(net_286), .ck(clk), .d(n3827) );
ms00f80  l0779 ( .o(net_6799), .ck(clk), .d(n3831) );
ms00f80  l0780 ( .o(_net_6419), .ck(clk), .d(n3836) );
ms00f80  l0781 ( .o(_net_7652), .ck(clk), .d(n3841) );
ms00f80  l0782 ( .o(_net_6158), .ck(clk), .d(n3846) );
ms00f80  l0783 ( .o(net_6829), .ck(clk), .d(n3851) );
ms00f80  l0784 ( .o(net_6595), .ck(clk), .d(n3855) );
ms00f80  l0785 ( .o(_net_7290), .ck(clk), .d(n3859) );
ms00f80  l0786 ( .o(net_6850), .ck(clk), .d(n3864) );
ms00f80  l0787 ( .o(net_6636), .ck(clk), .d(n3867) );
ms00f80  l0788 ( .o(_net_188), .ck(clk), .d(n3872) );
ms00f80  l0789 ( .o(_net_6065), .ck(clk), .d(n3877) );
ms00f80  l0790 ( .o(net_6899), .ck(clk), .d(n3881) );
ms00f80  l0791 ( .o(_net_7574), .ck(clk), .d(n3886) );
ms00f80  l0792 ( .o(_net_123), .ck(clk), .d(n3891) );
ms00f80  l0793 ( .o(net_6855), .ck(clk), .d(n3896) );
ms00f80  l0794 ( .o(net_7034), .ck(clk), .d(n3899) );
ms00f80  l0795 ( .o(net_7239), .ck(clk), .d(n3904) );
ms00f80  l0796 ( .o(net_223), .ck(clk), .d(n3908) );
ms00f80  l0797 ( .o(_net_7270), .ck(clk), .d(n3913) );
ms00f80  l0798 ( .o(net_7184), .ck(clk), .d(n3917) );
ms00f80  l0799 ( .o(_net_6116), .ck(clk), .d(n3922) );
ms00f80  l0800 ( .o(_net_7563), .ck(clk), .d(n3927) );
ms00f80  l0801 ( .o(_net_7418), .ck(clk), .d(n3932) );
ms00f80  l0802 ( .o(net_6685), .ck(clk), .d(n3936) );
ms00f80  l0803 ( .o(_net_7591), .ck(clk), .d(n3941) );
ms00f80  l0804 ( .o(net_369), .ck(clk), .d(n3945) );
ms00f80  l0805 ( .o(net_6819), .ck(clk), .d(n3949) );
ms00f80  l0806 ( .o(net_7185), .ck(clk), .d(n3953) );
ms00f80  l0807 ( .o(net_372), .ck(clk), .d(n3957) );
ms00f80  l0808 ( .o(net_6372), .ck(clk), .d(n3962) );
ms00f80  l0809 ( .o(_net_7510), .ck(clk), .d(n3967) );
ms00f80  l0810 ( .o(net_7537), .ck(clk), .d(n3972) );
ms00f80  l0811 ( .o(_net_6202), .ck(clk), .d(n3976) );
ms00f80  l0812 ( .o(_net_6112), .ck(clk), .d(n3981) );
ms00f80  l0813 ( .o(net_7050), .ck(clk), .d(n3985) );
ms00f80  l0814 ( .o(net_309), .ck(clk), .d(n3989) );
ms00f80  l0815 ( .o(net_7165), .ck(clk), .d(n3993) );
ms00f80  l0816 ( .o(_net_7095), .ck(clk), .d(n3998) );
ms00f80  l0817 ( .o(net_6949), .ck(clk), .d(n4002) );
ms00f80  l0818 ( .o(net_6852), .ck(clk), .d(n4007) );
ms00f80  l0819 ( .o(net_6279), .ck(clk), .d(n4011) );
ms00f80  l0820 ( .o(_net_7733), .ck(clk), .d(n4016) );
ms00f80  l0821 ( .o(net_6810), .ck(clk), .d(n4020) );
ms00f80  l0822 ( .o(net_141), .ck(clk), .d(n4024) );
ms00f80  l0823 ( .o(_net_7601), .ck(clk), .d(n4029) );
ms00f80  l0824 ( .o(net_7191), .ck(clk), .d(n4033) );
ms00f80  l0825 ( .o(net_6790), .ck(clk), .d(n4037) );
ms00f80  l0826 ( .o(_net_7633), .ck(clk), .d(n4042) );
ms00f80  l0827 ( .o(net_355), .ck(clk), .d(n4046) );
ms00f80  l0828 ( .o(net_6613), .ck(clk), .d(n4051) );
ms00f80  l0829 ( .o(net_7711), .ck(clk), .d(n4055) );
ms00f80  l0830 ( .o(net_7013), .ck(clk), .d(n4059) );
ms00f80  l0831 ( .o(_net_7329), .ck(clk), .d(n4063) );
ms00f80  l0832 ( .o(net_6444), .ck(clk), .d(n4068) );
ms00f80  l0833 ( .o(net_6541), .ck(clk), .d(n4071) );
ms00f80  l0834 ( .o(net_364), .ck(clk), .d(n4075) );
ms00f80  l0835 ( .o(net_7636), .ck(clk), .d(n4079) );
ms00f80  l0836 ( .o(_net_294), .ck(clk), .d(n4084) );
ms00f80  l0837 ( .o(_net_6411), .ck(clk), .d(n4089) );
ms00f80  l0838 ( .o(_net_7404), .ck(clk), .d(n4094) );
ms00f80  l0839 ( .o(net_6493), .ck(clk), .d(n4098) );
ms00f80  l0840 ( .o(net_6778), .ck(clk), .d(n4102) );
ms00f80  l0841 ( .o(_net_7719), .ck(clk), .d(n4107) );
ms00f80  l0842 ( .o(net_6867), .ck(clk), .d(n4112) );
ms00f80  l0843 ( .o(_net_7364), .ck(clk), .d(n4116) );
ms00f80  l0844 ( .o(_net_276), .ck(clk), .d(n4121) );
ms00f80  l0845 ( .o(_net_7227), .ck(clk), .d(n4126) );
ms00f80  l0846 ( .o(net_7400), .ck(clk), .d(n4131) );
ms00f80  l0847 ( .o(_net_7232), .ck(clk), .d(n4135) );
ms00f80  l0848 ( .o(_net_7347), .ck(clk), .d(n4140) );
ms00f80  l0849 ( .o(net_6592), .ck(clk), .d(n4145) );
ms00f80  l0850 ( .o(net_7028), .ck(clk), .d(n4148) );
ms00f80  l0851 ( .o(_net_6239), .ck(clk), .d(n4153) );
ms00f80  l0852 ( .o(net_6714), .ck(clk), .d(n4158) );
ms00f80  l0853 ( .o(net_367), .ck(clk), .d(n4161) );
ms00f80  l0854 ( .o(_net_7437), .ck(clk), .d(n4166) );
ms00f80  l0855 ( .o(_net_7784), .ck(clk), .d(n4171) );
ms00f80  l0856 ( .o(net_6263), .ck(clk), .d(n4176) );
ms00f80  l0857 ( .o(net_234), .ck(clk), .d(n4181) );
ms00f80  l0858 ( .o(_net_7321), .ck(clk), .d(n4186) );
ms00f80  l0859 ( .o(net_7123), .ck(clk), .d(n4191) );
ms00f80  l0860 ( .o(net_6684), .ck(clk), .d(n4194) );
ms00f80  l0861 ( .o(net_6447), .ck(clk), .d(n4199) );
ms00f80  l0862 ( .o(_net_277), .ck(clk), .d(n4203) );
ms00f80  l0863 ( .o(net_7178), .ck(clk), .d(n4207) );
ms00f80  l0864 ( .o(net_206), .ck(clk), .d(n4212) );
ms00f80  l0865 ( .o(_net_7630), .ck(clk), .d(n4217) );
ms00f80  l0866 ( .o(net_7049), .ck(clk), .d(n4221) );
ms00f80  l0867 ( .o(_net_5968), .ck(clk), .d(n4226) );
ms00f80  l0868 ( .o(net_5858), .ck(clk), .d(n4231) );
ms00f80  l0869 ( .o(net_6643), .ck(clk), .d(n4235) );
ms00f80  l0870 ( .o(_net_7635), .ck(clk), .d(n4240) );
ms00f80  l0871 ( .o(net_7398), .ck(clk), .d(n4245) );
ms00f80  l0872 ( .o(_net_6152), .ck(clk), .d(n4249) );
ms00f80  l0873 ( .o(net_376), .ck(clk), .d(n4253) );
ms00f80  l0874 ( .o(net_296), .ck(clk), .d(n4258) );
ms00f80  l0875 ( .o(net_7338), .ck(clk), .d(n4263) );
ms00f80  l0876 ( .o(net_7031), .ck(clk), .d(n4267) );
ms00f80  l0877 ( .o(net_312), .ck(clk), .d(n4271) );
ms00f80  l0878 ( .o(_net_5981), .ck(clk), .d(n4276) );
ms00f80  l0879 ( .o(net_6926), .ck(clk), .d(n4280) );
ms00f80  l0880 ( .o(_net_7810), .ck(clk), .d(n4284) );
ms00f80  l0881 ( .o(_net_229), .ck(clk), .d(n4289) );
ms00f80  l0882 ( .o(_net_7318), .ck(clk), .d(n4294) );
ms00f80  l0883 ( .o(_net_6128), .ck(clk), .d(n4299) );
ms00f80  l0884 ( .o(_net_7688), .ck(clk), .d(n4304) );
ms00f80  l0885 ( .o(net_6753), .ck(clk), .d(n4309) );
ms00f80  l0886 ( .o(_net_6422), .ck(clk), .d(n4313) );
ms00f80  l0887 ( .o(net_6471), .ck(clk), .d(n4318) );
ms00f80  l0888 ( .o(_net_6050), .ck(clk), .d(n4322) );
ms00f80  l0889 ( .o(net_6388), .ck(clk), .d(n4326) );
ms00f80  l0890 ( .o(net_6978), .ck(clk), .d(n4330) );
ms00f80  l0891 ( .o(net_7641), .ck(clk), .d(n4333) );
ms00f80  l0892 ( .o(net_6805), .ck(clk), .d(n4338) );
ms00f80  l0893 ( .o(net_7771), .ck(clk), .d(n4343) );
ms00f80  l0894 ( .o(_net_7505), .ck(clk), .d(n4348) );
ms00f80  l0895 ( .o(net_7646), .ck(clk), .d(n4352) );
ms00f80  l0896 ( .o(_net_6009), .ck(clk), .d(n4357) );
ms00f80  l0897 ( .o(net_6863), .ck(clk), .d(n4362) );
ms00f80  l0898 ( .o(net_6762), .ck(clk), .d(n4365) );
ms00f80  l0899 ( .o(net_6641), .ck(clk), .d(n4370) );
ms00f80  l0900 ( .o(net_6950), .ck(clk), .d(n4374) );
ms00f80  l0901 ( .o(_net_7278), .ck(clk), .d(n4379) );
ms00f80  l0902 ( .o(net_6974), .ck(clk), .d(n4384) );
ms00f80  l0903 ( .o(net_6431), .ck(clk), .d(n4388) );
ms00f80  l0904 ( .o(_net_7301), .ck(clk), .d(n4392) );
ms00f80  l0905 ( .o(net_6564), .ck(clk), .d(n4397) );
ms00f80  l0906 ( .o(net_7162), .ck(clk), .d(n4401) );
ms00f80  l0907 ( .o(_net_265), .ck(clk), .d(n4405) );
ms00f80  l0908 ( .o(net_7111), .ck(clk), .d(n4410) );
ms00f80  l0909 ( .o(_net_7718), .ck(clk), .d(n4414) );
ms00f80  l0910 ( .o(net_6347), .ck(clk), .d(n4419) );
ms00f80  l0911 ( .o(_net_6045), .ck(clk), .d(n4424) );
ms00f80  l0912 ( .o(net_7366), .ck(clk), .d(n4428) );
ms00f80  l0913 ( .o(_net_7332), .ck(clk), .d(n4433) );
ms00f80  l0914 ( .o(_net_7403), .ck(clk), .d(n4438) );
ms00f80  l0915 ( .o(_net_6206), .ck(clk), .d(n4443) );
ms00f80  l0916 ( .o(net_6886), .ck(clk), .d(n4448) );
ms00f80  l0917 ( .o(net_7374), .ck(clk), .d(n4451) );
ms00f80  l0918 ( .o(x179), .ck(clk), .d(n4456) );
ms00f80  l0919 ( .o(net_7741), .ck(clk), .d(n4459) );
ms00f80  l0920 ( .o(_net_7323), .ck(clk), .d(n4464) );
ms00f80  l0921 ( .o(net_6343), .ck(clk), .d(n4469) );
ms00f80  l0922 ( .o(net_7199), .ck(clk), .d(n4473) );
ms00f80  l0923 ( .o(net_6448), .ck(clk), .d(n4478) );
ms00f80  l0924 ( .o(_net_6148), .ck(clk), .d(n4482) );
ms00f80  l0925 ( .o(net_7129), .ck(clk), .d(n4487) );
ms00f80  l0926 ( .o(_net_6018), .ck(clk), .d(n4491) );
ms00f80  l0927 ( .o(net_389), .ck(clk), .d(n4496) );
ms00f80  l0928 ( .o(net_155), .ck(clk), .d(n4501) );
ms00f80  l0929 ( .o(net_7075), .ck(clk), .d(n4505) );
ms00f80  l0930 ( .o(_net_7469), .ck(clk), .d(n4510) );
ms00f80  l0931 ( .o(_net_6173), .ck(clk), .d(n4515) );
ms00f80  l0932 ( .o(net_246), .ck(clk), .d(n4520) );
ms00f80  l0933 ( .o(net_138), .ck(clk), .d(n4524) );
ms00f80  l0934 ( .o(_net_6189), .ck(clk), .d(n4529) );
ms00f80  l0935 ( .o(net_6195), .ck(clk), .d(n4534) );
ms00f80  l0936 ( .o(_net_6172), .ck(clk), .d(n4539) );
ms00f80  l0937 ( .o(_net_7480), .ck(clk), .d(n4544) );
ms00f80  l0938 ( .o(net_6489), .ck(clk), .d(n4548) );
ms00f80  l0939 ( .o(_net_6165), .ck(clk), .d(n4553) );
ms00f80  l0940 ( .o(net_146), .ck(clk), .d(n4558) );
ms00f80  l0941 ( .o(net_6761), .ck(clk), .d(n4562) );
ms00f80  l0942 ( .o(net_6225), .ck(clk), .d(n4567) );
ms00f80  l0943 ( .o(_net_7475), .ck(clk), .d(n4572) );
ms00f80  l0944 ( .o(net_6305), .ck(clk), .d(n4577) );
ms00f80  l0945 ( .o(net_7079), .ck(clk), .d(n4581) );
ms00f80  l0946 ( .o(_net_6297), .ck(clk), .d(n4586) );
ms00f80  l0947 ( .o(_net_7233), .ck(clk), .d(n4591) );
ms00f80  l0948 ( .o(_net_7413), .ck(clk), .d(n4596) );
ms00f80  l0949 ( .o(net_7068), .ck(clk), .d(n4600) );
ms00f80  l0950 ( .o(net_6635), .ck(clk), .d(n4604) );
ms00f80  l0951 ( .o(_net_7586), .ck(clk), .d(n4609) );
ms00f80  l0952 ( .o(net_6776), .ck(clk), .d(n4613) );
ms00f80  l0953 ( .o(net_6637), .ck(clk), .d(n4617) );
ms00f80  l0954 ( .o(net_6273), .ck(clk), .d(n4622) );
ms00f80  l0955 ( .o(_net_7346), .ck(clk), .d(n4627) );
ms00f80  l0956 ( .o(net_6786), .ck(clk), .d(n4631) );
ms00f80  l0957 ( .o(net_253), .ck(clk), .d(n4636) );
ms00f80  l0958 ( .o(_net_6064), .ck(clk), .d(n4641) );
ms00f80  l0959 ( .o(_net_7269), .ck(clk), .d(n4646) );
ms00f80  l0960 ( .o(net_6367), .ck(clk), .d(n4651) );
ms00f80  l0961 ( .o(_net_7288), .ck(clk), .d(n4656) );
ms00f80  l0962 ( .o(net_7197), .ck(clk), .d(n4660) );
ms00f80  l0963 ( .o(net_6736), .ck(clk), .d(n4665) );
ms00f80  l0964 ( .o(net_6581), .ck(clk), .d(n4669) );
ms00f80  l0965 ( .o(net_6055), .ck(clk), .d(n4673) );
ms00f80  l0966 ( .o(x744), .ck(clk), .d(n4678) );
ms00f80  l0967 ( .o(_net_7797), .ck(clk), .d(n4681) );
ms00f80  l0968 ( .o(net_378), .ck(clk), .d(n4686) );
ms00f80  l0969 ( .o(net_7370), .ck(clk), .d(n4690) );
ms00f80  l0970 ( .o(net_7493), .ck(clk), .d(n4694) );
ms00f80  l0971 ( .o(net_6993), .ck(clk), .d(n4699) );
ms00f80  l0972 ( .o(_net_7749), .ck(clk), .d(n4703) );
ms00f80  l0973 ( .o(_net_6073), .ck(clk), .d(n4708) );
ms00f80  l0974 ( .o(net_7142), .ck(clk), .d(n4713) );
ms00f80  l0975 ( .o(net_6544), .ck(clk), .d(n4717) );
ms00f80  l0976 ( .o(net_6271), .ck(clk), .d(n4722) );
ms00f80  l0977 ( .o(_net_7692), .ck(clk), .d(n4727) );
ms00f80  l0978 ( .o(_net_7286), .ck(clk), .d(n4732) );
ms00f80  l0979 ( .o(_net_7382), .ck(clk), .d(n4737) );
ms00f80  l0980 ( .o(net_6735), .ck(clk), .d(n4742) );
ms00f80  l0981 ( .o(net_6502), .ck(clk), .d(n4745) );
ms00f80  l0982 ( .o(net_6334), .ck(clk), .d(n4750) );
ms00f80  l0983 ( .o(net_6349), .ck(clk), .d(n4755) );
ms00f80  l0984 ( .o(_net_7706), .ck(clk), .d(n4760) );
ms00f80  l0985 ( .o(net_6231), .ck(clk), .d(n4765) );
ms00f80  l0986 ( .o(net_7455), .ck(clk), .d(n4769) );
ms00f80  l0987 ( .o(net_7545), .ck(clk), .d(n4774) );
ms00f80  l0988 ( .o(net_6449), .ck(clk), .d(n4778) );
ms00f80  l0989 ( .o(net_6352), .ck(clk), .d(n4782) );
ms00f80  l0990 ( .o(_net_7559), .ck(clk), .d(n4787) );
ms00f80  l0991 ( .o(net_6931), .ck(clk), .d(n4791) );
ms00f80  l0992 ( .o(net_6935), .ck(clk), .d(n4795) );
ms00f80  l0993 ( .o(_net_7452), .ck(clk), .d(n4800) );
ms00f80  l0994 ( .o(net_7014), .ck(clk), .d(n4805) );
ms00f80  l0995 ( .o(_net_7655), .ck(clk), .d(n4809) );
ms00f80  l0996 ( .o(net_7128), .ck(clk), .d(n4814) );
ms00f80  l0997 ( .o(_net_7624), .ck(clk), .d(n4818) );
ms00f80  l0998 ( .o(net_7304), .ck(clk), .d(n4822) );
ms00f80  l0999 ( .o(net_6567), .ck(clk), .d(n4827) );
ms00f80  l1000 ( .o(x234), .ck(clk), .d(n4831) );
ms00f80  l1001 ( .o(net_6650), .ck(clk), .d(n4834) );
ms00f80  l1002 ( .o(net_6509), .ck(clk), .d(n4838) );
ms00f80  l1003 ( .o(_net_6019), .ck(clk), .d(n4843) );
ms00f80  l1004 ( .o(net_6250), .ck(clk), .d(n4848) );
ms00f80  l1005 ( .o(net_6875), .ck(clk), .d(n4853) );
ms00f80  l1006 ( .o(_net_5975), .ck(clk), .d(n4857) );
ms00f80  l1007 ( .o(net_6403), .ck(clk), .d(n4862) );
ms00f80  l1008 ( .o(net_7189), .ck(clk), .d(n4867) );
ms00f80  l1009 ( .o(_net_284), .ck(clk), .d(n4872) );
ms00f80  l1010 ( .o(_net_6406), .ck(clk), .d(n4877) );
ms00f80  l1011 ( .o(net_349), .ck(clk), .d(n4881) );
ms00f80  l1012 ( .o(net_202), .ck(clk), .d(n4886) );
ms00f80  l1013 ( .o(net_7203), .ck(clk), .d(n4890) );
ms00f80  l1014 ( .o(net_7154), .ck(clk), .d(n4895) );
ms00f80  l1015 ( .o(net_6339), .ck(clk), .d(n4899) );
ms00f80  l1016 ( .o(net_7001), .ck(clk), .d(n4904) );
ms00f80  l1017 ( .o(_net_5967), .ck(clk), .d(n4908) );
ms00f80  l1018 ( .o(net_6573), .ck(clk), .d(n4913) );
ms00f80  l1019 ( .o(_net_6011), .ck(clk), .d(n4917) );
ms00f80  l1020 ( .o(_net_5970), .ck(clk), .d(n4922) );
ms00f80  l1021 ( .o(_net_7782), .ck(clk), .d(n4927) );
ms00f80  l1022 ( .o(net_6820), .ck(clk), .d(n4931) );
ms00f80  l1023 ( .o(_net_7659), .ck(clk), .d(n4936) );
ms00f80  l1024 ( .o(net_7047), .ck(clk), .d(n4940) );
ms00f80  l1025 ( .o(net_144), .ck(clk), .d(n4944) );
ms00f80  l1026 ( .o(net_7085), .ck(clk), .d(n4947) );
ms00f80  l1027 ( .o(_net_295), .ck(clk), .d(n4952) );
ms00f80  l1028 ( .o(net_6718), .ck(clk), .d(n4957) );
ms00f80  l1029 ( .o(_net_7651), .ck(clk), .d(n4961) );
ms00f80  l1030 ( .o(net_6923), .ck(clk), .d(n4965) );
ms00f80  l1031 ( .o(net_6808), .ck(clk), .d(n4969) );
ms00f80  l1032 ( .o(_net_6157), .ck(clk), .d(n4974) );
ms00f80  l1033 ( .o(net_6484), .ck(clk), .d(n4979) );
ms00f80  l1034 ( .o(net_6858), .ck(clk), .d(n4983) );
ms00f80  l1035 ( .o(_net_7571), .ck(clk), .d(n4987) );
ms00f80  l1036 ( .o(x765), .ck(clk), .d(n4992) );
ms00f80  l1037 ( .o(net_6241), .ck(clk), .d(n4996) );
ms00f80  l1038 ( .o(net_6617), .ck(clk), .d(n5001) );
ms00f80  l1039 ( .o(net_6854), .ck(clk), .d(n5005) );
ms00f80  l1040 ( .o(net_331), .ck(clk), .d(n5008) );
ms00f80  l1041 ( .o(_net_7727), .ck(clk), .d(n5013) );
ms00f80  l1042 ( .o(_net_6693), .ck(clk), .d(n5018) );
ms00f80  l1043 ( .o(net_7539), .ck(clk), .d(n5023) );
ms00f80  l1044 ( .o(net_7518), .ck(clk), .d(n5027) );
ms00f80  l1045 ( .o(net_6546), .ck(clk), .d(n5031) );
ms00f80  l1046 ( .o(net_7219), .ck(clk), .d(n5035) );
ms00f80  l1047 ( .o(_net_6034), .ck(clk), .d(n5040) );
ms00f80  l1048 ( .o(net_7399), .ck(clk), .d(n5045) );
ms00f80  l1049 ( .o(net_7614), .ck(clk), .d(n5048) );
ms00f80  l1050 ( .o(net_6970), .ck(clk), .d(n5053) );
ms00f80  l1051 ( .o(net_7376), .ck(clk), .d(n5056) );
ms00f80  l1052 ( .o(_net_7507), .ck(clk), .d(n5061) );
ms00f80  l1053 ( .o(net_6311), .ck(clk), .d(n5066) );
ms00f80  l1054 ( .o(net_6663), .ck(clk), .d(n5070) );
ms00f80  l1055 ( .o(_net_7508), .ck(clk), .d(n5075) );
ms00f80  l1056 ( .o(_net_7514), .ck(clk), .d(n5080) );
ms00f80  l1057 ( .o(net_6057), .ck(clk), .d(n5085) );
ms00f80  l1058 ( .o(net_7011), .ck(clk), .d(n5090) );
ms00f80  l1059 ( .o(_net_7433), .ck(clk), .d(n5094) );
ms00f80  l1060 ( .o(net_324), .ck(clk), .d(n5098) );
ms00f80  l1061 ( .o(x379), .ck(clk), .d(n5103) );
ms00f80  l1062 ( .o(net_208), .ck(clk), .d(n5107) );
ms00f80  l1063 ( .o(_net_6415), .ck(clk), .d(n5112) );
ms00f80  l1064 ( .o(_net_227), .ck(clk), .d(n5117) );
ms00f80  l1065 ( .o(net_308), .ck(clk), .d(n5121) );
ms00f80  l1066 ( .o(net_6589), .ck(clk), .d(n5126) );
ms00f80  l1067 ( .o(x149), .ck(clk), .d(n5130) );
ms00f80  l1068 ( .o(net_218), .ck(clk), .d(n5134) );
ms00f80  l1069 ( .o(net_6985), .ck(clk), .d(n5139) );
ms00f80  l1070 ( .o(_net_7272), .ck(clk), .d(n5143) );
ms00f80  l1071 ( .o(net_6572), .ck(clk), .d(n5148) );
ms00f80  l1072 ( .o(net_6516), .ck(clk), .d(n5151) );
ms00f80  l1073 ( .o(net_6428), .ck(clk), .d(n5156) );
ms00f80  l1074 ( .o(net_130), .ck(clk), .d(n5159) );
ms00f80  l1075 ( .o(_net_271), .ck(clk), .d(n5164) );
ms00f80  l1076 ( .o(_net_7435), .ck(clk), .d(n5169) );
ms00f80  l1077 ( .o(net_6940), .ck(clk), .d(n5173) );
ms00f80  l1078 ( .o(net_6841), .ck(clk), .d(n5178) );
ms00f80  l1079 ( .o(_net_7803), .ck(clk), .d(n5181) );
ms00f80  l1080 ( .o(net_7691), .ck(clk), .d(n5186) );
ms00f80  l1081 ( .o(net_6656), .ck(clk), .d(n5189) );
ms00f80  l1082 ( .o(net_7037), .ck(clk), .d(n5193) );
ms00f80  l1083 ( .o(_net_6084), .ck(clk), .d(n5198) );
ms00f80  l1084 ( .o(net_6506), .ck(clk), .d(n5202) );
ms00f80  l1085 ( .o(_net_7686), .ck(clk), .d(n5207) );
ms00f80  l1086 ( .o(_net_6114), .ck(clk), .d(n5212) );
ms00f80  l1087 ( .o(net_6569), .ck(clk), .d(n5217) );
ms00f80  l1088 ( .o(net_6857), .ck(clk), .d(n5221) );
ms00f80  l1089 ( .o(_net_7593), .ck(clk), .d(n5225) );
ms00f80  l1090 ( .o(_net_7422), .ck(clk), .d(n5230) );
ms00f80  l1091 ( .o(net_7176), .ck(clk), .d(n5234) );
ms00f80  l1092 ( .o(net_6487), .ck(clk), .d(n5239) );
ms00f80  l1093 ( .o(net_6676), .ck(clk), .d(n5242) );
ms00f80  l1094 ( .o(net_6897), .ck(clk), .d(n5246) );
ms00f80  l1095 ( .o(_net_7297), .ck(clk), .d(n5251) );
ms00f80  l1096 ( .o(_net_7567), .ck(clk), .d(n5256) );
ms00f80  l1097 ( .o(net_6843), .ck(clk), .d(n5261) );
ms00f80  l1098 ( .o(_net_7416), .ck(clk), .d(n5265) );
ms00f80  l1099 ( .o(net_7168), .ck(clk), .d(n5269) );
ms00f80  l1100 ( .o(_net_7292), .ck(clk), .d(n5274) );
ms00f80  l1101 ( .o(_net_7731), .ck(clk), .d(n5279) );
ms00f80  l1102 ( .o(_net_6284), .ck(clk), .d(n5284) );
ms00f80  l1103 ( .o(net_320), .ck(clk), .d(n5288) );
ms00f80  l1104 ( .o(_net_7599), .ck(clk), .d(n5293) );
ms00f80  l1105 ( .o(net_6965), .ck(clk), .d(n5298) );
ms00f80  l1106 ( .o(net_6324), .ck(clk), .d(n5302) );
ms00f80  l1107 ( .o(_net_7411), .ck(clk), .d(n5307) );
ms00f80  l1108 ( .o(net_7006), .ck(clk), .d(n5312) );
ms00f80  l1109 ( .o(net_6061), .ck(clk), .d(n5316) );
ms00f80  l1110 ( .o(_net_7684), .ck(clk), .d(n5321) );
ms00f80  l1111 ( .o(net_6844), .ck(clk), .d(n5326) );
ms00f80  l1112 ( .o(_net_7662), .ck(clk), .d(n5330) );
ms00f80  l1113 ( .o(net_7002), .ck(clk), .d(n5335) );
ms00f80  l1114 ( .o(net_6357), .ck(clk), .d(n5339) );
ms00f80  l1115 ( .o(_net_6420), .ck(clk), .d(n5344) );
ms00f80  l1116 ( .o(net_6987), .ck(clk), .d(n5349) );
ms00f80  l1117 ( .o(_net_7280), .ck(clk), .d(n5353) );
ms00f80  l1118 ( .o(net_6454), .ck(clk), .d(n5358) );
ms00f80  l1119 ( .o(net_6460), .ck(clk), .d(n5362) );
ms00f80  l1120 ( .o(net_6860), .ck(clk), .d(n5366) );
ms00f80  l1121 ( .o(_net_7657), .ck(clk), .d(n5370) );
ms00f80  l1122 ( .o(net_6237), .ck(clk), .d(n5375) );
ms00f80  l1123 ( .o(net_6729), .ck(clk), .d(n5380) );
ms00f80  l1124 ( .o(net_6816), .ck(clk), .d(n5383) );
ms00f80  l1125 ( .o(_net_6096), .ck(clk), .d(n5388) );
ms00f80  l1126 ( .o(net_7021), .ck(clk), .d(n5393) );
ms00f80  l1127 ( .o(net_159), .ck(clk), .d(n5397) );
ms00f80  l1128 ( .o(net_7151), .ck(clk), .d(n5402) );
ms00f80  l1129 ( .o(_net_7429), .ck(clk), .d(n5406) );
ms00f80  l1130 ( .o(_net_7631), .ck(clk), .d(n5411) );
ms00f80  l1131 ( .o(net_7206), .ck(clk), .d(n5415) );
ms00f80  l1132 ( .o(_net_7295), .ck(clk), .d(n5420) );
ms00f80  l1133 ( .o(net_7167), .ck(clk), .d(n5424) );
ms00f80  l1134 ( .o(_net_6030), .ck(clk), .d(n5429) );
ms00f80  l1135 ( .o(net_6766), .ck(clk), .d(n5433) );
ms00f80  l1136 ( .o(net_380), .ck(clk), .d(n5437) );
ms00f80  l1137 ( .o(net_6551), .ck(clk), .d(n5441) );
ms00f80  l1138 ( .o(_net_119), .ck(clk), .d(n5446) );
ms00f80  l1139 ( .o(net_6436), .ck(clk), .d(n5451) );
ms00f80  l1140 ( .o(_net_5987), .ck(clk), .d(n5455) );
ms00f80  l1141 ( .o(net_6251), .ck(clk), .d(n5460) );
ms00f80  l1142 ( .o(net_7335), .ck(clk), .d(n5464) );
ms00f80  l1143 ( .o(net_6610), .ck(clk), .d(n5469) );
ms00f80  l1144 ( .o(net_7610), .ck(clk), .d(n5472) );
ms00f80  l1145 ( .o(_net_7587), .ck(clk), .d(n5477) );
ms00f80  l1146 ( .o(net_6915), .ck(clk), .d(n5481) );
ms00f80  l1147 ( .o(net_390), .ck(clk), .d(n5486) );
ms00f80  l1148 ( .o(_net_7513), .ck(clk), .d(n5490) );
ms00f80  l1149 ( .o(_net_270), .ck(clk), .d(n5495) );
ms00f80  l1150 ( .o(net_6575), .ck(clk), .d(n5500) );
ms00f80  l1151 ( .o(net_7100), .ck(clk), .d(n5504) );
ms00f80  l1152 ( .o(_net_7467), .ck(clk), .d(n5508) );
ms00f80  l1153 ( .o(net_6024), .ck(clk), .d(n5513) );
ms00f80  l1154 ( .o(x390), .ck(clk), .d(n5517) );
ms00f80  l1155 ( .o(net_7018), .ck(clk), .d(n5521) );
ms00f80  l1156 ( .o(x172), .ck(clk), .d(n5525) );
ms00f80  l1157 ( .o(net_7780), .ck(clk), .d(n5529) );
ms00f80  l1158 ( .o(_net_7721), .ck(clk), .d(n5534) );
ms00f80  l1159 ( .o(net_6839), .ck(clk), .d(n5539) );
ms00f80  l1160 ( .o(_net_7577), .ck(clk), .d(n5543) );
ms00f80  l1161 ( .o(net_6670), .ck(clk), .d(n5547) );
ms00f80  l1162 ( .o(net_7528), .ck(clk), .d(n5552) );
ms00f80  l1163 ( .o(net_343), .ck(clk), .d(n5556) );
ms00f80  l1164 ( .o(net_6789), .ck(clk), .d(n5560) );
ms00f80  l1165 ( .o(_net_7430), .ck(clk), .d(n5565) );
ms00f80  l1166 ( .o(_net_7502), .ck(clk), .d(n5570) );
ms00f80  l1167 ( .o(net_6620), .ck(clk), .d(n5575) );
ms00f80  l1168 ( .o(_net_7622), .ck(clk), .d(n5579) );
ms00f80  l1169 ( .o(net_7546), .ck(clk), .d(n5584) );
ms00f80  l1170 ( .o(net_7235), .ck(clk), .d(n5588) );
ms00f80  l1171 ( .o(net_7640), .ck(clk), .d(n5591) );
ms00f80  l1172 ( .o(_net_6162), .ck(clk), .d(n5596) );
ms00f80  l1173 ( .o(_net_7420), .ck(clk), .d(n5601) );
ms00f80  l1174 ( .o(net_6368), .ck(clk), .d(n5606) );
ms00f80  l1175 ( .o(net_133), .ck(clk), .d(n5610) );
ms00f80  l1176 ( .o(net_7080), .ck(clk), .d(n5613) );
ms00f80  l1177 ( .o(net_6243), .ck(clk), .d(n5618) );
ms00f80  l1178 ( .o(_net_6138), .ck(clk), .d(n5623) );
ms00f80  l1179 ( .o(net_7647), .ck(clk), .d(n5628) );
ms00f80  l1180 ( .o(_net_7736), .ck(clk), .d(n5633) );
ms00f80  l1181 ( .o(_net_6205), .ck(clk), .d(n5638) );
ms00f80  l1182 ( .o(_net_7634), .ck(clk), .d(n5643) );
ms00f80  l1183 ( .o(net_6983), .ck(clk), .d(n5648) );
ms00f80  l1184 ( .o(net_7202), .ck(clk), .d(n5651) );
ms00f80  l1185 ( .o(net_6490), .ck(clk), .d(n5655) );
ms00f80  l1186 ( .o(net_5849), .ck(clk), .d(n5660) );
ms00f80  l1187 ( .o(net_7215), .ck(clk), .d(n5664) );
ms00f80  l1188 ( .o(_net_7380), .ck(clk), .d(n5669) );
ms00f80  l1189 ( .o(_net_7564), .ck(clk), .d(n5674) );
ms00f80  l1190 ( .o(net_6727), .ck(clk), .d(n5679) );
ms00f80  l1191 ( .o(net_7030), .ck(clk), .d(n5682) );
ms00f80  l1192 ( .o(_net_7822), .ck(clk), .d(n5686) );
ms00f80  l1193 ( .o(_net_6283), .ck(clk), .d(n5691) );
ms00f80  l1194 ( .o(net_6609), .ck(clk), .d(n5696) );
ms00f80  l1195 ( .o(net_169), .ck(clk), .d(n5700) );
ms00f80  l1196 ( .o(net_6942), .ck(clk), .d(n5704) );
ms00f80  l1197 ( .o(net_6412), .ck(clk), .d(n5709) );
ms00f80  l1198 ( .o(net_6668), .ck(clk), .d(n5713) );
ms00f80  l1199 ( .o(net_6523), .ck(clk), .d(n5717) );
ms00f80  l1200 ( .o(_net_269), .ck(clk), .d(n5722) );
ms00f80  l1201 ( .o(net_6598), .ck(clk), .d(n5727) );
ms00f80  l1202 ( .o(net_7107), .ck(clk), .d(n5731) );
ms00f80  l1203 ( .o(net_7026), .ck(clk), .d(n5735) );
ms00f80  l1204 ( .o(_net_5998), .ck(clk), .d(n5739) );
ms00f80  l1205 ( .o(net_7244), .ck(clk), .d(n5744) );
ms00f80  l1206 ( .o(_net_6825), .ck(clk), .d(n5748) );
ms00f80  l1207 ( .o(_net_6414), .ck(clk), .d(n5753) );
ms00f80  l1208 ( .o(net_6327), .ck(clk), .d(n5758) );
ms00f80  l1209 ( .o(net_6560), .ck(clk), .d(n5763) );
ms00f80  l1210 ( .o(net_6590), .ck(clk), .d(n5767) );
ms00f80  l1211 ( .o(net_6480), .ck(clk), .d(n5771) );
ms00f80  l1212 ( .o(_net_6154), .ck(clk), .d(n5775) );
ms00f80  l1213 ( .o(net_6642), .ck(clk), .d(n5779) );
ms00f80  l1214 ( .o(net_373), .ck(clk), .d(n5783) );
ms00f80  l1215 ( .o(net_6779), .ck(clk), .d(n5787) );
ms00f80  l1216 ( .o(net_7529), .ck(clk), .d(n5792) );
ms00f80  l1217 ( .o(net_6632), .ck(clk), .d(n5796) );
ms00f80  l1218 ( .o(net_7012), .ck(clk), .d(n5801) );
ms00f80  l1219 ( .o(net_6437), .ck(clk), .d(n5805) );
ms00f80  l1220 ( .o(_net_7561), .ck(clk), .d(n5809) );
ms00f80  l1221 ( .o(net_7676), .ck(clk), .d(n5814) );
ms00f80  l1222 ( .o(net_247), .ck(clk), .d(n5819) );
ms00f80  l1223 ( .o(net_7113), .ck(clk), .d(n5824) );
ms00f80  l1224 ( .o(net_164), .ck(clk), .d(n5828) );
ms00f80  l1225 ( .o(net_6878), .ck(clk), .d(n5833) );
ms00f80  l1226 ( .o(net_6934), .ck(clk), .d(n5836) );
ms00f80  l1227 ( .o(net_6925), .ck(clk), .d(n5840) );
ms00f80  l1228 ( .o(net_259), .ck(clk), .d(n5845) );
ms00f80  l1229 ( .o(_net_7734), .ck(clk), .d(n5850) );
ms00f80  l1230 ( .o(net_6416), .ck(clk), .d(n5855) );
ms00f80  l1231 ( .o(net_6479), .ck(clk), .d(n5860) );
ms00f80  l1232 ( .o(net_7102), .ck(clk), .d(n5864) );
ms00f80  l1233 ( .o(net_7306), .ck(clk), .d(n5867) );
ms00f80  l1234 ( .o(net_6340), .ck(clk), .d(n5872) );
ms00f80  l1235 ( .o(net_6954), .ck(clk), .d(n5876) );
ms00f80  l1236 ( .o(net_6720), .ck(clk), .d(n5881) );
ms00f80  l1237 ( .o(_net_5982), .ck(clk), .d(n5885) );
ms00f80  l1238 ( .o(_net_283), .ck(clk), .d(n5890) );
ms00f80  l1239 ( .o(net_356), .ck(clk), .d(n5894) );
ms00f80  l1240 ( .o(_net_7407), .ck(clk), .d(n5899) );
ms00f80  l1241 ( .o(net_7792), .ck(clk), .d(n5903) );
ms00f80  l1242 ( .o(net_6376), .ck(clk), .d(n5908) );
ms00f80  l1243 ( .o(net_6538), .ck(clk), .d(n5912) );
ms00f80  l1244 ( .o(net_6971), .ck(clk), .d(n5917) );
ms00f80  l1245 ( .o(net_6927), .ck(clk), .d(n5920) );
ms00f80  l1246 ( .o(_net_6040), .ck(clk), .d(n5925) );
ms00f80  l1247 ( .o(net_6580), .ck(clk), .d(n5930) );
ms00f80  l1248 ( .o(net_7127), .ck(clk), .d(n5934) );
ms00f80  l1249 ( .o(_net_7553), .ck(clk), .d(n5938) );
ms00f80  l1250 ( .o(net_6887), .ck(clk), .d(n5943) );
ms00f80  l1251 ( .o(net_6562), .ck(clk), .d(n5947) );
ms00f80  l1252 ( .o(net_6973), .ck(clk), .d(n5951) );
ms00f80  l1253 ( .o(net_6255), .ck(clk), .d(n5955) );
ms00f80  l1254 ( .o(_net_6006), .ck(clk), .d(n5960) );
ms00f80  l1255 ( .o(_net_7798), .ck(clk), .d(n5964) );
ms00f80  l1256 ( .o(net_7056), .ck(clk), .d(n5968) );
ms00f80  l1257 ( .o(_net_7360), .ck(clk), .d(n5973) );
ms00f80  l1258 ( .o(net_6618), .ck(clk), .d(n5978) );
ms00f80  l1259 ( .o(_net_6689), .ck(clk), .d(n5982) );
ms00f80  l1260 ( .o(_net_6410), .ck(clk), .d(n5987) );
ms00f80  l1261 ( .o(_net_7357), .ck(clk), .d(n5992) );
ms00f80  l1262 ( .o(_net_6066), .ck(clk), .d(n5997) );
ms00f80  l1263 ( .o(net_7712), .ck(clk), .d(n6002) );
ms00f80  l1264 ( .o(net_7115), .ck(clk), .d(n6006) );
ms00f80  l1265 ( .o(net_6497), .ck(clk), .d(n6009) );
ms00f80  l1266 ( .o(net_5861), .ck(clk), .d(n6014) );
ms00f80  l1267 ( .o(net_6314), .ck(clk), .d(n6019) );
ms00f80  l1268 ( .o(_net_7596), .ck(clk), .d(n6024) );
ms00f80  l1269 ( .o(_net_6081), .ck(clk), .d(n6029) );
ms00f80  l1270 ( .o(net_7125), .ck(clk), .d(n6034) );
ms00f80  l1271 ( .o(net_251), .ck(clk), .d(n6038) );
ms00f80  l1272 ( .o(net_6733), .ck(clk), .d(n6043) );
ms00f80  l1273 ( .o(net_6362), .ck(clk), .d(n6047) );
ms00f80  l1274 ( .o(_net_6132), .ck(clk), .d(n6052) );
ms00f80  l1275 ( .o(net_6802), .ck(clk), .d(n6056) );
ms00f80  l1276 ( .o(_net_7482), .ck(clk), .d(n6061) );
ms00f80  l1277 ( .o(net_6466), .ck(clk), .d(n6066) );
ms00f80  l1278 ( .o(net_6630), .ck(clk), .d(n6069) );
ms00f80  l1279 ( .o(_net_6558), .ck(clk), .d(n6074) );
ms00f80  l1280 ( .o(_net_7796), .ck(clk), .d(n6078) );
ms00f80  l1281 ( .o(net_261), .ck(clk), .d(n6083) );
ms00f80  l1282 ( .o(net_6054), .ck(clk), .d(n6088) );
ms00f80  l1283 ( .o(_net_7405), .ck(clk), .d(n6093) );
ms00f80  l1284 ( .o(net_6335), .ck(clk), .d(n6098) );
ms00f80  l1285 ( .o(net_6763), .ck(clk), .d(n6102) );
ms00f80  l1286 ( .o(net_6686), .ck(clk), .d(n6106) );
ms00f80  l1287 ( .o(net_7372), .ck(clk), .d(n6110) );
ms00f80  l1288 ( .o(net_6804), .ck(clk), .d(n6114) );
ms00f80  l1289 ( .o(_net_6181), .ck(clk), .d(n6119) );
ms00f80  l1290 ( .o(_net_7729), .ck(clk), .d(n6124) );
ms00f80  l1291 ( .o(net_7038), .ck(clk), .d(n6128) );
ms00f80  l1292 ( .o(_net_7808), .ck(clk), .d(n6132) );
ms00f80  l1293 ( .o(net_6385), .ck(clk), .d(n6136) );
ms00f80  l1294 ( .o(_net_7681), .ck(clk), .d(n6140) );
ms00f80  l1295 ( .o(net_6594), .ck(clk), .d(n6145) );
ms00f80  l1296 ( .o(net_274), .ck(clk), .d(n6148) );
ms00f80  l1297 ( .o(_net_6293), .ck(clk), .d(n6153) );
ms00f80  l1298 ( .o(net_6892), .ck(clk), .d(n6158) );
ms00f80  l1299 ( .o(net_7083), .ck(clk), .d(n6161) );
ms00f80  l1300 ( .o(_net_6209), .ck(clk), .d(n6166) );
ms00f80  l1301 ( .o(_net_6071), .ck(clk), .d(n6171) );
ms00f80  l1302 ( .o(net_6301), .ck(clk), .d(n6176) );
ms00f80  l1303 ( .o(net_6309), .ck(clk), .d(n6181) );
ms00f80  l1304 ( .o(_net_6124), .ck(clk), .d(n6186) );
ms00f80  l1305 ( .o(_net_6149), .ck(clk), .d(n6191) );
ms00f80  l1306 ( .o(net_6508), .ck(clk), .d(n6195) );
ms00f80  l1307 ( .o(_net_7693), .ck(clk), .d(n6200) );
ms00f80  l1308 ( .o(net_382), .ck(clk), .d(n6204) );
ms00f80  l1309 ( .o(_net_7254), .ck(clk), .d(n6209) );
ms00f80  l1310 ( .o(net_7385), .ck(clk), .d(n6214) );
ms00f80  l1311 ( .o(_net_6099), .ck(clk), .d(n6218) );
ms00f80  l1312 ( .o(net_7679), .ck(clk), .d(n6222) );
ms00f80  l1313 ( .o(net_186), .ck(clk), .d(n6227) );
ms00f80  l1314 ( .o(net_7739), .ck(clk), .d(n6231) );
ms00f80  l1315 ( .o(net_6629), .ck(clk), .d(n6235) );
ms00f80  l1316 ( .o(net_385), .ck(clk), .d(n6239) );
ms00f80  l1317 ( .o(_net_210), .ck(clk), .d(n6244) );
ms00f80  l1318 ( .o(_net_201), .ck(clk), .d(n6249) );
ms00f80  l1319 ( .o(net_6697), .ck(clk), .d(n6254) );
ms00f80  l1320 ( .o(net_6750), .ck(clk), .d(n6258) );
ms00f80  l1321 ( .o(_net_7801), .ck(clk), .d(n6261) );
ms00f80  l1322 ( .o(_net_7434), .ck(clk), .d(n6266) );
ms00f80  l1323 ( .o(net_167), .ck(clk), .d(n6271) );
ms00f80  l1324 ( .o(net_7752), .ck(clk), .d(n6276) );
ms00f80  l1325 ( .o(_net_174), .ck(clk), .d(n6281) );
ms00f80  l1326 ( .o(net_6212), .ck(clk), .d(n6285) );
ms00f80  l1327 ( .o(x718), .ck(clk), .d(n6290) );
ms00f80  l1328 ( .o(_net_7789), .ck(clk), .d(n6294) );
ms00f80  l1329 ( .o(net_7130), .ck(clk), .d(n6299) );
ms00f80  l1330 ( .o(net_7454), .ck(clk), .d(n6302) );
ms00f80  l1331 ( .o(net_302), .ck(clk), .d(n6306) );
ms00f80  l1332 ( .o(_net_5994), .ck(clk), .d(n6311) );
ms00f80  l1333 ( .o(net_7770), .ck(clk), .d(n6316) );
ms00f80  l1334 ( .o(_net_5922), .ck(clk), .d(n6319) );
ms00f80  l1335 ( .o(_net_6001), .ck(clk), .d(n6324) );
ms00f80  l1336 ( .o(net_7161), .ck(clk), .d(n6329) );
ms00f80  l1337 ( .o(net_381), .ck(clk), .d(n6332) );
ms00f80  l1338 ( .o(_net_6074), .ck(clk), .d(n6337) );
ms00f80  l1339 ( .o(net_6469), .ck(clk), .d(n6342) );
ms00f80  l1340 ( .o(_net_7353), .ck(clk), .d(n6346) );
ms00f80  l1341 ( .o(net_131), .ck(clk), .d(n6350) );
ms00f80  l1342 ( .o(net_6747), .ck(clk), .d(n6354) );
ms00f80  l1343 ( .o(net_6679), .ck(clk), .d(n6357) );
ms00f80  l1344 ( .o(_net_7440), .ck(clk), .d(n6362) );
ms00f80  l1345 ( .o(net_6439), .ck(clk), .d(n6367) );
ms00f80  l1346 ( .o(_net_7098), .ck(clk), .d(n6371) );
ms00f80  l1347 ( .o(net_7341), .ck(clk), .d(n6376) );
ms00f80  l1348 ( .o(_net_7661), .ck(clk), .d(n6381) );
ms00f80  l1349 ( .o(net_7117), .ck(clk), .d(n6386) );
ms00f80  l1350 ( .o(net_6361), .ck(clk), .d(n6390) );
ms00f80  l1351 ( .o(_net_6101), .ck(clk), .d(n6395) );
ms00f80  l1352 ( .o(net_6399), .ck(clk), .d(n6399) );
ms00f80  l1353 ( .o(net_6738), .ck(clk), .d(n6403) );
ms00f80  l1354 ( .o(net_6481), .ck(clk), .d(n6407) );
ms00f80  l1355 ( .o(_net_7438), .ck(clk), .d(n6411) );
ms00f80  l1356 ( .o(net_7208), .ck(clk), .d(n6415) );
ms00f80  l1357 ( .o(net_6625), .ck(clk), .d(n6419) );
ms00f80  l1358 ( .o(net_6383), .ck(clk), .d(n6423) );
ms00f80  l1359 ( .o(net_6826), .ck(clk), .d(n6427) );
ms00f80  l1360 ( .o(net_156), .ck(clk), .d(n6432) );
ms00f80  l1361 ( .o(net_7462), .ck(clk), .d(n6437) );
ms00f80  l1362 ( .o(net_7069), .ck(clk), .d(n6441) );
ms00f80  l1363 ( .o(net_6702), .ck(clk), .d(n6446) );
ms00f80  l1364 ( .o(_net_6692), .ck(clk), .d(n6450) );
ms00f80  l1365 ( .o(_net_7257), .ck(clk), .d(n6455) );
ms00f80  l1366 ( .o(net_6348), .ck(clk), .d(n6460) );
ms00f80  l1367 ( .o(net_6647), .ck(clk), .d(n6464) );
ms00f80  l1368 ( .o(net_6980), .ck(clk), .d(n6469) );
ms00f80  l1369 ( .o(net_6777), .ck(clk), .d(n6472) );
ms00f80  l1370 ( .o(net_7148), .ck(clk), .d(n6477) );
ms00f80  l1371 ( .o(net_6626), .ck(clk), .d(n6480) );
ms00f80  l1372 ( .o(net_6462), .ck(clk), .d(n6485) );
ms00f80  l1373 ( .o(net_7242), .ck(clk), .d(n6489) );
ms00f80  l1374 ( .o(net_205), .ck(clk), .d(n6493) );
ms00f80  l1375 ( .o(net_6355), .ck(clk), .d(n6498) );
ms00f80  l1376 ( .o(net_7074), .ck(clk), .d(n6502) );
ms00f80  l1377 ( .o(net_6563), .ck(clk), .d(n6507) );
ms00f80  l1378 ( .o(net_6604), .ck(clk), .d(n6511) );
ms00f80  l1379 ( .o(net_6836), .ck(clk), .d(n6515) );
ms00f80  l1380 ( .o(net_6866), .ck(clk), .d(n6519) );
ms00f80  l1381 ( .o(_net_7805), .ck(clk), .d(n6522) );
ms00f80  l1382 ( .o(_net_5857), .ck(clk), .d(n6527) );
ms00f80  l1383 ( .o(net_330), .ck(clk), .d(n6531) );
ms00f80  l1384 ( .o(net_7606), .ck(clk), .d(n6535) );
ms00f80  l1385 ( .o(_net_6126), .ck(clk), .d(n6540) );
ms00f80  l1386 ( .o(_net_118), .ck(clk), .d(n6545) );
ms00f80  l1387 ( .o(net_7397), .ck(clk), .d(n6550) );
ms00f80  l1388 ( .o(net_6713), .ck(clk), .d(n6554) );
ms00f80  l1389 ( .o(_net_7654), .ck(clk), .d(n6558) );
ms00f80  l1390 ( .o(net_6846), .ck(clk), .d(n6563) );
ms00f80  l1391 ( .o(net_6382), .ck(clk), .d(n6566) );
ms00f80  l1392 ( .o(_net_6146), .ck(clk), .d(n6570) );
ms00f80  l1393 ( .o(net_7485), .ck(clk), .d(n6574) );
ms00f80  l1394 ( .o(net_6226), .ck(clk), .d(n6578) );
ms00f80  l1395 ( .o(net_386), .ck(clk), .d(n6583) );
ms00f80  l1396 ( .o(net_6814), .ck(clk), .d(n6586) );
ms00f80  l1397 ( .o(net_157), .ck(clk), .d(n6591) );
ms00f80  l1398 ( .o(_net_6119), .ck(clk), .d(n6596) );
ms00f80  l1399 ( .o(_net_7448), .ck(clk), .d(n6601) );
ms00f80  l1400 ( .o(_net_5976), .ck(clk), .d(n6606) );
ms00f80  l1401 ( .o(net_6272), .ck(clk), .d(n6611) );
ms00f80  l1402 ( .o(net_6917), .ck(clk), .d(n6615) );
ms00f80  l1403 ( .o(net_7163), .ck(clk), .d(n6619) );
ms00f80  l1404 ( .o(net_168), .ck(clk), .d(n6624) );
ms00f80  l1405 ( .o(net_6261), .ck(clk), .d(n6629) );
ms00f80  l1406 ( .o(_net_6170), .ck(clk), .d(n6634) );
ms00f80  l1407 ( .o(net_7187), .ck(clk), .d(n6638) );
ms00f80  l1408 ( .o(net_6003), .ck(clk), .d(n6643) );
ms00f80  l1409 ( .o(net_7145), .ck(clk), .d(n6648) );
ms00f80  l1410 ( .o(_net_124), .ck(clk), .d(n6652) );
ms00f80  l1411 ( .o(net_7638), .ck(clk), .d(n6656) );
ms00f80  l1412 ( .o(net_6424), .ck(clk), .d(n6661) );
ms00f80  l1413 ( .o(_net_6129), .ck(clk), .d(n6665) );
ms00f80  l1414 ( .o(net_315), .ck(clk), .d(n6669) );
ms00f80  l1415 ( .o(net_6834), .ck(clk), .d(n6674) );
ms00f80  l1416 ( .o(net_6708), .ck(clk), .d(n6678) );
ms00f80  l1417 ( .o(_net_278), .ck(clk), .d(n6682) );
ms00f80  l1418 ( .o(net_6997), .ck(clk), .d(n6687) );
ms00f80  l1419 ( .o(x681), .ck(clk), .d(n6691) );
ms00f80  l1420 ( .o(_net_7623), .ck(clk), .d(n6695) );
ms00f80  l1421 ( .o(net_6353), .ck(clk), .d(n6700) );
ms00f80  l1422 ( .o(net_7029), .ck(clk), .d(n6704) );
ms00f80  l1423 ( .o(_net_7279), .ck(clk), .d(n6709) );
ms00f80  l1424 ( .o(net_6655), .ck(clk), .d(n6713) );
ms00f80  l1425 ( .o(net_6793), .ck(clk), .d(n6717) );
ms00f80  l1426 ( .o(net_7345), .ck(clk), .d(n6722) );
ms00f80  l1427 ( .o(_net_6113), .ck(clk), .d(n6727) );
ms00f80  l1428 ( .o(net_7180), .ck(clk), .d(n6732) );
ms00f80  l1429 ( .o(net_136), .ck(clk), .d(n6736) );
ms00f80  l1430 ( .o(_net_7620), .ck(clk), .d(n6741) );
ms00f80  l1431 ( .o(net_7549), .ck(clk), .d(n6746) );
ms00f80  l1432 ( .o(net_147), .ck(clk), .d(n6749) );
ms00f80  l1433 ( .o(net_6894), .ck(clk), .d(n6752) );
ms00f80  l1434 ( .o(net_314), .ck(clk), .d(n6756) );
ms00f80  l1435 ( .o(net_6728), .ck(clk), .d(n6761) );
ms00f80  l1436 ( .o(_net_6136), .ck(clk), .d(n6765) );
ms00f80  l1437 ( .o(net_6830), .ck(clk), .d(n6770) );
ms00f80  l1438 ( .o(_net_6117), .ck(clk), .d(n6774) );
ms00f80  l1439 ( .o(_net_7723), .ck(clk), .d(n6779) );
ms00f80  l1440 ( .o(net_6519), .ck(clk), .d(n6783) );
ms00f80  l1441 ( .o(_net_7446), .ck(clk), .d(n6788) );
ms00f80  l1442 ( .o(net_7394), .ck(clk), .d(n6793) );
ms00f80  l1443 ( .o(net_6933), .ck(clk), .d(n6796) );
ms00f80  l1444 ( .o(_net_7258), .ck(clk), .d(n6801) );
ms00f80  l1445 ( .o(net_6990), .ck(clk), .d(n6806) );
ms00f80  l1446 ( .o(net_6526), .ck(clk), .d(n6809) );
ms00f80  l1447 ( .o(net_7033), .ck(clk), .d(n6813) );
ms00f80  l1448 ( .o(_net_7700), .ck(clk), .d(n6818) );
ms00f80  l1449 ( .o(net_301), .ck(clk), .d(n6822) );
ms00f80  l1450 ( .o(net_7044), .ck(clk), .d(n6826) );
ms00f80  l1451 ( .o(_net_7584), .ck(clk), .d(n6831) );
ms00f80  l1452 ( .o(net_7025), .ck(clk), .d(n6836) );
ms00f80  l1453 ( .o(_net_5993), .ck(clk), .d(n6840) );
ms00f80  l1454 ( .o(_net_7325), .ck(clk), .d(n6845) );
ms00f80  l1455 ( .o(net_240), .ck(clk), .d(n6850) );
ms00f80  l1456 ( .o(_net_5990), .ck(clk), .d(n6855) );
ms00f80  l1457 ( .o(net_6470), .ck(clk), .d(n6860) );
ms00f80  l1458 ( .o(net_7166), .ck(clk), .d(n6863) );
ms00f80  l1459 ( .o(net_7193), .ck(clk), .d(n6867) );
ms00f80  l1460 ( .o(net_216), .ck(clk), .d(n6872) );
ms00f80  l1461 ( .o(net_7209), .ck(clk), .d(n6876) );
ms00f80  l1462 ( .o(_net_6161), .ck(clk), .d(n6881) );
ms00f80  l1463 ( .o(net_6712), .ck(clk), .d(n6886) );
ms00f80  l1464 ( .o(_net_7427), .ck(clk), .d(n6890) );
ms00f80  l1465 ( .o(net_7009), .ck(clk), .d(n6895) );
ms00f80  l1466 ( .o(net_6607), .ck(clk), .d(n6899) );
ms00f80  l1467 ( .o(net_340), .ck(clk), .d(n6902) );
ms00f80  l1468 ( .o(net_6904), .ck(clk), .d(n6906) );
ms00f80  l1469 ( .o(net_7053), .ck(clk), .d(n6910) );
ms00f80  l1470 ( .o(_net_215), .ck(clk), .d(n6915) );
ms00f80  l1471 ( .o(net_7309), .ck(clk), .d(n6919) );
ms00f80  l1472 ( .o(_net_7443), .ck(clk), .d(n6924) );
ms00f80  l1473 ( .o(net_244), .ck(clk), .d(n6929) );
ms00f80  l1474 ( .o(net_7150), .ck(clk), .d(n6934) );
ms00f80  l1475 ( .o(_net_114), .ck(clk), .d(n6938) );
ms00f80  l1476 ( .o(_net_7589), .ck(clk), .d(n6943) );
ms00f80  l1477 ( .o(net_375), .ck(clk), .d(n6947) );
ms00f80  l1478 ( .o(_net_7500), .ck(clk), .d(n6952) );
ms00f80  l1479 ( .o(net_6587), .ck(clk), .d(n6957) );
ms00f80  l1480 ( .o(net_149), .ck(clk), .d(n6960) );
ms00f80  l1481 ( .o(_net_6098), .ck(clk), .d(n6964) );
ms00f80  l1482 ( .o(net_194), .ck(clk), .d(n6969) );
ms00f80  l1483 ( .o(net_7245), .ck(clk), .d(n6974) );
ms00f80  l1484 ( .o(net_7051), .ck(clk), .d(n6977) );
ms00f80  l1485 ( .o(net_6342), .ck(clk), .d(n6982) );
ms00f80  l1486 ( .o(net_7172), .ck(clk), .d(n6986) );
ms00f80  l1487 ( .o(net_6495), .ck(clk), .d(n6990) );
ms00f80  l1488 ( .o(_net_7256), .ck(clk), .d(n6995) );
ms00f80  l1489 ( .o(_net_281), .ck(clk), .d(n7000) );
ms00f80  l1490 ( .o(net_6621), .ck(clk), .d(n7005) );
ms00f80  l1491 ( .o(net_6597), .ck(clk), .d(n7009) );
ms00f80  l1492 ( .o(_net_7408), .ck(clk), .d(n7013) );
ms00f80  l1493 ( .o(_net_6140), .ck(clk), .d(n7018) );
ms00f80  l1494 ( .o(net_222), .ck(clk), .d(n7023) );
ms00f80  l1495 ( .o(net_6902), .ck(clk), .d(n7027) );
ms00f80  l1496 ( .o(_net_7298), .ck(clk), .d(n7032) );
ms00f80  l1497 ( .o(net_306), .ck(clk), .d(n7036) );
ms00f80  l1498 ( .o(net_6889), .ck(clk), .d(n7041) );
ms00f80  l1499 ( .o(net_6378), .ck(clk), .d(n7045) );
ms00f80  l1500 ( .o(net_6394), .ck(clk), .d(n7049) );
ms00f80  l1501 ( .o(_net_7579), .ck(clk), .d(n7053) );
ms00f80  l1502 ( .o(_net_7268), .ck(clk), .d(n7058) );
ms00f80  l1503 ( .o(net_6769), .ck(clk), .d(n7062) );
ms00f80  l1504 ( .o(_net_6122), .ck(clk), .d(n7067) );
ms00f80  l1505 ( .o(_net_7761), .ck(clk), .d(n7072) );
ms00f80  l1506 ( .o(_net_6285), .ck(clk), .d(n7077) );
ms00f80  l1507 ( .o(net_6872), .ck(clk), .d(n7082) );
ms00f80  l1508 ( .o(net_7460), .ck(clk), .d(n7085) );
ms00f80  l1509 ( .o(net_6673), .ck(clk), .d(n7089) );
ms00f80  l1510 ( .o(net_383), .ck(clk), .d(n7093) );
ms00f80  l1511 ( .o(net_7152), .ck(clk), .d(n7098) );
ms00f80  l1512 ( .o(_net_193), .ck(clk), .d(n7102) );
ms00f80  l1513 ( .o(net_7769), .ck(clk), .d(n7107) );
ms00f80  l1514 ( .o(net_7088), .ck(clk), .d(n7111) );
ms00f80  l1515 ( .o(net_6329), .ck(clk), .d(n7116) );
ms00f80  l1516 ( .o(net_6498), .ck(clk), .d(n7120) );
ms00f80  l1517 ( .o(net_6561), .ck(clk), .d(n7125) );
ms00f80  l1518 ( .o(net_6660), .ck(clk), .d(n7128) );
ms00f80  l1519 ( .o(_net_7705), .ck(clk), .d(n7133) );
ms00f80  l1520 ( .o(_net_5848), .ck(clk), .d(n7138) );
ms00f80  l1521 ( .o(net_7496), .ck(clk), .d(n7142) );
ms00f80  l1522 ( .o(net_6249), .ck(clk), .d(n7147) );
ms00f80  l1523 ( .o(net_6948), .ck(clk), .d(n7151) );
ms00f80  l1524 ( .o(net_7226), .ck(clk), .d(n7155) );
ms00f80  l1525 ( .o(net_6862), .ck(clk), .d(n7160) );
ms00f80  l1526 ( .o(x195), .ck(clk), .d(n7164) );
ms00f80  l1527 ( .o(net_6235), .ck(clk), .d(n7167) );
ms00f80  l1528 ( .o(_net_5979), .ck(clk), .d(n7172) );
ms00f80  l1529 ( .o(net_161), .ck(clk), .d(n7177) );
ms00f80  l1530 ( .o(net_7543), .ck(clk), .d(n7182) );
ms00f80  l1531 ( .o(net_7307), .ck(clk), .d(n7185) );
ms00f80  l1532 ( .o(net_6430), .ck(clk), .d(n7190) );
ms00f80  l1533 ( .o(_net_6554), .ck(clk), .d(n7194) );
ms00f80  l1534 ( .o(net_7238), .ck(clk), .d(n7199) );
ms00f80  l1535 ( .o(net_6477), .ck(clk), .d(n7203) );
ms00f80  l1536 ( .o(_net_6080), .ck(clk), .d(n7207) );
ms00f80  l1537 ( .o(net_6559), .ck(clk), .d(n7212) );
ms00f80  l1538 ( .o(_net_7361), .ck(clk), .d(n7216) );
ms00f80  l1539 ( .o(net_6211), .ck(clk), .d(n7221) );
ms00f80  l1540 ( .o(_net_6200), .ck(clk), .d(n7226) );
ms00f80  l1541 ( .o(net_7090), .ck(clk), .d(n7230) );
ms00f80  l1542 ( .o(_net_6295), .ck(clk), .d(n7235) );
ms00f80  l1543 ( .o(_net_6145), .ck(clk), .d(n7240) );
ms00f80  l1544 ( .o(_net_6423), .ck(clk), .d(n7245) );
ms00f80  l1545 ( .o(net_7807), .ck(clk), .d(n7249) );
ms00f80  l1546 ( .o(net_6801), .ck(clk), .d(n7252) );
ms00f80  l1547 ( .o(_net_7791), .ck(clk), .d(n7256) );
ms00f80  l1548 ( .o(net_6627), .ck(clk), .d(n7260) );
ms00f80  l1549 ( .o(_net_6402), .ck(clk), .d(n7265) );
ms00f80  l1550 ( .o(_net_6151), .ck(clk), .d(n7270) );
ms00f80  l1551 ( .o(_net_6291), .ck(clk), .d(n7275) );
ms00f80  l1552 ( .o(_net_6026), .ck(clk), .d(n7280) );
ms00f80  l1553 ( .o(net_6511), .ck(clk), .d(n7284) );
ms00f80  l1554 ( .o(net_342), .ck(clk), .d(n7288) );
ms00f80  l1555 ( .o(_net_7816), .ck(clk), .d(n7292) );
ms00f80  l1556 ( .o(_net_6028), .ck(clk), .d(n7297) );
ms00f80  l1557 ( .o(_net_6288), .ck(clk), .d(n7302) );
ms00f80  l1558 ( .o(_net_7697), .ck(clk), .d(n7307) );
ms00f80  l1559 ( .o(net_6869), .ck(clk), .d(n7312) );
ms00f80  l1560 ( .o(net_6374), .ck(clk), .d(n7316) );
ms00f80  l1561 ( .o(_net_7365), .ck(clk), .d(n7321) );
ms00f80  l1562 ( .o(net_6715), .ck(clk), .d(n7326) );
ms00f80  l1563 ( .o(net_6264), .ck(clk), .d(n7330) );
ms00f80  l1564 ( .o(net_5860), .ck(clk), .d(n7335) );
ms00f80  l1565 ( .o(_net_6179), .ck(clk), .d(n7340) );
ms00f80  l1566 ( .o(net_7173), .ck(clk), .d(n7344) );
ms00f80  l1567 ( .o(net_6193), .ck(clk), .d(n7349) );
ms00f80  l1568 ( .o(net_250), .ck(clk), .d(n7354) );
ms00f80  l1569 ( .o(net_7008), .ck(clk), .d(n7359) );
ms00f80  l1570 ( .o(net_185), .ck(clk), .d(n7363) );
ms00f80  l1571 ( .o(net_6317), .ck(clk), .d(n7368) );
ms00f80  l1572 ( .o(net_7065), .ck(clk), .d(n7372) );
ms00f80  l1573 ( .o(net_6228), .ck(clk), .d(n7376) );
ms00f80  l1574 ( .o(_net_7666), .ck(clk), .d(n7381) );
ms00f80  l1575 ( .o(_net_6105), .ck(clk), .d(n7386) );
ms00f80  l1576 ( .o(net_7118), .ck(clk), .d(n7391) );
ms00f80  l1577 ( .o(_net_117), .ck(clk), .d(n7395) );
ms00f80  l1578 ( .o(_net_7473), .ck(clk), .d(n7400) );
ms00f80  l1579 ( .o(net_6503), .ck(clk), .d(n7404) );
ms00f80  l1580 ( .o(net_7054), .ck(clk), .d(n7408) );
ms00f80  l1581 ( .o(net_6994), .ck(clk), .d(n7413) );
ms00f80  l1582 ( .o(net_6257), .ck(clk), .d(n7417) );
ms00f80  l1583 ( .o(_net_6957), .ck(clk), .d(n7422) );
ms00f80  l1584 ( .o(net_6345), .ck(clk), .d(n7427) );
ms00f80  l1585 ( .o(_net_7757), .ck(clk), .d(n7432) );
ms00f80  l1586 ( .o(_net_6069), .ck(clk), .d(n7437) );
ms00f80  l1587 ( .o(net_6700), .ck(clk), .d(n7442) );
ms00f80  l1588 ( .o(net_6696), .ck(clk), .d(n7446) );
ms00f80  l1589 ( .o(net_6740), .ck(clk), .d(n7450) );
ms00f80  l1590 ( .o(_net_6007), .ck(clk), .d(n7454) );
ms00f80  l1591 ( .o(_net_7263), .ck(clk), .d(n7459) );
ms00f80  l1592 ( .o(net_7216), .ck(clk), .d(n7463) );
ms00f80  l1593 ( .o(net_6337), .ck(clk), .d(n7468) );
ms00f80  l1594 ( .o(_net_6222), .ck(clk), .d(n7473) );
ms00f80  l1595 ( .o(_net_7351), .ck(clk), .d(n7478) );
ms00f80  l1596 ( .o(net_7077), .ck(clk), .d(n7482) );
ms00f80  l1597 ( .o(_net_6962), .ck(clk), .d(n7487) );
ms00f80  l1598 ( .o(net_6726), .ck(clk), .d(n7492) );
ms00f80  l1599 ( .o(_net_6068), .ck(clk), .d(n7496) );
ms00f80  l1600 ( .o(_net_264), .ck(clk), .d(n7501) );
ms00f80  l1601 ( .o(net_348), .ck(clk), .d(n7505) );
ms00f80  l1602 ( .o(net_6774), .ck(clk), .d(n7509) );
ms00f80  l1603 ( .o(net_6550), .ck(clk), .d(n7513) );
ms00f80  l1604 ( .o(_net_7471), .ck(clk), .d(n7518) );
ms00f80  l1605 ( .o(net_7211), .ck(clk), .d(n7522) );
ms00f80  l1606 ( .o(net_6451), .ck(clk), .d(n7527) );
ms00f80  l1607 ( .o(net_7210), .ck(clk), .d(n7530) );
ms00f80  l1608 ( .o(net_6757), .ck(clk), .d(n7535) );
ms00f80  l1609 ( .o(x476), .ck(clk), .d(n7539) );
ms00f80  l1610 ( .o(_net_177), .ck(clk), .d(n7543) );
ms00f80  l1611 ( .o(net_243), .ck(clk), .d(n7548) );
ms00f80  l1612 ( .o(net_6266), .ck(clk), .d(n7553) );
ms00f80  l1613 ( .o(_net_7381), .ck(clk), .d(n7558) );
ms00f80  l1614 ( .o(_net_7293), .ck(clk), .d(n7563) );
ms00f80  l1615 ( .o(_net_7824), .ck(clk), .d(n7567) );
ms00f80  l1616 ( .o(_net_6127), .ck(clk), .d(n7572) );
ms00f80  l1617 ( .o(_net_6319), .ck(clk), .d(n7577) );
ms00f80  l1618 ( .o(net_6811), .ck(clk), .d(n7581) );
ms00f80  l1619 ( .o(_net_6033), .ck(clk), .d(n7586) );
ms00f80  l1620 ( .o(_net_127), .ck(clk), .d(n7591) );
ms00f80  l1621 ( .o(x187), .ck(clk), .d(n7596) );
ms00f80  l1622 ( .o(net_7494), .ck(clk), .d(n7599) );
ms00f80  l1623 ( .o(net_6716), .ck(clk), .d(n7604) );
ms00f80  l1624 ( .o(_net_6959), .ck(clk), .d(n7608) );
ms00f80  l1625 ( .o(net_199), .ck(clk), .d(n7613) );
ms00f80  l1626 ( .o(net_7392), .ck(clk), .d(n7618) );
ms00f80  l1627 ( .o(_net_6207), .ck(clk), .d(n7622) );
ms00f80  l1628 ( .o(net_7489), .ck(clk), .d(n7626) );
ms00f80  l1629 ( .o(_net_7331), .ck(clk), .d(n7631) );
ms00f80  l1630 ( .o(net_7668), .ck(clk), .d(n7635) );
ms00f80  l1631 ( .o(_net_5999), .ck(clk), .d(n7640) );
ms00f80  l1632 ( .o(net_341), .ck(clk), .d(n7644) );
ms00f80  l1633 ( .o(net_6299), .ck(clk), .d(n7649) );
ms00f80  l1634 ( .o(net_7139), .ck(clk), .d(n7654) );
ms00f80  l1635 ( .o(net_6467), .ck(clk), .d(n7658) );
ms00f80  l1636 ( .o(net_7486), .ck(clk), .d(n7661) );
ms00f80  l1637 ( .o(_net_7228), .ck(clk), .d(n7666) );
ms00f80  l1638 ( .o(_net_6091), .ck(clk), .d(n7671) );
ms00f80  l1639 ( .o(_net_6103), .ck(clk), .d(n7676) );
ms00f80  l1640 ( .o(_net_125), .ck(clk), .d(n7681) );
ms00f80  l1641 ( .o(net_231), .ck(clk), .d(n7686) );
ms00f80  l1642 ( .o(x38), .ck(clk), .d(n7691) );
ms00f80  l1643 ( .o(_net_5995), .ck(clk), .d(n7695) );
ms00f80  l1644 ( .o(net_6748), .ck(clk), .d(n7700) );
ms00f80  l1645 ( .o(net_6304), .ck(clk), .d(n7704) );
ms00f80  l1646 ( .o(net_6047), .ck(clk), .d(n7709) );
ms00f80  l1647 ( .o(net_7764), .ck(clk), .d(n7714) );
ms00f80  l1648 ( .o(net_6837), .ck(clk), .d(n7719) );
ms00f80  l1649 ( .o(_net_7273), .ck(clk), .d(n7723) );
ms00f80  l1650 ( .o(_net_7289), .ck(clk), .d(n7728) );
ms00f80  l1651 ( .o(net_7526), .ck(clk), .d(n7732) );
ms00f80  l1652 ( .o(x522), .ck(clk), .d(n7737) );
ms00f80  l1653 ( .o(_net_392), .ck(clk), .d(n7741) );
ms00f80  l1654 ( .o(_net_6828), .ck(clk), .d(n7746) );
ms00f80  l1655 ( .o(_net_7555), .ck(clk), .d(n7751) );
ms00f80  l1656 ( .o(net_6441), .ck(clk), .d(n7756) );
ms00f80  l1657 ( .o(net_7143), .ck(clk), .d(n7760) );
ms00f80  l1658 ( .o(net_7160), .ck(clk), .d(n7764) );
ms00f80  l1659 ( .o(_net_7699), .ck(clk), .d(n7768) );
ms00f80  l1660 ( .o(x420), .ck(clk), .d(n7773) );
ms00f80  l1661 ( .o(net_6397), .ck(clk), .d(n7776) );
ms00f80  l1662 ( .o(net_7059), .ck(clk), .d(n7779) );
ms00f80  l1663 ( .o(net_6710), .ck(clk), .d(n7784) );
ms00f80  l1664 ( .o(_net_6093), .ck(clk), .d(n7788) );
ms00f80  l1665 ( .o(_net_6049), .ck(clk), .d(n7793) );
ms00f80  l1666 ( .o(_net_7442), .ck(clk), .d(n7798) );
ms00f80  l1667 ( .o(net_6797), .ck(clk), .d(n7802) );
ms00f80  l1668 ( .o(net_6947), .ck(clk), .d(n7806) );
ms00f80  l1669 ( .o(net_6659), .ck(clk), .d(n7810) );
ms00f80  l1670 ( .o(net_6734), .ck(clk), .d(n7815) );
ms00f80  l1671 ( .o(net_6387), .ck(clk), .d(n7818) );
ms00f80  l1672 ( .o(_net_5974), .ck(clk), .d(n7822) );
ms00f80  l1673 ( .o(net_6528), .ck(clk), .d(n7826) );
ms00f80  l1674 ( .o(net_6566), .ck(clk), .d(n7831) );
ms00f80  l1675 ( .o(_net_7276), .ck(clk), .d(n7835) );
ms00f80  l1676 ( .o(net_6331), .ck(clk), .d(n7840) );
ms00f80  l1677 ( .o(x264), .ck(clk), .d(n7845) );
ms00f80  l1678 ( .o(net_327), .ck(clk), .d(n7848) );
ms00f80  l1679 ( .o(net_200), .ck(clk), .d(n7853) );
ms00f80  l1680 ( .o(_net_5971), .ck(clk), .d(n7858) );
ms00f80  l1681 ( .o(_net_6409), .ck(clk), .d(n7863) );
ms00f80  l1682 ( .o(net_358), .ck(clk), .d(n7867) );
ms00f80  l1683 ( .o(net_137), .ck(clk), .d(n7871) );
ms00f80  l1684 ( .o(net_6874), .ck(clk), .d(n7875) );
ms00f80  l1685 ( .o(net_7673), .ck(clk), .d(n7878) );
ms00f80  l1686 ( .o(net_6344), .ck(clk), .d(n7883) );
ms00f80  l1687 ( .o(_net_7484), .ck(clk), .d(n7888) );
ms00f80  l1688 ( .o(net_7249), .ck(clk), .d(n7893) );
ms00f80  l1689 ( .o(_net_5850), .ck(clk), .d(n7897) );
ms00f80  l1690 ( .o(_net_6031), .ck(clk), .d(n7902) );
ms00f80  l1691 ( .o(net_7192), .ck(clk), .d(n7906) );
ms00f80  l1692 ( .o(_net_6552), .ck(clk), .d(n7911) );
ms00f80  l1693 ( .o(net_6363), .ck(clk), .d(n7916) );
ms00f80  l1694 ( .o(net_311), .ck(clk), .d(n7920) );
ms00f80  l1695 ( .o(net_7456), .ck(clk), .d(n7924) );
ms00f80  l1696 ( .o(net_6568), .ck(clk), .d(n7929) );
ms00f80  l1697 ( .o(net_237), .ck(clk), .d(n7933) );
ms00f80  l1698 ( .o(net_6930), .ck(clk), .d(n7937) );
ms00f80  l1699 ( .o(net_7540), .ck(clk), .d(n7942) );
ms00f80  l1700 ( .o(net_335), .ck(clk), .d(n7945) );
ms00f80  l1701 ( .o(net_6056), .ck(clk), .d(n7950) );
ms00f80  l1702 ( .o(net_6724), .ck(clk), .d(n7955) );
ms00f80  l1703 ( .o(net_6232), .ck(clk), .d(n7958) );
ms00f80  l1704 ( .o(net_7078), .ck(clk), .d(n7962) );
ms00f80  l1705 ( .o(net_6992), .ck(clk), .d(n7967) );
ms00f80  l1706 ( .o(net_7491), .ck(clk), .d(n7970) );
ms00f80  l1707 ( .o(_net_5855), .ck(clk), .d(n7975) );
ms00f80  l1708 ( .o(net_158), .ck(clk), .d(n7980) );
ms00f80  l1709 ( .o(_net_7425), .ck(clk), .d(n7985) );
ms00f80  l1710 ( .o(net_6651), .ck(clk), .d(n7989) );
ms00f80  l1711 ( .o(net_6585), .ck(clk), .d(n7994) );
ms00f80  l1712 ( .o(net_7087), .ck(clk), .d(n7997) );
ms00f80  l1713 ( .o(net_6975), .ck(clk), .d(n8002) );
ms00f80  l1714 ( .o(net_379), .ck(clk), .d(n8005) );
ms00f80  l1715 ( .o(_net_5852), .ck(clk), .d(n8010) );
ms00f80  l1716 ( .o(net_7131), .ck(clk), .d(n8015) );
ms00f80  l1717 ( .o(_net_291), .ck(clk), .d(n8019) );
ms00f80  l1718 ( .o(_net_6287), .ck(clk), .d(n8024) );
ms00f80  l1719 ( .o(net_6542), .ck(clk), .d(n8028) );
ms00f80  l1720 ( .o(_net_6072), .ck(clk), .d(n8033) );
ms00f80  l1721 ( .o(net_7680), .ck(clk), .d(n8038) );
ms00f80  l1722 ( .o(net_7744), .ck(clk), .d(n8042) );
ms00f80  l1723 ( .o(net_6365), .ck(clk), .d(n8047) );
ms00f80  l1724 ( .o(net_344), .ck(clk), .d(n8051) );
ms00f80  l1725 ( .o(net_6988), .ck(clk), .d(n8056) );
ms00f80  l1726 ( .o(net_6919), .ck(clk), .d(n8059) );
ms00f80  l1727 ( .o(net_6968), .ck(clk), .d(n8064) );
ms00f80  l1728 ( .o(net_6675), .ck(clk), .d(n8067) );
ms00f80  l1729 ( .o(net_6614), .ck(clk), .d(n8072) );
ms00f80  l1730 ( .o(net_6924), .ck(clk), .d(n8075) );
ms00f80  l1731 ( .o(_net_7262), .ck(clk), .d(n8080) );
ms00f80  l1732 ( .o(net_6596), .ck(clk), .d(n8085) );
ms00f80  l1733 ( .o(net_285), .ck(clk), .d(n8088) );
ms00f80  l1734 ( .o(net_7036), .ck(clk), .d(n8092) );
ms00f80  l1735 ( .o(_net_7573), .ck(clk), .d(n8097) );
ms00f80  l1736 ( .o(_net_7499), .ck(clk), .d(n8102) );
ms00f80  l1737 ( .o(_net_7417), .ck(clk), .d(n8107) );
ms00f80  l1738 ( .o(_net_6115), .ck(clk), .d(n8112) );
ms00f80  l1739 ( .o(net_6798), .ck(clk), .d(n8116) );
ms00f80  l1740 ( .o(_net_7562), .ck(clk), .d(n8121) );
ms00f80  l1741 ( .o(net_6895), .ck(clk), .d(n8125) );
ms00f80  l1742 ( .o(_net_7291), .ck(clk), .d(n8130) );
ms00f80  l1743 ( .o(_net_7592), .ck(clk), .d(n8135) );
ms00f80  l1744 ( .o(net_7141), .ck(clk), .d(n8140) );
ms00f80  l1745 ( .o(net_6571), .ck(clk), .d(n8144) );
ms00f80  l1746 ( .o(net_6638), .ck(clk), .d(n8147) );
ms00f80  l1747 ( .o(_net_262), .ck(clk), .d(n8152) );
ms00f80  l1748 ( .o(net_7339), .ck(clk), .d(n8156) );
ms00f80  l1749 ( .o(net_242), .ck(clk), .d(n8161) );
ms00f80  l1750 ( .o(net_7715), .ck(clk), .d(n8166) );
ms00f80  l1751 ( .o(_net_221), .ck(clk), .d(n8170) );
ms00f80  l1752 ( .o(net_6682), .ck(clk), .d(n8174) );
ms00f80  l1753 ( .o(_net_180), .ck(clk), .d(n8179) );
ms00f80  l1754 ( .o(net_6767), .ck(clk), .d(n8183) );
ms00f80  l1755 ( .o(net_6835), .ck(clk), .d(n8188) );
ms00f80  l1756 ( .o(_net_7275), .ck(clk), .d(n8192) );
ms00f80  l1757 ( .o(net_275), .ck(clk), .d(n8197) );
ms00f80  l1758 ( .o(_net_6159), .ck(clk), .d(n8202) );
ms00f80  l1759 ( .o(net_6678), .ck(clk), .d(n8206) );
ms00f80  l1760 ( .o(net_7772), .ck(clk), .d(n8211) );
ms00f80  l1761 ( .o(_net_7702), .ck(clk), .d(n8216) );
ms00f80  l1762 ( .o(net_6390), .ck(clk), .d(n8220) );
ms00f80  l1763 ( .o(_net_7755), .ck(clk), .d(n8224) );
ms00f80  l1764 ( .o(net_6910), .ck(clk), .d(n8228) );
ms00f80  l1765 ( .o(net_7177), .ck(clk), .d(n8232) );
ms00f80  l1766 ( .o(_net_7580), .ck(clk), .d(n8237) );
ms00f80  l1767 ( .o(net_370), .ck(clk), .d(n8241) );
ms00f80  l1768 ( .o(net_6494), .ck(clk), .d(n8245) );
ms00f80  l1769 ( .o(net_6389), .ck(clk), .d(n8249) );
ms00f80  l1770 ( .o(_net_7432), .ck(clk), .d(n8253) );
ms00f80  l1771 ( .o(net_196), .ck(clk), .d(n8258) );
ms00f80  l1772 ( .o(net_7615), .ck(clk), .d(n8262) );
ms00f80  l1773 ( .o(net_7169), .ck(clk), .d(n8266) );
ms00f80  l1774 ( .o(net_6312), .ck(clk), .d(n8271) );
ms00f80  l1775 ( .o(net_6615), .ck(clk), .d(n8276) );
ms00f80  l1776 ( .o(net_7538), .ck(clk), .d(n8280) );
ms00f80  l1777 ( .o(_net_6413), .ck(clk), .d(n8284) );
ms00f80  l1778 ( .o(net_6321), .ck(clk), .d(n8289) );
ms00f80  l1779 ( .o(_net_7648), .ck(clk), .d(n8294) );
ms00f80  l1780 ( .o(_net_6020), .ck(clk), .d(n8299) );
ms00f80  l1781 ( .o(net_7045), .ck(clk), .d(n8303) );
ms00f80  l1782 ( .o(net_7181), .ck(clk), .d(n8307) );
ms00f80  l1783 ( .o(net_7186), .ck(clk), .d(n8311) );
ms00f80  l1784 ( .o(net_6853), .ck(clk), .d(n8316) );
ms00f80  l1785 ( .o(net_7138), .ck(clk), .d(n8320) );
ms00f80  l1786 ( .o(_net_6201), .ck(clk), .d(n8324) );
ms00f80  l1787 ( .o(net_6276), .ck(clk), .d(n8329) );
ms00f80  l1788 ( .o(net_6851), .ck(clk), .d(n8334) );
ms00f80  l1789 ( .o(net_143), .ck(clk), .d(n8337) );
ms00f80  l1790 ( .o(net_6809), .ck(clk), .d(n8340) );
ms00f80  l1791 ( .o(_net_6123), .ck(clk), .d(n8345) );
ms00f80  l1792 ( .o(net_7023), .ck(clk), .d(n8350) );
ms00f80  l1793 ( .o(_net_6823), .ck(clk), .d(n8354) );
ms00f80  l1794 ( .o(net_6427), .ck(clk), .d(n8359) );
ms00f80  l1795 ( .o(net_7605), .ck(clk), .d(n8362) );
ms00f80  l1796 ( .o(_net_189), .ck(clk), .d(n8367) );
ms00f80  l1797 ( .o(_net_7685), .ck(clk), .d(n8372) );
ms00f80  l1798 ( .o(_net_7735), .ck(clk), .d(n8377) );
ms00f80  l1799 ( .o(_net_7602), .ck(clk), .d(n8382) );
ms00f80  l1800 ( .o(_net_6027), .ck(clk), .d(n8387) );
ms00f80  l1801 ( .o(net_6425), .ck(clk), .d(n8392) );
ms00f80  l1802 ( .o(_net_7568), .ck(clk), .d(n8396) );
ms00f80  l1803 ( .o(net_7104), .ck(clk), .d(n8401) );
ms00f80  l1804 ( .o(_net_6958), .ck(clk), .d(n8405) );
ms00f80  l1805 ( .o(_net_7333), .ck(clk), .d(n8410) );
ms00f80  l1806 ( .o(net_7137), .ck(clk), .d(n8415) );
ms00f80  l1807 ( .o(net_6393), .ck(clk), .d(n8418) );
ms00f80  l1808 ( .o(net_7237), .ck(clk), .d(n8422) );
ms00f80  l1809 ( .o(_net_6089), .ck(clk), .d(n8426) );
ms00f80  l1810 ( .o(net_332), .ck(clk), .d(n8430) );
ms00f80  l1811 ( .o(x342), .ck(clk), .d(n8435) );
ms00f80  l1812 ( .o(_net_5924), .ck(clk), .d(n8438) );
ms00f80  l1813 ( .o(_net_7687), .ck(clk), .d(n8443) );
ms00f80  l1814 ( .o(net_7375), .ck(clk), .d(n8447) );
ms00f80  l1815 ( .o(net_7459), .ck(clk), .d(n8451) );
ms00f80  l1816 ( .o(net_6945), .ck(clk), .d(n8455) );
ms00f80  l1817 ( .o(net_6518), .ck(clk), .d(n8459) );
ms00f80  l1818 ( .o(net_6742), .ck(clk), .d(n8464) );
ms00f80  l1819 ( .o(net_7039), .ck(clk), .d(n8467) );
ms00f80  l1820 ( .o(_net_5961), .ck(clk), .d(n8472) );
ms00f80  l1821 ( .o(net_6754), .ck(clk), .d(n8477) );
ms00f80  l1822 ( .o(_net_7450), .ck(clk), .d(n8481) );
ms00f80  l1823 ( .o(_net_6178), .ck(clk), .d(n8486) );
ms00f80  l1824 ( .o(net_7020), .ck(clk), .d(n8491) );
ms00f80  l1825 ( .o(net_7212), .ck(clk), .d(n8494) );
ms00f80  l1826 ( .o(_net_6039), .ck(clk), .d(n8499) );
ms00f80  l1827 ( .o(net_6622), .ck(clk), .d(n8504) );
ms00f80  l1828 ( .o(_net_6557), .ck(clk), .d(n8508) );
ms00f80  l1829 ( .o(net_6744), .ck(clk), .d(n8513) );
ms00f80  l1830 ( .o(_net_7575), .ck(clk), .d(n8517) );
ms00f80  l1831 ( .o(net_6838), .ck(clk), .d(n8522) );
ms00f80  l1832 ( .o(_net_7349), .ck(clk), .d(n8526) );
ms00f80  l1833 ( .o(_net_7284), .ck(clk), .d(n8531) );
ms00f80  l1834 ( .o(net_6771), .ck(clk), .d(n8535) );
ms00f80  l1835 ( .o(net_239), .ck(clk), .d(n8540) );
ms00f80  l1836 ( .o(net_6499), .ck(clk), .d(n8544) );
ms00f80  l1837 ( .o(net_6707), .ck(clk), .d(n8549) );
ms00f80  l1838 ( .o(net_6792), .ck(clk), .d(n8552) );
ms00f80  l1839 ( .o(net_166), .ck(clk), .d(n8557) );
ms00f80  l1840 ( .o(net_6956), .ck(clk), .d(n8561) );
ms00f80  l1841 ( .o(net_6794), .ck(clk), .d(n8565) );
ms00f80  l1842 ( .o(_net_122), .ck(clk), .d(n8570) );
ms00f80  l1843 ( .o(net_6475), .ck(clk), .d(n8575) );
ms00f80  l1844 ( .o(net_350), .ck(clk), .d(n8578) );
ms00f80  l1845 ( .o(_net_6282), .ck(clk), .d(n8583) );
ms00f80  l1846 ( .o(net_7778), .ck(clk), .d(n8588) );
ms00f80  l1847 ( .o(_net_7695), .ck(clk), .d(n8593) );
ms00f80  l1848 ( .o(net_6695), .ck(clk), .d(n8598) );
ms00f80  l1849 ( .o(_net_7319), .ck(clk), .d(n8602) );
ms00f80  l1850 ( .o(net_181), .ck(clk), .d(n8607) );
ms00f80  l1851 ( .o(net_6463), .ck(clk), .d(n8612) );
ms00f80  l1852 ( .o(net_6360), .ck(clk), .d(n8616) );
ms00f80  l1853 ( .o(net_6831), .ck(clk), .d(n8621) );
ms00f80  l1854 ( .o(net_388), .ck(clk), .d(n8625) );
ms00f80  l1855 ( .o(net_151), .ck(clk), .d(n8628) );
ms00f80  l1856 ( .o(net_6683), .ck(clk), .d(n8632) );
ms00f80  l1857 ( .o(net_6013), .ck(clk), .d(n8637) );
ms00f80  l1858 ( .o(net_6756), .ck(clk), .d(n8641) );
ms00f80  l1859 ( .o(_net_6141), .ck(clk), .d(n8645) );
ms00f80  l1860 ( .o(net_6865), .ck(clk), .d(n8650) );
ms00f80  l1861 ( .o(net_6577), .ck(clk), .d(n8654) );
ms00f80  l1862 ( .o(net_6600), .ck(clk), .d(n8658) );
ms00f80  l1863 ( .o(net_198), .ck(clk), .d(n8662) );
ms00f80  l1864 ( .o(net_7373), .ck(clk), .d(n8666) );
ms00f80  l1865 ( .o(_net_7267), .ck(clk), .d(n8671) );
ms00f80  l1866 ( .o(_net_6418), .ck(clk), .d(n8676) );
ms00f80  l1867 ( .o(net_6891), .ck(clk), .d(n8681) );
ms00f80  l1868 ( .o(net_6722), .ck(clk), .d(n8685) );
ms00f80  l1869 ( .o(_net_7627), .ck(clk), .d(n8689) );
ms00f80  l1870 ( .o(_net_6144), .ck(clk), .d(n8694) );
ms00f80  l1871 ( .o(_net_7811), .ck(clk), .d(n8698) );
ms00f80  l1872 ( .o(_net_6010), .ck(clk), .d(n8703) );
ms00f80  l1873 ( .o(x538), .ck(clk), .d(n8708) );
ms00f80  l1874 ( .o(net_7521), .ck(clk), .d(n8711) );
ms00f80  l1875 ( .o(net_333), .ck(clk), .d(n8715) );
ms00f80  l1876 ( .o(_net_7477), .ck(clk), .d(n8720) );
ms00f80  l1877 ( .o(_net_6824), .ck(clk), .d(n8725) );
ms00f80  l1878 ( .o(_net_6109), .ck(clk), .d(n8730) );
ms00f80  l1879 ( .o(net_7340), .ck(clk), .d(n8734) );
ms00f80  l1880 ( .o(net_7389), .ck(clk), .d(n8739) );
ms00f80  l1881 ( .o(_net_6043), .ck(clk), .d(n8743) );
ms00f80  l1882 ( .o(_net_7476), .ck(clk), .d(n8748) );
ms00f80  l1883 ( .o(_net_7585), .ck(clk), .d(n8753) );
ms00f80  l1884 ( .o(net_6234), .ck(clk), .d(n8757) );
ms00f80  l1885 ( .o(_net_6289), .ck(clk), .d(n8762) );
ms00f80  l1886 ( .o(net_7110), .ck(clk), .d(n8767) );
ms00f80  l1887 ( .o(net_387), .ck(clk), .d(n8771) );
ms00f80  l1888 ( .o(_net_7230), .ck(clk), .d(n8775) );
ms00f80  l1889 ( .o(_net_7265), .ck(clk), .d(n8780) );
ms00f80  l1890 ( .o(_net_7818), .ck(clk), .d(n8784) );
ms00f80  l1891 ( .o(net_6046), .ck(clk), .d(n8788) );
ms00f80  l1892 ( .o(net_6882), .ck(clk), .d(n8793) );
ms00f80  l1893 ( .o(net_6457), .ck(clk), .d(n8797) );
ms00f80  l1894 ( .o(net_7043), .ck(clk), .d(n8800) );
ms00f80  l1895 ( .o(net_6982), .ck(clk), .d(n8805) );
ms00f80  l1896 ( .o(net_6417), .ck(clk), .d(n8809) );
ms00f80  l1897 ( .o(net_7064), .ck(clk), .d(n8813) );
ms00f80  l1898 ( .o(_net_7409), .ck(clk), .d(n8818) );
ms00f80  l1899 ( .o(net_7542), .ck(clk), .d(n8823) );
ms00f80  l1900 ( .o(net_6787), .ck(clk), .d(n8826) );
ms00f80  l1901 ( .o(net_195), .ck(clk), .d(n8831) );
ms00f80  l1902 ( .o(net_7046), .ck(clk), .d(n8835) );
ms00f80  l1903 ( .o(_net_7664), .ck(clk), .d(n8840) );
ms00f80  l1904 ( .o(_net_6048), .ck(clk), .d(n8845) );
ms00f80  l1905 ( .o(_net_228), .ck(clk), .d(n8850) );
ms00f80  l1906 ( .o(_net_7363), .ck(clk), .d(n8855) );
ms00f80  l1907 ( .o(_net_7625), .ck(clk), .d(n8860) );
ms00f80  l1908 ( .o(_net_7806), .ck(clk), .d(n8864) );
ms00f80  l1909 ( .o(_net_6186), .ck(clk), .d(n8869) );
ms00f80  l1910 ( .o(net_6217), .ck(clk), .d(n8873) );
ms00f80  l1911 ( .o(net_307), .ck(clk), .d(n8877) );
ms00f80  l1912 ( .o(net_6196), .ck(clk), .d(n8882) );
ms00f80  l1913 ( .o(net_7086), .ck(clk), .d(n8886) );
ms00f80  l1914 ( .o(net_7132), .ck(clk), .d(n8891) );
ms00f80  l1915 ( .o(_net_6298), .ck(clk), .d(n8895) );
ms00f80  l1916 ( .o(net_7302), .ck(clk), .d(n8899) );
ms00f80  l1917 ( .o(net_6549), .ck(clk), .d(n8903) );
ms00f80  l1918 ( .o(net_6315), .ck(clk), .d(n8908) );
ms00f80  l1919 ( .o(net_6531), .ck(clk), .d(n8912) );
ms00f80  l1920 ( .o(_net_6166), .ck(clk), .d(n8917) );
ms00f80  l1921 ( .o(_net_7787), .ck(clk), .d(n8922) );
ms00f80  l1922 ( .o(net_6504), .ck(clk), .d(n8926) );
ms00f80  l1923 ( .o(net_7243), .ck(clk), .d(n8931) );
ms00f80  l1924 ( .o(net_7368), .ck(clk), .d(n8934) );
ms00f80  l1925 ( .o(net_6458), .ck(clk), .d(n8939) );
ms00f80  l1926 ( .o(net_6262), .ck(clk), .d(n8943) );
ms00f80  l1927 ( .o(_net_7322), .ck(clk), .d(n8948) );
ms00f80  l1928 ( .o(_net_7451), .ck(clk), .d(n8953) );
ms00f80  l1929 ( .o(net_6326), .ck(clk), .d(n8958) );
ms00f80  l1930 ( .o(net_7544), .ck(clk), .d(n8963) );
ms00f80  l1931 ( .o(_net_209), .ck(clk), .d(n8967) );
ms00f80  l1932 ( .o(net_6534), .ck(clk), .d(n8971) );
ms00f80  l1933 ( .o(_net_7466), .ck(clk), .d(n8976) );
ms00f80  l1934 ( .o(net_6350), .ck(clk), .d(n8981) );
ms00f80  l1935 ( .o(_net_7581), .ck(clk), .d(n8986) );
ms00f80  l1936 ( .o(net_304), .ck(clk), .d(n8990) );
ms00f80  l1937 ( .o(_net_293), .ck(clk), .d(n8995) );
ms00f80  l1938 ( .o(_net_268), .ck(clk), .d(n9000) );
ms00f80  l1939 ( .o(_net_7783), .ck(clk), .d(n9005) );
ms00f80  l1940 ( .o(net_6582), .ck(clk), .d(n9010) );
ms00f80  l1941 ( .o(net_7017), .ck(clk), .d(n9014) );
ms00f80  l1942 ( .o(net_6230), .ck(clk), .d(n9017) );
ms00f80  l1943 ( .o(net_6445), .ck(clk), .d(n9022) );
ms00f80  l1944 ( .o(net_6932), .ck(clk), .d(n9025) );
ms00f80  l1945 ( .o(x249), .ck(clk), .d(n9030) );
ms00f80  l1946 ( .o(net_6864), .ck(clk), .d(n9034) );
ms00f80  l1947 ( .o(net_6937), .ck(clk), .d(n9037) );
ms00f80  l1948 ( .o(net_230), .ck(clk), .d(n9042) );
ms00f80  l1949 ( .o(net_7762), .ck(clk), .d(n9047) );
ms00f80  l1950 ( .o(_net_7423), .ck(clk), .d(n9052) );
ms00f80  l1951 ( .o(net_6966), .ck(clk), .d(n9057) );
ms00f80  l1952 ( .o(net_7305), .ck(clk), .d(n9060) );
ms00f80  l1953 ( .o(net_6984), .ck(clk), .d(n9065) );
ms00f80  l1954 ( .o(net_6306), .ck(clk), .d(n9069) );
ms00f80  l1955 ( .o(_net_115), .ck(clk), .d(n9074) );
ms00f80  l1956 ( .o(net_7101), .ck(clk), .d(n9079) );
ms00f80  l1957 ( .o(net_7084), .ck(clk), .d(n9082) );
ms00f80  l1958 ( .o(net_6649), .ck(clk), .d(n9086) );
ms00f80  l1959 ( .o(net_6270), .ck(clk), .d(n9091) );
ms00f80  l1960 ( .o(net_256), .ck(clk), .d(n9096) );
ms00f80  l1961 ( .o(_net_289), .ck(clk), .d(n9101) );
ms00f80  l1962 ( .o(_net_7716), .ck(clk), .d(n9106) );
ms00f80  l1963 ( .o(_net_7804), .ck(clk), .d(n9110) );
ms00f80  l1964 ( .o(_net_292), .ck(clk), .d(n9115) );
ms00f80  l1965 ( .o(net_7155), .ck(clk), .d(n9120) );
ms00f80  l1966 ( .o(_net_7558), .ck(clk), .d(n9124) );
ms00f80  l1967 ( .o(_net_7660), .ck(clk), .d(n9129) );
ms00f80  l1968 ( .o(net_6333), .ck(clk), .d(n9134) );
ms00f80  l1969 ( .o(net_6520), .ck(clk), .d(n9138) );
ms00f80  l1970 ( .o(net_6876), .ck(clk), .d(n9143) );
ms00f80  l1971 ( .o(net_6665), .ck(clk), .d(n9146) );
ms00f80  l1972 ( .o(net_162), .ck(clk), .d(n9151) );
ms00f80  l1973 ( .o(_net_7259), .ck(clk), .d(n9156) );
ms00f80  l1974 ( .o(net_318), .ck(clk), .d(n9160) );
ms00f80  l1975 ( .o(net_6911), .ck(clk), .d(n9164) );
ms00f80  l1976 ( .o(net_6565), .ck(clk), .d(n9169) );
ms00f80  l1977 ( .o(_net_6188), .ck(clk), .d(n9173) );
ms00f80  l1978 ( .o(net_6253), .ck(clk), .d(n9178) );
ms00f80  l1979 ( .o(net_6492), .ck(clk), .d(n9182) );
ms00f80  l1980 ( .o(_net_7260), .ck(clk), .d(n9187) );
ms00f80  l1981 ( .o(_net_172), .ck(clk), .d(n9192) );
ms00f80  l1982 ( .o(net_328), .ck(clk), .d(n9196) );
ms00f80  l1983 ( .o(_net_7682), .ck(clk), .d(n9201) );
ms00f80  l1984 ( .o(_net_5986), .ck(clk), .d(n9206) );
ms00f80  l1985 ( .o(net_7776), .ck(clk), .d(n9211) );
ms00f80  l1986 ( .o(net_7367), .ck(clk), .d(n9215) );
ms00f80  l1987 ( .o(_net_6094), .ck(clk), .d(n9220) );
ms00f80  l1988 ( .o(net_7156), .ck(clk), .d(n9225) );
ms00f80  l1989 ( .o(net_7463), .ck(clk), .d(n9228) );
ms00f80  l1990 ( .o(_net_7701), .ck(clk), .d(n9233) );
ms00f80  l1991 ( .o(net_6705), .ck(clk), .d(n9238) );
ms00f80  l1992 ( .o(net_6483), .ck(clk), .d(n9242) );
ms00f80  l1993 ( .o(net_6527), .ck(clk), .d(n9245) );
ms00f80  l1994 ( .o(net_6701), .ck(clk), .d(n9250) );
ms00f80  l1995 ( .o(net_7103), .ck(clk), .d(n9254) );
ms00f80  l1996 ( .o(_net_6405), .ck(clk), .d(n9258) );
ms00f80  l1997 ( .o(_net_7515), .ck(clk), .d(n9263) );
ms00f80  l1998 ( .o(net_6669), .ck(clk), .d(n9267) );
ms00f80  l1999 ( .o(_net_7530), .ck(clk), .d(n9272) );
ms00f80  l2000 ( .o(_net_6106), .ck(clk), .d(n9277) );
ms00f80  l2001 ( .o(_net_6137), .ck(clk), .d(n9282) );
ms00f80  l2002 ( .o(net_6848), .ck(clk), .d(n9287) );
ms00f80  l2003 ( .o(net_7190), .ck(clk), .d(n9290) );
ms00f80  l2004 ( .o(net_7218), .ck(clk), .d(n9294) );
ms00f80  l2005 ( .o(net_7612), .ck(clk), .d(n9298) );
ms00f80  l2006 ( .o(net_7519), .ck(clk), .d(n9302) );
ms00f80  l2007 ( .o(_net_7516), .ck(clk), .d(n9307) );
ms00f80  l2008 ( .o(_net_7726), .ck(clk), .d(n9312) );
ms00f80  l2009 ( .o(net_7377), .ck(clk), .d(n9316) );
ms00f80  l2010 ( .o(net_219), .ck(clk), .d(n9321) );
ms00f80  l2011 ( .o(net_6749), .ck(clk), .d(n9326) );
ms00f80  l2012 ( .o(_net_5983), .ck(clk), .d(n9330) );
ms00f80  l2013 ( .o(_net_7725), .ck(clk), .d(n9335) );
ms00f80  l2014 ( .o(net_6662), .ck(clk), .d(n9339) );
ms00f80  l2015 ( .o(net_6535), .ck(clk), .d(n9343) );
ms00f80  l2016 ( .o(net_7541), .ck(clk), .d(n9348) );
ms00f80  l2017 ( .o(_net_7504), .ck(clk), .d(n9352) );
ms00f80  l2018 ( .o(net_7164), .ck(clk), .d(n9356) );
ms00f80  l2019 ( .o(net_6464), .ck(clk), .d(n9361) );
ms00f80  l2020 ( .o(net_6265), .ck(clk), .d(n9365) );
ms00f80  l2021 ( .o(net_7099), .ck(clk), .d(n9370) );
ms00f80  l2022 ( .o(net_6640), .ck(clk), .d(n9373) );
ms00f80  l2023 ( .o(net_6817), .ck(clk), .d(n9377) );
ms00f80  l2024 ( .o(net_6921), .ck(clk), .d(n9381) );
ms00f80  l2025 ( .o(net_7072), .ck(clk), .d(n9385) );
ms00f80  l2026 ( .o(net_6601), .ck(clk), .d(n9390) );
ms00f80  l2027 ( .o(net_6936), .ck(clk), .d(n9393) );
ms00f80  l2028 ( .o(net_6278), .ck(clk), .d(n9398) );
ms00f80  l2029 ( .o(x0), .ck(clk), .d(n9402) );
ms00f80  l2030 ( .o(net_6908), .ck(clk), .d(n9405) );
ms00f80  l2031 ( .o(_net_7569), .ck(clk), .d(n9410) );
ms00f80  l2032 ( .o(_net_6085), .ck(clk), .d(n9415) );
ms00f80  l2033 ( .o(_net_7317), .ck(clk), .d(n9420) );
ms00f80  l2034 ( .o(net_6459), .ck(clk), .d(n9425) );
ms00f80  l2035 ( .o(net_145), .ck(clk), .d(n9428) );
ms00f80  l2036 ( .o(net_6775), .ck(clk), .d(n9431) );
ms00f80  l2037 ( .o(_net_7745), .ck(clk), .d(n9436) );
ms00f80  l2038 ( .o(x638), .ck(clk), .d(n9441) );
ms00f80  l2039 ( .o(net_6731), .ck(clk), .d(n9445) );
ms00f80  l2040 ( .o(_net_6280), .ck(clk), .d(n9449) );
ms00f80  l2041 ( .o(_net_6005), .ck(clk), .d(n9454) );
ms00f80  l2042 ( .o(net_7709), .ck(clk), .d(n9459) );
ms00f80  l2043 ( .o(net_6916), .ck(clk), .d(n9462) );
ms00f80  l2044 ( .o(net_6972), .ck(clk), .d(n9467) );
ms00f80  l2045 ( .o(net_359), .ck(clk), .d(n9470) );
ms00f80  l2046 ( .o(net_6842), .ck(clk), .d(n9475) );
ms00f80  l2047 ( .o(net_7464), .ck(clk), .d(n9478) );
ms00f80  l2048 ( .o(net_6611), .ck(clk), .d(n9483) );
ms00f80  l2049 ( .o(_net_7415), .ck(clk), .d(n9487) );
ms00f80  l2050 ( .o(_net_7282), .ck(clk), .d(n9492) );
ms00f80  l2051 ( .o(_net_7597), .ck(clk), .d(n9497) );
ms00f80  l2052 ( .o(net_6359), .ck(clk), .d(n9502) );
ms00f80  l2053 ( .o(_net_7617), .ck(clk), .d(n9507) );
ms00f80  l2054 ( .o(_net_7616), .ck(clk), .d(n9512) );
ms00f80  l2055 ( .o(net_6871), .ck(clk), .d(n9517) );
ms00f80  l2056 ( .o(net_316), .ck(clk), .d(n9520) );
ms00f80  l2057 ( .o(net_7015), .ck(clk), .d(n9525) );
ms00f80  l2058 ( .o(net_6667), .ck(clk), .d(n9528) );
ms00f80  l2059 ( .o(_net_217), .ck(clk), .d(n9533) );
ms00f80  l2060 ( .o(net_6782), .ck(clk), .d(n9537) );
ms00f80  l2061 ( .o(net_7183), .ck(clk), .d(n9541) );
ms00f80  l2062 ( .o(x138), .ck(clk), .d(n9546) );
ms00f80  l2063 ( .o(net_7524), .ck(clk), .d(n9549) );
ms00f80  l2064 ( .o(net_6058), .ck(clk), .d(n9554) );
ms00f80  l2065 ( .o(_net_190), .ck(clk), .d(n9559) );
ms00f80  l2066 ( .o(_net_6021), .ck(clk), .d(n9564) );
ms00f80  l2067 ( .o(_net_7509), .ck(clk), .d(n9569) );
ms00f80  l2068 ( .o(net_297), .ck(clk), .d(n9574) );
ms00f80  l2069 ( .o(net_6840), .ck(clk), .d(n9579) );
ms00f80  l2070 ( .o(_net_7506), .ck(clk), .d(n9583) );
ms00f80  l2071 ( .o(net_6455), .ck(clk), .d(n9588) );
ms00f80  l2072 ( .o(net_6036), .ck(clk), .d(n9592) );
ms00f80  l2073 ( .o(_net_6153), .ck(clk), .d(n9597) );
ms00f80  l2074 ( .o(_net_7324), .ck(clk), .d(n9602) );
ms00f80  l2075 ( .o(net_6818), .ck(clk), .d(n9606) );
ms00f80  l2076 ( .o(net_6307), .ck(clk), .d(n9611) );
ms00f80  l2077 ( .o(_net_6052), .ck(clk), .d(n9616) );
ms00f80  l2078 ( .o(net_6785), .ck(clk), .d(n9620) );
ms00f80  l2079 ( .o(net_7205), .ck(clk), .d(n9624) );
ms00f80  l2080 ( .o(_net_6219), .ck(clk), .d(n9628) );
ms00f80  l2081 ( .o(_net_7436), .ck(clk), .d(n9633) );
ms00f80  l2082 ( .o(_net_7414), .ck(clk), .d(n9638) );
ms00f80  l2083 ( .o(net_6644), .ck(clk), .d(n9642) );
ms00f80  l2084 ( .o(net_7386), .ck(clk), .d(n9647) );
ms00f80  l2085 ( .o(net_7548), .ck(clk), .d(n9651) );
ms00f80  l2086 ( .o(_net_7327), .ck(clk), .d(n9655) );
ms00f80  l2087 ( .o(net_7005), .ck(clk), .d(n9660) );
ms00f80  l2088 ( .o(_net_7656), .ck(clk), .d(n9664) );
ms00f80  l2089 ( .o(net_368), .ck(clk), .d(n9668) );
ms00f80  l2090 ( .o(_net_7588), .ck(clk), .d(n9673) );
ms00f80  l2091 ( .o(_net_225), .ck(clk), .d(n9678) );
ms00f80  l2092 ( .o(_net_7560), .ck(clk), .d(n9683) );
ms00f80  l2093 ( .o(net_317), .ck(clk), .d(n9687) );
ms00f80  l2094 ( .o(net_6703), .ck(clk), .d(n9692) );
ms00f80  l2095 ( .o(net_366), .ck(clk), .d(n9695) );
ms00f80  l2096 ( .o(_net_5964), .ck(clk), .d(n9700) );
ms00f80  l2097 ( .o(net_6634), .ck(clk), .d(n9704) );
ms00f80  l2098 ( .o(_net_6051), .ck(clk), .d(n9709) );
ms00f80  l2099 ( .o(_net_6143), .ck(clk), .d(n9714) );
ms00f80  l2100 ( .o(_net_6174), .ck(clk), .d(n9719) );
ms00f80  l2101 ( .o(net_6358), .ck(clk), .d(n9724) );
ms00f80  l2102 ( .o(net_6472), .ck(clk), .d(n9729) );
ms00f80  l2103 ( .o(_net_192), .ck(clk), .d(n9733) );
ms00f80  l2104 ( .o(_net_7817), .ck(clk), .d(n9737) );
ms00f80  l2105 ( .o(net_170), .ck(clk), .d(n9742) );
ms00f80  l2106 ( .o(net_7214), .ck(clk), .d(n9746) );
ms00f80  l2107 ( .o(net_6657), .ck(clk), .d(n9750) );
ms00f80  l2108 ( .o(net_7522), .ck(clk), .d(n9754) );
ms00f80  l2109 ( .o(net_7669), .ck(clk), .d(n9758) );
ms00f80  l2110 ( .o(_net_7576), .ck(clk), .d(n9763) );
ms00f80  l2111 ( .o(_net_7283), .ck(clk), .d(n9768) );
ms00f80  l2112 ( .o(_net_6002), .ck(clk), .d(n9773) );
ms00f80  l2113 ( .o(_net_5973), .ck(clk), .d(n9778) );
ms00f80  l2114 ( .o(net_7027), .ck(clk), .d(n9783) );
ms00f80  l2115 ( .o(_net_7566), .ck(clk), .d(n9787) );
ms00f80  l2116 ( .o(_net_5989), .ck(clk), .d(n9792) );
ms00f80  l2117 ( .o(net_6807), .ck(clk), .d(n9796) );
ms00f80  l2118 ( .o(_net_7384), .ck(clk), .d(n9801) );
ms00f80  l2119 ( .o(net_384), .ck(clk), .d(n9805) );
ms00f80  l2120 ( .o(net_313), .ck(clk), .d(n9809) );
ms00f80  l2121 ( .o(_net_5859), .ck(clk), .d(n9814) );
ms00f80  l2122 ( .o(_net_7533), .ck(clk), .d(n9819) );
ms00f80  l2123 ( .o(_net_7383), .ck(clk), .d(n9824) );
ms00f80  l2124 ( .o(net_7674), .ck(clk), .d(n9828) );
ms00f80  l2125 ( .o(net_7135), .ck(clk), .d(n9833) );
ms00f80  l2126 ( .o(net_7122), .ck(clk), .d(n9837) );
ms00f80  l2127 ( .o(net_321), .ck(clk), .d(n9840) );
ms00f80  l2128 ( .o(net_305), .ck(clk), .d(n9844) );
ms00f80  l2129 ( .o(_net_7421), .ck(clk), .d(n9849) );
ms00f80  l2130 ( .o(net_7644), .ck(clk), .d(n9853) );
ms00f80  l2131 ( .o(_net_6407), .ck(clk), .d(n9858) );
ms00f80  l2132 ( .o(_net_7097), .ck(clk), .d(n9863) );
ms00f80  l2133 ( .o(net_6943), .ck(clk), .d(n9867) );
ms00f80  l2134 ( .o(net_6929), .ck(clk), .d(n9871) );
ms00f80  l2135 ( .o(net_6533), .ck(clk), .d(n9875) );
ms00f80  l2136 ( .o(_net_6421), .ck(clk), .d(n9880) );
ms00f80  l2137 ( .o(net_7109), .ck(clk), .d(n9885) );
ms00f80  l2138 ( .o(_net_6111), .ck(clk), .d(n9889) );
ms00f80  l2139 ( .o(_net_287), .ck(clk), .d(n9894) );
ms00f80  l2140 ( .o(net_6752), .ck(clk), .d(n9899) );
ms00f80  l2141 ( .o(net_6795), .ck(clk), .d(n9902) );
ms00f80  l2142 ( .o(x361), .ck(clk), .d(n9907) );
ms00f80  l2143 ( .o(net_6446), .ck(clk), .d(n9911) );
ms00f80  l2144 ( .o(net_7221), .ck(clk), .d(n9914) );
ms00f80  l2145 ( .o(_net_7795), .ck(clk), .d(n9918) );
ms00f80  l2146 ( .o(net_6719), .ck(clk), .d(n9923) );
ms00f80  l2147 ( .o(net_374), .ck(clk), .d(n9926) );
ms00f80  l2148 ( .o(net_338), .ck(clk), .d(n9930) );
ms00f80  l2149 ( .o(net_6465), .ck(clk), .d(n9935) );
ms00f80  l2150 ( .o(_net_288), .ck(clk), .d(n9939) );
ms00f80  l2151 ( .o(net_6370), .ck(clk), .d(n9944) );
ms00f80  l2152 ( .o(_net_7348), .ck(clk), .d(n9949) );
ms00f80  l2153 ( .o(net_7740), .ck(clk), .d(n9953) );
ms00f80  l2154 ( .o(net_354), .ck(clk), .d(n9957) );
ms00f80  l2155 ( .o(net_7071), .ck(clk), .d(n9961) );
ms00f80  l2156 ( .o(_net_7402), .ck(clk), .d(n9966) );
ms00f80  l2157 ( .o(_net_6076), .ck(clk), .d(n9971) );
ms00f80  l2158 ( .o(net_6192), .ck(clk), .d(n9976) );
ms00f80  l2159 ( .o(_net_7788), .ck(clk), .d(n9981) );
ms00f80  l2160 ( .o(net_6381), .ck(clk), .d(n9985) );
ms00f80  l2161 ( .o(net_6905), .ck(clk), .d(n9988) );
ms00f80  l2162 ( .o(net_7175), .ck(clk), .d(n9992) );
ms00f80  l2163 ( .o(_net_7717), .ck(clk), .d(n9997) );
ms00f80  l2164 ( .o(net_6507), .ck(clk), .d(n10001) );
ms00f80  l2165 ( .o(net_6198), .ck(clk), .d(n10006) );
ms00f80  l2166 ( .o(net_6529), .ck(clk), .d(n10010) );
ms00f80  l2167 ( .o(_net_7823), .ck(clk), .d(n10014) );
ms00f80  l2168 ( .o(_net_267), .ck(clk), .d(n10019) );
ms00f80  l2169 ( .o(net_6224), .ck(clk), .d(n10023) );
ms00f80  l2170 ( .o(net_6879), .ck(clk), .d(n10028) );
ms00f80  l2171 ( .o(_net_7582), .ck(clk), .d(n10032) );
ms00f80  l2172 ( .o(_net_6017), .ck(clk), .d(n10037) );
ms00f80  l2173 ( .o(_net_6203), .ck(clk), .d(n10042) );
ms00f80  l2174 ( .o(net_6351), .ck(clk), .d(n10047) );
ms00f80  l2175 ( .o(_net_7287), .ck(clk), .d(n10052) );
ms00f80  l2176 ( .o(net_7677), .ck(clk), .d(n10056) );
ms00f80  l2177 ( .o(net_7773), .ck(clk), .d(n10061) );
ms00f80  l2178 ( .o(x620), .ck(clk), .d(n10066) );
ms00f80  l2179 ( .o(net_6884), .ck(clk), .d(n10070) );
ms00f80  l2180 ( .o(_net_7251), .ck(clk), .d(n10074) );
ms00f80  l2181 ( .o(_net_6555), .ck(clk), .d(n10079) );
ms00f80  l2182 ( .o(_net_6131), .ck(clk), .d(n10084) );
ms00f80  l2183 ( .o(_net_6183), .ck(clk), .d(n10089) );
ms00f80  l2184 ( .o(_net_7264), .ck(clk), .d(n10094) );
ms00f80  l2185 ( .o(_net_7479), .ck(clk), .d(n10099) );
ms00f80  l2186 ( .o(net_6645), .ck(clk), .d(n10103) );
ms00f80  l2187 ( .o(net_6648), .ck(clk), .d(n10107) );
ms00f80  l2188 ( .o(net_7112), .ck(clk), .d(n10112) );
ms00f80  l2189 ( .o(net_248), .ck(clk), .d(n10116) );
ms00f80  l2190 ( .o(net_6780), .ck(clk), .d(n10120) );
ms00f80  l2191 ( .o(net_148), .ck(clk), .d(n10124) );
ms00f80  l2192 ( .o(_net_7356), .ck(clk), .d(n10128) );
ms00f80  l2193 ( .o(net_6532), .ck(clk), .d(n10132) );
ms00f80  l2194 ( .o(_net_6176), .ck(clk), .d(n10137) );
ms00f80  l2195 ( .o(_net_7793), .ck(clk), .d(n10141) );
ms00f80  l2196 ( .o(net_7313), .ck(clk), .d(n10145) );
ms00f80  l2197 ( .o(_net_6164), .ck(clk), .d(n10150) );
ms00f80  l2198 ( .o(net_6772), .ck(clk), .d(n10154) );
ms00f80  l2199 ( .o(net_7041), .ck(clk), .d(n10158) );
vcc      t0 ( .o(n7265) );

endmodule
