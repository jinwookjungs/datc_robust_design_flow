VERSION 5.7 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS	2000 ;
END UNITS

MANUFACTURINGGRID	0.0025 ;

SITE core
  SIZE 0.19 BY 1.71 ;
  CLASS CORE ;
END core

LAYER metal1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.19 ;
  WIDTH 0.065 ;
END metal1

LAYER metal2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.19 ;
  WIDTH 0.07 ;
END metal2

LAYER metal3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.19 ;
  WIDTH 0.07 ;
END metal3

LAYER metal4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.285 ;
  WIDTH 0.14 ;
END metal4

LAYER metal5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.285 ;
  WIDTH 0.14 ;
END metal5

LAYER metal6
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.285 ;
  WIDTH 0.14 ;
END metal6

LAYER metal7
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.38 ;
  WIDTH 0.21 ;
END metal7

LAYER metal8
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.38 ;
  WIDTH 0.21 ;
END metal8

LAYER metal9
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.38 ;
  WIDTH 0.21 ;
END metal9

MACRO in01s01
    CLASS CORE ;
    FOREIGN in01s01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.760 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.465 0.150 0.53 1.255 ;
        RECT 0.415 0.150 0.61 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.210 0.340 0.34 0.405 ;
        END
    END a
END in01s01

MACRO in01s02
    CLASS CORE ;
    FOREIGN in01s02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.925 0.150 1.12 1.255 ;
        RECT 0.835 0.150 1.225 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.420 0.340 0.68 0.405 ;
        END
    END a
END in01s02

MACRO in01s03
    CLASS CORE ;
    FOREIGN in01s03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.900 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.160 0.150 1.355 1.255 ;
        RECT 1.040 0.150 1.495 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.525 0.340 0.85 0.405 ;
        END
    END a
END in01s03

MACRO in01s04
    CLASS CORE ;
    FOREIGN in01s04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.900 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.160 0.150 1.355 1.255 ;
        RECT 1.040 0.150 1.495 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.525 0.340 0.85 0.405 ;
        END
    END a
END in01s04

MACRO in01s06
    CLASS CORE ;
    FOREIGN in01s06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.280 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.150 1.65 1.255 ;
        RECT 1.250 0.150 1.77 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.630 0.340 1.02 0.405 ;
        END
    END a
END in01s06

MACRO in01s08
    CLASS CORE ;
    FOREIGN in01s08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.620 0.150 1.945 1.255 ;
        RECT 1.460 0.150 2.11 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.735 0.340 1.19 0.405 ;
        END
    END a
END in01s08

MACRO in01s10
    CLASS CORE ;
    FOREIGN in01s10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.620 0.150 1.945 1.255 ;
        RECT 1.460 0.150 2.11 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.735 0.340 1.19 0.405 ;
        END
    END a
END in01s10

MACRO in01s20
    CLASS CORE ;
    FOREIGN in01s20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.315 0.150 2.77 1.255 ;
        RECT 2.085 0.150 2.995 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.050 0.340 1.7 0.405 ;
        END
    END a
END in01s20

MACRO in01s40
    CLASS CORE ;
    FOREIGN in01s40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.940 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.010 0.150 3.595 1.255 ;
        RECT 2.710 0.150 3.88 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.365 0.340 2.21 0.405 ;
        END
    END a
END in01s40

MACRO in01s80
    CLASS CORE ;
    FOREIGN in01s80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.840 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.170 0.150 4.95 1.255 ;
        RECT 3.750 0.150 5.375 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.890 0.340 3.06 0.405 ;
        END
    END a
END in01s80

MACRO in01m01
    CLASS CORE ;
    FOREIGN in01m01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.760 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.465 0.150 0.53 1.255 ;
        RECT 0.415 0.150 0.61 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.210 0.340 0.34 0.405 ;
        END
    END a
END in01m01

MACRO in01m02
    CLASS CORE ;
    FOREIGN in01m02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.925 0.150 1.12 1.255 ;
        RECT 0.835 0.150 1.225 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.420 0.340 0.68 0.405 ;
        END
    END a
END in01m02

MACRO in01m03
    CLASS CORE ;
    FOREIGN in01m03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.900 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.160 0.150 1.355 1.255 ;
        RECT 1.040 0.150 1.495 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.525 0.340 0.85 0.405 ;
        END
    END a
END in01m03

MACRO in01m04
    CLASS CORE ;
    FOREIGN in01m04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.900 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.160 0.150 1.355 1.255 ;
        RECT 1.040 0.150 1.495 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.525 0.340 0.85 0.405 ;
        END
    END a
END in01m04

MACRO in01m06
    CLASS CORE ;
    FOREIGN in01m06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.280 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.150 1.65 1.255 ;
        RECT 1.250 0.150 1.77 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.630 0.340 1.02 0.405 ;
        END
    END a
END in01m06

MACRO in01m08
    CLASS CORE ;
    FOREIGN in01m08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.620 0.150 1.945 1.255 ;
        RECT 1.460 0.150 2.11 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.735 0.340 1.19 0.405 ;
        END
    END a
END in01m08

MACRO in01m10
    CLASS CORE ;
    FOREIGN in01m10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.620 0.150 1.945 1.255 ;
        RECT 1.460 0.150 2.11 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.735 0.340 1.19 0.405 ;
        END
    END a
END in01m10

MACRO in01m20
    CLASS CORE ;
    FOREIGN in01m20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.315 0.150 2.77 1.255 ;
        RECT 2.085 0.150 2.995 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.050 0.340 1.7 0.405 ;
        END
    END a
END in01m20

MACRO in01m40
    CLASS CORE ;
    FOREIGN in01m40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.940 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.010 0.150 3.595 1.255 ;
        RECT 2.710 0.150 3.88 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.365 0.340 2.21 0.405 ;
        END
    END a
END in01m40

MACRO in01m80
    CLASS CORE ;
    FOREIGN in01m80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.840 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.170 0.150 4.95 1.255 ;
        RECT 3.750 0.150 5.375 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.890 0.340 3.06 0.405 ;
        END
    END a
END in01m80

MACRO in01f01
    CLASS CORE ;
    FOREIGN in01f01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.760 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.465 0.150 0.53 1.255 ;
        RECT 0.415 0.150 0.61 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.210 0.340 0.34 0.405 ;
        END
    END a
END in01f01

MACRO in01f02
    CLASS CORE ;
    FOREIGN in01f02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.925 0.150 1.12 1.255 ;
        RECT 0.835 0.150 1.225 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.420 0.340 0.68 0.405 ;
        END
    END a
END in01f02

MACRO in01f03
    CLASS CORE ;
    FOREIGN in01f03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.900 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.160 0.150 1.355 1.255 ;
        RECT 1.040 0.150 1.495 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.525 0.340 0.85 0.405 ;
        END
    END a
END in01f03

MACRO in01f04
    CLASS CORE ;
    FOREIGN in01f04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.900 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.160 0.150 1.355 1.255 ;
        RECT 1.040 0.150 1.495 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.525 0.340 0.85 0.405 ;
        END
    END a
END in01f04

MACRO in01f06
    CLASS CORE ;
    FOREIGN in01f06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.280 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.150 1.65 1.255 ;
        RECT 1.250 0.150 1.77 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.630 0.340 1.02 0.405 ;
        END
    END a
END in01f06

MACRO in01f08
    CLASS CORE ;
    FOREIGN in01f08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.620 0.150 1.945 1.255 ;
        RECT 1.460 0.150 2.11 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.735 0.340 1.19 0.405 ;
        END
    END a
END in01f08

MACRO in01f10
    CLASS CORE ;
    FOREIGN in01f10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.620 0.150 1.945 1.255 ;
        RECT 1.460 0.150 2.11 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.735 0.340 1.19 0.405 ;
        END
    END a
END in01f10

MACRO in01f20
    CLASS CORE ;
    FOREIGN in01f20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.315 0.150 2.77 1.255 ;
        RECT 2.085 0.150 2.995 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.050 0.340 1.7 0.405 ;
        END
    END a
END in01f20

MACRO in01f40
    CLASS CORE ;
    FOREIGN in01f40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.940 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.010 0.150 3.595 1.255 ;
        RECT 2.710 0.150 3.88 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.365 0.340 2.21 0.405 ;
        END
    END a
END in01f40

MACRO in01f80
    CLASS CORE ;
    FOREIGN in01f80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.840 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.170 0.150 4.95 1.255 ;
        RECT 3.750 0.150 5.375 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.890 0.340 3.06 0.405 ;
        END
    END a
END in01f80

MACRO na02s01
    CLASS CORE ;
    FOREIGN na02s01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.140 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.450 0.110 0.58 1.215 ;
        RECT 0.430 0.725 0.625 1.245 ;
        RECT 0.450 0.110 0.905 0.175 ;
        RECT 0.805 0.110 0.935 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.070 0.535 0.33 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.645 0.540 0.905 0.67 ;
        END
    END b
END na02s01

MACRO na02s02
    CLASS CORE ;
    FOREIGN na02s02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.050 0.110 1.31 1.215 ;
        RECT 1.000 0.725 1.455 1.245 ;
        RECT 1.050 0.110 2.09 0.175 ;
        RECT 1.875 0.110 2.135 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.160 0.535 0.81 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.505 0.540 2.09 0.67 ;
        END
    END b
END na02s02

MACRO na02s03
    CLASS CORE ;
    FOREIGN na02s03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.420 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.350 0.110 1.675 1.215 ;
        RECT 1.285 0.725 1.87 1.245 ;
        RECT 1.350 0.110 2.715 0.175 ;
        RECT 2.410 0.110 2.735 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.205 0.535 1.05 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.935 0.540 2.715 0.67 ;
        END
    END b
END na02s03

MACRO na02s04
    CLASS CORE ;
    FOREIGN na02s04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.500 0.110 1.825 1.215 ;
        RECT 1.425 0.725 2.075 1.245 ;
        RECT 1.500 0.110 2.995 0.175 ;
        RECT 2.675 0.110 3.0 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.225 0.535 1.2 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.150 0.540 2.995 0.67 ;
        END
    END b
END na02s04

MACRO na02s06
    CLASS CORE ;
    FOREIGN na02s06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.800 0.110 2.19 1.215 ;
        RECT 1.710 0.725 2.49 1.245 ;
        RECT 1.800 0.110 3.62 0.175 ;
        RECT 3.210 0.110 3.6 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.270 0.535 1.44 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.580 0.540 3.62 0.67 ;
        END
    END b
END na02s06

MACRO na02s08
    CLASS CORE ;
    FOREIGN na02s08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.940 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.950 0.110 2.405 1.215 ;
        RECT 1.855 0.725 2.7 1.245 ;
        RECT 1.950 0.110 3.9 0.175 ;
        RECT 3.480 0.110 3.935 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.290 0.535 1.525 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.795 0.540 3.9 0.67 ;
        END
    END b
END na02s08

MACRO na02s10
    CLASS CORE ;
    FOREIGN na02s10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.700 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.250 0.110 2.77 1.215 ;
        RECT 2.140 0.725 3.18 1.245 ;
        RECT 2.250 0.110 4.525 0.175 ;
        RECT 4.015 0.110 4.535 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.340 0.535 1.77 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.225 0.540 4.525 0.67 ;
        END
    END b
END na02s10

MACRO na02s20
    CLASS CORE ;
    FOREIGN na02s20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.000 0.110 3.65 1.215 ;
        RECT 2.850 0.725 4.215 1.245 ;
        RECT 3.000 0.110 5.99 0.175 ;
        RECT 5.350 0.110 6.0 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.450 0.535 2.335 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.300 0.540 6.055 0.67 ;
        END
    END b
END na02s20

MACRO na02s40
    CLASS CORE ;
    FOREIGN na02s40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.200 0.110 5.11 1.215 ;
        RECT 3.990 0.725 5.875 1.245 ;
        RECT 4.200 0.110 8.425 0.175 ;
        RECT 7.490 0.110 8.4 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.630 0.535 3.295 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.020 0.540 8.425 0.67 ;
        END
    END b
END na02s40

MACRO na02s80
    CLASS CORE ;
    FOREIGN na02s80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.440 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.700 0.110 6.935 1.215 ;
        RECT 5.415 0.725 7.95 1.245 ;
        RECT 5.700 0.110 11.42 0.175 ;
        RECT 10.165 0.110 11.4 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.855 0.535 4.495 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.170 0.540 11.42 0.67 ;
        END
    END b
END na02s80

MACRO na02m01
    CLASS CORE ;
    FOREIGN na02m01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.140 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.450 0.110 0.58 1.215 ;
        RECT 0.430 0.725 0.625 1.245 ;
        RECT 0.450 0.110 0.905 0.175 ;
        RECT 0.805 0.110 0.935 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.070 0.535 0.33 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.645 0.540 0.905 0.67 ;
        END
    END b
END na02m01

MACRO na02m02
    CLASS CORE ;
    FOREIGN na02m02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.050 0.110 1.31 1.215 ;
        RECT 1.000 0.725 1.455 1.245 ;
        RECT 1.050 0.110 2.09 0.175 ;
        RECT 1.875 0.110 2.135 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.160 0.535 0.81 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.505 0.540 2.09 0.67 ;
        END
    END b
END na02m02

MACRO na02m03
    CLASS CORE ;
    FOREIGN na02m03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.420 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.350 0.110 1.675 1.215 ;
        RECT 1.285 0.725 1.87 1.245 ;
        RECT 1.350 0.110 2.715 0.175 ;
        RECT 2.410 0.110 2.735 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.205 0.535 1.05 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.935 0.540 2.715 0.67 ;
        END
    END b
END na02m03

MACRO na02m04
    CLASS CORE ;
    FOREIGN na02m04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.500 0.110 1.825 1.215 ;
        RECT 1.425 0.725 2.075 1.245 ;
        RECT 1.500 0.110 2.995 0.175 ;
        RECT 2.675 0.110 3.0 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.225 0.535 1.2 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.150 0.540 2.995 0.67 ;
        END
    END b
END na02m04

MACRO na02m06
    CLASS CORE ;
    FOREIGN na02m06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.800 0.110 2.19 1.215 ;
        RECT 1.710 0.725 2.49 1.245 ;
        RECT 1.800 0.110 3.62 0.175 ;
        RECT 3.210 0.110 3.6 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.270 0.535 1.44 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.580 0.540 3.62 0.67 ;
        END
    END b
END na02m06

MACRO na02m08
    CLASS CORE ;
    FOREIGN na02m08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.940 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.950 0.110 2.405 1.215 ;
        RECT 1.855 0.725 2.7 1.245 ;
        RECT 1.950 0.110 3.9 0.175 ;
        RECT 3.480 0.110 3.935 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.290 0.535 1.525 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.795 0.540 3.9 0.67 ;
        END
    END b
END na02m08

MACRO na02m10
    CLASS CORE ;
    FOREIGN na02m10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.700 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.250 0.110 2.77 1.215 ;
        RECT 2.140 0.725 3.18 1.245 ;
        RECT 2.250 0.110 4.525 0.175 ;
        RECT 4.015 0.110 4.535 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.340 0.535 1.77 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.225 0.540 4.525 0.67 ;
        END
    END b
END na02m10

MACRO na02m20
    CLASS CORE ;
    FOREIGN na02m20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.000 0.110 3.65 1.215 ;
        RECT 2.850 0.725 4.215 1.245 ;
        RECT 3.000 0.110 5.99 0.175 ;
        RECT 5.350 0.110 6.0 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.450 0.535 2.335 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.300 0.540 6.055 0.67 ;
        END
    END b
END na02m20

MACRO na02m40
    CLASS CORE ;
    FOREIGN na02m40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.200 0.110 5.11 1.215 ;
        RECT 3.990 0.725 5.875 1.245 ;
        RECT 4.200 0.110 8.425 0.175 ;
        RECT 7.490 0.110 8.4 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.630 0.535 3.295 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.020 0.540 8.425 0.67 ;
        END
    END b
END na02m40

MACRO na02m80
    CLASS CORE ;
    FOREIGN na02m80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.440 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.700 0.110 6.935 1.215 ;
        RECT 5.415 0.725 7.95 1.245 ;
        RECT 5.700 0.110 11.42 0.175 ;
        RECT 10.165 0.110 11.4 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.855 0.535 4.495 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.170 0.540 11.42 0.67 ;
        END
    END b
END na02m80

MACRO na02f01
    CLASS CORE ;
    FOREIGN na02f01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.140 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.450 0.110 0.58 1.215 ;
        RECT 0.430 0.725 0.625 1.245 ;
        RECT 0.450 0.110 0.905 0.175 ;
        RECT 0.805 0.110 0.935 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.070 0.535 0.33 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.645 0.540 0.905 0.67 ;
        END
    END b
END na02f01

MACRO na02f02
    CLASS CORE ;
    FOREIGN na02f02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.050 0.110 1.31 1.215 ;
        RECT 1.000 0.725 1.455 1.245 ;
        RECT 1.050 0.110 2.09 0.175 ;
        RECT 1.875 0.110 2.135 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.160 0.535 0.81 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.505 0.540 2.09 0.67 ;
        END
    END b
END na02f02

MACRO na02f03
    CLASS CORE ;
    FOREIGN na02f03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.420 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.350 0.110 1.675 1.215 ;
        RECT 1.285 0.725 1.87 1.245 ;
        RECT 1.350 0.110 2.715 0.175 ;
        RECT 2.410 0.110 2.735 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.205 0.535 1.05 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.935 0.540 2.715 0.67 ;
        END
    END b
END na02f03

MACRO na02f04
    CLASS CORE ;
    FOREIGN na02f04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.500 0.110 1.825 1.215 ;
        RECT 1.425 0.725 2.075 1.245 ;
        RECT 1.500 0.110 2.995 0.175 ;
        RECT 2.675 0.110 3.0 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.225 0.535 1.2 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.150 0.540 2.995 0.67 ;
        END
    END b
END na02f04

MACRO na02f06
    CLASS CORE ;
    FOREIGN na02f06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.800 0.110 2.19 1.215 ;
        RECT 1.710 0.725 2.49 1.245 ;
        RECT 1.800 0.110 3.62 0.175 ;
        RECT 3.210 0.110 3.6 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.270 0.535 1.44 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.580 0.540 3.62 0.67 ;
        END
    END b
END na02f06

MACRO na02f08
    CLASS CORE ;
    FOREIGN na02f08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.940 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.950 0.110 2.405 1.215 ;
        RECT 1.855 0.725 2.7 1.245 ;
        RECT 1.950 0.110 3.9 0.175 ;
        RECT 3.480 0.110 3.935 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.290 0.535 1.525 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.795 0.540 3.9 0.67 ;
        END
    END b
END na02f08

MACRO na02f10
    CLASS CORE ;
    FOREIGN na02f10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.700 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.250 0.110 2.77 1.215 ;
        RECT 2.140 0.725 3.18 1.245 ;
        RECT 2.250 0.110 4.525 0.175 ;
        RECT 4.015 0.110 4.535 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.340 0.535 1.77 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.225 0.540 4.525 0.67 ;
        END
    END b
END na02f10

MACRO na02f20
    CLASS CORE ;
    FOREIGN na02f20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.000 0.110 3.65 1.215 ;
        RECT 2.850 0.725 4.215 1.245 ;
        RECT 3.000 0.110 5.99 0.175 ;
        RECT 5.350 0.110 6.0 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.450 0.535 2.335 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.300 0.540 6.055 0.67 ;
        END
    END b
END na02f20

MACRO na02f40
    CLASS CORE ;
    FOREIGN na02f40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.200 0.110 5.11 1.215 ;
        RECT 3.990 0.725 5.875 1.245 ;
        RECT 4.200 0.110 8.425 0.175 ;
        RECT 7.490 0.110 8.4 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.630 0.535 3.295 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.020 0.540 8.425 0.67 ;
        END
    END b
END na02f40

MACRO na02f80
    CLASS CORE ;
    FOREIGN na02f80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.440 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.700 0.110 6.935 1.215 ;
        RECT 5.415 0.725 7.95 1.245 ;
        RECT 5.700 0.110 11.42 0.175 ;
        RECT 10.165 0.110 11.4 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.855 0.535 4.495 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.170 0.540 11.42 0.67 ;
        END
    END b
END na02f80

MACRO na03s01
    CLASS CORE ;
    FOREIGN na03s01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.140 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.415 0.805 0.48 1.26 ;
        RECT 0.415 0.805 0.935 0.87 ;
        RECT 0.875 0.090 0.94 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.040 0.630 0.3 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.350 0.090 0.545 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.640 0.090 0.77 0.74 ;
        END
    END c
END na03s01

MACRO na03s02
    CLASS CORE ;
    FOREIGN na03s02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.975 0.805 1.17 1.26 ;
        RECT 0.975 0.805 2.21 0.87 ;
        RECT 2.035 0.090 2.23 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.090 0.630 0.61 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.820 0.090 1.34 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.490 0.090 1.815 0.74 ;
        END
    END c
END na03s02

MACRO na03s03
    CLASS CORE ;
    FOREIGN na03s03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.420 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.250 0.805 1.51 1.26 ;
        RECT 1.250 0.805 2.875 0.87 ;
        RECT 2.620 0.090 2.88 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.115 0.630 0.83 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.055 0.090 1.705 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.915 0.090 2.37 0.74 ;
        END
    END c
END na03s03

MACRO na03s04
    CLASS CORE ;
    FOREIGN na03s04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.805 1.65 1.26 ;
        RECT 1.390 0.805 3.145 0.87 ;
        RECT 2.910 0.090 3.17 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.130 0.630 0.91 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.170 0.090 1.885 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.130 0.090 2.65 0.74 ;
        END
    END c
END na03s04

MACRO na03s06
    CLASS CORE ;
    FOREIGN na03s06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.670 0.805 1.995 1.26 ;
        RECT 1.670 0.805 3.815 0.87 ;
        RECT 3.490 0.090 3.815 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.155 0.630 1.065 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.405 0.090 2.25 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.555 0.090 3.14 0.74 ;
        END
    END c
END na03s06

MACRO na03s08
    CLASS CORE ;
    FOREIGN na03s08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.940 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.805 0.805 2.13 1.26 ;
        RECT 1.805 0.805 4.145 0.87 ;
        RECT 3.785 0.090 4.11 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.170 0.630 1.145 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.520 0.090 2.43 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.770 0.090 3.42 0.74 ;
        END
    END c
END na03s08

MACRO na03s10
    CLASS CORE ;
    FOREIGN na03s10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.700 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.085 0.805 2.475 1.26 ;
        RECT 2.085 0.805 4.75 0.87 ;
        RECT 4.365 0.090 4.755 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.195 0.630 1.365 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.755 0.090 2.795 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.195 0.090 3.975 0.74 ;
        END
    END c
END na03s10

MACRO na03s20
    CLASS CORE ;
    FOREIGN na03s20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.780 0.805 3.3 1.26 ;
        RECT 2.780 0.805 6.355 0.87 ;
        RECT 5.820 0.090 6.34 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.260 0.630 1.755 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.340 0.090 3.77 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.260 0.090 5.235 0.74 ;
        END
    END c
END na03s20

MACRO na03s40
    CLASS CORE ;
    FOREIGN na03s40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.890 0.805 4.605 1.26 ;
        RECT 3.890 0.805 8.895 0.87 ;
        RECT 8.150 0.090 8.865 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.365 0.630 2.51 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.275 0.090 5.225 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.965 0.090 7.395 0.74 ;
        END
    END c
END na03s40

MACRO na03s80
    CLASS CORE ;
    FOREIGN na03s80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.440 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.280 0.805 6.255 1.26 ;
        RECT 5.280 0.805 12.04 0.87 ;
        RECT 11.060 0.090 12.035 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.495 0.630 3.355 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.445 0.090 7.11 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.095 0.090 9.98 0.74 ;
        END
    END c
END na03s80

MACRO na03m01
    CLASS CORE ;
    FOREIGN na03m01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.140 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.415 0.805 0.48 1.26 ;
        RECT 0.415 0.805 0.935 0.87 ;
        RECT 0.875 0.090 0.94 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.040 0.630 0.3 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.350 0.090 0.545 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.640 0.090 0.77 0.74 ;
        END
    END c
END na03m01

MACRO na03m02
    CLASS CORE ;
    FOREIGN na03m02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.975 0.805 1.17 1.26 ;
        RECT 0.975 0.805 2.21 0.87 ;
        RECT 2.035 0.090 2.23 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.090 0.630 0.61 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.820 0.090 1.34 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.490 0.090 1.815 0.74 ;
        END
    END c
END na03m02

MACRO na03m03
    CLASS CORE ;
    FOREIGN na03m03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.420 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.250 0.805 1.51 1.26 ;
        RECT 1.250 0.805 2.875 0.87 ;
        RECT 2.620 0.090 2.88 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.115 0.630 0.83 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.055 0.090 1.705 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.915 0.090 2.37 0.74 ;
        END
    END c
END na03m03

MACRO na03m04
    CLASS CORE ;
    FOREIGN na03m04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.805 1.65 1.26 ;
        RECT 1.390 0.805 3.145 0.87 ;
        RECT 2.910 0.090 3.17 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.130 0.630 0.91 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.170 0.090 1.885 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.130 0.090 2.65 0.74 ;
        END
    END c
END na03m04

MACRO na03m06
    CLASS CORE ;
    FOREIGN na03m06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.670 0.805 1.995 1.26 ;
        RECT 1.670 0.805 3.815 0.87 ;
        RECT 3.490 0.090 3.815 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.155 0.630 1.065 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.405 0.090 2.25 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.555 0.090 3.14 0.74 ;
        END
    END c
END na03m06

MACRO na03m08
    CLASS CORE ;
    FOREIGN na03m08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.940 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.805 0.805 2.13 1.26 ;
        RECT 1.805 0.805 4.145 0.87 ;
        RECT 3.785 0.090 4.11 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.170 0.630 1.145 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.520 0.090 2.43 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.770 0.090 3.42 0.74 ;
        END
    END c
END na03m08

MACRO na03m10
    CLASS CORE ;
    FOREIGN na03m10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.700 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.085 0.805 2.475 1.26 ;
        RECT 2.085 0.805 4.75 0.87 ;
        RECT 4.365 0.090 4.755 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.195 0.630 1.365 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.755 0.090 2.795 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.195 0.090 3.975 0.74 ;
        END
    END c
END na03m10

MACRO na03m20
    CLASS CORE ;
    FOREIGN na03m20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.780 0.805 3.3 1.26 ;
        RECT 2.780 0.805 6.355 0.87 ;
        RECT 5.820 0.090 6.34 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.260 0.630 1.755 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.340 0.090 3.77 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.260 0.090 5.235 0.74 ;
        END
    END c
END na03m20

MACRO na03m40
    CLASS CORE ;
    FOREIGN na03m40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.890 0.805 4.605 1.26 ;
        RECT 3.890 0.805 8.895 0.87 ;
        RECT 8.150 0.090 8.865 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.365 0.630 2.51 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.275 0.090 5.225 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.965 0.090 7.395 0.74 ;
        END
    END c
END na03m40

MACRO na03m80
    CLASS CORE ;
    FOREIGN na03m80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.440 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.280 0.805 6.255 1.26 ;
        RECT 5.280 0.805 12.04 0.87 ;
        RECT 11.060 0.090 12.035 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.495 0.630 3.355 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.445 0.090 7.11 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.095 0.090 9.98 0.74 ;
        END
    END c
END na03m80

MACRO na03f01
    CLASS CORE ;
    FOREIGN na03f01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.140 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.415 0.805 0.48 1.26 ;
        RECT 0.415 0.805 0.935 0.87 ;
        RECT 0.875 0.090 0.94 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.040 0.630 0.3 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.350 0.090 0.545 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.640 0.090 0.77 0.74 ;
        END
    END c
END na03f01

MACRO na03f02
    CLASS CORE ;
    FOREIGN na03f02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.975 0.805 1.17 1.26 ;
        RECT 0.975 0.805 2.21 0.87 ;
        RECT 2.035 0.090 2.23 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.090 0.630 0.61 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.820 0.090 1.34 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.490 0.090 1.815 0.74 ;
        END
    END c
END na03f02

MACRO na03f03
    CLASS CORE ;
    FOREIGN na03f03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.420 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.250 0.805 1.51 1.26 ;
        RECT 1.250 0.805 2.875 0.87 ;
        RECT 2.620 0.090 2.88 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.115 0.630 0.83 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.055 0.090 1.705 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.915 0.090 2.37 0.74 ;
        END
    END c
END na03f03

MACRO na03f04
    CLASS CORE ;
    FOREIGN na03f04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.805 1.65 1.26 ;
        RECT 1.390 0.805 3.145 0.87 ;
        RECT 2.910 0.090 3.17 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.130 0.630 0.91 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.170 0.090 1.885 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.130 0.090 2.65 0.74 ;
        END
    END c
END na03f04

MACRO na03f06
    CLASS CORE ;
    FOREIGN na03f06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.670 0.805 1.995 1.26 ;
        RECT 1.670 0.805 3.815 0.87 ;
        RECT 3.490 0.090 3.815 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.155 0.630 1.065 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.405 0.090 2.25 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.555 0.090 3.14 0.74 ;
        END
    END c
END na03f06

MACRO na03f08
    CLASS CORE ;
    FOREIGN na03f08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.940 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.805 0.805 2.13 1.26 ;
        RECT 1.805 0.805 4.145 0.87 ;
        RECT 3.785 0.090 4.11 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.170 0.630 1.145 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.520 0.090 2.43 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.770 0.090 3.42 0.74 ;
        END
    END c
END na03f08

MACRO na03f10
    CLASS CORE ;
    FOREIGN na03f10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.700 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.085 0.805 2.475 1.26 ;
        RECT 2.085 0.805 4.75 0.87 ;
        RECT 4.365 0.090 4.755 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.195 0.630 1.365 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.755 0.090 2.795 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.195 0.090 3.975 0.74 ;
        END
    END c
END na03f10

MACRO na03f20
    CLASS CORE ;
    FOREIGN na03f20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.780 0.805 3.3 1.26 ;
        RECT 2.780 0.805 6.355 0.87 ;
        RECT 5.820 0.090 6.34 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.260 0.630 1.755 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.340 0.090 3.77 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.260 0.090 5.235 0.74 ;
        END
    END c
END na03f20

MACRO na03f40
    CLASS CORE ;
    FOREIGN na03f40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.890 0.805 4.605 1.26 ;
        RECT 3.890 0.805 8.895 0.87 ;
        RECT 8.150 0.090 8.865 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.365 0.630 2.51 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.275 0.090 5.225 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.965 0.090 7.395 0.74 ;
        END
    END c
END na03f40

MACRO na03f80
    CLASS CORE ;
    FOREIGN na03f80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.440 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.280 0.805 6.255 1.26 ;
        RECT 5.280 0.805 12.04 0.87 ;
        RECT 11.060 0.090 12.035 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.495 0.630 3.355 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.445 0.090 7.11 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.095 0.090 9.98 0.74 ;
        END
    END c
END na03f80

MACRO na04s01
    CLASS CORE ;
    FOREIGN na04s01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.465 0.210 0.53 0.925 ;
        RECT 0.465 0.870 0.79 0.935 ;
        RECT 0.715 0.870 0.78 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.145 0.725 1.34 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.890 0.725 1.085 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.210 0.635 0.405 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.635 0.725 0.83 0.79 ;
        END
    END d
END na04s01

MACRO na04s02
    CLASS CORE ;
    FOREIGN na04s02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.040 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.925 0.210 1.12 0.925 ;
        RECT 0.925 0.870 1.575 0.935 ;
        RECT 1.435 0.870 1.63 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.285 0.725 2.61 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.780 0.725 2.105 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.420 0.635 0.745 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.275 0.725 1.6 0.79 ;
        END
    END d
END na04s02

MACRO na04s03
    CLASS CORE ;
    FOREIGN na04s03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.160 0.210 1.355 0.925 ;
        RECT 1.160 0.870 2.005 0.935 ;
        RECT 1.790 0.870 1.985 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.860 0.725 3.25 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.225 0.725 2.615 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.525 0.635 0.915 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.590 0.725 1.98 0.79 ;
        END
    END d
END na04s03

MACRO na04s04
    CLASS CORE ;
    FOREIGN na04s04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.210 1.65 0.925 ;
        RECT 1.390 0.870 2.43 0.935 ;
        RECT 2.150 0.870 2.41 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.430 0.725 3.95 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.670 0.725 3.19 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.630 0.635 1.15 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.910 0.725 2.43 0.79 ;
        END
    END d
END na04s04

MACRO na04s06
    CLASS CORE ;
    FOREIGN na04s06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.620 0.210 1.945 0.925 ;
        RECT 1.620 0.870 2.79 0.935 ;
        RECT 2.510 0.870 2.835 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.000 0.725 4.585 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.115 0.725 3.7 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.735 0.635 1.32 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.230 0.725 2.815 0.79 ;
        END
    END d
END na04s06

MACRO na04s08
    CLASS CORE ;
    FOREIGN na04s08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.080 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.855 0.210 2.18 0.925 ;
        RECT 1.855 0.870 3.22 0.935 ;
        RECT 2.865 0.870 3.19 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.575 0.725 5.225 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.560 0.725 4.21 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.840 0.635 1.49 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.545 0.725 3.195 0.79 ;
        END
    END d
END na04s08

MACRO na04s10
    CLASS CORE ;
    FOREIGN na04s10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.460 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.970 0.210 2.36 0.925 ;
        RECT 1.970 0.870 3.4 0.935 ;
        RECT 3.045 0.870 3.435 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.860 0.725 5.575 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.785 0.725 4.5 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.895 0.635 1.61 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.705 0.725 3.42 0.79 ;
        END
    END d
END na04s10

MACRO na04s20
    CLASS CORE ;
    FOREIGN na04s20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.740 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.665 0.210 3.185 0.925 ;
        RECT 2.665 0.870 4.615 0.935 ;
        RECT 4.120 0.870 4.64 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.575 0.725 7.55 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.115 0.725 6.09 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.210 0.635 2.185 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.660 0.725 4.635 0.79 ;
        END
    END d
END na04s20

MACRO na04s40
    CLASS CORE ;
    FOREIGN na04s40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.780 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.590 0.210 4.24 0.925 ;
        RECT 3.590 0.870 6.255 0.935 ;
        RECT 5.555 0.870 6.205 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.860 0.725 10.16 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.895 0.725 8.195 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.625 0.635 2.925 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.935 0.725 6.235 0.79 ;
        END
    END d
END na04s40

MACRO na04s80
    CLASS CORE ;
    FOREIGN na04s80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.340 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.980 0.210 5.89 0.925 ;
        RECT 4.980 0.870 8.62 0.935 ;
        RECT 7.705 0.870 8.615 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 12.290 0.725 14.11 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 9.565 0.725 11.385 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.255 0.635 4.075 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.845 0.725 8.665 0.79 ;
        END
    END d
END na04s80

MACRO na04m01
    CLASS CORE ;
    FOREIGN na04m01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.465 0.210 0.53 0.925 ;
        RECT 0.465 0.870 0.79 0.935 ;
        RECT 0.715 0.870 0.78 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.145 0.725 1.34 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.890 0.725 1.085 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.210 0.635 0.405 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.635 0.725 0.83 0.79 ;
        END
    END d
END na04m01

MACRO na04m02
    CLASS CORE ;
    FOREIGN na04m02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.040 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.925 0.210 1.12 0.925 ;
        RECT 0.925 0.870 1.575 0.935 ;
        RECT 1.435 0.870 1.63 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.285 0.725 2.61 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.780 0.725 2.105 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.420 0.635 0.745 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.275 0.725 1.6 0.79 ;
        END
    END d
END na04m02

MACRO na04m03
    CLASS CORE ;
    FOREIGN na04m03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.160 0.210 1.355 0.925 ;
        RECT 1.160 0.870 2.005 0.935 ;
        RECT 1.790 0.870 1.985 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.860 0.725 3.25 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.225 0.725 2.615 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.525 0.635 0.915 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.590 0.725 1.98 0.79 ;
        END
    END d
END na04m03

MACRO na04m04
    CLASS CORE ;
    FOREIGN na04m04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.210 1.65 0.925 ;
        RECT 1.390 0.870 2.43 0.935 ;
        RECT 2.150 0.870 2.41 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.430 0.725 3.95 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.670 0.725 3.19 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.630 0.635 1.15 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.910 0.725 2.43 0.79 ;
        END
    END d
END na04m04

MACRO na04m06
    CLASS CORE ;
    FOREIGN na04m06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.620 0.210 1.945 0.925 ;
        RECT 1.620 0.870 2.79 0.935 ;
        RECT 2.510 0.870 2.835 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.000 0.725 4.585 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.115 0.725 3.7 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.735 0.635 1.32 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.230 0.725 2.815 0.79 ;
        END
    END d
END na04m06

MACRO na04m08
    CLASS CORE ;
    FOREIGN na04m08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.080 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.855 0.210 2.18 0.925 ;
        RECT 1.855 0.870 3.22 0.935 ;
        RECT 2.865 0.870 3.19 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.575 0.725 5.225 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.560 0.725 4.21 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.840 0.635 1.49 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.545 0.725 3.195 0.79 ;
        END
    END d
END na04m08

MACRO na04m10
    CLASS CORE ;
    FOREIGN na04m10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.460 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.970 0.210 2.36 0.925 ;
        RECT 1.970 0.870 3.4 0.935 ;
        RECT 3.045 0.870 3.435 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.860 0.725 5.575 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.785 0.725 4.5 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.895 0.635 1.61 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.705 0.725 3.42 0.79 ;
        END
    END d
END na04m10

MACRO na04m20
    CLASS CORE ;
    FOREIGN na04m20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.740 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.665 0.210 3.185 0.925 ;
        RECT 2.665 0.870 4.615 0.935 ;
        RECT 4.120 0.870 4.64 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.575 0.725 7.55 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.115 0.725 6.09 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.210 0.635 2.185 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.660 0.725 4.635 0.79 ;
        END
    END d
END na04m20

MACRO na04m40
    CLASS CORE ;
    FOREIGN na04m40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.780 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.590 0.210 4.24 0.925 ;
        RECT 3.590 0.870 6.255 0.935 ;
        RECT 5.555 0.870 6.205 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.860 0.725 10.16 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.895 0.725 8.195 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.625 0.635 2.925 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.935 0.725 6.235 0.79 ;
        END
    END d
END na04m40

MACRO na04m80
    CLASS CORE ;
    FOREIGN na04m80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.340 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.980 0.210 5.89 0.925 ;
        RECT 4.980 0.870 8.62 0.935 ;
        RECT 7.705 0.870 8.615 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 12.290 0.725 14.11 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 9.565 0.725 11.385 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.255 0.635 4.075 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.845 0.725 8.665 0.79 ;
        END
    END d
END na04m80

MACRO na04f01
    CLASS CORE ;
    FOREIGN na04f01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.465 0.210 0.53 0.925 ;
        RECT 0.465 0.870 0.79 0.935 ;
        RECT 0.715 0.870 0.78 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.145 0.725 1.34 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.890 0.725 1.085 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.210 0.635 0.405 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.635 0.725 0.83 0.79 ;
        END
    END d
END na04f01

MACRO na04f02
    CLASS CORE ;
    FOREIGN na04f02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.040 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.925 0.210 1.12 0.925 ;
        RECT 0.925 0.870 1.575 0.935 ;
        RECT 1.435 0.870 1.63 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.285 0.725 2.61 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.780 0.725 2.105 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.420 0.635 0.745 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.275 0.725 1.6 0.79 ;
        END
    END d
END na04f02

MACRO na04f03
    CLASS CORE ;
    FOREIGN na04f03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.160 0.210 1.355 0.925 ;
        RECT 1.160 0.870 2.005 0.935 ;
        RECT 1.790 0.870 1.985 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.860 0.725 3.25 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.225 0.725 2.615 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.525 0.635 0.915 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.590 0.725 1.98 0.79 ;
        END
    END d
END na04f03

MACRO na04f04
    CLASS CORE ;
    FOREIGN na04f04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.210 1.65 0.925 ;
        RECT 1.390 0.870 2.43 0.935 ;
        RECT 2.150 0.870 2.41 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.430 0.725 3.95 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.670 0.725 3.19 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.630 0.635 1.15 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.910 0.725 2.43 0.79 ;
        END
    END d
END na04f04

MACRO na04f06
    CLASS CORE ;
    FOREIGN na04f06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.620 0.210 1.945 0.925 ;
        RECT 1.620 0.870 2.79 0.935 ;
        RECT 2.510 0.870 2.835 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.000 0.725 4.585 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.115 0.725 3.7 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.735 0.635 1.32 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.230 0.725 2.815 0.79 ;
        END
    END d
END na04f06

MACRO na04f08
    CLASS CORE ;
    FOREIGN na04f08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.080 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.855 0.210 2.18 0.925 ;
        RECT 1.855 0.870 3.22 0.935 ;
        RECT 2.865 0.870 3.19 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.575 0.725 5.225 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.560 0.725 4.21 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.840 0.635 1.49 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.545 0.725 3.195 0.79 ;
        END
    END d
END na04f08

MACRO na04f10
    CLASS CORE ;
    FOREIGN na04f10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.460 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.970 0.210 2.36 0.925 ;
        RECT 1.970 0.870 3.4 0.935 ;
        RECT 3.045 0.870 3.435 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.860 0.725 5.575 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.785 0.725 4.5 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.895 0.635 1.61 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.705 0.725 3.42 0.79 ;
        END
    END d
END na04f10

MACRO na04f20
    CLASS CORE ;
    FOREIGN na04f20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.740 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.665 0.210 3.185 0.925 ;
        RECT 2.665 0.870 4.615 0.935 ;
        RECT 4.120 0.870 4.64 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.575 0.725 7.55 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.115 0.725 6.09 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.210 0.635 2.185 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.660 0.725 4.635 0.79 ;
        END
    END d
END na04f20

MACRO na04f40
    CLASS CORE ;
    FOREIGN na04f40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.780 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.590 0.210 4.24 0.925 ;
        RECT 3.590 0.870 6.255 0.935 ;
        RECT 5.555 0.870 6.205 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.860 0.725 10.16 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.895 0.725 8.195 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.625 0.635 2.925 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.935 0.725 6.235 0.79 ;
        END
    END d
END na04f40

MACRO na04f80
    CLASS CORE ;
    FOREIGN na04f80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.340 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.980 0.210 5.89 0.925 ;
        RECT 4.980 0.870 8.62 0.935 ;
        RECT 7.705 0.870 8.615 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 12.290 0.725 14.11 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 9.565 0.725 11.385 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.255 0.635 4.075 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.845 0.725 8.665 0.79 ;
        END
    END d
END na04f80

MACRO no02s01
    CLASS CORE ;
    FOREIGN no02s01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.140 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.520 0.150 0.65 0.54 ;
        RECT 0.465 0.150 0.66 0.28 ;
        RECT 0.520 0.505 0.91 0.57 ;
        RECT 0.805 0.505 0.935 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.235 0.340 0.43 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.715 0.340 0.91 0.405 ;
        END
    END b
END no02s01

MACRO no02s02
    CLASS CORE ;
    FOREIGN no02s02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.215 0.150 1.475 0.54 ;
        RECT 1.085 0.150 1.54 0.28 ;
        RECT 1.215 0.505 2.125 0.57 ;
        RECT 1.875 0.505 2.135 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.550 0.340 1.005 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.670 0.340 2.125 0.405 ;
        END
    END b
END no02s02

MACRO no02s03
    CLASS CORE ;
    FOREIGN no02s03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.420 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.565 0.150 1.89 0.54 ;
        RECT 1.395 0.150 1.98 0.28 ;
        RECT 1.565 0.505 2.67 0.57 ;
        RECT 2.410 0.505 2.735 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.710 0.340 1.295 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.150 0.340 2.735 0.405 ;
        END
    END b
END no02s03

MACRO no02s04
    CLASS CORE ;
    FOREIGN no02s04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.740 0.150 2.065 0.54 ;
        RECT 1.550 0.150 2.2 0.28 ;
        RECT 1.740 0.505 2.975 0.57 ;
        RECT 2.675 0.505 3.0 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.790 0.340 1.44 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.390 0.340 3.04 0.405 ;
        END
    END b
END no02s04

MACRO no02s06
    CLASS CORE ;
    FOREIGN no02s06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.085 0.150 2.475 0.54 ;
        RECT 1.860 0.150 2.64 0.28 ;
        RECT 2.085 0.505 3.58 0.57 ;
        RECT 3.210 0.505 3.6 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.945 0.340 1.725 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.865 0.340 3.645 0.405 ;
        END
    END b
END no02s06

MACRO no02s08
    CLASS CORE ;
    FOREIGN no02s08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.940 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.260 0.150 2.715 0.54 ;
        RECT 2.015 0.150 2.86 0.28 ;
        RECT 2.260 0.505 3.885 0.57 ;
        RECT 3.480 0.505 3.935 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.025 0.340 1.87 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.105 0.340 3.95 0.405 ;
        END
    END b
END no02s08

MACRO no02s10
    CLASS CORE ;
    FOREIGN no02s10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.700 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.605 0.150 3.125 0.54 ;
        RECT 2.325 0.150 3.365 0.28 ;
        RECT 2.605 0.505 4.49 0.57 ;
        RECT 4.015 0.505 4.535 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.180 0.340 2.09 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.580 0.340 4.49 0.405 ;
        END
    END b
END no02s10

MACRO no02s20
    CLASS CORE ;
    FOREIGN no02s20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.475 0.150 4.125 0.54 ;
        RECT 3.100 0.150 4.465 0.28 ;
        RECT 3.475 0.505 6.01 0.57 ;
        RECT 5.350 0.505 6.0 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.575 0.340 2.81 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.775 0.340 6.01 0.405 ;
        END
    END b
END no02s20

MACRO no02s40
    CLASS CORE ;
    FOREIGN no02s40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.865 0.150 5.775 0.54 ;
        RECT 4.340 0.150 6.225 0.28 ;
        RECT 4.865 0.505 8.375 0.57 ;
        RECT 7.490 0.505 8.4 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.205 0.340 3.96 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.685 0.340 8.44 0.405 ;
        END
    END b
END no02s40

MACRO no02s80
    CLASS CORE ;
    FOREIGN no02s80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.440 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.605 0.150 7.84 0.54 ;
        RECT 5.890 0.150 8.425 0.28 ;
        RECT 6.605 0.505 11.415 0.57 ;
        RECT 10.165 0.505 11.4 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.995 0.340 5.4 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 9.075 0.340 11.48 0.405 ;
        END
    END b
END no02s80

MACRO no02m01
    CLASS CORE ;
    FOREIGN no02m01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.140 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.520 0.150 0.65 0.54 ;
        RECT 0.465 0.150 0.66 0.28 ;
        RECT 0.520 0.505 0.91 0.57 ;
        RECT 0.805 0.505 0.935 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.235 0.340 0.43 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.715 0.340 0.91 0.405 ;
        END
    END b
END no02m01

MACRO no02m02
    CLASS CORE ;
    FOREIGN no02m02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.215 0.150 1.475 0.54 ;
        RECT 1.085 0.150 1.54 0.28 ;
        RECT 1.215 0.505 2.125 0.57 ;
        RECT 1.875 0.505 2.135 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.550 0.340 1.005 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.670 0.340 2.125 0.405 ;
        END
    END b
END no02m02

MACRO no02m03
    CLASS CORE ;
    FOREIGN no02m03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.420 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.565 0.150 1.89 0.54 ;
        RECT 1.395 0.150 1.98 0.28 ;
        RECT 1.565 0.505 2.67 0.57 ;
        RECT 2.410 0.505 2.735 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.710 0.340 1.295 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.150 0.340 2.735 0.405 ;
        END
    END b
END no02m03

MACRO no02m04
    CLASS CORE ;
    FOREIGN no02m04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.740 0.150 2.065 0.54 ;
        RECT 1.550 0.150 2.2 0.28 ;
        RECT 1.740 0.505 2.975 0.57 ;
        RECT 2.675 0.505 3.0 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.790 0.340 1.44 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.390 0.340 3.04 0.405 ;
        END
    END b
END no02m04

MACRO no02m06
    CLASS CORE ;
    FOREIGN no02m06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.085 0.150 2.475 0.54 ;
        RECT 1.860 0.150 2.64 0.28 ;
        RECT 2.085 0.505 3.58 0.57 ;
        RECT 3.210 0.505 3.6 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.945 0.340 1.725 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.865 0.340 3.645 0.405 ;
        END
    END b
END no02m06

MACRO no02m08
    CLASS CORE ;
    FOREIGN no02m08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.940 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.260 0.150 2.715 0.54 ;
        RECT 2.015 0.150 2.86 0.28 ;
        RECT 2.260 0.505 3.885 0.57 ;
        RECT 3.480 0.505 3.935 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.025 0.340 1.87 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.105 0.340 3.95 0.405 ;
        END
    END b
END no02m08

MACRO no02m10
    CLASS CORE ;
    FOREIGN no02m10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.700 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.605 0.150 3.125 0.54 ;
        RECT 2.325 0.150 3.365 0.28 ;
        RECT 2.605 0.505 4.49 0.57 ;
        RECT 4.015 0.505 4.535 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.180 0.340 2.09 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.580 0.340 4.49 0.405 ;
        END
    END b
END no02m10

MACRO no02m20
    CLASS CORE ;
    FOREIGN no02m20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.475 0.150 4.125 0.54 ;
        RECT 3.100 0.150 4.465 0.28 ;
        RECT 3.475 0.505 6.01 0.57 ;
        RECT 5.350 0.505 6.0 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.575 0.340 2.81 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.775 0.340 6.01 0.405 ;
        END
    END b
END no02m20

MACRO no02m40
    CLASS CORE ;
    FOREIGN no02m40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.865 0.150 5.775 0.54 ;
        RECT 4.340 0.150 6.225 0.28 ;
        RECT 4.865 0.505 8.375 0.57 ;
        RECT 7.490 0.505 8.4 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.205 0.340 3.96 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.685 0.340 8.44 0.405 ;
        END
    END b
END no02m40

MACRO no02m80
    CLASS CORE ;
    FOREIGN no02m80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.440 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.605 0.150 7.84 0.54 ;
        RECT 5.890 0.150 8.425 0.28 ;
        RECT 6.605 0.505 11.415 0.57 ;
        RECT 10.165 0.505 11.4 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.995 0.340 5.4 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 9.075 0.340 11.48 0.405 ;
        END
    END b
END no02m80

MACRO no02f01
    CLASS CORE ;
    FOREIGN no02f01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.140 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.520 0.150 0.65 0.54 ;
        RECT 0.465 0.150 0.66 0.28 ;
        RECT 0.520 0.505 0.91 0.57 ;
        RECT 0.805 0.505 0.935 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.235 0.340 0.43 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.715 0.340 0.91 0.405 ;
        END
    END b
END no02f01

MACRO no02f02
    CLASS CORE ;
    FOREIGN no02f02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.215 0.150 1.475 0.54 ;
        RECT 1.085 0.150 1.54 0.28 ;
        RECT 1.215 0.505 2.125 0.57 ;
        RECT 1.875 0.505 2.135 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.550 0.340 1.005 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.670 0.340 2.125 0.405 ;
        END
    END b
END no02f02

MACRO no02f03
    CLASS CORE ;
    FOREIGN no02f03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.420 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.565 0.150 1.89 0.54 ;
        RECT 1.395 0.150 1.98 0.28 ;
        RECT 1.565 0.505 2.67 0.57 ;
        RECT 2.410 0.505 2.735 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.710 0.340 1.295 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.150 0.340 2.735 0.405 ;
        END
    END b
END no02f03

MACRO no02f04
    CLASS CORE ;
    FOREIGN no02f04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.740 0.150 2.065 0.54 ;
        RECT 1.550 0.150 2.2 0.28 ;
        RECT 1.740 0.505 2.975 0.57 ;
        RECT 2.675 0.505 3.0 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.790 0.340 1.44 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.390 0.340 3.04 0.405 ;
        END
    END b
END no02f04

MACRO no02f06
    CLASS CORE ;
    FOREIGN no02f06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.085 0.150 2.475 0.54 ;
        RECT 1.860 0.150 2.64 0.28 ;
        RECT 2.085 0.505 3.58 0.57 ;
        RECT 3.210 0.505 3.6 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.945 0.340 1.725 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.865 0.340 3.645 0.405 ;
        END
    END b
END no02f06

MACRO no02f08
    CLASS CORE ;
    FOREIGN no02f08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.940 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.260 0.150 2.715 0.54 ;
        RECT 2.015 0.150 2.86 0.28 ;
        RECT 2.260 0.505 3.885 0.57 ;
        RECT 3.480 0.505 3.935 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.025 0.340 1.87 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.105 0.340 3.95 0.405 ;
        END
    END b
END no02f08

MACRO no02f10
    CLASS CORE ;
    FOREIGN no02f10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.700 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.605 0.150 3.125 0.54 ;
        RECT 2.325 0.150 3.365 0.28 ;
        RECT 2.605 0.505 4.49 0.57 ;
        RECT 4.015 0.505 4.535 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.180 0.340 2.09 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.580 0.340 4.49 0.405 ;
        END
    END b
END no02f10

MACRO no02f20
    CLASS CORE ;
    FOREIGN no02f20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.475 0.150 4.125 0.54 ;
        RECT 3.100 0.150 4.465 0.28 ;
        RECT 3.475 0.505 6.01 0.57 ;
        RECT 5.350 0.505 6.0 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.575 0.340 2.81 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.775 0.340 6.01 0.405 ;
        END
    END b
END no02f20

MACRO no02f40
    CLASS CORE ;
    FOREIGN no02f40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.865 0.150 5.775 0.54 ;
        RECT 4.340 0.150 6.225 0.28 ;
        RECT 4.865 0.505 8.375 0.57 ;
        RECT 7.490 0.505 8.4 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.205 0.340 3.96 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.685 0.340 8.44 0.405 ;
        END
    END b
END no02f40

MACRO no02f80
    CLASS CORE ;
    FOREIGN no02f80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.440 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.605 0.150 7.84 0.54 ;
        RECT 5.890 0.150 8.425 0.28 ;
        RECT 6.605 0.505 11.415 0.57 ;
        RECT 10.165 0.505 11.4 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.995 0.340 5.4 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 9.075 0.340 11.48 0.405 ;
        END
    END b
END no02f80

MACRO no03s01
    CLASS CORE ;
    FOREIGN no03s01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.140 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.420 0.130 0.485 0.39 ;
        RECT 0.420 0.340 0.94 0.405 ;
        RECT 0.870 0.130 0.935 1.625 ;
        RECT 0.870 0.545 0.935 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.085 0.365 0.28 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.415 0.430 0.545 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.645 0.430 0.775 0.56 ;
        END
    END c
END no03s01

MACRO no03s02
    CLASS CORE ;
    FOREIGN no03s02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.980 0.130 1.175 0.39 ;
        RECT 0.980 0.340 2.215 0.405 ;
        RECT 2.030 0.130 2.225 1.625 ;
        RECT 2.030 0.545 2.225 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.195 0.365 0.65 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.975 0.430 1.3 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.505 0.430 1.83 0.56 ;
        END
    END c
END no03s02

MACRO no03s03
    CLASS CORE ;
    FOREIGN no03s03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.420 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.260 0.130 1.52 0.39 ;
        RECT 1.260 0.340 2.82 0.405 ;
        RECT 2.610 0.130 2.87 1.625 ;
        RECT 2.610 0.545 2.87 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.250 0.365 0.77 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.250 0.430 1.705 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.935 0.430 2.39 0.56 ;
        END
    END c
END no03s03

MACRO no03s04
    CLASS CORE ;
    FOREIGN no03s04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.400 0.130 1.66 0.39 ;
        RECT 1.400 0.340 3.155 0.405 ;
        RECT 2.900 0.130 3.16 1.625 ;
        RECT 2.900 0.545 3.16 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.280 0.365 0.865 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.430 1.845 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.150 0.430 2.67 0.56 ;
        END
    END c
END no03s04

MACRO no03s06
    CLASS CORE ;
    FOREIGN no03s06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.680 0.130 2.005 0.39 ;
        RECT 1.680 0.340 3.76 0.405 ;
        RECT 3.480 0.130 3.805 1.625 ;
        RECT 3.480 0.545 3.805 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.335 0.365 1.05 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.670 0.430 2.255 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.580 0.430 3.165 0.56 ;
        END
    END c
END no03s06

MACRO no03s08
    CLASS CORE ;
    FOREIGN no03s08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.940 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.820 0.130 2.145 0.39 ;
        RECT 1.820 0.340 4.095 0.405 ;
        RECT 3.770 0.130 4.095 1.625 ;
        RECT 3.770 0.545 4.095 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.365 0.365 1.145 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.805 0.430 2.39 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.795 0.430 3.445 0.56 ;
        END
    END c
END no03s08

MACRO no03s10
    CLASS CORE ;
    FOREIGN no03s10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.700 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.100 0.130 2.49 0.39 ;
        RECT 2.100 0.340 4.765 0.405 ;
        RECT 4.350 0.130 4.74 1.625 ;
        RECT 4.350 0.545 4.74 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.420 0.365 1.33 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.085 0.430 2.8 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.225 0.430 3.94 0.56 ;
        END
    END c
END no03s10

MACRO no03s20
    CLASS CORE ;
    FOREIGN no03s20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.800 0.130 3.32 0.39 ;
        RECT 2.800 0.340 6.31 0.405 ;
        RECT 5.800 0.130 6.32 1.625 ;
        RECT 5.800 0.545 6.32 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.560 0.365 1.795 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.780 0.430 3.69 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.300 0.430 5.275 0.56 ;
        END
    END c
END no03s20

MACRO no03s40
    CLASS CORE ;
    FOREIGN no03s40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.920 0.130 4.635 0.39 ;
        RECT 3.920 0.340 8.86 0.405 ;
        RECT 8.120 0.130 8.835 1.625 ;
        RECT 8.120 0.545 8.9 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.785 0.365 2.475 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.890 0.430 5.19 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.020 0.430 7.385 0.56 ;
        END
    END c
END no03s40

MACRO no03s80
    CLASS CORE ;
    FOREIGN no03s80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.440 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.320 0.130 6.295 0.39 ;
        RECT 5.320 0.340 12.015 0.405 ;
        RECT 11.020 0.130 11.995 1.625 ;
        RECT 11.020 0.545 12.06 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.065 0.365 3.405 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.280 0.430 7.035 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.170 0.430 10.055 0.56 ;
        END
    END c
END no03s80

MACRO no03m01
    CLASS CORE ;
    FOREIGN no03m01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.140 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.420 0.130 0.485 0.39 ;
        RECT 0.420 0.340 0.94 0.405 ;
        RECT 0.870 0.130 0.935 1.625 ;
        RECT 0.870 0.545 0.935 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.085 0.365 0.28 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.415 0.430 0.545 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.645 0.430 0.775 0.56 ;
        END
    END c
END no03m01

MACRO no03m02
    CLASS CORE ;
    FOREIGN no03m02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.980 0.130 1.175 0.39 ;
        RECT 0.980 0.340 2.215 0.405 ;
        RECT 2.030 0.130 2.225 1.625 ;
        RECT 2.030 0.545 2.225 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.195 0.365 0.65 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.975 0.430 1.3 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.505 0.430 1.83 0.56 ;
        END
    END c
END no03m02

MACRO no03m03
    CLASS CORE ;
    FOREIGN no03m03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.420 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.260 0.130 1.52 0.39 ;
        RECT 1.260 0.340 2.82 0.405 ;
        RECT 2.610 0.130 2.87 1.625 ;
        RECT 2.610 0.545 2.87 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.250 0.365 0.77 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.250 0.430 1.705 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.935 0.430 2.39 0.56 ;
        END
    END c
END no03m03

MACRO no03m04
    CLASS CORE ;
    FOREIGN no03m04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.400 0.130 1.66 0.39 ;
        RECT 1.400 0.340 3.155 0.405 ;
        RECT 2.900 0.130 3.16 1.625 ;
        RECT 2.900 0.545 3.16 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.280 0.365 0.865 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.430 1.845 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.150 0.430 2.67 0.56 ;
        END
    END c
END no03m04

MACRO no03m06
    CLASS CORE ;
    FOREIGN no03m06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.680 0.130 2.005 0.39 ;
        RECT 1.680 0.340 3.76 0.405 ;
        RECT 3.480 0.130 3.805 1.625 ;
        RECT 3.480 0.545 3.805 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.335 0.365 1.05 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.670 0.430 2.255 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.580 0.430 3.165 0.56 ;
        END
    END c
END no03m06

MACRO no03m08
    CLASS CORE ;
    FOREIGN no03m08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.940 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.820 0.130 2.145 0.39 ;
        RECT 1.820 0.340 4.095 0.405 ;
        RECT 3.770 0.130 4.095 1.625 ;
        RECT 3.770 0.545 4.095 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.365 0.365 1.145 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.805 0.430 2.39 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.795 0.430 3.445 0.56 ;
        END
    END c
END no03m08

MACRO no03m10
    CLASS CORE ;
    FOREIGN no03m10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.700 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.100 0.130 2.49 0.39 ;
        RECT 2.100 0.340 4.765 0.405 ;
        RECT 4.350 0.130 4.74 1.625 ;
        RECT 4.350 0.545 4.74 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.420 0.365 1.33 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.085 0.430 2.8 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.225 0.430 3.94 0.56 ;
        END
    END c
END no03m10

MACRO no03m20
    CLASS CORE ;
    FOREIGN no03m20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.800 0.130 3.32 0.39 ;
        RECT 2.800 0.340 6.31 0.405 ;
        RECT 5.800 0.130 6.32 1.625 ;
        RECT 5.800 0.545 6.32 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.560 0.365 1.795 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.780 0.430 3.69 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.300 0.430 5.275 0.56 ;
        END
    END c
END no03m20

MACRO no03m40
    CLASS CORE ;
    FOREIGN no03m40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.920 0.130 4.635 0.39 ;
        RECT 3.920 0.340 8.86 0.405 ;
        RECT 8.120 0.130 8.835 1.625 ;
        RECT 8.120 0.545 8.9 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.785 0.365 2.475 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.890 0.430 5.19 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.020 0.430 7.385 0.56 ;
        END
    END c
END no03m40

MACRO no03m80
    CLASS CORE ;
    FOREIGN no03m80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.440 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.320 0.130 6.295 0.39 ;
        RECT 5.320 0.340 12.015 0.405 ;
        RECT 11.020 0.130 11.995 1.625 ;
        RECT 11.020 0.545 12.06 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.065 0.365 3.405 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.280 0.430 7.035 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.170 0.430 10.055 0.56 ;
        END
    END c
END no03m80

MACRO no03f01
    CLASS CORE ;
    FOREIGN no03f01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.140 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.420 0.130 0.485 0.39 ;
        RECT 0.420 0.340 0.94 0.405 ;
        RECT 0.870 0.130 0.935 1.625 ;
        RECT 0.870 0.545 0.935 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.085 0.365 0.28 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.415 0.430 0.545 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.645 0.430 0.775 0.56 ;
        END
    END c
END no03f01

MACRO no03f02
    CLASS CORE ;
    FOREIGN no03f02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.980 0.130 1.175 0.39 ;
        RECT 0.980 0.340 2.215 0.405 ;
        RECT 2.030 0.130 2.225 1.625 ;
        RECT 2.030 0.545 2.225 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.195 0.365 0.65 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.975 0.430 1.3 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.505 0.430 1.83 0.56 ;
        END
    END c
END no03f02

MACRO no03f03
    CLASS CORE ;
    FOREIGN no03f03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.420 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.260 0.130 1.52 0.39 ;
        RECT 1.260 0.340 2.82 0.405 ;
        RECT 2.610 0.130 2.87 1.625 ;
        RECT 2.610 0.545 2.87 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.250 0.365 0.77 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.250 0.430 1.705 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.935 0.430 2.39 0.56 ;
        END
    END c
END no03f03

MACRO no03f04
    CLASS CORE ;
    FOREIGN no03f04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.400 0.130 1.66 0.39 ;
        RECT 1.400 0.340 3.155 0.405 ;
        RECT 2.900 0.130 3.16 1.625 ;
        RECT 2.900 0.545 3.16 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.280 0.365 0.865 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.430 1.845 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.150 0.430 2.67 0.56 ;
        END
    END c
END no03f04

MACRO no03f06
    CLASS CORE ;
    FOREIGN no03f06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.680 0.130 2.005 0.39 ;
        RECT 1.680 0.340 3.76 0.405 ;
        RECT 3.480 0.130 3.805 1.625 ;
        RECT 3.480 0.545 3.805 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.335 0.365 1.05 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.670 0.430 2.255 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.580 0.430 3.165 0.56 ;
        END
    END c
END no03f06

MACRO no03f08
    CLASS CORE ;
    FOREIGN no03f08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.940 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.820 0.130 2.145 0.39 ;
        RECT 1.820 0.340 4.095 0.405 ;
        RECT 3.770 0.130 4.095 1.625 ;
        RECT 3.770 0.545 4.095 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.365 0.365 1.145 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.805 0.430 2.39 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.795 0.430 3.445 0.56 ;
        END
    END c
END no03f08

MACRO no03f10
    CLASS CORE ;
    FOREIGN no03f10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.700 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.100 0.130 2.49 0.39 ;
        RECT 2.100 0.340 4.765 0.405 ;
        RECT 4.350 0.130 4.74 1.625 ;
        RECT 4.350 0.545 4.74 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.420 0.365 1.33 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.085 0.430 2.8 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.225 0.430 3.94 0.56 ;
        END
    END c
END no03f10

MACRO no03f20
    CLASS CORE ;
    FOREIGN no03f20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.800 0.130 3.32 0.39 ;
        RECT 2.800 0.340 6.31 0.405 ;
        RECT 5.800 0.130 6.32 1.625 ;
        RECT 5.800 0.545 6.32 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.560 0.365 1.795 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.780 0.430 3.69 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.300 0.430 5.275 0.56 ;
        END
    END c
END no03f20

MACRO no03f40
    CLASS CORE ;
    FOREIGN no03f40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.920 0.130 4.635 0.39 ;
        RECT 3.920 0.340 8.86 0.405 ;
        RECT 8.120 0.130 8.835 1.625 ;
        RECT 8.120 0.545 8.9 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.785 0.365 2.475 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.890 0.430 5.19 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.020 0.430 7.385 0.56 ;
        END
    END c
END no03f40

MACRO no03f80
    CLASS CORE ;
    FOREIGN no03f80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.440 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.320 0.130 6.295 0.39 ;
        RECT 5.320 0.340 12.015 0.405 ;
        RECT 11.020 0.130 11.995 1.625 ;
        RECT 11.020 0.545 12.06 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.065 0.365 3.405 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.280 0.430 7.035 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.170 0.430 10.055 0.56 ;
        END
    END c
END no03f80

MACRO no04s01
    CLASS CORE ;
    FOREIGN no04s01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.465 0.090 0.53 1.455 ;
        RECT 0.465 0.090 0.79 0.155 ;
        RECT 0.715 0.090 0.78 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.145 0.530 1.34 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.890 0.530 1.085 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.045 0.530 0.305 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.635 0.530 0.83 0.66 ;
        END
    END d
END no04s01

MACRO no04s02
    CLASS CORE ;
    FOREIGN no04s02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.040 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.925 0.090 1.12 1.455 ;
        RECT 0.925 0.090 1.575 0.155 ;
        RECT 1.425 0.090 1.62 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.285 0.530 2.61 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.780 0.530 2.105 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.085 0.530 0.605 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.275 0.530 1.6 0.66 ;
        END
    END d
END no04s02

MACRO no04s03
    CLASS CORE ;
    FOREIGN no04s03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.160 0.090 1.355 1.455 ;
        RECT 1.160 0.090 2.005 0.155 ;
        RECT 1.785 0.090 1.98 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.860 0.530 3.25 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.225 0.530 2.615 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.110 0.530 0.76 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.590 0.530 1.98 0.66 ;
        END
    END d
END no04s03

MACRO no04s04
    CLASS CORE ;
    FOREIGN no04s04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.090 1.65 1.455 ;
        RECT 1.390 0.090 2.43 0.155 ;
        RECT 2.140 0.090 2.4 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.430 0.530 3.95 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.670 0.530 3.19 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.130 0.530 0.91 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.910 0.530 2.43 0.66 ;
        END
    END d
END no04s04

MACRO no04s06
    CLASS CORE ;
    FOREIGN no04s06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.620 0.090 1.945 1.455 ;
        RECT 1.620 0.090 2.79 0.155 ;
        RECT 2.495 0.090 2.82 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.000 0.530 4.585 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.115 0.530 3.7 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.150 0.530 1.06 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.230 0.530 2.815 0.66 ;
        END
    END d
END no04s06

MACRO no04s08
    CLASS CORE ;
    FOREIGN no04s08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.080 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.855 0.090 2.18 1.455 ;
        RECT 1.855 0.090 3.22 0.155 ;
        RECT 2.855 0.090 3.18 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.575 0.530 5.225 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.560 0.530 4.21 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.175 0.530 1.215 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.545 0.530 3.195 0.66 ;
        END
    END d
END no04s08

MACRO no04s10
    CLASS CORE ;
    FOREIGN no04s10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.460 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.970 0.090 2.36 1.455 ;
        RECT 1.970 0.090 3.4 0.155 ;
        RECT 3.030 0.090 3.42 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.860 0.530 5.575 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.785 0.530 4.5 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.185 0.530 1.29 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.705 0.530 3.42 0.66 ;
        END
    END d
END no04s10

MACRO no04s20
    CLASS CORE ;
    FOREIGN no04s20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.740 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.665 0.090 3.185 1.455 ;
        RECT 2.665 0.090 4.615 0.155 ;
        RECT 4.100 0.090 4.62 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.575 0.530 7.55 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.115 0.530 6.09 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.250 0.530 1.68 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.660 0.530 4.635 0.66 ;
        END
    END d
END no04s20

MACRO no04s40
    CLASS CORE ;
    FOREIGN no04s40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.780 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.590 0.090 4.24 1.455 ;
        RECT 3.590 0.090 6.19 0.155 ;
        RECT 5.530 0.090 6.18 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.860 0.530 10.16 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.895 0.530 8.195 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.335 0.530 2.285 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.935 0.530 6.235 0.66 ;
        END
    END d
END no04s40

MACRO no04s80
    CLASS CORE ;
    FOREIGN no04s80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.340 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.980 0.090 5.89 1.455 ;
        RECT 4.980 0.090 8.62 0.155 ;
        RECT 7.670 0.090 8.58 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 12.290 0.530 14.11 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 9.565 0.530 11.385 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.465 0.530 3.195 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.845 0.530 8.665 0.66 ;
        END
    END d
END no04s80

MACRO no04m01
    CLASS CORE ;
    FOREIGN no04m01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.465 0.090 0.53 1.455 ;
        RECT 0.465 0.090 0.79 0.155 ;
        RECT 0.715 0.090 0.78 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.145 0.530 1.34 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.890 0.530 1.085 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.045 0.530 0.305 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.635 0.530 0.83 0.66 ;
        END
    END d
END no04m01

MACRO no04m02
    CLASS CORE ;
    FOREIGN no04m02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.040 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.925 0.090 1.12 1.455 ;
        RECT 0.925 0.090 1.575 0.155 ;
        RECT 1.425 0.090 1.62 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.285 0.530 2.61 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.780 0.530 2.105 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.085 0.530 0.605 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.275 0.530 1.6 0.66 ;
        END
    END d
END no04m02

MACRO no04m03
    CLASS CORE ;
    FOREIGN no04m03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.160 0.090 1.355 1.455 ;
        RECT 1.160 0.090 2.005 0.155 ;
        RECT 1.785 0.090 1.98 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.860 0.530 3.25 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.225 0.530 2.615 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.110 0.530 0.76 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.590 0.530 1.98 0.66 ;
        END
    END d
END no04m03

MACRO no04m04
    CLASS CORE ;
    FOREIGN no04m04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.090 1.65 1.455 ;
        RECT 1.390 0.090 2.43 0.155 ;
        RECT 2.140 0.090 2.4 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.430 0.530 3.95 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.670 0.530 3.19 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.130 0.530 0.91 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.910 0.530 2.43 0.66 ;
        END
    END d
END no04m04

MACRO no04m06
    CLASS CORE ;
    FOREIGN no04m06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.620 0.090 1.945 1.455 ;
        RECT 1.620 0.090 2.79 0.155 ;
        RECT 2.495 0.090 2.82 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.000 0.530 4.585 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.115 0.530 3.7 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.150 0.530 1.06 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.230 0.530 2.815 0.66 ;
        END
    END d
END no04m06

MACRO no04m08
    CLASS CORE ;
    FOREIGN no04m08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.080 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.855 0.090 2.18 1.455 ;
        RECT 1.855 0.090 3.22 0.155 ;
        RECT 2.855 0.090 3.18 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.575 0.530 5.225 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.560 0.530 4.21 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.175 0.530 1.215 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.545 0.530 3.195 0.66 ;
        END
    END d
END no04m08

MACRO no04m10
    CLASS CORE ;
    FOREIGN no04m10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.460 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.970 0.090 2.36 1.455 ;
        RECT 1.970 0.090 3.4 0.155 ;
        RECT 3.030 0.090 3.42 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.860 0.530 5.575 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.785 0.530 4.5 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.185 0.530 1.29 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.705 0.530 3.42 0.66 ;
        END
    END d
END no04m10

MACRO no04m20
    CLASS CORE ;
    FOREIGN no04m20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.740 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.665 0.090 3.185 1.455 ;
        RECT 2.665 0.090 4.615 0.155 ;
        RECT 4.100 0.090 4.62 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.575 0.530 7.55 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.115 0.530 6.09 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.250 0.530 1.68 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.660 0.530 4.635 0.66 ;
        END
    END d
END no04m20

MACRO no04m40
    CLASS CORE ;
    FOREIGN no04m40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.780 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.590 0.090 4.24 1.455 ;
        RECT 3.590 0.090 6.19 0.155 ;
        RECT 5.530 0.090 6.18 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.860 0.530 10.16 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.895 0.530 8.195 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.335 0.530 2.285 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.935 0.530 6.235 0.66 ;
        END
    END d
END no04m40

MACRO no04m80
    CLASS CORE ;
    FOREIGN no04m80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.340 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.980 0.090 5.89 1.455 ;
        RECT 4.980 0.090 8.62 0.155 ;
        RECT 7.670 0.090 8.58 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 12.290 0.530 14.11 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 9.565 0.530 11.385 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.465 0.530 3.195 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.845 0.530 8.665 0.66 ;
        END
    END d
END no04m80

MACRO no04f01
    CLASS CORE ;
    FOREIGN no04f01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.465 0.090 0.53 1.455 ;
        RECT 0.465 0.090 0.79 0.155 ;
        RECT 0.715 0.090 0.78 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.145 0.530 1.34 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.890 0.530 1.085 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.045 0.530 0.305 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.635 0.530 0.83 0.66 ;
        END
    END d
END no04f01

MACRO no04f02
    CLASS CORE ;
    FOREIGN no04f02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.040 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.925 0.090 1.12 1.455 ;
        RECT 0.925 0.090 1.575 0.155 ;
        RECT 1.425 0.090 1.62 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.285 0.530 2.61 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.780 0.530 2.105 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.085 0.530 0.605 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.275 0.530 1.6 0.66 ;
        END
    END d
END no04f02

MACRO no04f03
    CLASS CORE ;
    FOREIGN no04f03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.160 0.090 1.355 1.455 ;
        RECT 1.160 0.090 2.005 0.155 ;
        RECT 1.785 0.090 1.98 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.860 0.530 3.25 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.225 0.530 2.615 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.110 0.530 0.76 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.590 0.530 1.98 0.66 ;
        END
    END d
END no04f03

MACRO no04f04
    CLASS CORE ;
    FOREIGN no04f04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.090 1.65 1.455 ;
        RECT 1.390 0.090 2.43 0.155 ;
        RECT 2.140 0.090 2.4 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.430 0.530 3.95 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.670 0.530 3.19 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.130 0.530 0.91 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.910 0.530 2.43 0.66 ;
        END
    END d
END no04f04

MACRO no04f06
    CLASS CORE ;
    FOREIGN no04f06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.620 0.090 1.945 1.455 ;
        RECT 1.620 0.090 2.79 0.155 ;
        RECT 2.495 0.090 2.82 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.000 0.530 4.585 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.115 0.530 3.7 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.150 0.530 1.06 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.230 0.530 2.815 0.66 ;
        END
    END d
END no04f06

MACRO no04f08
    CLASS CORE ;
    FOREIGN no04f08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.080 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.855 0.090 2.18 1.455 ;
        RECT 1.855 0.090 3.22 0.155 ;
        RECT 2.855 0.090 3.18 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.575 0.530 5.225 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.560 0.530 4.21 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.175 0.530 1.215 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.545 0.530 3.195 0.66 ;
        END
    END d
END no04f08

MACRO no04f10
    CLASS CORE ;
    FOREIGN no04f10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.460 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.970 0.090 2.36 1.455 ;
        RECT 1.970 0.090 3.4 0.155 ;
        RECT 3.030 0.090 3.42 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.860 0.530 5.575 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.785 0.530 4.5 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.185 0.530 1.29 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.705 0.530 3.42 0.66 ;
        END
    END d
END no04f10

MACRO no04f20
    CLASS CORE ;
    FOREIGN no04f20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.740 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.665 0.090 3.185 1.455 ;
        RECT 2.665 0.090 4.615 0.155 ;
        RECT 4.100 0.090 4.62 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.575 0.530 7.55 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.115 0.530 6.09 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.250 0.530 1.68 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.660 0.530 4.635 0.66 ;
        END
    END d
END no04f20

MACRO no04f40
    CLASS CORE ;
    FOREIGN no04f40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.780 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.590 0.090 4.24 1.455 ;
        RECT 3.590 0.090 6.19 0.155 ;
        RECT 5.530 0.090 6.18 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.860 0.530 10.16 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.895 0.530 8.195 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.335 0.530 2.285 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.935 0.530 6.235 0.66 ;
        END
    END d
END no04f40

MACRO no04f80
    CLASS CORE ;
    FOREIGN no04f80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.340 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.980 0.090 5.89 1.455 ;
        RECT 4.980 0.090 8.62 0.155 ;
        RECT 7.670 0.090 8.58 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 12.290 0.530 14.11 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 9.565 0.530 11.385 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.465 0.530 3.195 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.845 0.530 8.665 0.66 ;
        END
    END d
END no04f80

MACRO  bf01s01
    CLASS CORE ;
    FOREIGN bf01s01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.060 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.660 0.150 0.725 1.255 ;
        RECT  0.615 0.150 0.810 0.280 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.320 0.340 0.450 0.405 ;
        END
    END a
END bf01s01

MACRO  bf01s02
    CLASS CORE ;
    FOREIGN bf01s02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.125 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.330 0.150 1.525 1.255 ;
        RECT  1.240 0.150 1.635 0.280 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.640 0.340 0.900 0.405 ;
        END
    END a
END bf01s02

MACRO  bf01s03
    CLASS CORE ;
    FOREIGN bf01s03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.655 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.660 0.150 1.855 1.255 ;
        RECT  1.540 0.150 1.995 0.280 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.795 0.340 1.120 0.405 ;
        END
    END a
END bf01s03

MACRO  bf01s04
    CLASS CORE ;
    FOREIGN bf01s04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.655 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.660 0.150 1.855 1.255 ;
        RECT  1.540 0.150 1.995 0.280 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.795 0.340 1.120 0.405 ;
        END
    END a
END bf01s04

MACRO  bf01s06
    CLASS CORE ;
    FOREIGN bf01s06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.190 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.995 0.150 2.250 1.255 ;
        RECT  1.845 0.150 2.370 0.280 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.955 0.340 1.345 0.405 ;
        END
    END a
END bf01s06

MACRO  bf01s08
    CLASS CORE ;
    FOREIGN bf01s08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.720 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.330 0.150 2.655 1.255 ;
        RECT  2.170 0.150 2.820 0.280 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.115 0.340 1.570 0.405 ;
        END
    END a
END bf01s08

MACRO  bf01s10
    CLASS CORE ;
    FOREIGN bf01s10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.720 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.330 0.150 2.655 1.255 ;
        RECT  2.170 0.150 2.820 0.280 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.115 0.340 1.570 0.405 ;
        END
    END a
END bf01s10

MACRO  bf01s20
    CLASS CORE ;
    FOREIGN bf01s20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.315 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.325 0.150 3.780 1.255 ;
        RECT  3.100 0.150 4.005 0.280 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.595 0.340 2.245 0.405 ;
        END
    END a
END bf01s20

MACRO  bf01s40
    CLASS CORE ;
    FOREIGN bf01s40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.915 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.325 0.150 4.910 1.255 ;
        RECT  4.025 0.150 5.195 0.280 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.075 0.340 2.920 0.405 ;
        END
    END a
END bf01s40

MACRO  bf01s80
    CLASS CORE ;
    FOREIGN bf01s80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.575 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.990 0.150 6.770 1.255 ;
        RECT  5.570 0.150 7.195 0.280 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.880 0.340 4.050 0.405 ;
        END
    END a
END bf01s80

MACRO  bf01m01
    CLASS CORE ;
    FOREIGN bf01m01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.060 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.660 0.150 0.725 1.255 ;
        RECT  0.615 0.150 0.810 0.280 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.320 0.340 0.450 0.405 ;
        END
    END a
END bf01m01

MACRO  bf01m02
    CLASS CORE ;
    FOREIGN bf01m02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.125 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.330 0.150 1.525 1.255 ;
        RECT  1.240 0.150 1.635 0.280 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.640 0.340 0.900 0.405 ;
        END
    END a
END bf01m02

MACRO  bf01m03
    CLASS CORE ;
    FOREIGN bf01m03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.655 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.660 0.150 1.855 1.255 ;
        RECT  1.540 0.150 1.995 0.280 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.795 0.340 1.120 0.405 ;
        END
    END a
END bf01m03

MACRO  bf01m04
    CLASS CORE ;
    FOREIGN bf01m04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.655 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.660 0.150 1.855 1.255 ;
        RECT  1.540 0.150 1.995 0.280 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.795 0.340 1.120 0.405 ;
        END
    END a
END bf01m04

MACRO  bf01m06
    CLASS CORE ;
    FOREIGN bf01m06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.190 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.995 0.150 2.250 1.255 ;
        RECT  1.845 0.150 2.370 0.280 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.955 0.340 1.345 0.405 ;
        END
    END a
END bf01m06

MACRO  bf01m08
    CLASS CORE ;
    FOREIGN bf01m08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.720 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.330 0.150 2.655 1.255 ;
        RECT  2.170 0.150 2.820 0.280 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.115 0.340 1.570 0.405 ;
        END
    END a
END bf01m08

MACRO  bf01m10
    CLASS CORE ;
    FOREIGN bf01m10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.720 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.330 0.150 2.655 1.255 ;
        RECT  2.170 0.150 2.820 0.280 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.115 0.340 1.570 0.405 ;
        END
    END a
END bf01m10

MACRO  bf01m20
    CLASS CORE ;
    FOREIGN bf01m20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.315 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.325 0.150 3.780 1.255 ;
        RECT  3.100 0.150 4.005 0.280 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.595 0.340 2.245 0.405 ;
        END
    END a
END bf01m20

MACRO  bf01m40
    CLASS CORE ;
    FOREIGN bf01m40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.915 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.325 0.150 4.910 1.255 ;
        RECT  4.025 0.150 5.195 0.280 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.075 0.340 2.920 0.405 ;
        END
    END a
END bf01m40

MACRO  bf01m80
    CLASS CORE ;
    FOREIGN bf01m80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.575 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.990 0.150 6.770 1.255 ;
        RECT  5.570 0.150 7.195 0.280 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.880 0.340 4.050 0.405 ;
        END
    END a
END bf01m80

MACRO  bf01f01
    CLASS CORE ;
    FOREIGN bf01f01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.060 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.660 0.150 0.725 1.255 ;
        RECT  0.615 0.150 0.810 0.280 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.320 0.340 0.450 0.405 ;
        END
    END a
END bf01f01

MACRO  bf01f02
    CLASS CORE ;
    FOREIGN bf01f02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.125 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.330 0.150 1.525 1.255 ;
        RECT  1.240 0.150 1.635 0.280 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.640 0.340 0.900 0.405 ;
        END
    END a
END bf01f02

MACRO  bf01f03
    CLASS CORE ;
    FOREIGN bf01f03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.655 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.660 0.150 1.855 1.255 ;
        RECT  1.540 0.150 1.995 0.280 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.795 0.340 1.120 0.405 ;
        END
    END a
END bf01f03

MACRO  bf01f04
    CLASS CORE ;
    FOREIGN bf01f04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.655 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.660 0.150 1.855 1.255 ;
        RECT  1.540 0.150 1.995 0.280 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.795 0.340 1.120 0.405 ;
        END
    END a
END bf01f04

MACRO  bf01f06
    CLASS CORE ;
    FOREIGN bf01f06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.190 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.995 0.150 2.250 1.255 ;
        RECT  1.845 0.150 2.370 0.280 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.955 0.340 1.345 0.405 ;
        END
    END a
END bf01f06

MACRO  bf01f08
    CLASS CORE ;
    FOREIGN bf01f08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.720 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.330 0.150 2.655 1.255 ;
        RECT  2.170 0.150 2.820 0.280 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.115 0.340 1.570 0.405 ;
        END
    END a
END bf01f08

MACRO  bf01f10
    CLASS CORE ;
    FOREIGN bf01f10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.720 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.330 0.150 2.655 1.255 ;
        RECT  2.170 0.150 2.820 0.280 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.115 0.340 1.570 0.405 ;
        END
    END a
END bf01f10

MACRO  bf01f20
    CLASS CORE ;
    FOREIGN bf01f20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.315 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.325 0.150 3.780 1.255 ;
        RECT  3.100 0.150 4.005 0.280 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.595 0.340 2.245 0.405 ;
        END
    END a
END bf01f20

MACRO  bf01f40
    CLASS CORE ;
    FOREIGN bf01f40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.915 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.325 0.150 4.910 1.255 ;
        RECT  4.025 0.150 5.195 0.280 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.075 0.340 2.920 0.405 ;
        END
    END a
END bf01f40

MACRO  bf01f80
    CLASS CORE ;
    FOREIGN bf01f80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.575 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.990 0.150 6.770 1.255 ;
        RECT  5.570 0.150 7.195 0.280 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.880 0.340 4.050 0.405 ;
        END
    END a
END bf01f80

MACRO ao12s01
    CLASS CORE ;
    FOREIGN ao12s01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.010 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.520 0.100 0.645 0.685 ;
        RECT  0.550 0.635 0.675 0.765 ;
        RECT  0.505 0.750 0.895 0.815 ;
        RECT  0.725 0.750 0.855 1.530 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.130 0.585 0.325 0.650 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.345 0.505 0.475 0.570 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.675 0.585 0.870 0.650 ;
        END
    END c
END ao12s01

MACRO ao12s02
    CLASS CORE ;
    FOREIGN ao12s02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.530 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.315 0.100 1.580 0.685 ;
        RECT  1.390 0.635 1.650 0.765 ;
        RECT  1.280 0.750 2.190 0.815 ;
        RECT  1.830 0.750 2.085 1.530 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.330 0.585 0.845 0.650 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.855 0.505 1.250 0.570 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.690 0.585 2.210 0.650 ;
        END
    END c
END ao12s02

MACRO ao12s03
    CLASS CORE ;
    FOREIGN ao12s03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.035 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.580 0.100 1.905 0.685 ;
        RECT  1.660 0.635 1.985 0.765 ;
        RECT  1.530 0.750 2.635 0.815 ;
        RECT  2.190 0.750 2.515 1.530 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.400 0.585 0.985 0.650 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.030 0.505 1.485 0.570 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.035 0.585 2.620 0.650 ;
        END
    END c
END ao12s03

MACRO ao12s04
    CLASS CORE ;
    FOREIGN ao12s04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.545 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.845 0.100 2.230 0.685 ;
        RECT  1.940 0.635 2.330 0.765 ;
        RECT  1.790 0.750 3.090 0.815 ;
        RECT  2.550 0.750 2.945 1.530 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.465 0.585 1.180 0.650 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.195 0.505 1.780 0.570 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.370 0.585 3.085 0.650 ;
        END
    END c
END ao12s04

MACRO ao12s06
    CLASS CORE ;
    FOREIGN ao12s06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.305 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.245 0.100 2.700 0.685 ;
        RECT  2.355 0.635 2.810 0.765 ;
        RECT  2.170 0.750 3.735 0.815 ;
        RECT  3.105 0.750 3.560 1.530 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.570 0.585 1.415 0.650 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.465 0.505 2.115 0.570 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.880 0.585 3.725 0.650 ;
        END
    END c
END ao12s06

MACRO ao12s08
    CLASS CORE ;
    FOREIGN ao12s08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.065 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.645 0.100 3.165 0.685 ;
        RECT  2.780 0.635 3.300 0.765 ;
        RECT  2.560 0.750 4.380 0.815 ;
        RECT  3.660 0.750 4.175 1.530 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.675 0.585 1.650 0.650 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.715 0.505 2.500 0.570 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.395 0.585 4.370 0.650 ;
        END
    END c
END ao12s08

MACRO ao12s10
    CLASS CORE ;
    FOREIGN ao12s10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.570 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.905 0.100 3.490 0.685 ;
        RECT  3.050 0.635 3.635 0.765 ;
        RECT  2.815 0.750 4.830 0.815 ;
        RECT  4.020 0.750 4.605 1.530 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.735 0.585 1.840 0.650 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.880 0.505 2.795 0.570 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.730 0.585 4.835 0.650 ;
        END
    END c
END ao12s10

MACRO ao12s20
    CLASS CORE ;
    FOREIGN ao12s20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.970 0.100 4.750 0.685 ;
        RECT  4.160 0.635 4.945 0.765 ;
        RECT  3.845 0.750 6.570 0.815 ;
        RECT  5.485 0.750 6.270 1.530 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.005 0.585 2.500 0.650 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.585 0.505 3.755 0.570 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.085 0.585 6.580 0.650 ;
        END
    END c
END ao12s20

MACRO ao12s40
    CLASS CORE ;
    FOREIGN ao12s40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.385 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.430 0.100 6.470 0.685 ;
        RECT  5.695 0.635 6.740 0.765 ;
        RECT  5.240 0.750 9.015 0.815 ;
        RECT  7.505 0.750 8.545 1.530 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.375 0.585 3.455 0.650 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.525 0.505 5.150 0.570 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.945 0.585 9.025 0.650 ;
        END
    END c
END ao12s40

MACRO ao12s80
    CLASS CORE ;
    FOREIGN ao12s80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.440 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.535 0.100 9.030 0.685 ;
        RECT  7.915 0.635 9.410 0.765 ;
        RECT  7.285 0.750 12.550 0.815 ;
        RECT  10.425 0.750 11.920 1.530 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.915 0.585 4.775 0.650 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.900 0.505 7.175 0.570 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.670 0.585 12.525 0.650 ;
        END
    END c
END ao12s80

MACRO ao12m01
    CLASS CORE ;
    FOREIGN ao12m01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.010 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.520 0.100 0.645 0.685 ;
        RECT  0.550 0.635 0.675 0.765 ;
        RECT  0.505 0.750 0.895 0.815 ;
        RECT  0.725 0.750 0.855 1.530 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.130 0.585 0.325 0.650 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.345 0.505 0.475 0.570 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.675 0.585 0.870 0.650 ;
        END
    END c
END ao12m01

MACRO ao12m02
    CLASS CORE ;
    FOREIGN ao12m02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.530 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.315 0.100 1.580 0.685 ;
        RECT  1.390 0.635 1.650 0.765 ;
        RECT  1.280 0.750 2.190 0.815 ;
        RECT  1.830 0.750 2.085 1.530 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.330 0.585 0.845 0.650 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.855 0.505 1.250 0.570 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.690 0.585 2.210 0.650 ;
        END
    END c
END ao12m02

MACRO ao12m03
    CLASS CORE ;
    FOREIGN ao12m03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.035 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.580 0.100 1.905 0.685 ;
        RECT  1.660 0.635 1.985 0.765 ;
        RECT  1.530 0.750 2.635 0.815 ;
        RECT  2.190 0.750 2.515 1.530 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.400 0.585 0.985 0.650 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.030 0.505 1.485 0.570 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.035 0.585 2.620 0.650 ;
        END
    END c
END ao12m03

MACRO ao12m04
    CLASS CORE ;
    FOREIGN ao12m04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.545 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.845 0.100 2.230 0.685 ;
        RECT  1.940 0.635 2.330 0.765 ;
        RECT  1.790 0.750 3.090 0.815 ;
        RECT  2.550 0.750 2.945 1.530 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.465 0.585 1.180 0.650 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.195 0.505 1.780 0.570 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.370 0.585 3.085 0.650 ;
        END
    END c
END ao12m04

MACRO ao12m06
    CLASS CORE ;
    FOREIGN ao12m06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.305 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.245 0.100 2.700 0.685 ;
        RECT  2.355 0.635 2.810 0.765 ;
        RECT  2.170 0.750 3.735 0.815 ;
        RECT  3.105 0.750 3.560 1.530 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.570 0.585 1.415 0.650 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.465 0.505 2.115 0.570 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.880 0.585 3.725 0.650 ;
        END
    END c
END ao12m06

MACRO ao12m08
    CLASS CORE ;
    FOREIGN ao12m08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.065 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.645 0.100 3.165 0.685 ;
        RECT  2.780 0.635 3.300 0.765 ;
        RECT  2.560 0.750 4.380 0.815 ;
        RECT  3.660 0.750 4.175 1.530 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.675 0.585 1.650 0.650 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.715 0.505 2.500 0.570 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.395 0.585 4.370 0.650 ;
        END
    END c
END ao12m08

MACRO ao12m10
    CLASS CORE ;
    FOREIGN ao12m10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.570 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.905 0.100 3.490 0.685 ;
        RECT  3.050 0.635 3.635 0.765 ;
        RECT  2.815 0.750 4.830 0.815 ;
        RECT  4.020 0.750 4.605 1.530 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.735 0.585 1.840 0.650 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.880 0.505 2.795 0.570 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.730 0.585 4.835 0.650 ;
        END
    END c
END ao12m10

MACRO ao12m20
    CLASS CORE ;
    FOREIGN ao12m20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.970 0.100 4.750 0.685 ;
        RECT  4.160 0.635 4.945 0.765 ;
        RECT  3.845 0.750 6.570 0.815 ;
        RECT  5.485 0.750 6.270 1.530 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.005 0.585 2.500 0.650 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.585 0.505 3.755 0.570 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.085 0.585 6.580 0.650 ;
        END
    END c
END ao12m20

MACRO ao12m40
    CLASS CORE ;
    FOREIGN ao12m40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.385 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.430 0.100 6.470 0.685 ;
        RECT  5.695 0.635 6.740 0.765 ;
        RECT  5.240 0.750 9.015 0.815 ;
        RECT  7.505 0.750 8.545 1.530 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.375 0.585 3.455 0.650 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.525 0.505 5.150 0.570 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.945 0.585 9.025 0.650 ;
        END
    END c
END ao12m40

MACRO ao12m80
    CLASS CORE ;
    FOREIGN ao12m80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.440 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.535 0.100 9.030 0.685 ;
        RECT  7.915 0.635 9.410 0.765 ;
        RECT  7.285 0.750 12.550 0.815 ;
        RECT  10.425 0.750 11.920 1.530 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.915 0.585 4.775 0.650 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.900 0.505 7.175 0.570 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.670 0.585 12.525 0.650 ;
        END
    END c
END ao12m80

MACRO ao12f01
    CLASS CORE ;
    FOREIGN ao12f01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.010 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.520 0.100 0.645 0.685 ;
        RECT  0.550 0.635 0.675 0.765 ;
        RECT  0.505 0.750 0.895 0.815 ;
        RECT  0.725 0.750 0.855 1.530 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.130 0.585 0.325 0.650 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.345 0.505 0.475 0.570 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.675 0.585 0.870 0.650 ;
        END
    END c
END ao12f01

MACRO ao12f02
    CLASS CORE ;
    FOREIGN ao12f02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.530 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.315 0.100 1.580 0.685 ;
        RECT  1.390 0.635 1.650 0.765 ;
        RECT  1.280 0.750 2.190 0.815 ;
        RECT  1.830 0.750 2.085 1.530 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.330 0.585 0.845 0.650 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.855 0.505 1.250 0.570 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.690 0.585 2.210 0.650 ;
        END
    END c
END ao12f02

MACRO ao12f03
    CLASS CORE ;
    FOREIGN ao12f03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.035 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.580 0.100 1.905 0.685 ;
        RECT  1.660 0.635 1.985 0.765 ;
        RECT  1.530 0.750 2.635 0.815 ;
        RECT  2.190 0.750 2.515 1.530 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.400 0.585 0.985 0.650 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.030 0.505 1.485 0.570 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.035 0.585 2.620 0.650 ;
        END
    END c
END ao12f03

MACRO ao12f04
    CLASS CORE ;
    FOREIGN ao12f04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.545 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.845 0.100 2.230 0.685 ;
        RECT  1.940 0.635 2.330 0.765 ;
        RECT  1.790 0.750 3.090 0.815 ;
        RECT  2.550 0.750 2.945 1.530 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.465 0.585 1.180 0.650 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.195 0.505 1.780 0.570 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.370 0.585 3.085 0.650 ;
        END
    END c
END ao12f04

MACRO ao12f06
    CLASS CORE ;
    FOREIGN ao12f06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.305 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.245 0.100 2.700 0.685 ;
        RECT  2.355 0.635 2.810 0.765 ;
        RECT  2.170 0.750 3.735 0.815 ;
        RECT  3.105 0.750 3.560 1.530 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.570 0.585 1.415 0.650 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.465 0.505 2.115 0.570 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.880 0.585 3.725 0.650 ;
        END
    END c
END ao12f06

MACRO ao12f08
    CLASS CORE ;
    FOREIGN ao12f08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.065 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.645 0.100 3.165 0.685 ;
        RECT  2.780 0.635 3.300 0.765 ;
        RECT  2.560 0.750 4.380 0.815 ;
        RECT  3.660 0.750 4.175 1.530 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.675 0.585 1.650 0.650 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.715 0.505 2.500 0.570 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.395 0.585 4.370 0.650 ;
        END
    END c
END ao12f08

MACRO ao12f10
    CLASS CORE ;
    FOREIGN ao12f10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.570 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.905 0.100 3.490 0.685 ;
        RECT  3.050 0.635 3.635 0.765 ;
        RECT  2.815 0.750 4.830 0.815 ;
        RECT  4.020 0.750 4.605 1.530 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.735 0.585 1.840 0.650 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.880 0.505 2.795 0.570 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.730 0.585 4.835 0.650 ;
        END
    END c
END ao12f10

MACRO ao12f20
    CLASS CORE ;
    FOREIGN ao12f20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.970 0.100 4.750 0.685 ;
        RECT  4.160 0.635 4.945 0.765 ;
        RECT  3.845 0.750 6.570 0.815 ;
        RECT  5.485 0.750 6.270 1.530 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.005 0.585 2.500 0.650 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.585 0.505 3.755 0.570 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.085 0.585 6.580 0.650 ;
        END
    END c
END ao12f20

MACRO ao12f40
    CLASS CORE ;
    FOREIGN ao12f40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.385 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.430 0.100 6.470 0.685 ;
        RECT  5.695 0.635 6.740 0.765 ;
        RECT  5.240 0.750 9.015 0.815 ;
        RECT  7.505 0.750 8.545 1.530 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.375 0.585 3.455 0.650 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.525 0.505 5.150 0.570 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.945 0.585 9.025 0.650 ;
        END
    END c
END ao12f40

MACRO ao12f80
    CLASS CORE ;
    FOREIGN ao12f80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.440 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.535 0.100 9.030 0.685 ;
        RECT  7.915 0.635 9.410 0.765 ;
        RECT  7.285 0.750 12.550 0.815 ;
        RECT  10.425 0.750 11.920 1.530 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.915 0.585 4.775 0.650 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.900 0.505 7.175 0.570 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.670 0.585 12.525 0.650 ;
        END
    END c
END ao12f80

MACRO ao22s01
    CLASS CORE ;
    FOREIGN ao22s01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.010 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.295 0.090 0.360 1.455 ;
        RECT  0.250 0.090 0.575 0.155 ;
        RECT  0.460 0.090 0.525 0.480 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.725 0.530 0.920 0.660 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.555 0.530 0.750 0.660 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  -0.015 0.530 0.245 0.660 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.385 0.530 0.580 0.660 ;
        END
    END d
END ao22s01

MACRO ao22s02
    CLASS CORE ;
    FOREIGN ao22s02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.785 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.805 0.090 1.060 1.455 ;
        RECT  0.695 0.090 1.605 0.155 ;
        RECT  1.260 0.090 1.520 0.480 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.015 0.530 2.470 0.660 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.550 0.530 2.005 0.660 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  -0.040 0.530 0.670 0.660 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.085 0.530 1.540 0.660 ;
        END
    END d
END ao22s02

MACRO ao22s03
    CLASS CORE ;
    FOREIGN ao22s03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.545 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.020 0.090 1.345 1.455 ;
        RECT  0.885 0.090 2.050 0.155 ;
        RECT  1.605 0.090 1.930 0.480 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.565 0.530 3.150 0.660 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.975 0.530 2.560 0.660 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  -0.050 0.530 0.855 0.660 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.385 0.530 1.970 0.660 ;
        END
    END d
END ao22s03

MACRO ao22s04
    CLASS CORE ;
    FOREIGN ao22s04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.050 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.180 0.090 1.505 1.455 ;
        RECT  1.005 0.090 2.370 0.155 ;
        RECT  1.845 0.090 2.170 0.480 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.940 0.530 3.590 0.660 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.260 0.530 2.915 0.660 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  -0.060 0.530 0.980 0.660 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.585 0.530 2.235 0.660 ;
        END
    END d
END ao22s04

MACRO ao22s06
    CLASS CORE ;
    FOREIGN ao22s06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.810 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.400 0.090 1.785 1.455 ;
        RECT  1.190 0.090 2.815 0.155 ;
        RECT  2.195 0.090 2.585 0.480 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.485 0.530 4.265 0.660 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.690 0.530 3.465 0.660 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  -0.070 0.530 1.160 0.660 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.880 0.530 2.665 0.660 ;
        END
    END d
END ao22s06

MACRO ao22s08
    CLASS CORE ;
    FOREIGN ao22s08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.570 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.620 0.090 2.075 1.455 ;
        RECT  1.395 0.090 3.215 0.155 ;
        RECT  2.535 0.090 2.990 0.480 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.040 0.530 4.950 0.660 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.110 0.530 4.015 0.660 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  -0.065 0.530 1.295 0.660 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.180 0.530 3.090 0.660 ;
        END
    END d
END ao22s08

MACRO ao22s10
    CLASS CORE ;
    FOREIGN ao22s10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.075 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.765 0.090 2.285 1.455 ;
        RECT  1.515 0.090 3.530 0.155 ;
        RECT  2.765 0.090 3.280 0.480 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.405 0.530 5.380 0.660 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.395 0.530 4.370 0.660 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  -0.075 0.530 1.415 0.660 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.380 0.530 3.355 0.660 ;
        END
    END d
END ao22s10

MACRO ao22s20
    CLASS CORE ;
    FOREIGN ao22s20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.610 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.505 0.090 3.220 1.455 ;
        RECT  2.150 0.090 5.005 0.155 ;
        RECT  3.920 0.090 4.635 0.480 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.240 0.530 7.670 0.660 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.805 0.530 6.230 0.660 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  -0.110 0.530 2.030 0.660 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.365 0.530 4.795 0.660 ;
        END
    END d
END ao22s20

MACRO ao22s40
    CLASS CORE ;
    FOREIGN ao22s40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.650 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.385 0.090 4.360 1.455 ;
        RECT  2.900 0.090 6.800 0.155 ;
        RECT  5.300 0.090 6.275 0.480 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.450 0.530 10.335 0.660 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.505 0.530 8.390 0.660 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  -0.155 0.530 2.765 0.660 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.560 0.530 6.445 0.660 ;
        END
    END d
END ao22s40

MACRO ao22s80
    CLASS CORE ;
    FOREIGN ao22s80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.210 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.710 0.090 6.075 1.455 ;
        RECT  4.040 0.090 9.435 0.155 ;
        RECT  7.375 0.090 8.740 0.480 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.750 0.530 14.415 0.660 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.045 0.530 11.710 0.660 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  -0.205 0.530 3.815 0.660 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.340 0.530 9.005 0.660 ;
        END
    END d
END ao22s80

MACRO ao22m01
    CLASS CORE ;
    FOREIGN ao22m01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.010 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.295 0.090 0.360 1.455 ;
        RECT  0.250 0.090 0.575 0.155 ;
        RECT  0.460 0.090 0.525 0.480 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.725 0.530 0.920 0.660 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.555 0.530 0.750 0.660 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  -0.015 0.530 0.245 0.660 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.385 0.530 0.580 0.660 ;
        END
    END d
END ao22m01

MACRO ao22m02
    CLASS CORE ;
    FOREIGN ao22m02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.785 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.805 0.090 1.060 1.455 ;
        RECT  0.695 0.090 1.605 0.155 ;
        RECT  1.260 0.090 1.520 0.480 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.015 0.530 2.470 0.660 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.550 0.530 2.005 0.660 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  -0.040 0.530 0.670 0.660 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.085 0.530 1.540 0.660 ;
        END
    END d
END ao22m02

MACRO ao22m03
    CLASS CORE ;
    FOREIGN ao22m03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.545 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.020 0.090 1.345 1.455 ;
        RECT  0.885 0.090 2.050 0.155 ;
        RECT  1.605 0.090 1.930 0.480 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.565 0.530 3.150 0.660 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.975 0.530 2.560 0.660 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  -0.050 0.530 0.855 0.660 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.385 0.530 1.970 0.660 ;
        END
    END d
END ao22m03

MACRO ao22m04
    CLASS CORE ;
    FOREIGN ao22m04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.050 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.180 0.090 1.505 1.455 ;
        RECT  1.005 0.090 2.370 0.155 ;
        RECT  1.845 0.090 2.170 0.480 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.940 0.530 3.590 0.660 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.260 0.530 2.915 0.660 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  -0.060 0.530 0.980 0.660 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.585 0.530 2.235 0.660 ;
        END
    END d
END ao22m04

MACRO ao22m06
    CLASS CORE ;
    FOREIGN ao22m06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.810 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.400 0.090 1.785 1.455 ;
        RECT  1.190 0.090 2.815 0.155 ;
        RECT  2.195 0.090 2.585 0.480 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.485 0.530 4.265 0.660 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.690 0.530 3.465 0.660 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  -0.070 0.530 1.160 0.660 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.880 0.530 2.665 0.660 ;
        END
    END d
END ao22m06

MACRO ao22m08
    CLASS CORE ;
    FOREIGN ao22m08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.570 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.620 0.090 2.075 1.455 ;
        RECT  1.395 0.090 3.215 0.155 ;
        RECT  2.535 0.090 2.990 0.480 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.040 0.530 4.950 0.660 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.110 0.530 4.015 0.660 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  -0.065 0.530 1.295 0.660 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.180 0.530 3.090 0.660 ;
        END
    END d
END ao22m08

MACRO ao22m10
    CLASS CORE ;
    FOREIGN ao22m10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.075 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.765 0.090 2.285 1.455 ;
        RECT  1.515 0.090 3.530 0.155 ;
        RECT  2.765 0.090 3.280 0.480 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.405 0.530 5.380 0.660 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.395 0.530 4.370 0.660 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  -0.075 0.530 1.415 0.660 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.380 0.530 3.355 0.660 ;
        END
    END d
END ao22m10

MACRO ao22m20
    CLASS CORE ;
    FOREIGN ao22m20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.610 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.505 0.090 3.220 1.455 ;
        RECT  2.150 0.090 5.005 0.155 ;
        RECT  3.920 0.090 4.635 0.480 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.240 0.530 7.670 0.660 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.805 0.530 6.230 0.660 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  -0.110 0.530 2.030 0.660 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.365 0.530 4.795 0.660 ;
        END
    END d
END ao22m20

MACRO ao22m40
    CLASS CORE ;
    FOREIGN ao22m40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.650 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.385 0.090 4.360 1.455 ;
        RECT  2.900 0.090 6.800 0.155 ;
        RECT  5.300 0.090 6.275 0.480 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.450 0.530 10.335 0.660 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.505 0.530 8.390 0.660 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  -0.155 0.530 2.765 0.660 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.560 0.530 6.445 0.660 ;
        END
    END d
END ao22m40

MACRO ao22m80
    CLASS CORE ;
    FOREIGN ao22m80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.210 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.710 0.090 6.075 1.455 ;
        RECT  4.040 0.090 9.435 0.155 ;
        RECT  7.375 0.090 8.740 0.480 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.750 0.530 14.415 0.660 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.045 0.530 11.710 0.660 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  -0.205 0.530 3.815 0.660 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.340 0.530 9.005 0.660 ;
        END
    END d
END ao22m80

MACRO ao22f01
    CLASS CORE ;
    FOREIGN ao22f01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.010 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.295 0.090 0.360 1.455 ;
        RECT  0.250 0.090 0.575 0.155 ;
        RECT  0.460 0.090 0.525 0.480 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.725 0.530 0.920 0.660 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.555 0.530 0.750 0.660 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  -0.015 0.530 0.245 0.660 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.385 0.530 0.580 0.660 ;
        END
    END d
END ao22f01

MACRO ao22f02
    CLASS CORE ;
    FOREIGN ao22f02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.785 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.805 0.090 1.060 1.455 ;
        RECT  0.695 0.090 1.605 0.155 ;
        RECT  1.260 0.090 1.520 0.480 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.015 0.530 2.470 0.660 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.550 0.530 2.005 0.660 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  -0.040 0.530 0.670 0.660 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.085 0.530 1.540 0.660 ;
        END
    END d
END ao22f02

MACRO ao22f03
    CLASS CORE ;
    FOREIGN ao22f03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.545 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.020 0.090 1.345 1.455 ;
        RECT  0.885 0.090 2.050 0.155 ;
        RECT  1.605 0.090 1.930 0.480 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.565 0.530 3.150 0.660 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.975 0.530 2.560 0.660 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  -0.050 0.530 0.855 0.660 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.385 0.530 1.970 0.660 ;
        END
    END d
END ao22f03

MACRO ao22f04
    CLASS CORE ;
    FOREIGN ao22f04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.050 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.180 0.090 1.505 1.455 ;
        RECT  1.005 0.090 2.370 0.155 ;
        RECT  1.845 0.090 2.170 0.480 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.940 0.530 3.590 0.660 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.260 0.530 2.915 0.660 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  -0.060 0.530 0.980 0.660 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.585 0.530 2.235 0.660 ;
        END
    END d
END ao22f04

MACRO ao22f06
    CLASS CORE ;
    FOREIGN ao22f06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.810 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.400 0.090 1.785 1.455 ;
        RECT  1.190 0.090 2.815 0.155 ;
        RECT  2.195 0.090 2.585 0.480 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.485 0.530 4.265 0.660 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.690 0.530 3.465 0.660 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  -0.070 0.530 1.160 0.660 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.880 0.530 2.665 0.660 ;
        END
    END d
END ao22f06

MACRO ao22f08
    CLASS CORE ;
    FOREIGN ao22f08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.570 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.620 0.090 2.075 1.455 ;
        RECT  1.395 0.090 3.215 0.155 ;
        RECT  2.535 0.090 2.990 0.480 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.040 0.530 4.950 0.660 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.110 0.530 4.015 0.660 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  -0.065 0.530 1.295 0.660 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.180 0.530 3.090 0.660 ;
        END
    END d
END ao22f08

MACRO ao22f10
    CLASS CORE ;
    FOREIGN ao22f10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.075 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.765 0.090 2.285 1.455 ;
        RECT  1.515 0.090 3.530 0.155 ;
        RECT  2.765 0.090 3.280 0.480 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.405 0.530 5.380 0.660 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.395 0.530 4.370 0.660 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  -0.075 0.530 1.415 0.660 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.380 0.530 3.355 0.660 ;
        END
    END d
END ao22f10

MACRO ao22f20
    CLASS CORE ;
    FOREIGN ao22f20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.610 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.505 0.090 3.220 1.455 ;
        RECT  2.150 0.090 5.005 0.155 ;
        RECT  3.920 0.090 4.635 0.480 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.240 0.530 7.670 0.660 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.805 0.530 6.230 0.660 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  -0.110 0.530 2.030 0.660 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.365 0.530 4.795 0.660 ;
        END
    END d
END ao22f20

MACRO ao22f40
    CLASS CORE ;
    FOREIGN ao22f40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.650 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.385 0.090 4.360 1.455 ;
        RECT  2.900 0.090 6.800 0.155 ;
        RECT  5.300 0.090 6.275 0.480 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.450 0.530 10.335 0.660 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.505 0.530 8.390 0.660 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  -0.155 0.530 2.765 0.660 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.560 0.530 6.445 0.660 ;
        END
    END d
END ao22f40

MACRO ao22f80
    CLASS CORE ;
    FOREIGN ao22f80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.210 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.710 0.090 6.075 1.455 ;
        RECT  4.040 0.090 9.435 0.155 ;
        RECT  7.375 0.090 8.740 0.480 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.750 0.530 14.415 0.660 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.045 0.530 11.710 0.660 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  -0.205 0.530 3.815 0.660 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.340 0.530 9.005 0.660 ;
        END
    END d
END ao22f80

MACRO oa12s01
    CLASS CORE ;
    FOREIGN oa12s01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.010 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.550 0.650 0.675 1.235 ;
        RECT  0.460 0.900 0.655 1.225 ;
        RECT  0.710 0.135 0.840 0.720 ;
        RECT  0.515 0.650 0.840 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.130 0.720 0.325 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.345 0.720 0.475 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.675 0.740 0.870 0.805 ;
        END
    END c
END oa12s01

MACRO oa12s02
    CLASS CORE ;
    FOREIGN oa12s02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.530 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.390 0.650 1.650 1.235 ;
        RECT  1.155 0.900 1.680 1.225 ;
        RECT  1.790 0.135 2.045 0.720 ;
        RECT  1.285 0.650 2.130 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.340 0.720 0.795 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.865 0.720 1.190 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.690 0.740 2.210 0.805 ;
        END
    END c
END oa12s02

MACRO oa12s03
    CLASS CORE ;
    FOREIGN oa12s03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.035 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.660 0.650 1.985 1.235 ;
        RECT  1.385 0.900 2.035 1.225 ;
        RECT  2.140 0.135 2.465 0.720 ;
        RECT  1.545 0.650 2.585 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.415 0.720 0.935 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.040 0.720 1.435 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.035 0.740 2.620 0.805 ;
        END
    END c
END oa12s03

MACRO oa12s04
    CLASS CORE ;
    FOREIGN oa12s04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.545 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.940 0.650 2.330 1.235 ;
        RECT  1.615 0.900 2.390 1.225 ;
        RECT  2.500 0.135 2.885 0.720 ;
        RECT  1.795 0.650 3.030 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.485 0.720 1.070 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.215 0.720 1.670 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.370 0.740 3.085 0.805 ;
        END
    END c
END oa12s04

MACRO oa12s06
    CLASS CORE ;
    FOREIGN oa12s06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.305 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.355 0.650 2.810 1.235 ;
        RECT  1.965 0.900 2.875 1.225 ;
        RECT  3.035 0.135 3.490 0.720 ;
        RECT  2.195 0.650 3.625 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.575 0.720 1.355 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.490 0.720 2.005 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.880 0.740 3.725 0.805 ;
        END
    END c
END oa12s06

MACRO oa12s08
    CLASS CORE ;
    FOREIGN oa12s08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.065 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.780 0.650 3.300 1.235 ;
        RECT  2.305 0.900 3.410 1.225 ;
        RECT  3.580 0.135 4.095 0.720 ;
        RECT  2.580 0.650 4.270 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.685 0.720 1.595 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.735 0.720 2.390 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.395 0.740 4.370 0.805 ;
        END
    END c
END oa12s08

MACRO oa12s10
    CLASS CORE ;
    FOREIGN oa12s10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.570 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.050 0.650 3.635 1.235 ;
        RECT  2.545 0.900 3.715 1.225 ;
        RECT  3.930 0.135 4.515 0.720 ;
        RECT  2.835 0.650 4.720 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.755 0.720 1.730 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.915 0.720 2.630 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.730 0.740 4.835 0.805 ;
        END
    END c
END oa12s10

MACRO oa12s20
    CLASS CORE ;
    FOREIGN oa12s20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.160 0.650 4.945 1.235 ;
        RECT  3.465 0.900 5.090 1.225 ;
        RECT  5.370 0.135 6.145 0.720 ;
        RECT  3.860 0.650 6.465 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.040 0.720 2.335 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.615 0.720 3.590 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.085 0.740 6.580 0.805 ;
        END
    END c
END oa12s20

MACRO oa12s40
    CLASS CORE ;
    FOREIGN oa12s40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.385 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.695 0.650 6.740 1.235 ;
        RECT  4.740 0.900 6.945 1.225 ;
        RECT  7.340 0.135 8.375 0.720 ;
        RECT  5.290 0.650 8.800 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.420 0.720 3.240 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.580 0.720 4.880 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.945 0.740 9.025 0.805 ;
        END
    END c
END oa12s40

MACRO oa12s80
    CLASS CORE ;
    FOREIGN oa12s80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.440 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.915 0.650 9.410 1.235 ;
        RECT  6.595 0.900 9.650 1.225 ;
        RECT  10.195 0.135 11.690 0.720 ;
        RECT  7.355 0.650 12.230 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.965 0.720 4.500 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.980 0.720 6.795 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.670 0.740 12.525 0.805 ;
        END
    END c
END oa12s80

MACRO oa12m01
    CLASS CORE ;
    FOREIGN oa12m01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.010 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.550 0.650 0.675 1.235 ;
        RECT  0.460 0.900 0.655 1.225 ;
        RECT  0.710 0.135 0.840 0.720 ;
        RECT  0.515 0.650 0.840 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.130 0.720 0.325 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.345 0.720 0.475 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.675 0.740 0.870 0.805 ;
        END
    END c
END oa12m01

MACRO oa12m02
    CLASS CORE ;
    FOREIGN oa12m02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.530 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.390 0.650 1.650 1.235 ;
        RECT  1.155 0.900 1.680 1.225 ;
        RECT  1.790 0.135 2.045 0.720 ;
        RECT  1.285 0.650 2.130 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.340 0.720 0.795 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.865 0.720 1.190 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.690 0.740 2.210 0.805 ;
        END
    END c
END oa12m02

MACRO oa12m03
    CLASS CORE ;
    FOREIGN oa12m03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.035 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.660 0.650 1.985 1.235 ;
        RECT  1.385 0.900 2.035 1.225 ;
        RECT  2.140 0.135 2.465 0.720 ;
        RECT  1.545 0.650 2.585 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.415 0.720 0.935 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.040 0.720 1.435 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.035 0.740 2.620 0.805 ;
        END
    END c
END oa12m03

MACRO oa12m04
    CLASS CORE ;
    FOREIGN oa12m04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.545 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.940 0.650 2.330 1.235 ;
        RECT  1.615 0.900 2.390 1.225 ;
        RECT  2.500 0.135 2.885 0.720 ;
        RECT  1.795 0.650 3.030 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.485 0.720 1.070 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.215 0.720 1.670 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.370 0.740 3.085 0.805 ;
        END
    END c
END oa12m04

MACRO oa12m06
    CLASS CORE ;
    FOREIGN oa12m06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.305 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.355 0.650 2.810 1.235 ;
        RECT  1.965 0.900 2.875 1.225 ;
        RECT  3.035 0.135 3.490 0.720 ;
        RECT  2.195 0.650 3.625 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.575 0.720 1.355 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.490 0.720 2.005 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.880 0.740 3.725 0.805 ;
        END
    END c
END oa12m06

MACRO oa12m08
    CLASS CORE ;
    FOREIGN oa12m08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.065 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.780 0.650 3.300 1.235 ;
        RECT  2.305 0.900 3.410 1.225 ;
        RECT  3.580 0.135 4.095 0.720 ;
        RECT  2.580 0.650 4.270 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.685 0.720 1.595 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.735 0.720 2.390 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.395 0.740 4.370 0.805 ;
        END
    END c
END oa12m08

MACRO oa12m10
    CLASS CORE ;
    FOREIGN oa12m10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.570 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.050 0.650 3.635 1.235 ;
        RECT  2.545 0.900 3.715 1.225 ;
        RECT  3.930 0.135 4.515 0.720 ;
        RECT  2.835 0.650 4.720 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.755 0.720 1.730 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.915 0.720 2.630 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.730 0.740 4.835 0.805 ;
        END
    END c
END oa12m10

MACRO oa12m20
    CLASS CORE ;
    FOREIGN oa12m20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.160 0.650 4.945 1.235 ;
        RECT  3.465 0.900 5.090 1.225 ;
        RECT  5.370 0.135 6.145 0.720 ;
        RECT  3.860 0.650 6.465 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.040 0.720 2.335 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.615 0.720 3.590 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.085 0.740 6.580 0.805 ;
        END
    END c
END oa12m20

MACRO oa12m40
    CLASS CORE ;
    FOREIGN oa12m40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.385 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.695 0.650 6.740 1.235 ;
        RECT  4.740 0.900 6.945 1.225 ;
        RECT  7.340 0.135 8.375 0.720 ;
        RECT  5.290 0.650 8.800 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.420 0.720 3.240 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.580 0.720 4.880 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.945 0.740 9.025 0.805 ;
        END
    END c
END oa12m40

MACRO oa12m80
    CLASS CORE ;
    FOREIGN oa12m80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.440 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.915 0.650 9.410 1.235 ;
        RECT  6.595 0.900 9.650 1.225 ;
        RECT  10.195 0.135 11.690 0.720 ;
        RECT  7.355 0.650 12.230 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.965 0.720 4.500 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.980 0.720 6.795 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.670 0.740 12.525 0.805 ;
        END
    END c
END oa12m80

MACRO oa12f01
    CLASS CORE ;
    FOREIGN oa12f01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.010 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.550 0.650 0.675 1.235 ;
        RECT  0.460 0.900 0.655 1.225 ;
        RECT  0.710 0.135 0.840 0.720 ;
        RECT  0.515 0.650 0.840 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.130 0.720 0.325 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.345 0.720 0.475 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.675 0.740 0.870 0.805 ;
        END
    END c
END oa12f01

MACRO oa12f02
    CLASS CORE ;
    FOREIGN oa12f02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.530 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.390 0.650 1.650 1.235 ;
        RECT  1.155 0.900 1.680 1.225 ;
        RECT  1.790 0.135 2.045 0.720 ;
        RECT  1.285 0.650 2.130 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.340 0.720 0.795 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.865 0.720 1.190 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.690 0.740 2.210 0.805 ;
        END
    END c
END oa12f02

MACRO oa12f03
    CLASS CORE ;
    FOREIGN oa12f03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.035 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.660 0.650 1.985 1.235 ;
        RECT  1.385 0.900 2.035 1.225 ;
        RECT  2.140 0.135 2.465 0.720 ;
        RECT  1.545 0.650 2.585 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.415 0.720 0.935 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.040 0.720 1.435 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.035 0.740 2.620 0.805 ;
        END
    END c
END oa12f03

MACRO oa12f04
    CLASS CORE ;
    FOREIGN oa12f04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.545 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.940 0.650 2.330 1.235 ;
        RECT  1.615 0.900 2.390 1.225 ;
        RECT  2.500 0.135 2.885 0.720 ;
        RECT  1.795 0.650 3.030 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.485 0.720 1.070 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.215 0.720 1.670 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.370 0.740 3.085 0.805 ;
        END
    END c
END oa12f04

MACRO oa12f06
    CLASS CORE ;
    FOREIGN oa12f06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.305 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.355 0.650 2.810 1.235 ;
        RECT  1.965 0.900 2.875 1.225 ;
        RECT  3.035 0.135 3.490 0.720 ;
        RECT  2.195 0.650 3.625 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.575 0.720 1.355 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.490 0.720 2.005 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.880 0.740 3.725 0.805 ;
        END
    END c
END oa12f06

MACRO oa12f08
    CLASS CORE ;
    FOREIGN oa12f08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.065 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.780 0.650 3.300 1.235 ;
        RECT  2.305 0.900 3.410 1.225 ;
        RECT  3.580 0.135 4.095 0.720 ;
        RECT  2.580 0.650 4.270 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.685 0.720 1.595 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.735 0.720 2.390 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.395 0.740 4.370 0.805 ;
        END
    END c
END oa12f08

MACRO oa12f10
    CLASS CORE ;
    FOREIGN oa12f10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.570 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.050 0.650 3.635 1.235 ;
        RECT  2.545 0.900 3.715 1.225 ;
        RECT  3.930 0.135 4.515 0.720 ;
        RECT  2.835 0.650 4.720 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.755 0.720 1.730 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.915 0.720 2.630 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.730 0.740 4.835 0.805 ;
        END
    END c
END oa12f10

MACRO oa12f20
    CLASS CORE ;
    FOREIGN oa12f20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.160 0.650 4.945 1.235 ;
        RECT  3.465 0.900 5.090 1.225 ;
        RECT  5.370 0.135 6.145 0.720 ;
        RECT  3.860 0.650 6.465 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.040 0.720 2.335 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.615 0.720 3.590 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.085 0.740 6.580 0.805 ;
        END
    END c
END oa12f20

MACRO oa12f40
    CLASS CORE ;
    FOREIGN oa12f40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.385 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.695 0.650 6.740 1.235 ;
        RECT  4.740 0.900 6.945 1.225 ;
        RECT  7.340 0.135 8.375 0.720 ;
        RECT  5.290 0.650 8.800 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.420 0.720 3.240 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.580 0.720 4.880 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.945 0.740 9.025 0.805 ;
        END
    END c
END oa12f40

MACRO oa12f80
    CLASS CORE ;
    FOREIGN oa12f80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.440 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.915 0.650 9.410 1.235 ;
        RECT  6.595 0.900 9.650 1.225 ;
        RECT  10.195 0.135 11.690 0.720 ;
        RECT  7.355 0.650 12.230 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.965 0.720 4.500 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.980 0.720 6.795 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.670 0.740 12.525 0.805 ;
        END
    END c
END oa12f80

MACRO oa22s01
    CLASS CORE ;
    FOREIGN oa22s01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.010 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.295 0.210 0.360 0.925 ;
        RECT  0.250 0.870 0.575 0.935 ;
        RECT  0.460 0.870 0.525 1.520 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.725 0.725 0.920 0.790 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.555 0.725 0.750 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.105 0.635 0.300 0.700 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.385 0.725 0.580 0.790 ;
        END
    END d
END oa22s01

MACRO oa22s02
    CLASS CORE ;
    FOREIGN oa22s02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.785 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.805 0.210 1.060 0.925 ;
        RECT  0.695 0.870 1.605 0.935 ;
        RECT  1.270 0.870 1.530 1.520 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.015 0.725 2.470 0.790 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.550 0.725 2.005 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.305 0.635 0.760 0.700 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.085 0.725 1.540 0.790 ;
        END
    END d
END oa22s02

MACRO oa22s03
    CLASS CORE ;
    FOREIGN oa22s03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.545 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.020 0.210 1.345 0.925 ;
        RECT  0.885 0.870 2.050 0.935 ;
        RECT  1.615 0.870 1.940 1.520 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.565 0.725 3.150 0.790 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.975 0.725 2.560 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.390 0.635 0.975 0.700 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.385 0.725 1.970 0.790 ;
        END
    END d
END oa22s03

MACRO oa22s04
    CLASS CORE ;
    FOREIGN oa22s04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.050 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.180 0.210 1.505 0.925 ;
        RECT  1.005 0.870 2.370 0.935 ;
        RECT  1.850 0.870 2.175 1.520 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.940 0.725 3.590 0.790 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.260 0.725 2.915 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.450 0.635 1.100 0.700 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.585 0.725 2.235 0.790 ;
        END
    END d
END oa22s04

MACRO oa22s06
    CLASS CORE ;
    FOREIGN oa22s06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.810 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.400 0.210 1.785 0.925 ;
        RECT  1.190 0.870 2.815 0.935 ;
        RECT  2.205 0.870 2.590 1.520 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.485 0.725 4.265 0.790 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.690 0.725 3.465 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.530 0.635 1.310 0.700 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.880 0.725 2.665 0.790 ;
        END
    END d
END oa22s06

MACRO oa22s08
    CLASS CORE ;
    FOREIGN oa22s08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.570 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.620 0.210 2.075 0.925 ;
        RECT  1.380 0.870 3.265 0.935 ;
        RECT  2.545 0.870 3.000 1.520 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.040 0.725 4.950 0.790 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.110 0.725 4.015 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.615 0.635 1.525 0.700 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.180 0.725 3.090 0.790 ;
        END
    END d
END oa22s08

MACRO oa22s10
    CLASS CORE ;
    FOREIGN oa22s10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.075 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.765 0.210 2.285 0.925 ;
        RECT  1.515 0.870 3.530 0.935 ;
        RECT  2.780 0.870 3.300 1.520 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.405 0.725 5.380 0.790 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.395 0.725 4.370 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.675 0.635 1.650 0.700 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.380 0.725 3.355 0.790 ;
        END
    END d
END oa22s10

MACRO oa22s20
    CLASS CORE ;
    FOREIGN oa22s20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.610 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.505 0.210 3.220 0.925 ;
        RECT  2.150 0.870 5.005 0.935 ;
        RECT  3.935 0.870 4.650 1.520 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.240 0.725 7.670 0.790 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.805 0.725 6.230 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.950 0.635 2.375 0.700 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.365 0.725 4.795 0.790 ;
        END
    END d
END oa22s20

MACRO oa22s40
    CLASS CORE ;
    FOREIGN oa22s40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.650 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.385 0.210 4.360 0.925 ;
        RECT  2.900 0.870 6.800 0.935 ;
        RECT  5.325 0.870 6.300 1.520 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.450 0.725 10.335 0.790 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.505 0.725 8.390 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.290 0.635 3.175 0.700 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.560 0.725 6.445 0.790 ;
        END
    END d
END oa22s40

MACRO oa22s80
    CLASS CORE ;
    FOREIGN oa22s80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.210 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.710 0.210 6.075 0.925 ;
        RECT  4.025 0.870 9.490 0.935 ;
        RECT  7.410 0.870 8.775 1.520 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.750 0.725 14.415 0.790 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.045 0.725 11.710 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.790 0.635 4.455 0.700 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.340 0.725 9.005 0.790 ;
        END
    END d
END oa22s80

MACRO oa22m01
    CLASS CORE ;
    FOREIGN oa22m01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.010 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.295 0.210 0.360 0.925 ;
        RECT  0.250 0.870 0.575 0.935 ;
        RECT  0.460 0.870 0.525 1.520 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.725 0.725 0.920 0.790 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.555 0.725 0.750 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.105 0.635 0.300 0.700 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.385 0.725 0.580 0.790 ;
        END
    END d
END oa22m01

MACRO oa22m02
    CLASS CORE ;
    FOREIGN oa22m02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.785 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.805 0.210 1.060 0.925 ;
        RECT  0.695 0.870 1.605 0.935 ;
        RECT  1.270 0.870 1.530 1.520 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.015 0.725 2.470 0.790 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.550 0.725 2.005 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.305 0.635 0.760 0.700 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.085 0.725 1.540 0.790 ;
        END
    END d
END oa22m02

MACRO oa22m03
    CLASS CORE ;
    FOREIGN oa22m03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.545 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.020 0.210 1.345 0.925 ;
        RECT  0.885 0.870 2.050 0.935 ;
        RECT  1.615 0.870 1.940 1.520 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.565 0.725 3.150 0.790 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.975 0.725 2.560 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.390 0.635 0.975 0.700 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.385 0.725 1.970 0.790 ;
        END
    END d
END oa22m03

MACRO oa22m04
    CLASS CORE ;
    FOREIGN oa22m04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.050 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.180 0.210 1.505 0.925 ;
        RECT  1.005 0.870 2.370 0.935 ;
        RECT  1.850 0.870 2.175 1.520 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.940 0.725 3.590 0.790 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.260 0.725 2.915 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.450 0.635 1.100 0.700 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.585 0.725 2.235 0.790 ;
        END
    END d
END oa22m04

MACRO oa22m06
    CLASS CORE ;
    FOREIGN oa22m06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.810 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.400 0.210 1.785 0.925 ;
        RECT  1.190 0.870 2.815 0.935 ;
        RECT  2.205 0.870 2.590 1.520 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.485 0.725 4.265 0.790 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.690 0.725 3.465 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.530 0.635 1.310 0.700 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.880 0.725 2.665 0.790 ;
        END
    END d
END oa22m06

MACRO oa22m08
    CLASS CORE ;
    FOREIGN oa22m08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.570 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.620 0.210 2.075 0.925 ;
        RECT  1.380 0.870 3.265 0.935 ;
        RECT  2.545 0.870 3.000 1.520 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.040 0.725 4.950 0.790 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.110 0.725 4.015 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.615 0.635 1.525 0.700 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.180 0.725 3.090 0.790 ;
        END
    END d
END oa22m08

MACRO oa22m10
    CLASS CORE ;
    FOREIGN oa22m10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.075 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.765 0.210 2.285 0.925 ;
        RECT  1.515 0.870 3.530 0.935 ;
        RECT  2.780 0.870 3.300 1.520 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.405 0.725 5.380 0.790 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.395 0.725 4.370 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.675 0.635 1.650 0.700 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.380 0.725 3.355 0.790 ;
        END
    END d
END oa22m10

MACRO oa22m20
    CLASS CORE ;
    FOREIGN oa22m20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.610 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.505 0.210 3.220 0.925 ;
        RECT  2.150 0.870 5.005 0.935 ;
        RECT  3.935 0.870 4.650 1.520 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.240 0.725 7.670 0.790 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.805 0.725 6.230 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.950 0.635 2.375 0.700 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.365 0.725 4.795 0.790 ;
        END
    END d
END oa22m20

MACRO oa22m40
    CLASS CORE ;
    FOREIGN oa22m40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.650 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.385 0.210 4.360 0.925 ;
        RECT  2.900 0.870 6.800 0.935 ;
        RECT  5.325 0.870 6.300 1.520 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.450 0.725 10.335 0.790 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.505 0.725 8.390 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.290 0.635 3.175 0.700 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.560 0.725 6.445 0.790 ;
        END
    END d
END oa22m40

MACRO oa22m80
    CLASS CORE ;
    FOREIGN oa22m80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.210 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.710 0.210 6.075 0.925 ;
        RECT  4.025 0.870 9.490 0.935 ;
        RECT  7.410 0.870 8.775 1.520 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.750 0.725 14.415 0.790 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.045 0.725 11.710 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.790 0.635 4.455 0.700 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.340 0.725 9.005 0.790 ;
        END
    END d
END oa22m80

MACRO oa22f01
    CLASS CORE ;
    FOREIGN oa22f01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.010 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.295 0.210 0.360 0.925 ;
        RECT  0.250 0.870 0.575 0.935 ;
        RECT  0.460 0.870 0.525 1.520 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.725 0.725 0.920 0.790 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.555 0.725 0.750 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.105 0.635 0.300 0.700 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.385 0.725 0.580 0.790 ;
        END
    END d
END oa22f01

MACRO oa22f02
    CLASS CORE ;
    FOREIGN oa22f02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.785 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.805 0.210 1.060 0.925 ;
        RECT  0.695 0.870 1.605 0.935 ;
        RECT  1.270 0.870 1.530 1.520 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.015 0.725 2.470 0.790 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.550 0.725 2.005 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.305 0.635 0.760 0.700 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.085 0.725 1.540 0.790 ;
        END
    END d
END oa22f02

MACRO oa22f03
    CLASS CORE ;
    FOREIGN oa22f03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.545 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.020 0.210 1.345 0.925 ;
        RECT  0.885 0.870 2.050 0.935 ;
        RECT  1.615 0.870 1.940 1.520 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.565 0.725 3.150 0.790 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.975 0.725 2.560 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.390 0.635 0.975 0.700 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.385 0.725 1.970 0.790 ;
        END
    END d
END oa22f03

MACRO oa22f04
    CLASS CORE ;
    FOREIGN oa22f04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.050 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.180 0.210 1.505 0.925 ;
        RECT  1.005 0.870 2.370 0.935 ;
        RECT  1.850 0.870 2.175 1.520 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.940 0.725 3.590 0.790 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.260 0.725 2.915 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.450 0.635 1.100 0.700 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.585 0.725 2.235 0.790 ;
        END
    END d
END oa22f04

MACRO oa22f06
    CLASS CORE ;
    FOREIGN oa22f06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.810 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.400 0.210 1.785 0.925 ;
        RECT  1.190 0.870 2.815 0.935 ;
        RECT  2.205 0.870 2.590 1.520 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.485 0.725 4.265 0.790 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.690 0.725 3.465 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.530 0.635 1.310 0.700 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.880 0.725 2.665 0.790 ;
        END
    END d
END oa22f06

MACRO oa22f08
    CLASS CORE ;
    FOREIGN oa22f08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.570 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.620 0.210 2.075 0.925 ;
        RECT  1.380 0.870 3.265 0.935 ;
        RECT  2.545 0.870 3.000 1.520 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.040 0.725 4.950 0.790 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.110 0.725 4.015 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.615 0.635 1.525 0.700 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.180 0.725 3.090 0.790 ;
        END
    END d
END oa22f08

MACRO oa22f10
    CLASS CORE ;
    FOREIGN oa22f10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.075 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.765 0.210 2.285 0.925 ;
        RECT  1.515 0.870 3.530 0.935 ;
        RECT  2.780 0.870 3.300 1.520 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.405 0.725 5.380 0.790 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.395 0.725 4.370 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.675 0.635 1.650 0.700 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.380 0.725 3.355 0.790 ;
        END
    END d
END oa22f10

MACRO oa22f20
    CLASS CORE ;
    FOREIGN oa22f20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.610 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.505 0.210 3.220 0.925 ;
        RECT  2.150 0.870 5.005 0.935 ;
        RECT  3.935 0.870 4.650 1.520 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.240 0.725 7.670 0.790 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.805 0.725 6.230 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.950 0.635 2.375 0.700 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.365 0.725 4.795 0.790 ;
        END
    END d
END oa22f20

MACRO oa22f40
    CLASS CORE ;
    FOREIGN oa22f40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.650 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.385 0.210 4.360 0.925 ;
        RECT  2.900 0.870 6.800 0.935 ;
        RECT  5.325 0.870 6.300 1.520 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.450 0.725 10.335 0.790 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.505 0.725 8.390 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.290 0.635 3.175 0.700 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.560 0.725 6.445 0.790 ;
        END
    END d
END oa22f40

MACRO oa22f80
    CLASS CORE ;
    FOREIGN oa22f80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.210 BY 1.710 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.710 0.210 6.075 0.925 ;
        RECT  4.025 0.870 9.490 0.935 ;
        RECT  7.410 0.870 8.775 1.520 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.750 0.725 14.415 0.790 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.045 0.725 11.710 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.790 0.635 4.455 0.700 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.340 0.725 9.005 0.790 ;
        END
    END d
END oa22f80

MACRO ms00f20
    CLASS CORE ;
    FOREIGN ms00f20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.75 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.19 0.15 0.45 1.58 ;
        RECT 0.19 0.635 0.775 0.7 ;
        RECT 0.19 1.14 1.62 1.205 ;
        END
    END o
    PIN ck
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.6375 0.99 2.8975 1.38 ;
        RECT 2.635 0.705 2.895 1.03 ;
        RECT 2.63 1.47 4.055 1.535 ;
        RECT 3.8 0.775 4.06 1.49 ;
        RECT 3.5 0.775 4.02 0.84 ;
        RECT 2.6375 1.29 2.8975 1.485 ;
        RECT 2.6375 1.315 2.8975 1.38 ;
        RECT 1.3525 0.78 1.8075 0.845 ;
        RECT 1.6025 0.64 1.8625 0.835 ;
        RECT 1.6025 0.64 2.895 0.705 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.36 0.72 4.62 0.785 ;
        END
    END d
END ms00f20

MACRO ms00f40
    CLASS CORE ;
    FOREIGN ms00f40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.84 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.19 0.15 0.45 1.58 ;
        RECT 0.19 0.635 0.775 0.7 ;
        RECT 0.19 1.14 1.62 1.205 ;
        END
    END o
    PIN ck
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.7125 0.99 3.9725 1.38 ;
        RECT 3.71 0.705 3.97 1.03 ;
        RECT 3.705 1.47 5.13 1.535 ;
        RECT 4.875 0.775 5.135 1.49 ;
        RECT 4.575 0.775 5.095 0.84 ;
        RECT 3.7125 1.29 3.9725 1.485 ;
        RECT 3.7125 1.315 3.9725 1.38 ;
        RECT 2.0325 0.78 2.4875 0.845 ;
        RECT 2.2825 0.64 2.5425 0.835 ;
        RECT 2.2825 0.64 3.9725 0.705 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.0325 0.72 6.2925 0.785 ;
        END
    END d
END ms00f40

MACRO ms00f80
    CLASS CORE ;
    FOREIGN ms00f80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.500 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.190 0.150 0.45 1.58 ;
        RECT 0.190 0.635 0.775 0.7 ;
        RECT 0.190 1.140 1.62 1.205 ;
        END
    END o
    PIN ck
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.240 0.990 5.5 1.38 ;
        RECT 5.240 0.990 5.565 1.185 ;
        RECT 1.815 0.640 2.075 0.835 ;
        RECT 1.565 0.780 2.02 0.845 ;
        RECT 1.815 0.640 3.505 0.705 ;
        RECT 2.815 0.640 3.53 0.835 ;
        RECT 4.330 0.705 4.785 0.835 ;
        RECT 2.815 0.790 4.83 0.855 ;
        RECT 4.580 0.705 4.84 1.03 ;
        RECT 4.580 1.015 5.685 1.08 ;
        RECT 5.190 1.015 5.645 1.145 ;
        RECT 5.240 1.290 5.5 1.485 ;
        RECT 7.940 0.775 8.46 0.84 ;
        RECT 8.240 0.775 8.5 1.49 ;
        RECT 5.240 1.470 8.49 1.535 ;
        RECT 5.240 1.315 5.5 1.38 ;
        RECT 5.315 1.110 5.575 1.175 ;
        RECT 5.315 1.015 5.575 1.08 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.705 0.720 8.965 0.785 ;
        END
    END d
END ms00f80

MACRO vcc
    CLASS CORE ;
    FOREIGN vcc 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
				USE SIGNAL ;
        PORT
        LAYER metal1 ;
        RECT 0.925 0.150 1.12 1.255 ;
        RECT 0.835 0.150 1.225 0.28 ;
        END
    END o
END vcc

MACRO vss
    CLASS CORE ;
    FOREIGN vss 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.140 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
				USE SIGNAL ;
        PORT
        LAYER metal1 ;
        RECT 0.695 0.150 0.84 1.255 ;
        RECT 0.625 0.150 0.915 0.28 ;
        END
    END o
END vss

MACRO BLK_NETCARD_TYPE1
  CLASS BLOCK ;
	SIZE 190 BY 598.5 ;
	ORIGIN 0 0 ;
	SITE core ;
END BLK_NETCARD_TYPE1

MACRO BLK_NETCARD_TYPE2
  CLASS BLOCK ;
	SIZE 95 BY 598.5 ;
	ORIGIN 0 0 ;
	SITE core ;
END BLK_NETCARD_TYPE2

MACRO BLK_NETCARD_TYPE3
  CLASS BLOCK ;
	SIZE 190 BY 171 ;
	ORIGIN 0 0 ;
	SITE core ;
END BLK_NETCARD_TYPE3

MACRO BLK_MGC_TYPE1
  CLASS BLOCK ;
	SIZE 38 BY 68.4 ;
	ORIGIN 0 0 ;
	SITE core ;
END BLK_MGC_TYPE1

MACRO BLK_MGC_TYPE2
  CLASS BLOCK ;
	SIZE 38 BY 171 ;
	ORIGIN 0 0 ;
	SITE core ;
END BLK_MGC_TYPE2

END LIBRARY
