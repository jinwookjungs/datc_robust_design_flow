module usb_funct (
x185140,
x6157,
x5961,
x5143,
x3360,
x3320,
x2767,
x5850,
x185135,
x3300,
x3849,
x3613,
x5722,
x3022,
x6102,
x2098,
x3133,
x2214,
x5077,
x2400,
x3558,
x3249,
x185132,
x3653,
x3338,
x6327,
x1459,
x3314,
x6303,
x4851,
x185138,
x3606,
x6282,
x4359,
x6028,
x1418,
x3889,
x3599,
x2890,
x2278,
x5647,
x5548,
x3534,
x4781,
x2648,
x2531,
x6577,
x3307,
x2333,
x5003,
x3949,
x5225,
x1865,
x185141,
x185137,
x6599,
x4117,
x3588,
x1598,
x185130,
x3638,
x1974,
x4041,
x185133,
x6351,
x4285,
x1792,
x3327,
x5790,
x3867,
x4587,
x4937,
x1503,
x185134,
x6445,
x185142,
x6401,
x185136,
x2826,
x3733,
x5601,
x185131,
x5901,
x3645,
x2165,
x3772,
x1660,
x6198,
x2968,
x6186,
x3349,
x3621,
x3683,
x4694,
x2707,
x3828,
x6252,
x6220,
x3574,
x5427,
x2027,
x3675,
x185129,
x4209,
x6531,
x185139,
x5289,
x1911,
x3194,
x2589,
x6264,
x6241,
x3071,
x5498,
x5364,
x3565,
x3858,
x1743,
x4520,
x4449,
x1547,
x3507,
x3698,
x6496,
x2477,
x185128,
x3632,
x3390,
x19,
x715,
x916,
x465,
x91,
x329,
x293,
x86,
x1161,
x507,
x936,
x962,
x355,
x39,
x1329,
x381,
x143,
x348,
x257,
x1192,
x480,
x1215,
x1113,
x277,
x447,
x948,
x316,
x1290,
x1134,
x1121,
x111,
x420,
x921,
x1248,
x101,
x1262,
x784,
x33,
x682,
x957,
x427,
x1074,
x1402,
x1384,
x1274,
x1153,
x906,
x472,
x1357,
x1240,
x1104,
x454,
x244,
x941,
x494,
x401,
x769,
x73,
x297,
x589,
x268,
x1343,
x126,
x341,
x1029,
x926,
x1231,
x1197,
x132,
x1170,
x1066,
x871,
x198,
x374,
x121,
x304,
x813,
x1298,
x798,
x1142,
x80,
x1010,
x747,
x182,
x911,
x555,
x157,
x1313,
x637,
x1370,
x898,
x223,
x65,
x116,
x46,
x1223,
x233,
x285,
x0,
x413,
x166,
x57,
x1129,
x106,
x366,
x1187,
x987,
x27,
x1282,
x1095,
x208,
x890,
x461,
x389,
x526,
x931,
x1058,
x1206,
x1179,
x437,
x732);

// Start PIs
input x185140;
input x6157;
input x5961;
input x5143;
input x3360;
input x3320;
input x2767;
input x5850;
input x185135;
input x3300;
input x3849;
input x3613;
input x5722;
input x3022;
input x6102;
input x2098;
input x3133;
input x2214;
input x5077;
input x2400;
input x3558;
input x3249;
input x185132;
input x3653;
input x3338;
input x6327;
input x1459;
input x3314;
input x6303;
input x4851;
input x185138;
input x3606;
input x6282;
input x4359;
input x6028;
input x1418;
input x3889;
input x3599;
input x2890;
input x2278;
input x5647;
input x5548;
input x3534;
input x4781;
input x2648;
input x2531;
input x6577;
input x3307;
input x2333;
input x5003;
input x3949;
input x5225;
input x1865;
input x185141;
input x185137;
input x6599;
input x4117;
input x3588;
input x1598;
input x185130;
input x3638;
input x1974;
input x4041;
input x185133;
input x6351;
input x4285;
input x1792;
input x3327;
input x5790;
input x3867;
input x4587;
input x4937;
input x1503;
input x185134;
input x6445;
input x185142;
input x6401;
input x185136;
input x2826;
input x3733;
input x5601;
input x185131;
input x5901;
input x3645;
input x2165;
input x3772;
input x1660;
input x6198;
input x2968;
input x6186;
input x3349;
input x3621;
input x3683;
input x4694;
input x2707;
input x3828;
input x6252;
input x6220;
input x3574;
input x5427;
input x2027;
input x3675;
input x185129;
input x4209;
input x6531;
input x185139;
input x5289;
input x1911;
input x3194;
input x2589;
input x6264;
input x6241;
input x3071;
input x5498;
input x5364;
input x3565;
input x3858;
input x1743;
input x4520;
input x4449;
input x1547;
input x3507;
input x3698;
input x6496;
input x2477;
input x185128;
input x3632;
input x3390;

// Start POs
output x19;
output x715;
output x916;
output x465;
output x91;
output x329;
output x293;
output x86;
output x1161;
output x507;
output x936;
output x962;
output x355;
output x39;
output x1329;
output x381;
output x143;
output x348;
output x257;
output x1192;
output x480;
output x1215;
output x1113;
output x277;
output x447;
output x948;
output x316;
output x1290;
output x1134;
output x1121;
output x111;
output x420;
output x921;
output x1248;
output x101;
output x1262;
output x784;
output x33;
output x682;
output x957;
output x427;
output x1074;
output x1402;
output x1384;
output x1274;
output x1153;
output x906;
output x472;
output x1357;
output x1240;
output x1104;
output x454;
output x244;
output x941;
output x494;
output x401;
output x769;
output x73;
output x297;
output x589;
output x268;
output x1343;
output x126;
output x341;
output x1029;
output x926;
output x1231;
output x1197;
output x132;
output x1170;
output x1066;
output x871;
output x198;
output x374;
output x121;
output x304;
output x813;
output x1298;
output x798;
output x1142;
output x80;
output x1010;
output x747;
output x182;
output x911;
output x555;
output x157;
output x1313;
output x637;
output x1370;
output x898;
output x223;
output x65;
output x116;
output x46;
output x1223;
output x233;
output x285;
output x0;
output x413;
output x166;
output x57;
output x1129;
output x106;
output x366;
output x1187;
output x987;
output x27;
output x1282;
output x1095;
output x208;
output x890;
output x461;
output x389;
output x526;
output x931;
output x1058;
output x1206;
output x1179;
output x437;
output x732;

// Start wires
wire net_8298;
wire net_8631;
wire net_4065;
wire net_11968;
wire net_4854;
wire net_2418;
wire net_14672;
wire net_14199;
wire net_7279;
wire net_943;
wire net_11788;
wire net_10413;
wire net_4598;
wire net_4392;
wire net_11330;
wire net_12833;
wire net_1897;
wire net_9435;
wire net_980;
wire net_13088;
wire net_5499;
wire net_9803;
wire net_2542;
wire net_12029;
wire net_7081;
wire net_10629;
wire net_11370;
wire net_5515;
wire net_3996;
wire x2278;
wire net_11996;
wire net_7594;
wire net_15044;
wire net_6241;
wire net_7298;
wire net_4382;
wire net_13988;
wire net_12537;
wire net_13226;
wire net_12501;
wire net_8105;
wire net_4934;
wire net_2256;
wire net_4306;
wire net_264;
wire net_12959;
wire net_11178;
wire net_12809;
wire net_3904;
wire net_4122;
wire net_4315;
wire net_8914;
wire net_11757;
wire net_9072;
wire net_2769;
wire net_8503;
wire net_11190;
wire net_4996;
wire net_14016;
wire net_3707;
wire net_1064;
wire net_14405;
wire net_2082;
wire net_10165;
wire net_6227;
wire net_7173;
wire net_5035;
wire x5790;
wire net_15734;
wire net_12907;
wire net_4832;
wire net_4464;
wire net_8577;
wire net_9784;
wire net_12704;
wire net_13544;
wire net_10988;
wire net_7191;
wire net_703;
wire x5901;
wire net_5330;
wire net_193;
wire net_11377;
wire net_9989;
wire net_12447;
wire net_6037;
wire net_14381;
wire net_10554;
wire net_6773;
wire net_5273;
wire net_12413;
wire net_7283;
wire net_14609;
wire x1313;
wire net_5627;
wire net_2942;
wire net_3817;
wire net_9441;
wire net_13993;
wire net_3281;
wire net_13916;
wire net_10659;
wire net_4442;
wire net_3949;
wire net_3134;
wire net_13458;
wire net_8185;
wire net_10215;
wire net_5523;
wire net_1720;
wire net_14164;
wire net_13885;
wire net_8191;
wire net_6231;
wire net_3818;
wire net_3434;
wire net_15098;
wire net_6104;
wire net_2060;
wire net_2051;
wire net_6087;
wire net_4535;
wire net_9464;
wire net_3756;
wire net_6426;
wire net_593;
wire net_5563;
wire x5961;
wire net_10156;
wire net_6238;
wire net_4169;
wire net_2765;
wire net_15665;
wire net_15085;
wire net_13451;
wire net_7845;
wire net_9957;
wire net_11979;
wire net_742;
wire net_8341;
wire net_5139;
wire net_6384;
wire net_11044;
wire net_12976;
wire net_9597;
wire net_7092;
wire net_10343;
wire net_2830;
wire net_15449;
wire net_10320;
wire net_4509;
wire net_1198;
wire net_3975;
wire net_2862;
wire net_8100;
wire net_2457;
wire net_8260;
wire net_883;
wire net_13476;
wire net_11605;
wire net_8124;
wire net_4108;
wire net_9970;
wire net_5533;
wire net_2957;
wire net_446;
wire net_1516;
wire net_1712;
wire net_6782;
wire net_6473;
wire net_3063;
wire net_1083;
wire net_3423;
wire net_1499;
wire net_964;
wire net_2913;
wire net_8242;
wire net_3295;
wire net_15060;
wire net_13729;
wire net_6402;
wire net_14985;
wire net_11003;
wire net_4379;
wire net_2268;
wire net_10000;
wire net_15141;
wire net_6114;
wire net_14352;
wire net_2846;
wire net_2303;
wire net_13331;
wire net_11685;
wire net_9479;
wire net_4369;
wire net_1735;
wire net_2210;
wire net_8249;
wire net_2176;
wire net_13191;
wire net_11933;
wire net_8563;
wire net_997;
wire net_12243;
wire net_10837;
wire net_6401;
wire x116;
wire net_11060;
wire net_10007;
wire net_256;
wire net_8762;
wire net_4929;
wire net_3959;
wire net_4309;
wire net_8873;
wire net_12393;
wire net_11226;
wire net_6573;
wire net_1140;
wire net_2764;
wire net_1464;
wire net_7490;
wire net_10931;
wire net_5797;
wire net_11985;
wire net_4973;
wire net_12891;
wire net_3196;
wire net_14740;
wire net_5962;
wire net_515;
wire net_4835;
wire net_10620;
wire net_5342;
wire net_13216;
wire net_11124;
wire net_7463;
wire net_6806;
wire net_5121;
wire net_3987;
wire net_223;
wire net_6557;
wire net_15725;
wire net_7146;
wire net_2077;
wire net_15028;
wire net_8468;
wire net_7496;
wire net_2219;
wire net_2745;
wire net_7343;
wire net_11166;
wire net_15657;
wire net_5680;
wire net_13973;
wire net_5084;
wire net_3965;
wire net_13827;
wire net_15008;
wire net_7483;
wire net_1876;
wire net_13130;
wire net_15567;
wire net_6706;
wire net_14611;
wire net_130;
wire net_7212;
wire net_572;
wire net_9810;
wire net_5289;
wire net_15218;
wire net_10955;
wire net_9614;
wire net_5116;
wire net_369;
wire net_12709;
wire net_12051;
wire net_7850;
wire net_1662;
wire net_10396;
wire net_4358;
wire net_14615;
wire net_7543;
wire net_9835;
wire net_1079;
wire net_10495;
wire net_7959;
wire x5003;
wire net_3935;
wire net_15551;
wire net_11290;
wire net_10148;
wire net_6760;
wire net_15273;
wire net_5198;
wire net_2809;
wire net_14318;
wire net_3235;
wire net_780;
wire net_4938;
wire net_3586;
wire net_3184;
wire net_7099;
wire x244;
wire net_6812;
wire net_12226;
wire net_13261;
wire net_9272;
wire net_2391;
wire net_10095;
wire net_5263;
wire net_2802;
wire net_11350;
wire net_7965;
wire net_4614;
wire net_2906;
wire net_456;
wire net_155;
wire net_12555;
wire net_11357;
wire net_9301;
wire net_11299;
wire net_10636;
wire net_7238;
wire net_3850;
wire net_9153;
wire net_9023;
wire net_8222;
wire net_349;
wire net_12923;
wire net_8533;
wire net_14367;
wire net_8547;
wire net_3428;
wire net_1409;
wire net_12576;
wire net_14528;
wire net_2977;
wire net_493;
wire net_6374;
wire net_6080;
wire net_14306;
wire net_13140;
wire net_6506;
wire net_14629;
wire net_13679;
wire net_1428;
wire net_987;
wire net_14518;
wire net_15297;
wire net_13137;
wire net_6167;
wire net_5222;
wire net_3620;
wire net_10510;
wire net_14340;
wire net_7781;
wire net_13824;
wire net_4238;
wire net_5844;
wire net_8475;
wire net_2350;
wire net_6293;
wire net_3271;
wire net_13183;
wire net_11197;
wire net_10675;
wire net_13098;
wire net_12568;
wire net_10506;
wire net_5740;
wire net_14763;
wire net_12276;
wire net_12418;
wire net_721;
wire net_12366;
wire net_9033;
wire net_8950;
wire net_7779;
wire net_3226;
wire net_3143;
wire net_8164;
wire net_15590;
wire net_12127;
wire net_9819;
wire net_2757;
wire net_13634;
wire net_12776;
wire net_9531;
wire net_1018;
wire net_11085;
wire net_3629;
wire net_7315;
wire net_11701;
wire net_2369;
wire net_2038;
wire net_13289;
wire net_6591;
wire net_823;
wire net_9067;
wire net_12878;
wire net_9269;
wire net_1676;
wire net_7271;
wire net_4788;
wire x3653;
wire net_14230;
wire net_698;
wire net_12969;
wire net_11774;
wire net_9541;
wire net_7892;
wire net_14374;
wire net_11028;
wire net_5428;
wire net_1191;
wire net_13688;
wire net_5259;
wire net_8515;
wire net_2255;
wire net_4649;
wire net_4754;
wire net_2485;
wire net_13906;
wire net_6967;
wire net_3857;
wire net_8970;
wire net_7471;
wire net_12918;
wire net_749;
wire net_15053;
wire net_11729;
wire net_1019;
wire net_1948;
wire net_1616;
wire net_11500;
wire net_11898;
wire net_6180;
wire net_10348;
wire net_1006;
wire net_2781;
wire net_9415;
wire net_6767;
wire net_14181;
wire net_4342;
wire net_9724;
wire net_14695;
wire net_12863;
wire net_2969;
wire net_7839;
wire net_7518;
wire net_12522;
wire net_12351;
wire net_5490;
wire net_15253;
wire net_12960;
wire net_13167;
wire net_7544;
wire net_15078;
wire net_11406;
wire net_8886;
wire net_2985;
wire net_11551;
wire net_537;
wire net_3056;
wire net_14050;
wire net_12943;
wire net_11310;
wire net_10893;
wire net_8710;
wire net_12477;
wire net_3614;
wire net_7624;
wire net_13446;
wire net_13007;
wire net_5501;
wire net_12294;
wire net_3252;
wire net_6792;
wire net_5790;
wire net_5891;
wire net_513;
wire net_12020;
wire net_15600;
wire net_7950;
wire net_1576;
wire net_1421;
wire net_14991;
wire net_14282;
wire net_12462;
wire net_9525;
wire net_4496;
wire net_8737;
wire net_6067;
wire net_3407;
wire net_2736;
wire net_2127;
wire net_1280;
wire net_459;
wire net_12616;
wire net_9239;
wire net_8720;
wire net_13569;
wire net_3656;
wire net_737;
wire net_6590;
wire net_2284;
wire net_3412;
wire net_2113;
wire net_13305;
wire net_9397;
wire net_4793;
wire net_5865;
wire net_13372;
wire net_4760;
wire net_3915;
wire net_12737;
wire net_15623;
wire net_14424;
wire net_5957;
wire net_5606;
wire net_11722;
wire net_11541;
wire net_12375;
wire net_5201;
wire net_8063;
wire net_15127;
wire net_8353;
wire net_1156;
wire net_14127;
wire net_5150;
wire net_13641;
wire net_1966;
wire net_13049;
wire net_14299;
wire net_12188;
wire net_11718;
wire net_4571;
wire net_9212;
wire net_12713;
wire net_8176;
wire net_12873;
wire net_5977;
wire net_11493;
wire net_7709;
wire net_12672;
wire net_1659;
wire net_326;
wire net_2381;
wire net_589;
wire net_11012;
wire net_10286;
wire x1384;
wire net_15393;
wire net_9504;
wire net_1814;
wire net_5403;
wire net_11610;
wire net_5981;
wire net_10242;
wire net_6735;
wire net_6668;
wire net_3175;
wire net_14918;
wire net_10186;
wire net_10076;
wire x126;
wire net_7319;
wire net_2829;
wire net_10288;
wire net_8698;
wire net_724;
wire net_9826;
wire net_9123;
wire net_4815;
wire net_4099;
wire net_3142;
wire net_1219;
wire net_12826;
wire net_14410;
wire net_8058;
wire net_10886;
wire net_10871;
wire x5601;
wire net_13815;
wire net_2384;
wire net_3884;
wire net_7760;
wire net_8745;
wire net_3736;
wire net_2877;
wire net_5889;
wire net_2480;
wire net_9943;
wire net_12181;
wire net_9868;
wire net_9352;
wire net_874;
wire net_8334;
wire net_13706;
wire net_1632;
wire net_3796;
wire net_15264;
wire net_1661;
wire net_11399;
wire net_1236;
wire net_13627;
wire net_4277;
wire net_13771;
wire net_8987;
wire net_7907;
wire net_12107;
wire net_3674;
wire net_7555;
wire net_2700;
wire net_7996;
wire net_7868;
wire net_10307;
wire net_9548;
wire net_6841;
wire net_6273;
wire net_1488;
wire net_6187;
wire net_4966;
wire net_2812;
wire net_15522;
wire net_14973;
wire net_5244;
wire net_15406;
wire net_12721;
wire net_10178;
wire net_5691;
wire net_352;
wire net_11182;
wire net_9320;
wire net_12857;
wire net_3920;
wire net_436;
wire net_2837;
wire net_7963;
wire net_7181;
wire net_5641;
wire net_11157;
wire net_2824;
wire net_6342;
wire net_1777;
wire net_12983;
wire net_8263;
wire net_7373;
wire net_15706;
wire net_13647;
wire net_7903;
wire net_1641;
wire net_7511;
wire net_12325;
wire net_7246;
wire net_12153;
wire net_12134;
wire net_5556;
wire net_4919;
wire net_1702;
wire net_1103;
wire net_4403;
wire net_767;
wire net_7974;
wire net_6358;
wire net_1838;
wire net_4557;
wire net_11365;
wire net_10857;
wire net_131;
wire net_9754;
wire net_5488;
wire net_358;
wire net_1973;
wire net_8693;
wire net_8748;
wire net_7564;
wire net_4292;
wire net_2016;
wire net_14169;
wire net_2934;
wire net_7702;
wire net_10486;
wire net_11427;
wire net_3125;
wire net_1285;
wire net_10364;
wire net_5912;
wire net_3112;
wire net_15320;
wire net_13952;
wire net_1175;
wire net_13207;
wire net_13118;
wire net_12544;
wire net_10962;
wire net_9453;
wire net_6550;
wire net_9101;
wire net_9934;
wire net_5722;
wire net_13021;
wire net_9312;
wire net_9191;
wire net_2922;
wire net_9022;
wire net_10043;
wire net_1742;
wire net_13321;
wire net_11884;
wire net_7526;
wire net_7641;
wire net_14815;
wire net_11823;
wire net_468;
wire net_9308;
wire net_6890;
wire net_9372;
wire net_9257;
wire net_11654;
wire net_9738;
wire net_8011;
wire net_15368;
wire net_13734;
wire net_3370;
wire net_7025;
wire net_15573;
wire x732;
wire net_13040;
wire net_9497;
wire net_3947;
wire net_3441;
wire net_179;
wire net_9665;
wire net_4947;
wire net_4015;
wire net_3662;
wire net_10171;
wire net_12730;
wire net_8677;
wire net_14871;
wire net_14722;
wire net_8729;
wire net_3261;
wire net_9187;
wire net_13441;
wire net_6349;
wire net_2289;
wire net_10756;
wire net_7300;
wire net_11244;
wire net_6759;
wire net_5919;
wire net_3539;
wire net_2031;
wire net_1868;
wire net_1560;
wire net_13942;
wire net_4414;
wire net_12451;
wire net_4409;
wire net_10110;
wire net_7205;
wire net_12160;
wire net_10453;
wire net_6754;
wire net_13690;
wire net_12684;
wire net_3863;
wire net_10538;
wire net_9856;
wire net_8538;
wire net_9684;
wire net_8715;
wire net_14227;
wire net_13111;
wire net_5778;
wire net_7724;
wire net_6489;
wire net_3382;
wire net_4257;
wire net_1545;
wire net_13756;
wire net_4662;
wire net_4872;
wire net_8204;
wire net_990;
wire net_10798;
wire net_13838;
wire net_11728;
wire net_11485;
wire net_7423;
wire net_10428;
wire net_10473;
wire net_11763;
wire net_2332;
wire net_3774;
wire net_12491;
wire net_2715;
wire net_1803;
wire net_13803;
wire net_1941;
wire net_14915;
wire net_8031;
wire net_13074;
wire net_1134;
wire net_13968;
wire net_14276;
wire net_3899;
wire net_363;
wire net_1319;
wire net_8757;
wire net_776;
wire net_4550;
wire net_3080;
wire net_11075;
wire net_15358;
wire net_2508;
wire net_15091;
wire net_12118;
wire net_9624;
wire net_10353;
wire net_8451;
wire net_1650;
wire net_1582;
wire net_15174;
wire net_13574;
wire net_12696;
wire net_10717;
wire net_3149;
wire net_11253;
wire net_6454;
wire net_1675;
wire net_4016;
wire net_2247;
wire net_6028;
wire net_13747;
wire net_2333;
wire net_6544;
wire net_6464;
wire net_8115;
wire net_1368;
wire net_1248;
wire net_6525;
wire net_2291;
wire net_11108;
wire net_10531;
wire net_2238;
wire net_845;
wire net_15220;
wire net_10745;
wire x2477;
wire net_8003;
wire net_10973;
wire net_15558;
wire net_11096;
wire net_9081;
wire net_8414;
wire net_695;
wire net_12404;
wire net_7692;
wire net_2525;
wire net_1201;
wire net_14086;
wire x3849;
wire net_12073;
wire net_2671;
wire net_9701;
wire net_6787;
wire net_6569;
wire net_14331;
wire net_5106;
wire x1161;
wire net_8074;
wire net_13852;
wire net_12761;
wire net_859;
wire net_7259;
wire net_1167;
wire net_5896;
wire net_12788;
wire net_8636;
wire net_15169;
wire net_12610;
wire net_14605;
wire net_2198;
wire net_9043;
wire net_1044;
wire net_5250;
wire net_6435;
wire net_6661;
wire net_4322;
wire net_10948;
wire net_2940;
wire net_10617;
wire net_8672;
wire net_2043;
wire net_6775;
wire net_5583;
wire net_2095;
wire net_4681;
wire net_6955;
wire net_5231;
wire net_10662;
wire net_9726;
wire net_2314;
wire net_9905;
wire net_5454;
wire net_2613;
wire net_15311;
wire net_9995;
wire net_3605;
wire net_14336;
wire net_12174;
wire net_10865;
wire net_6635;
wire net_9010;
wire net_8849;
wire net_11055;
wire net_7250;
wire net_4114;
wire net_14220;
wire net_11479;
wire net_10330;
wire net_865;
wire net_13500;
wire net_9896;
wire net_231;
wire net_10197;
wire net_13326;
wire net_2621;
wire net_13832;
wire net_3024;
wire net_1223;
wire net_4691;
wire net_2750;
wire net_5816;
wire net_11961;
wire net_926;
wire net_4623;
wire net_12381;
wire net_7264;
wire net_7403;
wire net_4223;
wire net_6153;
wire net_14656;
wire net_11321;
wire net_8642;
wire net_2297;
wire net_13052;
wire net_9439;
wire net_7188;
wire net_3325;
wire net_12868;
wire net_10595;
wire net_9185;
wire net_6466;
wire net_6171;
wire net_2048;
wire net_582;
wire net_12485;
wire net_4481;
wire x461;
wire net_15331;
wire net_7419;
wire net_2341;
wire net_661;
wire net_3633;
wire net_3360;
wire net_13537;
wire net_15648;
wire net_11854;
wire net_7337;
wire net_7036;
wire x6157;
wire net_14705;
wire net_9086;
wire net_3561;
wire net_1543;
wire net_1295;
wire net_10006;
wire net_13692;
wire net_10993;
wire net_9429;
wire net_5661;
wire net_9460;
wire net_2071;
wire net_1923;
wire net_1275;
wire net_210;
wire net_13481;
wire net_11031;
wire net_916;
wire net_13463;
wire net_3395;
wire net_11641;
wire net_940;
wire net_4335;
wire net_851;
wire net_9924;
wire net_4411;
wire net_14865;
wire net_4857;
wire net_3719;
wire net_15681;
wire net_10572;
wire net_13247;
wire net_2426;
wire net_6061;
wire net_8311;
wire net_5350;
wire net_7405;
wire net_14329;
wire net_12330;
wire net_12237;
wire net_9627;
wire net_3310;
wire net_671;
wire net_8817;
wire net_8846;
wire net_13631;
wire x6599;
wire net_14425;
wire net_12849;
wire net_5335;
wire net_12431;
wire net_6830;
wire net_6965;
wire net_12438;
wire net_10133;
wire net_8734;
wire net_9485;
wire net_12978;
wire net_9054;
wire net_1454;
wire net_15473;
wire net_307;
wire net_6949;
wire net_3342;
wire net_13938;
wire net_3547;
wire net_14711;
wire net_14497;
wire net_1550;
wire net_3543;
wire net_11470;
wire net_10069;
wire net_9642;
wire net_15298;
wire net_5104;
wire net_15248;
wire net_14774;
wire net_6069;
wire net_233;
wire net_5138;
wire net_3459;
wire net_2656;
wire net_13411;
wire net_1268;
wire net_11127;
wire net_6326;
wire net_3922;
wire net_3212;
wire net_13783;
wire net_3780;
wire net_6530;
wire net_4051;
wire net_1115;
wire net_11465;
wire net_9632;
wire net_1764;
wire net_6641;
wire net_14067;
wire net_961;
wire net_9643;
wire net_3513;
wire net_9968;
wire net_13290;
wire net_4042;
wire net_2106;
wire net_9691;
wire net_3335;
wire net_14691;
wire net_5377;
wire net_3682;
wire net_6456;
wire net_5175;
wire net_14196;
wire net_11909;
wire net_4894;
wire net_12245;
wire net_5655;
wire net_9424;
wire net_7856;
wire net_9480;
wire net_3327;
wire net_5091;
wire net_13719;
wire net_2667;
wire net_13700;
wire net_3456;
wire net_12818;
wire net_7627;
wire net_13220;
wire net_12453;
wire net_12250;
wire net_5431;
wire net_9907;
wire net_4407;
wire net_13713;
wire net_8443;
wire net_1586;
wire net_14113;
wire net_5354;
wire net_480;
wire net_7662;
wire net_13284;
wire net_216;
wire net_4507;
wire net_10727;
wire net_4986;
wire net_2897;
wire net_5810;
wire net_2881;
wire net_836;
wire net_13817;
wire net_12630;
wire net_2161;
wire net_4602;
wire net_15556;
wire net_12075;
wire net_12057;
wire net_10671;
wire net_5635;
wire net_9495;
wire net_6568;
wire net_8408;
wire net_6059;
wire net_370;
wire net_8806;
wire net_8379;
wire net_11237;
wire net_13429;
wire net_12520;
wire net_9097;
wire net_6443;
wire net_5881;
wire net_1120;
wire net_2848;
wire net_7126;
wire net_1169;
wire net_973;
wire x472;
wire net_11832;
wire net_13416;
wire net_1139;
wire net_7057;
wire net_6998;
wire net_7013;
wire net_9337;
wire net_7394;
wire net_13677;
wire net_9238;
wire net_7389;
wire net_3902;
wire net_2206;
wire net_11206;
wire net_1392;
wire net_1574;
wire net_14575;
wire net_9008;
wire net_4842;
wire net_11576;
wire net_6121;
wire net_311;
wire net_2479;
wire net_10132;
wire net_8016;
wire net_154;
wire net_15453;
wire net_3699;
wire net_11119;
wire net_4469;
wire net_11452;
wire net_14598;
wire net_13847;
wire net_12527;
wire net_12056;
wire net_9986;
wire net_14946;
wire net_14075;
wire net_13210;
wire net_2520;
wire net_1478;
wire net_10166;
wire net_2179;
wire net_1696;
wire net_587;
wire net_1262;
wire net_10768;
wire net_9163;
wire net_10704;
wire net_4027;
wire net_14106;
wire net_6676;
wire net_8750;
wire net_4505;
wire net_4213;
wire net_2197;
wire x166;
wire net_10521;
wire net_5399;
wire net_10220;
wire net_4131;
wire net_12089;
wire net_10779;
wire net_9473;
wire net_7396;
wire net_14937;
wire net_14658;
wire net_11323;
wire net_2905;
wire net_1907;
wire net_10372;
wire net_200;
wire net_4435;
wire net_15420;
wire net_8612;
wire net_5220;
wire net_4164;
wire net_6312;
wire net_195;
wire net_5995;
wire net_14706;
wire net_10200;
wire net_1853;
wire net_9741;
wire net_10247;
wire net_10119;
wire net_10240;
wire net_2170;
wire net_6851;
wire net_10104;
wire net_15304;
wire net_15026;
wire net_8980;
wire net_2678;
wire net_11036;
wire net_8346;
wire net_13999;
wire net_9119;
wire x962;
wire net_9042;
wire net_8323;
wire net_7002;
wire net_10256;
wire net_9196;
wire net_8906;
wire net_3761;
wire net_6698;
wire net_13722;
wire net_11267;
wire x6028;
wire net_242;
wire net_7722;
wire net_7719;
wire net_7076;
wire net_10381;
wire net_15609;
wire net_7717;
wire net_6988;
wire net_9543;
wire net_6281;
wire net_6209;
wire net_2864;
wire net_8938;
wire net_1998;
wire net_11384;
wire net_9341;
wire net_13621;
wire net_11656;
wire net_8336;
wire net_13514;
wire net_2795;
wire net_1311;
wire net_13587;
wire net_5939;
wire net_5540;
wire net_13307;
wire net_11230;
wire net_7068;
wire net_1918;
wire net_12790;
wire net_10207;
wire net_15388;
wire net_10549;
wire net_5870;
wire net_11911;
wire net_7894;
wire net_5937;
wire net_8208;
wire net_3236;
wire net_5837;
wire net_12314;
wire net_3201;
wire net_11812;
wire net_11169;
wire net_9678;
wire net_3558;
wire x1298;
wire net_8147;
wire net_8096;
wire net_5613;
wire net_555;
wire net_9560;
wire net_8966;
wire net_13016;
wire net_7758;
wire net_7163;
wire net_1613;
wire net_15051;
wire net_8024;
wire net_6897;
wire net_12912;
wire net_11938;
wire net_790;
wire net_5300;
wire net_12359;
wire net_14665;
wire net_8926;
wire net_11466;
wire net_1417;
wire net_11520;
wire net_13423;
wire x3574;
wire x0;
wire net_11063;
wire net_2386;
wire net_2166;
wire net_5803;
wire net_5410;
wire net_14838;
wire net_3650;
wire net_8359;
wire net_2465;
wire net_15544;
wire net_5078;
wire net_11588;
wire net_5447;
wire net_12830;
wire net_12043;
wire net_15230;
wire net_14465;
wire net_10650;
wire net_8485;
wire net_10388;
wire net_7150;
wire net_13699;
wire net_7462;
wire net_9900;
wire net_6023;
wire net_13862;
wire net_898;
wire net_14855;
wire net_6136;
wire net_10416;
wire net_6537;
wire net_14873;
wire net_15548;
wire net_13023;
wire net_8364;
wire net_7229;
wire net_7045;
wire net_4416;
wire net_5015;
wire net_714;
wire net_8640;
wire net_2999;
wire net_1309;
wire net_9567;
wire net_683;
wire net_1771;
wire net_148;
wire net_1376;
wire net_12136;
wire net_5005;
wire net_4493;
wire net_13555;
wire net_13409;
wire net_8810;
wire net_6885;
wire net_7220;
wire net_6701;
wire net_1980;
wire net_13793;
wire net_9171;
wire net_10362;
wire net_9303;
wire net_7751;
wire net_7449;
wire net_1302;
wire net_244;
wire net_7341;
wire net_14504;
wire net_5547;
wire net_15411;
wire net_9361;
wire net_9149;
wire net_8687;
wire net_2395;
wire net_6012;
wire net_7353;
wire net_5616;
wire net_5347;
wire net_12117;
wire net_7113;
wire net_5439;
wire net_4002;
wire net_1989;
wire net_2855;
wire net_1795;
wire net_13310;
wire net_9247;
wire net_8588;
wire net_12186;
wire net_7740;
wire net_2403;
wire net_1539;
wire net_15173;
wire net_15582;
wire net_9626;
wire net_14147;
wire net_4261;
wire net_7913;
wire net_15238;
wire net_10123;
wire net_3490;
wire net_3035;
wire net_7646;
wire net_14417;
wire net_15191;
wire net_8550;
wire net_14761;
wire net_11483;
wire net_1548;
wire net_810;
wire net_92;
wire net_394;
wire net_13434;
wire net_3778;
wire net_1189;
wire net_6359;
wire net_12082;
wire net_11131;
wire net_7430;
wire net_409;
wire net_7183;
wire net_15366;
wire net_7437;
wire net_1469;
wire net_3470;
wire x1370;
wire net_11908;
wire net_15749;
wire net_11626;
wire net_4081;
wire net_15694;
wire net_13354;
wire net_2436;
wire net_8036;
wire net_11509;
wire net_15113;
wire net_10754;
wire net_3419;
wire net_10793;
wire net_1254;
wire net_10733;
wire net_14176;
wire net_11417;
wire net_11878;
wire net_621;
wire net_15616;
wire net_12793;
wire net_10018;
wire net_5153;
wire net_13316;
wire net_10375;
wire net_13171;
wire net_105;
wire net_10533;
wire net_11862;
wire net_7240;
wire net_12586;
wire net_7365;
wire net_7729;
wire net_5361;
wire net_15496;
wire net_8703;
wire net_5598;
wire net_12591;
wire net_11276;
wire net_3985;
wire net_14492;
wire net_14801;
wire net_12390;
wire net_9792;
wire net_9383;
wire net_9552;
wire net_10229;
wire net_9689;
wire net_12663;
wire net_9841;
wire net_4675;
wire net_8378;
wire net_327;
wire net_13032;
wire net_3877;
wire net_999;
wire net_8549;
wire net_353;
wire net_13799;
wire net_8052;
wire net_11730;
wire net_12322;
wire net_10888;
wire net_8838;
wire net_13924;
wire net_9584;
wire net_9752;
wire net_8552;
wire net_5730;
wire net_14209;
wire net_4994;
wire net_3588;
wire net_14140;
wire net_9151;
wire net_8770;
wire net_1480;
wire net_6927;
wire net_14759;
wire net_12628;
wire net_3046;
wire net_7700;
wire net_6019;
wire net_4952;
wire net_164;
wire net_377;
wire net_8836;
wire net_4702;
wire net_288;
wire net_7632;
wire net_15396;
wire net_2649;
wire net_3096;
wire net_14950;
wire net_8947;
wire net_1629;
wire net_1459;
wire net_12252;
wire net_7290;
wire net_5265;
wire net_14431;
wire net_11650;
wire net_11387;
wire net_3277;
wire net_805;
wire net_12032;
wire net_12093;
wire net_7749;
wire net_6740;
wire net_3741;
wire net_3590;
wire net_13257;
wire net_4470;
wire x747;
wire net_9168;
wire net_2151;
wire net_540;
wire net_8521;
wire net_2688;
wire net_2642;
wire net_14304;
wire net_6650;
wire net_1622;
wire net_891;
wire net_12899;
wire net_9388;
wire net_5224;
wire net_3065;
wire net_13392;
wire net_11664;
wire net_6299;
wire net_5149;
wire net_5821;
wire net_4167;
wire net_15011;
wire net_7796;
wire net_6746;
wire net_4711;
wire net_10236;
wire net_5868;
wire net_10358;
wire net_7815;
wire net_7453;
wire net_4802;
wire net_14793;
wire net_12998;
wire net_13420;
wire net_11744;
wire net_618;
wire net_12825;
wire net_2244;
wire net_9075;
wire net_3688;
wire net_5759;
wire net_12001;
wire net_11737;
wire net_7826;
wire net_12399;
wire net_8256;
wire net_783;
wire net_11955;
wire net_6970;
wire net_14907;
wire net_14255;
wire net_5945;
wire net_13686;
wire net_6148;
wire net_754;
wire net_10785;
wire net_9211;
wire net_11703;
wire net_6305;
wire net_9469;
wire net_2605;
wire net_7193;
wire net_921;
wire net_9875;
wire net_9113;
wire net_550;
wire net_7989;
wire net_11581;
wire net_4957;
wire net_10821;
wire net_14900;
wire net_12292;
wire net_5238;
wire net_3308;
wire net_12607;
wire net_10274;
wire net_9158;
wire net_5086;
wire net_3991;
wire net_2192;
wire net_1533;
wire net_10912;
wire net_14516;
wire net_8565;
wire net_7999;
wire net_461;
wire net_7681;
wire net_7778;
wire net_6879;
wire net_12962;
wire net_8524;
wire net_6657;
wire net_9284;
wire net_9138;
wire net_15525;
wire net_14185;
wire net_11158;
wire net_9884;
wire net_3502;
wire net_14014;
wire net_1512;
wire net_15370;
wire net_4827;
wire net_654;
wire net_14593;
wire net_330;
wire net_8047;
wire net_5025;
wire net_1330;
wire net_3506;
wire net_8082;
wire net_4275;
wire net_11011;
wire net_3015;
wire net_1785;
wire net_14538;
wire net_13507;
wire net_11077;
wire net_9116;
wire net_4771;
wire net_570;
wire net_444;
wire net_525;
wire net_10680;
wire net_3829;
wire net_3646;
wire net_1210;
wire net_1067;
wire net_15575;
wire net_9516;
wire net_6624;
wire net_5058;
wire net_6870;
wire net_14920;
wire net_5998;
wire net_9655;
wire net_7820;
wire net_5060;
wire net_14681;
wire net_12596;
wire net_6200;
wire net_5668;
wire net_10408;
wire net_6259;
wire net_15206;
wire net_4679;
wire net_985;
wire net_6719;
wire net_12190;
wire net_3933;
wire net_7061;
wire net_15494;
wire net_424;
wire net_11629;
wire net_6837;
wire net_1729;
wire net_12623;
wire net_3353;
wire net_9325;
wire x3071;
wire x5498;
wire net_4247;
wire net_4820;
wire net_5719;
wire net_13486;
wire net_10055;
wire net_7577;
wire net_14404;
wire net_3639;
wire net_8065;
wire net_12311;
wire net_12148;
wire net_11992;
wire net_3086;
wire net_4585;
wire net_11110;
wire net_9409;
wire net_2058;
wire net_12206;
wire net_9404;
wire net_3045;
wire net_1178;
wire net_9722;
wire net_5573;
wire net_4875;
wire x3133;
wire net_7098;
wire net_2018;
wire net_13100;
wire net_11731;
wire net_3825;
wire net_11142;
wire net_6218;
wire net_12380;
wire net_340;
wire net_6039;
wire net_2510;
wire net_15435;
wire net_9952;
wire net_2634;
wire net_434;
wire net_7881;
wire net_3808;
wire net_14631;
wire net_12941;
wire net_6915;
wire net_8434;
wire net_7024;
wire net_6936;
wire net_6243;
wire x5548;
wire net_14200;
wire net_7882;
wire net_1797;
wire net_6415;
wire net_9443;
wire net_14393;
wire net_11086;
wire net_9201;
wire net_14732;
wire net_4906;
wire net_4524;
wire net_6302;
wire net_8916;
wire net_339;
wire net_2279;
wire net_7686;
wire net_14048;
wire net_15633;
wire net_3447;
wire net_13105;
wire net_8401;
wire net_6174;
wire net_3468;
wire net_10443;
wire net_14588;
wire net_11775;
wire net_12753;
wire net_2710;
wire net_15722;
wire net_9267;
wire net_2660;
wire net_14486;
wire net_8624;
wire net_10083;
wire net_13893;
wire net_10826;
wire net_8087;
wire net_5389;
wire net_8497;
wire net_3671;
wire net_102;
wire net_8236;
wire net_8651;
wire net_10295;
wire net_3691;
wire net_7801;
wire net_3217;
wire net_6362;
wire net_4387;
wire net_1291;
wire net_1865;
wire net_13896;
wire net_678;
wire net_6076;
wire net_5168;
wire net_5329;
wire net_14541;
wire net_11631;
wire net_8979;
wire net_10985;
wire net_928;
wire net_15251;
wire net_10490;
wire net_8460;
wire net_5459;
wire net_13363;
wire net_2578;
wire net_208;
wire net_9225;
wire net_7878;
wire net_8658;
wire net_8215;
wire net_10462;
wire net_2744;
wire net_2377;
wire net_1433;
wire net_415;
wire net_116;
wire net_3251;
wire net_2786;
wire net_11672;
wire net_347;
wire net_13745;
wire net_15503;
wire net_14784;
wire net_13526;
wire net_11059;
wire net_3794;
wire net_12664;
wire net_14786;
wire net_8606;
wire net_7306;
wire net_5440;
wire net_9425;
wire net_1335;
wire net_5928;
wire net_2574;
wire net_15716;
wire net_14235;
wire net_15519;
wire net_3531;
wire net_12210;
wire net_5477;
wire net_3747;
wire net_2212;
wire net_5453;
wire net_11535;
wire net_7730;
wire net_12212;
wire net_5732;
wire net_8593;
wire net_3571;
wire net_4642;
wire net_610;
wire net_1844;
wire net_8130;
wire net_11512;
wire net_7870;
wire net_389;
wire net_902;
wire net_15187;
wire net_13981;
wire net_2344;
wire net_11287;
wire net_10588;
wire net_1323;
wire net_14130;
wire net_1506;
wire net_10470;
wire net_13386;
wire net_13237;
wire net_6496;
wire net_13193;
wire net_736;
wire net_8771;
wire net_539;
wire net_13068;
wire net_692;
wire net_5462;
wire net_5282;
wire net_4568;
wire net_6498;
wire net_8372;
wire net_10807;
wire net_15737;
wire net_6262;
wire net_4377;
wire net_15130;
wire net_14261;
wire net_7704;
wire net_13125;
wire net_15379;
wire net_15104;
wire net_10905;
wire net_10311;
wire net_12517;
wire net_1400;
wire net_14092;
wire net_885;
wire net_10034;
wire net_9202;
wire net_7249;
wire net_11698;
wire net_15152;
wire net_14320;
wire net_9918;
wire net_5717;
wire net_10770;
wire net_869;
wire net_12144;
wire net_6822;
wire net_3714;
wire net_8308;
wire net_11280;
wire net_4077;
wire net_11607;
wire net_2441;
wire net_6594;
wire net_3517;
wire net_496;
wire net_761;
wire net_11396;
wire net_6799;
wire net_5828;
wire net_4749;
wire net_1554;
wire net_7101;
wire net_8775;
wire net_13774;
wire net_12092;
wire net_2459;
wire net_15512;
wire net_10638;
wire net_4370;
wire net_10394;
wire net_4979;
wire net_14613;
wire net_12578;
wire net_2249;
wire net_14434;
wire net_5422;
wire net_6629;
wire net_5686;
wire net_6704;
wire net_15129;
wire net_739;
wire net_12395;
wire net_15329;
wire net_8760;
wire net_6508;
wire net_2548;
wire net_2075;
wire net_826;
wire net_15069;
wire net_1738;
wire net_10384;
wire net_10504;
wire net_14887;
wire net_3359;
wire net_5848;
wire x2648;
wire net_10085;
wire net_12296;
wire net_11644;
wire net_9069;
wire net_6716;
wire net_7548;
wire net_2624;
wire net_12889;
wire net_14866;
wire net_11761;
wire net_343;
wire net_6165;
wire net_4795;
wire net_511;
wire net_9263;
wire net_12759;
wire net_7313;
wire net_3967;
wire net_9672;
wire net_8456;
wire net_5236;
wire net_4424;
wire net_7541;
wire net_9615;
wire net_2654;
wire net_7451;
wire net_2487;
wire net_11791;
wire net_7803;
wire net_2911;
wire net_1819;
wire net_15509;
wire net_8258;
wire net_12821;
wire net_8227;
wire net_12763;
wire net_13132;
wire net_15674;
wire net_2975;
wire net_4625;
wire net_7236;
wire net_5257;
wire net_8220;
wire net_2779;
wire net_14187;
wire net_11552;
wire net_6392;
wire net_13181;
wire net_11379;
wire net_9031;
wire net_15158;
wire net_9346;
wire net_13661;
wire net_11352;
wire net_8169;
wire net_1490;
wire net_11083;
wire net_9274;
wire net_4282;
wire net_15216;
wire net_989;
wire net_11806;
wire x1282;
wire net_12774;
wire net_8446;
wire net_15565;
wire net_14765;
wire net_14342;
wire net_5742;
wire net_458;
wire net_4356;
wire net_11748;
wire net_685;
wire net_8466;
wire net_7442;
wire net_8322;
wire net_14471;
wire net_10998;
wire net_9030;
wire net_10957;
wire net_12349;
wire net_14183;
wire net_13333;
wire net_11843;
wire net_4052;
wire net_8513;
wire net_4616;
wire net_8681;
wire net_13096;
wire net_11408;
wire net_4786;
wire net_8616;
wire net_7872;
wire net_5893;
wire net_10542;
wire x5077;
wire net_13469;
wire net_10891;
wire net_10652;
wire net_7160;
wire net_12876;
wire net_4686;
wire net_3410;
wire net_2111;
wire net_1946;
wire net_2733;
wire net_14954;
wire net_8162;
wire net_5525;
wire net_12496;
wire net_14280;
wire net_6764;
wire net_14894;
wire net_13252;
wire net_5610;
wire net_14278;
wire net_6769;
wire net_3612;
wire net_11634;
wire net_1605;
wire net_12795;
wire net_13045;
wire net_2535;
wire net_13165;
wire net_3191;
wire net_5118;
wire net_15106;
wire net_14396;
wire net_13822;
wire net_747;
wire net_15597;
wire net_10355;
wire net_2305;
wire net_1653;
wire net_12865;
wire net_14125;
wire net_5842;
wire net_12125;
wire net_9817;
wire net_7377;
wire net_2983;
wire net_12916;
wire net_14617;
wire net_10024;
wire net_2258;
wire net_198;
wire net_1647;
wire net_12460;
wire net_11168;
wire net_12510;
wire net_14327;
wire net_10058;
wire net_7509;
wire net_4756;
wire net_15293;
wire net_13280;
wire net_6500;
wire net_5196;
wire net_2367;
wire net_14697;
wire net_4573;
wire net_4127;
wire net_2892;
wire net_13263;
wire net_15646;
wire net_2810;
wire net_13546;
wire net_13077;
wire net_1053;
wire net_4444;
wire net_11292;
wire net_1004;
wire net_848;
wire net_4921;
wire net_11716;
wire net_11359;
wire net_9550;
wire net_12022;
wire net_1080;
wire net_10641;
wire net_3232;
wire net_1890;
wire net_13356;
wire net_13648;
wire net_4498;
wire net_11293;
wire net_3228;
wire net_2282;
wire net_10029;
wire net_4501;
wire net_2357;
wire net_13319;
wire net_12449;
wire net_11114;
wire net_1546;
wire net_11772;
wire net_11367;
wire net_8542;
wire net_5492;
wire net_15695;
wire net_12383;
wire net_6042;
wire net_13654;
wire net_11372;
wire net_10199;
wire net_1046;
wire net_15728;
wire net_6536;
wire net_11502;
wire net_7417;
wire net_4363;
wire net_606;
wire net_10332;
wire net_4960;
wire net_3906;
wire net_623;
wire net_12503;
wire net_663;
wire net_1213;
wire net_1891;
wire net_2265;
wire net_8118;
wire net_10163;
wire net_5180;
wire net_3998;
wire net_579;
wire net_9490;
wire net_8597;
wire net_5795;
wire net_12812;
wire net_769;
wire net_1780;
wire net_2062;
wire net_13668;
wire net_13666;
wire net_9828;
wire x1134;
wire net_10844;
wire net_6418;
wire net_1025;
wire net_3758;
wire net_7296;
wire net_4834;
wire net_9317;
wire net_8061;
wire net_4067;
wire net_4717;
wire net_15062;
wire net_13157;
wire net_10403;
wire net_7502;
wire net_1518;
wire net_4618;
wire net_1089;
wire net_12169;
wire net_1194;
wire net_1437;
wire net_11998;
wire net_5517;
wire net_6770;
wire net_11923;
wire net_7587;
wire net_1664;
wire net_13651;
wire net_4528;
wire net_15718;
wire net_6233;
wire net_5625;
wire net_10326;
wire net_705;
wire net_4141;
wire net_2948;
wire net_10523;
wire net_14094;
wire net_12535;
wire net_10669;
wire net_1036;
wire net_6052;
wire net_5608;
wire net_11966;
wire net_7497;
wire net_5146;
wire net_4537;
wire net_8701;
wire net_1196;
wire net_6331;
wire net_3973;
wire net_5326;
wire net_12921;
wire net_4394;
wire net_9077;
wire net_6762;
wire net_15421;
wire net_5531;
wire net_5953;
wire net_12442;
wire net_11047;
wire net_12702;
wire net_9433;
wire net_6085;
wire net_10816;
wire net_6598;
wire net_14124;
wire net_13248;
wire net_5701;
wire net_11786;
wire net_3626;
wire net_12095;
wire net_5779;
wire net_14798;
wire net_3136;
wire net_12553;
wire net_6417;
wire net_4726;
wire net_4090;
wire net_15475;
wire net_14377;
wire net_13086;
wire net_9588;
wire net_14572;
wire net_6149;
wire net_10809;
wire net_9178;
wire net_5344;
wire net_3834;
wire net_7492;
wire net_12468;
wire net_5364;
wire net_10300;
wire net_13471;
wire net_8743;
wire net_3152;
wire net_6388;
wire x2098;
wire net_14311;
wire net_13478;
wire net_3648;
wire net_740;
wire net_1722;
wire net_4072;
wire net_6395;
wire net_2008;
wire net_11633;
wire net_11090;
wire net_5825;
wire net_3183;
wire net_2808;
wire net_3908;
wire net_8265;
wire net_4837;
wire net_730;
wire net_9055;
wire net_4150;
wire net_14008;
wire net_8049;
wire net_7094;
wire net_5405;
wire net_11931;
wire net_6575;
wire net_2105;
wire net_13918;
wire net_7226;
wire net_6432;
wire net_4707;
wire net_1127;
wire net_6381;
wire net_9458;
wire net_11243;
wire net_15667;
wire net_12771;
wire net_6420;
wire net_957;
wire net_1287;
wire net_13831;
wire net_10625;
wire net_7465;
wire net_14040;
wire net_9297;
wire net_2726;
wire net_15732;
wire net_4143;
wire net_12900;
wire net_8679;
wire net_7285;
wire net_1340;
wire net_5140;
wire net_7277;
wire net_3123;
wire net_2955;
wire net_7165;
wire net_9599;
wire net_12363;
wire net_771;
wire net_2844;
wire net_2301;
wire net_12415;
wire net_2978;
wire net_9977;
wire net_15033;
wire net_5538;
wire net_5185;
wire net_13139;
wire net_9941;
wire net_6804;
wire net_4852;
wire net_10341;
wire net_14361;
wire net_3950;
wire net_10435;
wire net_4437;
wire net_4028;
wire net_2860;
wire net_432;
wire net_6025;
wire net_4927;
wire net_1062;
wire net_6329;
wire net_14395;
wire net_10627;
wire net_4936;
wire net_3293;
wire net_1142;
wire net_14556;
wire net_4120;
wire net_9246;
wire net_7733;
wire net_3159;
wire net_14987;
wire net_5644;
wire net_6050;
wire net_14600;
wire net_2240;
wire net_2416;
wire net_13214;
wire net_12882;
wire net_6404;
wire net_5188;
wire net_4590;
wire net_8727;
wire net_14354;
wire net_6185;
wire net_6116;
wire net_9713;
wire net_1411;
wire net_12549;
wire net_505;
wire net_5383;
wire net_4088;
wire net_10471;
wire net_3723;
wire net_10540;
wire net_7487;
wire net_13520;
wire net_14724;
wire net_10493;
wire net_10426;
wire net_7152;
wire net_6527;
wire net_4013;
wire net_992;
wire net_11517;
wire net_7485;
wire net_9781;
wire net_6727;
wire x6102;
wire net_782;
wire net_2144;
wire net_2236;
wire net_10527;
wire net_13576;
wire net_11106;
wire net_11057;
wire net_3443;
wire net_6291;
wire net_4186;
wire net_13328;
wire net_4738;
wire net_3314;
wire net_7422;
wire net_3945;
wire net_2971;
wire net_5776;
wire net_8824;
wire net_13322;
wire net_11529;
wire net_10339;
wire net_14622;
wire net_8072;
wire net_8244;
wire net_2836;
wire net_1505;
wire net_10615;
wire net_5689;
wire net_7429;
wire net_1805;
wire net_4667;
wire net_13836;
wire net_11536;
wire net_8279;
wire net_3952;
wire net_3669;
wire net_13448;
wire net_10660;
wire net_1861;
wire net_3635;
wire net_9999;
wire net_4388;
wire net_11852;
wire net_13559;
wire net_5672;
wire net_221;
wire net_1594;
wire net_7120;
wire net_1110;
wire net_15356;
wire net_442;
wire net_14999;
wire net_542;
wire net_14218;
wire net_13026;
wire net_13789;
wire net_12483;
wire x1503;
wire net_6487;
wire net_7202;
wire net_4562;
wire net_9437;
wire net_3087;
wire net_2376;
wire net_14627;
wire net_6562;
wire net_1520;
wire net_6713;
wire net_13900;
wire net_1821;
wire net_8579;
wire net_9638;
wire net_11675;
wire net_7480;
wire net_3865;
wire net_1588;
wire net_15287;
wire net_9029;
wire net_4037;
wire net_8005;
wire net_3937;
wire net_1495;
wire net_2992;
wire net_12974;
wire net_3664;
wire net_5124;
wire net_3233;
wire net_14521;
wire net_9731;
wire net_3522;
wire net_7178;
wire net_10937;
wire net_668;
wire net_7601;
wire net_11814;
wire net_9649;
wire net_3079;
wire net_1584;
wire net_14203;
wire net_13539;
wire net_12612;
wire net_2330;
wire net_8040;
wire net_5814;
wire net_7890;
wire net_12707;
wire net_3397;
wire net_1070;
wire net_9777;
wire net_8878;
wire net_1225;
wire net_812;
wire net_5898;
wire net_6785;
wire net_7814;
wire net_4391;
wire net_11473;
wire net_14993;
wire net_13805;
wire net_9045;
wire net_6314;
wire net_12659;
wire net_6875;
wire net_6972;
wire net_2857;
wire net_1107;
wire net_8674;
wire net_2767;
wire net_9594;
wire net_6120;
wire net_11491;
wire net_11053;
wire net_15621;
wire net_3384;
wire net_12652;
wire net_6604;
wire net_1203;
wire net_13347;
wire net_825;
wire net_309;
wire net_15055;
wire net_1366;
wire net_13054;
wire net_2615;
wire net_14978;
wire net_9011;
wire net_12402;
wire net_12176;
wire net_10867;
wire net_10715;
wire net_14268;
wire net_5321;
wire net_11434;
wire net_9290;
wire net_7367;
wire net_12789;
wire net_8158;
wire net_1151;
wire net_5240;
wire net_5318;
wire net_9993;
wire net_11138;
wire net_8291;
wire net_15046;
wire net_5884;
wire net_3213;
wire net_2818;
wire net_863;
wire net_7131;
wire net_7690;
wire net_6468;
wire net_3164;
wire net_4173;
wire net_580;
wire net_14058;
wire net_13150;
wire net_9805;
wire net_2136;
wire net_904;
wire net_2339;
wire net_8884;
wire net_7699;
wire net_15580;
wire net_12850;
wire net_14226;
wire net_4157;
wire net_13552;
wire net_1879;
wire net_14821;
wire net_6777;
wire net_12286;
wire net_6663;
wire net_12122;
wire net_13224;
wire net_8202;
wire net_6633;
wire net_8126;
wire net_4941;
wire net_4221;
wire net_6092;
wire net_6732;
wire net_6559;
wire net_15553;
wire net_12524;
wire net_11360;
wire net_9183;
wire net_15688;
wire net_4845;
wire net_1160;
wire net_12683;
wire net_159;
wire net_11147;
wire net_9379;
wire net_3268;
wire net_11022;
wire net_5604;
wire net_11612;
wire net_5863;
wire net_8351;
wire net_11615;
wire net_9523;
wire net_10181;
wire net_4887;
wire x936;
wire net_9354;
wire net_13116;
wire net_14834;
wire net_2875;
wire net_763;
wire net_13704;
wire net_12952;
wire net_14088;
wire net_10213;
wire net_7762;
wire net_14495;
wire net_5639;
wire net_1740;
wire net_324;
wire net_6848;
wire net_11724;
wire net_10284;
wire net_10074;
wire net_13397;
wire net_9455;
wire net_5480;
wire net_14675;
wire net_10309;
wire net_7257;
wire net_872;
wire net_13047;
wire net_9706;
wire net_14248;
wire net_14103;
wire net_9125;
wire net_12647;
wire net_10964;
wire net_10502;
wire net_5046;
wire net_3066;
wire net_8251;
wire net_6270;
wire net_3880;
wire net_15385;
wire net_6275;
wire net_5581;
wire net_4333;
wire net_4181;
wire net_11285;
wire net_14776;
wire net_376;
wire net_5558;
wire net_7575;
wire net_2133;
wire net_13643;
wire net_4817;
wire net_4880;
wire net_13374;
wire net_2515;
wire net_1812;
wire net_8174;
wire net_3173;
wire net_12584;
wire net_8038;
wire net_4825;
wire net_10850;
wire net_3738;
wire net_8696;
wire net_7994;
wire net_15529;
wire net_4138;
wire net_5298;
wire net_5119;
wire net_3203;
wire net_422;
wire net_4290;
wire net_14739;
wire net_1345;
wire net_12811;
wire net_1450;
wire net_561;
wire net_12694;
wire net_11881;
wire net_4899;
wire net_12670;
wire net_7515;
wire net_2659;
wire net_2589;
wire net_12739;
wire net_591;
wire net_1700;
wire net_12985;
wire net_5955;
wire net_8501;
wire net_4299;
wire net_2290;
wire net_12741;
wire net_10188;
wire net_7557;
wire net_2851;
wire net_178;
wire net_11751;
wire net_8427;
wire net_15266;
wire net_14640;
wire net_9074;
wire net_2843;
wire net_14081;
wire net_14019;
wire net_6780;
wire net_7961;
wire net_15322;
wire net_10191;
wire net_3772;
wire net_7901;
wire net_3807;
wire net_4868;
wire net_10480;
wire net_2698;
wire net_809;
wire net_13995;
wire net_8393;
wire net_6552;
wire net_8453;
wire net_3450;
wire net_635;
wire net_4279;
wire net_266;
wire net_1235;
wire net_14412;
wire net_2691;
wire net_14813;
wire net_3528;
wire net_8559;
wire net_8610;
wire net_12600;
wire net_8956;
wire net_350;
wire net_6622;
wire net_4270;
wire net_15520;
wire net_8332;
wire net_6007;
wire net_13205;
wire net_13178;
wire net_10176;
wire net_7606;
wire net_6549;
wire net_13275;
wire net_6542;
wire net_13091;
wire net_3460;
wire net_12859;
wire net_3117;
wire net_14245;
wire net_11816;
wire net_3482;
wire net_6648;
wire net_3198;
wire net_8366;
wire net_5720;
wire net_1626;
wire net_2822;
wire net_7317;
wire net_8413;
wire net_1258;
wire net_7375;
wire net_15712;
wire net_12041;
wire net_3369;
wire net_9866;
wire net_9020;
wire net_1101;
wire net_994;
wire net_12828;
wire net_12268;
wire net_10231;
wire net_318;
wire net_6685;
wire net_3927;
wire net_11837;
wire net_10859;
wire net_1971;
wire net_8931;
wire net_4166;
wire net_2409;
wire net_4608;
wire net_3192;
wire net_1900;
wire net_1779;
wire net_2647;
wire net_5218;
wire net_15122;
wire net_3340;
wire net_8492;
wire net_4545;
wire net_3844;
wire net_1849;
wire net_7972;
wire net_10045;
wire net_228;
wire net_5486;
wire net_11886;
wire net_4737;
wire net_2640;
wire net_13011;
wire net_966;
wire net_7083;
wire net_13516;
wire net_4698;
wire net_3372;
wire net_14994;
wire net_14637;
wire net_11122;
wire net_6049;
wire net_2201;
wire net_1108;
wire net_2827;
wire net_2025;
wire net_8583;
wire net_7905;
wire net_2936;
wire net_5643;
wire net_9756;
wire net_9936;
wire net_1878;
wire net_13736;
wire net_5728;
wire net_13070;
wire net_9255;
wire net_11446;
wire net_8013;
wire net_3890;
wire net_5975;
wire net_133;
wire net_12425;
wire net_10702;
wire net_10366;
wire net_7528;
wire net_14297;
wire net_4025;
wire net_11414;
wire net_12444;
wire net_11265;
wire net_10920;
wire net_15024;
wire net_9194;
wire net_15459;
wire net_7078;
wire net_12529;
wire net_10579;
wire net_7008;
wire net_11957;
wire net_7997;
wire net_4522;
wire net_3882;
wire net_557;
wire net_3043;
wire net_11925;
wire x39;
wire net_15288;
wire net_14836;
wire net_8908;
wire net_7860;
wire net_8689;
wire net_6611;
wire net_3652;
wire net_6829;
wire net_2669;
wire net_13891;
wire net_11386;
wire net_4083;
wire net_12316;
wire net_1991;
wire net_1611;
wire net_1173;
wire net_14046;
wire net_1431;
wire net_1754;
wire net_2328;
wire net_7715;
wire net_11401;
wire net_8080;
wire net_1714;
wire net_5571;
wire net_15302;
wire net_13014;
wire net_11970;
wire net_10205;
wire net_5805;
wire net_8868;
wire net_240;
wire net_12792;
wire net_15115;
wire net_7254;
wire net_13623;
wire net_7684;
wire x268;
wire net_295;
wire net_8411;
wire net_12991;
wire net_10743;
wire net_14467;
wire net_13605;
wire net_13565;
wire net_13425;
wire net_9604;
wire net_9241;
wire net_6887;
wire net_9838;
wire net_15427;
wire net_15546;
wire net_4462;
wire net_5935;
wire net_11038;
wire net_13490;
wire net_1394;
wire net_7753;
wire net_2963;
wire net_5546;
wire net_5412;
wire net_15236;
wire net_14879;
wire net_12115;
wire net_7720;
wire net_6134;
wire net_9395;
wire net_1281;
wire net_2463;
wire net_11239;
wire net_9291;
wire net_12619;
wire net_6691;
wire net_8210;
wire net_12967;
wire net_278;
wire net_6864;
wire net_11258;
wire net_8995;
wire net_8367;
wire net_4058;
wire net_9063;
wire net_8432;
wire net_4874;
wire net_3509;
wire net_1162;
wire net_10090;
wire net_13856;
wire net_13309;
wire net_2443;
wire net_10736;
wire net_2472;
wire net_1307;
wire net_13589;
wire net_4514;
wire net_2790;
wire net_2742;
wire net_13120;
wire net_10738;
wire net_5007;
wire net_15386;
wire net_10318;
wire net_6940;
wire net_13795;
wire net_10434;
wire net_5591;
wire net_4810;
wire net_11902;
wire net_8360;
wire net_10269;
wire net_6521;
wire net_15413;
wire net_10561;
wire net_4418;
wire net_3320;
wire net_5221;
wire net_3657;
wire net_5550;
wire net_5385;
wire net_14145;
wire net_6099;
wire net_1353;
wire net_14683;
wire net_9786;
wire net_11652;
wire net_15165;
wire net_12679;
wire net_7630;
wire net_5303;
wire net_3581;
wire net_14961;
wire net_13854;
wire net_13712;
wire net_4049;
wire net_3776;
wire net_1300;
wire net_14322;
wire net_1252;
wire net_12131;
wire net_14419;
wire net_9173;
wire net_7739;
wire net_9095;
wire net_7784;
wire net_13432;
wire net_14026;
wire net_10941;
wire net_547;
wire net_1098;
wire net_10731;
wire net_507;
wire net_10097;
wire net_10049;
wire net_8981;
wire net_1902;
wire net_6683;
wire net_238;
wire net_3074;
wire net_7111;
wire net_8973;
wire net_5475;
wire net_11354;
wire net_7055;
wire net_7896;
wire net_2438;
wire net_2600;
wire net_1911;
wire net_6906;
wire net_5734;
wire net_3563;
wire net_12224;
wire net_8726;
wire net_6585;
wire net_649;
wire net_9565;
wire net_13597;
wire net_11936;
wire net_4491;
wire net_11543;
wire net_1374;
wire net_13887;
wire net_8282;
wire net_7538;
wire net_4843;
wire net_8959;
wire net_1962;
wire net_291;
wire net_9502;
wire net_7351;
wire net_1964;
wire net_2494;
wire net_857;
wire net_867;
wire net_15747;
wire net_5964;
wire net_11217;
wire net_15618;
wire net_6819;
wire net_396;
wire net_14811;
wire net_12274;
wire net_3700;
wire net_13349;
wire net_107;
wire net_14845;
wire net_10602;
wire net_8851;
wire net_10535;
wire net_530;
wire net_15155;
wire net_9140;
wire net_1541;
wire net_14966;
wire net_11839;
wire net_10529;
wire net_14216;
wire net_9748;
wire net_15683;
wire net_5177;
wire net_271;
wire net_3329;
wire net_10067;
wire net_10004;
wire net_6111;
wire net_673;
wire net_7022;
wire net_4268;
wire net_12247;
wire net_12208;
wire net_7029;
wire net_14693;
wire net_3611;
wire net_2064;
wire net_9966;
wire net_6256;
wire net_2797;
wire net_15274;
wire net_3846;
wire net_12261;
wire net_5333;
wire net_1925;
wire net_9790;
wire net_3549;
wire net_1445;
wire net_10227;
wire net_8581;
wire net_1909;
wire net_6729;
wire net_13807;
wire net_9922;
wire net_10126;
wire net_7639;
wire net_1410;
wire net_11454;
wire net_11583;
wire net_365;
wire net_13412;
wire net_5379;
wire net_13340;
wire net_3913;
wire net_11643;
wire net_9988;
wire net_3344;
wire net_12060;
wire net_8374;
wire net_3787;
wire net_10729;
wire net_4413;
wire net_1810;
wire net_10776;
wire net_1118;
wire net_13849;
wire net_8719;
wire net_4313;
wire net_11000;
wire net_12235;
wire net_6858;
wire net_372;
wire net_9882;
wire net_8313;
wire net_7086;
wire net_2990;
wire net_9339;
wire net_6324;
wire net_7128;
wire net_7915;
wire net_13723;
wire net_11749;
wire net_13730;
wire net_4892;
wire net_803;
wire net_10884;
wire net_3595;
wire net_13787;
wire net_10383;
wire net_8923;
wire net_2788;
wire net_14713;
wire net_10142;
wire net_6899;
wire net_14111;
wire net_14490;
wire net_7764;
wire net_6375;
wire net_1476;
wire net_15346;
wire net_3489;
wire net_1293;
wire net_14939;
wire net_11098;
wire net_11184;
wire net_13581;
wire net_2883;
wire net_8665;
wire net_563;
wire net_7854;
wire net_13979;
wire net_1147;
wire net_11742;
wire net_13388;
wire net_15242;
wire net_2681;
wire net_15193;
wire net_8815;
wire x2027;
wire x4209;
wire net_13452;
wire net_12159;
wire net_9629;
wire net_2158;
wire net_5136;
wire net_4855;
wire net_14668;
wire net_4366;
wire net_10234;
wire net_13936;
wire net_10175;
wire net_12254;
wire net_5009;
wire net_1266;
wire net_3684;
wire net_14677;
wire net_1452;
wire net_8418;
wire net_2773;
wire net_2428;
wire net_909;
wire net_4529;
wire net_10695;
wire net_4898;
wire net_152;
wire net_8652;
wire net_11575;
wire net_10814;
wire net_3105;
wire net_2895;
wire net_15488;
wire net_13299;
wire net_2138;
wire net_13418;
wire net_8238;
wire net_258;
wire net_12957;
wire net_11192;
wire net_2477;
wire net_10761;
wire net_12935;
wire x381;
wire net_12054;
wire net_9927;
wire net_5653;
wire net_13983;
wire net_13819;
wire net_7664;
wire net_5083;
wire net_2446;
wire net_7171;
wire net_11999;
wire net_15644;
wire net_4188;
wire net_15451;
wire net_7605;
wire net_585;
wire net_7611;
wire net_7809;
wire net_6146;
wire net_4040;
wire net_14823;
wire x6577;
wire net_11913;
wire net_11347;
wire net_12766;
wire net_5433;
wire net_12061;
wire net_10593;
wire net_3759;
wire net_14514;
wire net_3511;
wire net_12839;
wire net_374;
wire net_14069;
wire net_10293;
wire net_8755;
wire net_1987;
wire net_12816;
wire net_12632;
wire net_788;
wire net_12910;
wire net_9090;
wire net_214;
wire net_7011;
wire net_8113;
wire net_3602;
wire net_249;
wire net_13155;
wire net_13028;
wire net_9963;
wire net_8144;
wire net_3578;
wire net_12455;
wire net_5283;
wire net_13903;
wire net_8804;
wire net_9013;
wire net_8871;
wire net_6310;
wire net_6196;
wire net_13488;
wire net_10766;
wire net_4009;
wire net_7648;
wire net_5097;
wire net_13880;
wire net_8508;
wire net_7329;
wire net_5993;
wire net_4259;
wire net_2565;
wire net_8018;
wire net_2632;
wire net_2547;
wire net_8634;
wire net_5076;
wire net_13229;
wire net_9084;
wire net_6783;
wire net_5908;
wire net_2118;
wire net_463;
wire net_15440;
wire net_2295;
wire net_5831;
wire net_15281;
wire net_5628;
wire net_9487;
wire net_1817;
wire net_197;
wire net_2560;
wire net_11009;
wire net_9348;
wire net_1381;
wire net_9331;
wire net_6445;
wire net_5017;
wire net_3709;
wire net_202;
wire net_13596;
wire net_3312;
wire net_13085;
wire net_7325;
wire net_1756;
wire net_12803;
wire net_7588;
wire net_11468;
wire net_2208;
wire net_6475;
wire net_5352;
wire net_2595;
wire net_1383;
wire net_7302;
wire net_2751;
wire net_918;
wire net_11204;
wire net_7727;
wire net_9663;
wire net_9165;
wire net_5397;
wire net_9204;
wire net_4446;
wire net_14160;
wire net_10484;
wire net_6269;
wire net_6176;
wire net_5901;
wire net_14170;
wire net_13672;
wire net_13610;
wire net_11116;
wire net_13497;
wire net_1683;
wire net_12515;
wire x1329;
wire net_978;
wire net_15510;
wire net_9356;
wire net_1313;
wire net_10780;
wire net_1129;
wire net_11345;
wire net_7618;
wire net_3331;
wire net_1056;
wire net_14689;
wire net_4908;
wire net_14561;
wire net_11994;
wire net_13286;
wire net_10896;
wire net_5712;
wire net_14446;
wire net_10877;
wire net_8383;
wire net_4781;
wire net_2044;
wire net_9954;
wire net_7402;
wire net_6360;
wire net_2181;
wire net_8626;
wire net_6913;
wire net_14782;
wire net_1789;
wire net_14035;
wire x1248;
wire net_13142;
wire net_13940;
wire net_8406;
wire net_7379;
wire net_4530;
wire net_838;
wire net_3219;
wire net_10441;
wire net_6123;
wire net_7520;
wire net_14316;
wire net_11151;
wire net_14202;
wire net_4587;
wire net_11750;
wire net_5872;
wire net_7107;
wire net_4980;
wire net_2576;
wire net_15341;
wire net_11270;
wire net_3827;
wire net_2352;
wire net_1038;
wire net_8405;
wire net_12072;
wire net_6931;
wire net_4241;
wire net_9920;
wire net_8168;
wire net_5308;
wire net_5710;
wire net_5369;
wire net_3763;
wire net_15445;
wire net_3515;
wire x2165;
wire net_12747;
wire net_5033;
wire net_8085;
wire net_6333;
wire net_9720;
wire net_11338;
wire net_14662;
wire net_9223;
wire net_7697;
wire net_3398;
wire net_2277;
wire net_342;
wire net_13400;
wire net_6078;
wire net_975;
wire net_5421;
wire net_612;
wire net_892;
wire net_15538;
wire net_8098;
wire net_12871;
wire net_4650;
wire net_4198;
wire net_13061;
wire net_10423;
wire net_15735;
wire net_5434;
wire net_11144;
wire net_6160;
wire net_10848;
wire net_14488;
wire net_5874;
wire net_2006;
wire net_13570;
wire net_12639;
wire net_8344;
wire net_10060;
wire net_6511;
wire net_1331;
wire net_1537;
wire net_13051;
wire net_11105;
wire x5850;
wire net_12307;
wire net_13399;
wire net_15071;
wire net_5826;
wire net_4074;
wire net_4000;
wire net_13912;
wire net_14913;
wire net_2214;
wire net_3338;
wire net_5987;
wire net_15468;
wire net_8604;
wire net_2728;
wire net_13238;
wire net_9929;
wire net_4636;
wire net_417;
wire net_122;
wire net_6264;
wire net_13619;
wire net_12847;
wire net_11514;
wire net_10634;
wire net_10026;
wire net_5387;
wire x1192;
wire net_8217;
wire net_9262;
wire net_14752;
wire net_7467;
wire net_4092;
wire x447;
wire net_10758;
wire net_12300;
wire net_8595;
wire net_8287;
wire net_3337;
wire net_2662;
wire net_94;
wire net_11760;
wire net_10751;
wire net_15361;
wire net_3752;
wire net_4486;
wire net_9427;
wire net_9131;
wire net_482;
wire net_5144;
wire net_10805;
wire net_3258;
wire net_10942;
wire net_15437;
wire net_10983;
wire net_7262;
wire net_149;
wire net_387;
wire net_7790;
wire net_15327;
wire net_3275;
wire net_7447;
wire net_6297;
wire net_13107;
wire net_13127;
wire net_10828;
wire net_5291;
wire net_5160;
wire net_1893;
wire net_14137;
wire net_6494;
wire net_15355;
wire net_1932;
wire net_15035;
wire net_9639;
wire net_8896;
wire net_11620;
wire net_8268;
wire net_3836;
wire net_577;
wire net_13245;
wire net_3401;
wire net_10313;
wire net_14554;
wire net_2550;
wire net_797;
wire net_7747;
wire net_3545;
wire net_1957;
wire net_1799;
wire net_10150;
wire net_11224;
wire net_10102;
wire net_15132;
wire net_13743;
wire net_13231;
wire net_9368;
wire net_11859;
wire net_15377;
wire net_12909;
wire net_9218;
wire net_7581;
wire net_2572;
wire net_2414;
wire net_337;
wire net_10581;
wire net_1846;
wire net_13312;
wire net_4476;
wire net_690;
wire net_13381;
wire net_5667;
wire net_11222;
wire net_7933;
wire net_6820;
wire net_9662;
wire net_3743;
wire net_7888;
wire net_12475;
wire net_523;
wire net_11066;
wire net_13984;
wire net_11070;
wire net_4254;
wire net_13760;
wire net_6718;
wire net_3815;
wire net_3555;
wire net_7144;
wire net_5739;
wire net_2371;
wire net_3375;
wire net_6744;
wire net_9620;
wire net_6794;
wire net_14077;
wire net_4926;
wire net_3467;
wire net_9617;
wire net_13368;
wire net_8972;
wire net_11014;
wire net_9760;
wire net_8396;
wire net_12546;
wire net_9640;
wire net_7843;
wire net_7392;
wire net_4467;
wire net_3982;
wire net_1388;
wire net_12129;
wire net_5028;
wire net_4709;
wire net_14409;
wire net_4721;
wire net_14959;
wire net_5756;
wire net_9858;
wire net_3391;
wire net_15018;
wire net_2730;
wire net_4426;
wire net_1631;
wire net_1337;
wire net_6835;
wire net_5786;
wire net_14254;
wire net_13553;
wire net_1182;
wire net_4655;
wire net_1624;
wire net_7231;
wire net_6618;
wire net_12332;
wire net_13656;
wire net_1638;
wire net_14458;
wire net_1950;
wire net_15067;
wire net_9052;
wire net_7455;
wire net_3875;
wire net_12146;
wire net_9319;
wire net_9280;
wire net_14803;
wire net_7039;
wire net_14436;
wire net_10135;
wire net_2421;
wire net_5684;
wire net_5268;
wire net_11389;
wire net_4901;
wire net_4804;
wire net_880;
wire net_1402;
wire net_14980;
wire net_6335;
wire net_2153;
wire net_1939;
wire net_9582;
wire net_4100;
wire net_8781;
wire net_8474;
wire net_3098;
wire net_7242;
wire net_14190;
wire net_8535;
wire net_6288;
wire net_4673;
wire net_5762;
wire net_9061;
wire net_5151;
wire net_13922;
wire net_10249;
wire net_11876;
wire net_7828;
wire net_2901;
wire net_162;
wire net_15751;
wire net_14952;
wire net_8301;
wire net_13255;
wire net_4950;
wire net_7776;
wire net_4944;
wire net_653;
wire net_14301;
wire net_13160;
wire net_5066;
wire net_13919;
wire net_14718;
wire net_11735;
wire net_12661;
wire net_12030;
wire net_4847;
wire net_3052;
wire net_3145;
wire net_10906;
wire net_6652;
wire net_9558;
wire net_13694;
wire net_3694;
wire net_11554;
wire net_7295;
wire net_14880;
wire net_10262;
wire net_11592;
wire net_6368;
wire net_14889;
wire net_3855;
wire net_236;
wire net_12324;
wire net_487;
wire net_9286;
wire net_552;
wire net_10823;
wire net_8861;
wire net_8206;
wire net_7992;
wire net_1787;
wire net_3551;
wire net_6654;
wire net_7440;
wire net_14791;
wire net_13390;
wire net_5056;
wire net_9518;
wire net_756;
wire net_7067;
wire net_7735;
wire net_13636;
wire net_4765;
wire net_15143;
wire net_14234;
wire net_8329;
wire net_104;
wire net_12230;
wire net_10101;
wire net_7798;
wire net_14402;
wire net_11301;
wire net_5031;
wire net_15477;
wire net_3416;
wire net_7198;
wire net_5166;
wire net_11845;
wire net_14595;
wire net_4886;
wire net_9878;
wire net_3537;
wire net_15655;
wire net_10914;
wire net_14070;
wire net_12039;
wire net_8522;
wire net_6659;
wire net_15541;
wire net_12897;
wire net_12192;
wire net_6877;
wire net_711;
wire net_2225;
wire net_7659;
wire net_15257;
wire net_15635;
wire net_4741;
wire net_11687;
wire net_15720;
wire net_8618;
wire net_4700;
wire net_846;
wire net_10469;
wire net_9402;
wire net_12852;
wire net_3017;
wire x1343;
wire net_11864;
wire net_4677;
wire net_11420;
wire net_8033;
wire net_10996;
wire net_10038;
wire net_5768;
wire net_174;
wire net_2607;
wire net_7799;
wire net_15210;
wire net_7957;
wire net_10971;
wire net_7987;
wire net_14755;
wire net_7214;
wire net_15208;
wire net_11691;
wire net_8769;
wire net_6202;
wire net_1831;
wire net_1482;
wire net_13870;
wire x1660;
wire net_5023;
wire net_3291;
wire net_2168;
wire net_3306;
wire net_2928;
wire net_14573;
wire net_14460;
wire net_7563;
wire net_1885;
wire net_1030;
wire net_4129;
wire net_1485;
wire net_14357;
wire net_10272;
wire net_9236;
wire net_10406;
wire net_10053;
wire net_6929;
wire net_3245;
wire net_13300;
wire net_10682;
wire net_9385;
wire net_7473;
wire net_6920;
wire x208;
wire net_14742;
wire net_7335;
wire net_7387;
wire net_15498;
wire net_11987;
wire net_13407;
wire net_12740;
wire net_12711;
wire net_10787;
wire net_11498;
wire net_10031;
wire net_4773;
wire net_4201;
wire net_13929;
wire net_4273;
wire net_1969;
wire net_745;
wire net_14737;
wire net_9651;
wire net_7991;
wire net_15514;
wire net_12306;
wire net_8009;
wire net_7064;
wire net_14271;
wire net_933;
wire net_1244;
wire net_12532;
wire net_429;
wire net_12036;
wire net_10966;
wire net_10860;
wire net_3377;
wire net_373;
wire net_12593;
wire net_356;
wire net_13701;
wire net_452;
wire net_11432;
wire net_545;
wire net_3683;
wire net_11700;
wire net_1483;
wire net_2147;
wire net_10361;
wire net_8067;
wire net_560;
wire net_3031;
wire net_9253;
wire net_10098;
wire net_5148;
wire net_15120;
wire net_4603;
wire net_2645;
wire net_14017;
wire net_10433;
wire net_15586;
wire net_11951;
wire net_5510;
wire net_5356;
wire net_10500;
wire net_9359;
wire net_6709;
wire net_14386;
wire net_8078;
wire net_7310;
wire net_7674;
wire net_7386;
wire net_6684;
wire net_13151;
wire net_4278;
wire net_7522;
wire net_2674;
wire net_13801;
wire net_2872;
wire net_6833;
wire net_2432;
wire net_12780;
wire net_10193;
wire net_8934;
wire net_7059;
wire net_5401;
wire net_14428;
wire net_322;
wire net_1671;
wire net_4764;
wire x4285;
wire net_420;
wire net_665;
wire net_1746;
wire net_2222;
wire net_8944;
wire net_2322;
wire net_2825;
wire net_7209;
wire net_3670;
wire net_14647;
wire net_9109;
wire net_5940;
wire net_4344;
wire net_13376;
wire net_3341;
wire net_5985;
wire net_7925;
wire net_1072;
wire net_6606;
wire net_10182;
wire net_10376;
wire net_7136;
wire net_4861;
wire net_13738;
wire net_11666;
wire net_109;
wire net_1706;
wire net_15527;
wire net_4510;
wire net_11113;
wire net_3574;
wire net_6278;
wire net_5994;
wire net_1730;
wire net_10852;
wire net_2921;
wire x6252;
wire net_3289;
wire net_8829;
wire net_6311;
wire net_13501;
wire net_4575;
wire net_10225;
wire net_651;
wire net_14653;
wire net_12097;
wire net_2931;
wire net_3114;
wire net_3415;
wire net_6846;
wire net_10019;
wire net_744;
wire net_8276;
wire net_4967;
wire net_598;
wire net_15620;
wire net_7985;
wire net_4136;
wire net_2011;
wire net_3455;
wire net_6317;
wire net_12011;
wire net_15023;
wire net_10068;
wire net_777;
wire net_4806;
wire net_13203;
wire net_7185;
wire net_4818;
wire net_3157;
wire net_8690;
wire net_2820;
wire net_8348;
wire net_7532;
wire net_6091;
wire net_490;
wire net_4404;
wire net_14805;
wire net_11497;
wire net_3068;
wire net_12677;
wire net_8585;
wire net_5973;
wire net_12130;
wire net_3892;
wire net_13930;
wire net_7921;
wire net_6009;
wire net_3462;
wire net_7080;
wire net_6739;
wire net_5978;
wire net_5670;
wire net_632;
wire net_4439;
wire net_843;
wire net_3860;
wire net_15652;
wire net_15603;
wire net_5602;
wire net_12720;
wire net_7638;
wire net_2841;
wire net_10106;
wire net_10063;
wire net_11889;
wire net_5484;
wire net_7255;
wire net_5813;
wire net_1977;
wire net_11959;
wire net_2100;
wire net_2938;
wire net_14009;
wire net_2122;
wire net_14568;
wire x1402;
wire net_12572;
wire net_6617;
wire net_1171;
wire net_10691;
wire net_1540;
wire net_9680;
wire net_248;
wire net_3594;
wire net_6548;
wire net_5341;
wire net_11835;
wire net_9734;
wire net_10393;
wire net_1725;
wire net_14064;
wire net_13583;
wire net_3541;
wire net_15268;
wire net_5649;
wire net_13718;
wire net_3532;
wire net_12725;
wire net_5112;
wire net_1767;
wire net_4010;
wire net_7333;
wire net_11827;
wire net_1640;
wire net_12956;
wire x6186;
wire net_13788;
wire net_10303;
wire net_9750;
wire net_5190;
wire net_2724;
wire net_11916;
wire net_14712;
wire net_6554;
wire net_12090;
wire net_7504;
wire net_503;
wire net_1741;
wire net_10141;
wire net_13510;
wire net_4227;
wire net_5695;
wire net_11818;
wire net_1672;
wire net_2103;
wire net_996;
wire net_3091;
wire net_7550;
wire net_14165;
wire net_2994;
wire net_11617;
wire net_959;
wire net_5381;
wire net_10838;
wire net_8327;
wire net_11476;
wire net_7911;
wire net_3051;
wire net_8767;
wire net_4004;
wire net_7706;
wire net_2345;
wire net_12342;
wire net_9304;
wire net_2973;
wire net_6981;
wire net_6460;
wire net_3106;
wire net_13792;
wire net_2503;
wire net_9705;
wire net_6660;
wire net_2164;
wire net_15170;
wire net_11079;
wire net_6646;
wire net_5659;
wire net_11797;
wire net_13578;
wire net_6469;
wire net_3751;
wire net_8330;
wire net_9821;
wire net_6211;
wire net_5311;
wire net_4564;
wire net_13670;
wire net_2338;
wire net_15685;
wire net_10982;
wire net_10556;
wire net_4606;
wire net_3721;
wire net_2616;
wire net_8200;
wire net_8894;
wire net_282;
wire net_1596;
wire net_10804;
wire net_6572;
wire net_12397;
wire net_4296;
wire net_11677;
wire net_7416;
wire net_15064;
wire net_6901;
wire net_14726;
wire net_11857;
wire net_5051;
wire net_10688;
wire net_10908;
wire net_11693;
wire net_2370;
wire net_2047;
wire net_8320;
wire net_2469;
wire net_11214;
wire net_9647;
wire net_12733;
wire net_2693;
wire net_13115;
wire net_14819;
wire net_14824;
wire net_11212;
wire net_10458;
wire net_1012;
wire net_1404;
wire net_12765;
wire net_12185;
wire net_9621;
wire net_907;
wire net_14473;
wire net_3076;
wire net_8809;
wire net_5807;
wire net_4694;
wire net_15124;
wire net_395;
wire net_2036;
wire net_15448;
wire net_12988;
wire net_9182;
wire net_8070;
wire net_2719;
wire net_10219;
wire net_6343;
wire net_8623;
wire net_2323;
wire net_9688;
wire net_3867;
wire x1223;
wire net_3677;
wire net_641;
wire net_15088;
wire net_4811;
wire net_5451;
wire net_2798;
wire net_15336;
wire net_5071;
wire net_10977;
wire net_10599;
wire net_4972;
wire net_3869;
wire net_14335;
wire net_1152;
wire net_1226;
wire net_10459;
wire net_14212;
wire x890;
wire net_10525;
wire net_8429;
wire net_4890;
wire net_1901;
wire net_3021;
wire net_5315;
wire net_15533;
wire net_3711;
wire net_14976;
wire net_10257;
wire net_3805;
wire net_7580;
wire net_3942;
wire net_15352;
wire net_7836;
wire net_4580;
wire net_602;
wire net_12605;
wire net_8273;
wire net_2379;
wire net_13199;
wire net_1818;
wire net_12783;
wire net_11850;
wire net_13335;
wire net_12288;
wire net_10932;
wire net_8646;
wire net_2918;
wire net_11658;
wire net_9371;
wire net_1497;
wire net_1800;
wire net_14480;
wire net_4634;
wire net_279;
wire net_1523;
wire net_3347;
wire net_1656;
wire net_6522;
wire net_12281;
wire net_4039;
wire net_11326;
wire net_4030;
wire net_15179;
wire net_691;
wire net_10212;
wire net_6951;
wire net_15506;
wire net_10713;
wire net_6337;
wire net_14119;
wire net_5551;
wire net_3178;
wire net_2701;
wire net_14289;
wire net_10422;
wire net_4078;
wire net_1863;
wire net_2833;
wire x3307;
wire net_2561;
wire net_15108;
wire net_12170;
wire net_15224;
wire net_13775;
wire net_10774;
wire net_8399;
wire net_2519;
wire net_471;
wire net_1055;
wire net_3813;
wire net_3894;
wire net_878;
wire net_1531;
wire net_1159;
wire net_10666;
wire net_518;
wire net_10334;
wire net_861;
wire net_6755;
wire net_7217;
wire net_12645;
wire net_11136;
wire net_10172;
wire net_14523;
wire net_13533;
wire net_929;
wire net_6696;
wire net_12400;
wire net_11102;
wire net_2523;
wire net_4914;
wire net_11779;
wire net_4210;
wire net_3954;
wire net_12939;
wire net_11811;
wire net_5726;
wire net_1565;
wire net_10882;
wire net_8544;
wire net_5262;
wire net_14487;
wire net_169;
wire net_15347;
wire net_12951;
wire net_9948;
wire net_5213;
wire net_7696;
wire net_8567;
wire net_12986;
wire net_2234;
wire net_4552;
wire net_12120;
wire net_15629;
wire net_6828;
wire net_10481;
wire net_967;
wire net_1527;
wire net_13270;
wire net_13056;
wire net_4420;
wire net_11849;
wire net_8007;
wire net_268;
wire net_13861;
wire net_4318;
wire net_12358;
wire net_11475;
wire net_3386;
wire net_4134;
wire net_4910;
wire x526;
wire net_6631;
wire net_15627;
wire net_13324;
wire net_1645;
wire net_2962;
wire net_9406;
wire net_4365;
wire net_14536;
wire net_176;
wire net_3638;
wire net_2570;
wire net_12410;
wire net_5793;
wire net_15036;
wire net_13195;
wire net_3354;
wire net_9468;
wire net_614;
wire net_2712;
wire net_13976;
wire net_2005;
wire net_14827;
wire net_12505;
wire net_1123;
wire net_2771;
wire net_8293;
wire net_6040;
wire net_4897;
wire net_3194;
wire net_3572;
wire net_5537;
wire net_13911;
wire net_9343;
wire net_4740;
wire net_9980;
wire net_8338;
wire net_1192;
wire net_11241;
wire net_10697;
wire net_6857;
wire net_4838;
wire net_5958;
wire net_14368;
wire net_4542;
wire net_984;
wire net_3363;
wire net_11894;
wire net_11753;
wire net_11705;
wire net_6407;
wire net_5467;
wire net_15093;
wire net_10915;
wire net_7263;
wire net_13652;
wire net_8730;
wire net_4061;
wire net_1105;
wire net_12370;
wire net_12201;
wire net_2172;
wire net_3156;
wire net_12109;
wire net_2482;
wire net_13043;
wire net_11448;
wire net_7275;
wire net_707;
wire net_14023;
wire net_6534;
wire net_7491;
wire net_4457;
wire net_5039;
wire net_9519;
wire net_11174;
wire net_6867;
wire net_4850;
wire net_1856;
wire net_830;
wire net_13828;
wire net_4531;
wire net_14778;
wire net_575;
wire net_1279;
wire net_14642;
wire net_1047;
wire net_5833;
wire net_13003;
wire net_4715;
wire net_7169;
wire net_9475;
wire net_3697;
wire net_12642;
wire net_11374;
wire net_8439;
wire net_6394;
wire net_14810;
wire net_14553;
wire net_12582;
wire net_11425;
wire net_6193;
wire net_4688;
wire net_2631;
wire net_8101;
wire net_12386;
wire net_6431;
wire net_3618;
wire net_12926;
wire net_1467;
wire net_9156;
wire net_7562;
wire net_5623;
wire net_1061;
wire net_3181;
wire net_14012;
wire net_10842;
wire net_5951;
wire net_5512;
wire net_765;
wire net_1342;
wire net_2633;
wire net_1666;
wire net_3837;
wire net_9096;
wire net_4839;
wire net_2288;
wire net_14843;
wire net_4193;
wire net_15661;
wire net_8718;
wire net_13752;
wire net_8573;
wire net_8253;
wire net_11189;
wire net_15213;
wire net_2099;
wire net_15390;
wire net_5745;
wire net_6750;
wire net_5182;
wire net_7612;
wire net_13454;
wire net_9809;
wire net_10302;
wire net_8195;
wire net_5850;
wire net_5646;
wire net_2021;
wire net_11248;
wire net_1068;
wire net_15200;
wire net_186;
wire net_14378;
wire net_3983;
wire net_8121;
wire net_2495;
wire net_15229;
wire net_15730;
wire net_12823;
wire net_6672;
wire net_3814;
wire net_10534;
wire net_1050;
wire net_6266;
wire net_2072;
wire net_2760;
wire net_5914;
wire net_4751;
wire net_1872;
wire net_2271;
wire net_1716;
wire net_13926;
wire net_5327;
wire net_5003;
wire net_1607;
wire net_14083;
wire net_11768;
wire net_5247;
wire net_12164;
wire net_6125;
wire net_7143;
wire net_13472;
wire net_7983;
wire net_1263;
wire net_12331;
wire net_4591;
wire net_196;
wire net_3452;
wire net_14356;
wire net_11969;
wire net_10324;
wire net_8766;
wire net_2067;
wire net_14243;
wire net_8120;
wire net_3130;
wire net_8881;
wire net_8572;
wire net_15157;
wire net_5183;
wire x1792;
wire net_7200;
wire net_5704;
wire net_1639;
wire net_5267;
wire net_4126;
wire net_4289;
wire net_4549;
wire net_9775;
wire net_7284;
wire net_11431;
wire net_3625;
wire net_14435;
wire net_9510;
wire x813;
wire net_4145;
wire net_7604;
wire net_13806;
wire net_4712;
wire net_11340;
wire net_260;
wire net_15145;
wire net_2947;
wire net_15729;
wire net_12552;
wire net_11784;
wire net_3137;
wire net_11981;
wire net_732;
wire net_2152;
wire net_8649;
wire net_12880;
wire net_12423;
wire x6220;
wire net_5286;
wire net_1597;
wire net_8285;
wire net_6105;
wire net_7946;
wire net_2088;
wire net_13083;
wire net_8785;
wire net_7572;
wire net_6423;
wire net_13963;
wire net_10655;
wire net_7593;
wire net_4217;
wire net_2689;
wire net_3988;
wire net_2761;
wire net_6396;
wire net_8422;
wire net_3788;
wire net_15605;
wire net_4355;
wire net_11678;
wire net_15399;
wire net_11092;
wire net_10623;
wire net_1503;
wire net_3961;
wire net_13970;
wire net_8430;
wire net_4639;
wire net_8628;
wire net_11089;
wire net_449;
wire net_5494;
wire net_5234;
wire net_9299;
wire net_8225;
wire net_11523;
wire net_11928;
wire net_9574;
wire net_12638;
wire net_15697;
wire net_1087;
wire net_4234;
wire net_11064;
wire net_3995;
wire net_733;
wire net_8245;
wire net_887;
wire net_5856;
wire net_9606;
wire net_12362;
wire net_11409;
wire net_6098;
wire net_11975;
wire net_7537;
wire net_6595;
wire net_13663;
wire net_11653;
wire net_10491;
wire net_6151;
wire net_13866;
wire net_6301;
wire net_5443;
wire net_2308;
wire net_5211;
wire net_4731;
wire net_2989;
wire net_9105;
wire net_497;
wire net_6720;
wire net_4628;
wire net_12494;
wire net_2770;
wire net_7658;
wire net_15291;
wire net_1424;
wire net_2636;
wire net_8160;
wire net_1414;
wire net_4375;
wire net_4153;
wire net_4412;
wire net_11307;
wire net_10927;
wire net_9864;
wire net_300;
wire net_9287;
wire net_2652;
wire net_5526;
wire net_10149;
wire net_1233;
wire net_2720;
wire net_8167;
wire net_6351;
wire net_4280;
wire net_15058;
wire net_12917;
wire net_10347;
wire net_1834;
wire net_9563;
wire net_950;
wire net_6027;
wire net_4925;
wire net_13213;
wire net_15258;
wire net_13024;
wire net_13313;
wire net_15690;
wire net_11441;
wire net_11355;
wire net_5474;
wire net_14363;
wire net_9839;
wire net_9745;
wire net_2816;
wire net_6610;
wire net_7651;
wire net_14507;
wire net_8984;
wire net_14344;
wire net_12565;
wire net_1214;
wire net_9529;
wire net_3641;
wire net_13405;
wire net_12895;
wire net_10203;
wire net_866;
wire net_11946;
wire net_13603;
wire net_15705;
wire net_12700;
wire net_5194;
wire net_4220;
wire net_12025;
wire net_3150;
wire net_9596;
wire net_10681;
wire net_1032;
wire net_15563;
wire net_567;
wire net_13985;
wire net_3726;
wire net_3979;
wire net_5255;
wire net_5787;
wire net_272;
wire net_8822;
wire net_13345;
wire net_13384;
wire net_8458;
wire net_3939;
wire x3858;
wire net_14625;
wire net_12712;
wire net_12480;
wire net_1024;
wire net_1590;
wire net_14097;
wire net_1612;
wire net_839;
wire net_11121;
wire net_814;
wire net_13542;
wire net_11778;
wire net_13685;
wire net_7095;
wire net_8128;
wire net_5840;
wire net_6184;
wire net_12705;
wire net_4660;
wire net_12525;
wire net_14003;
wire net_10639;
wire net_4785;
wire net_3930;
wire x1459;
wire net_9815;
wire net_2586;
wire net_3299;
wire net_13013;
wire net_10290;
wire net_1655;
wire net_11294;
wire net_6963;
wire net_7805;
wire net_11313;
wire net_954;
wire net_2365;
wire net_13094;
wire net_4565;
wire net_9051;
wire net_9037;
wire net_4797;
wire net_15048;
wire net_8796;
wire net_11271;
wire net_8962;
wire net_10897;
wire net_9240;
wire net_10810;
wire net_2361;
wire net_2598;
wire net_14767;
wire net_11194;
wire net_2879;
wire net_10152;
wire net_1680;
wire net_15671;
wire net_14219;
wire net_3302;
wire net_13359;
wire net_13265;
wire net_14456;
wire net_9545;
wire net_10411;
wire net_15276;
wire net_7540;
wire net_12445;
wire net_11337;
wire net_11989;
wire net_4790;
wire net_3187;
wire x4937;
wire net_12048;
wire net_15250;
wire net_2622;
wire net_5363;
wire net_5966;
wire x6401;
wire net_7529;
wire net_10514;
wire net_8294;
wire net_10997;
wire net_8888;
wire net_6665;
wire net_4900;
wire net_14500;
wire net_9807;
wire net_13222;
wire net_2262;
wire net_7505;
wire net_6502;
wire net_14888;
wire net_14783;
wire net_7305;
wire net_6163;
wire net_3011;
wire net_13079;
wire net_10643;
wire net_2087;
wire net_13187;
wire net_10021;
wire net_1002;
wire net_12946;
wire net_6817;
wire net_6000;
wire net_9079;
wire net_8863;
wire net_14859;
wire net_7620;
wire net_11930;
wire net_7224;
wire net_6118;
wire net_13628;
wire net_3188;
wire net_12466;
wire net_9536;
wire net_13308;
wire net_12887;
wire net_1993;
wire net_8198;
wire net_3010;
wire net_11128;
wire net_881;
wire net_12657;
wire net_8724;
wire net_10544;
wire net_2805;
wire net_8683;
wire net_1397;
wire net_2903;
wire net_14619;
wire net_14231;
wire net_15182;
wire net_4474;
wire net_14623;
wire x916;
wire net_11623;
wire net_8392;
wire net_9556;
wire net_4128;
wire net_4923;
wire net_1954;
wire net_13036;
wire net_11866;
wire net_3873;
wire net_7615;
wire net_6015;
wire net_2155;
wire net_14294;
wire net_6741;
wire net_168;
wire net_15056;
wire net_14924;
wire net_2041;
wire net_13090;
wire net_11830;
wire net_10354;
wire net_385;
wire net_13253;
wire net_2609;
wire net_14179;
wire net_5736;
wire net_5365;
wire net_7937;
wire net_7930;
wire net_5404;
wire net_14890;
wire net_5044;
wire net_10260;
wire net_8657;
wire net_7196;
wire net_8139;
wire net_12197;
wire net_10468;
wire net_11220;
wire net_6236;
wire net_14143;
wire net_2423;
wire net_7660;
wire net_13675;
wire net_7535;
wire net_6723;
wire net_2380;
wire net_3393;
wire net_4548;
wire net_13875;
wire net_8231;
wire net_9323;
wire net_12379;
wire net_11283;
wire net_895;
wire net_10781;
wire net_14797;
wire net_6412;
wire net_14469;
wire net_11603;
wire net_5990;
wire x1197;
wire net_14358;
wire net_1412;
wire net_15202;
wire net_12006;
wire net_8240;
wire net_7048;
wire net_9715;
wire net_15402;
wire net_7767;
wire net_8831;
wire net_12394;
wire net_10683;
wire net_12965;
wire net_12327;
wire net_13357;
wire net_1255;
wire net_7358;
wire net_12603;
wire net_7211;
wire net_1250;
wire net_8247;
wire net_13928;
wire net_15176;
wire net_207;
wire net_3040;
wire net_13762;
wire net_10825;
wire net_3557;
wire net_10609;
wire net_3643;
wire net_15149;
wire net_8801;
wire net_3004;
wire net_13639;
wire net_12102;
wire x6264;
wire net_8014;
wire net_13382;
wire net_11874;
wire net_1689;
wire net_12624;
wire net_10345;
wire net_10271;
wire net_7244;
wire net_6186;
wire net_7981;
wire net_15466;
wire net_10315;
wire net_8569;
wire net_9757;
wire net_5698;
wire net_3830;
wire net_8464;
wire net_274;
wire net_13987;
wire net_1075;
wire net_12806;
wire net_12561;
wire net_9387;
wire net_10282;
wire net_13360;
wire net_14044;
wire net_6204;
wire net_833;
wire net_930;
wire net_2387;
wire net_12599;
wire net_99;
wire net_12744;
wire net_9316;
wire net_8358;
wire net_6656;
wire net_4723;
wire net_2267;
wire net_4758;
wire net_7323;
wire net_4249;
wire net_4769;
wire net_14757;
wire net_14512;
wire net_13590;
wire net_12931;
wire net_13681;
wire net_11349;
wire net_1399;
wire net_8529;
wire net_10016;
wire net_8667;
wire net_4888;
wire net_9539;
wire net_3350;
wire net_14636;
wire net_3553;
wire net_5161;
wire net_14489;
wire x1074;
wire net_7623;
wire net_3304;
wire net_15416;
wire net_15382;
wire net_12751;
wire net_2549;
wire net_11024;
wire net_8654;
wire net_1781;
wire net_14390;
wire net_3465;
wire net_6217;
wire net_7457;
wire net_3049;
wire net_10299;
wire net_6918;
wire net_637;
wire net_13062;
wire net_2514;
wire net_9250;
wire net_2390;
wire net_12183;
wire net_5436;
wire net_4775;
wire net_2686;
wire net_3474;
wire net_5577;
wire net_5472;
wire net_2013;
wire net_1509;
wire net_529;
wire net_7477;
wire net_13503;
wire net_9447;
wire net_3495;
wire net_11262;
wire net_9887;
wire net_97;
wire net_2028;
wire net_2553;
wire net_9758;
wire net_4881;
wire net_1889;
wire net_3766;
wire net_7361;
wire net_12065;
wire net_8717;
wire net_2981;
wire net_8506;
wire net_6477;
wire net_11303;
wire net_1164;
wire net_10817;
wire net_8912;
wire net_6810;
wire net_15528;
wire net_14449;
wire net_121;
wire net_5228;
wire net_6923;
wire net_11148;
wire net_7475;
wire net_15324;
wire net_12500;
wire net_2583;
wire net_9762;
wire net_15579;
wire net_5708;
wire net_3820;
wire net_3799;
wire net_8854;
wire net_4175;
wire net_10938;
wire net_5824;
wire net_4665;
wire net_9366;
wire net_2664;
wire net_14206;
wire net_2706;
wire net_11202;
wire net_5163;
wire net_849;
wire net_5580;
wire net_14161;
wire net_11842;
wire net_10577;
wire net_8304;
wire net_7470;
wire net_5294;
wire net_11681;
wire net_2602;
wire net_14545;
wire net_6366;
wire net_5751;
wire net_401;
wire net_8449;
wire net_8165;
wire net_10720;
wire net_4484;
wire net_3798;
wire net_14906;
wire net_2714;
wire net_2183;
wire net_2557;
wire net_14903;
wire net_440;
wire x1113;
wire net_14265;
wire net_9229;
wire net_11361;
wire net_8069;
wire net_8048;
wire net_758;
wire net_10866;
wire net_14955;
wire net_5664;
wire net_13754;
wire net_14747;
wire net_14558;
wire net_6874;
wire net_4652;
wire net_718;
wire net_14482;
wire net_10846;
wire net_7773;
wire net_6178;
wire net_13563;
wire net_7682;
wire net_14193;
wire net_8707;
wire net_5504;
wire net_12995;
wire net_5714;
wire net_15133;
wire net_13367;
wire net_5838;
wire net_4998;
wire net_3255;
wire net_13946;
wire net_12215;
wire net_12303;
wire net_14078;
wire net_13545;
wire net_9848;
wire net_6564;
wire x132;
wire net_4448;
wire net_9797;
wire net_9419;
wire net_336;
wire net_12973;
wire net_10946;
wire net_15598;
wire net_5306;
wire net_10404;
wire net_14033;
wire net_9577;
wire net_1578;
wire net_14584;
wire net_9938;
wire net_11539;
wire net_8417;
wire net_2917;
wire net_8404;
wire net_15630;
wire net_6711;
wire net_3221;
wire net_697;
wire net_2003;
wire net_7708;
wire net_605;
wire net_3411;
wire net_5053;
wire net_4987;
wire net_10447;
wire x1095;
wire net_3426;
wire net_9233;
wire net_13008;
wire net_15632;
wire net_5095;
wire net_9527;
wire net_924;
wire net_8883;
wire net_12255;
wire net_5469;
wire net_1333;
wire net_5325;
wire net_9205;
wire net_10980;
wire net_7829;
wire x465;
wire net_2348;
wire net_5924;
wire net_489;
wire net_14911;
wire net_5593;
wire net_5107;
wire net_14422;
wire net_3082;
wire net_5859;
wire net_11503;
wire net_10802;
wire net_5457;
wire net_13521;
wire net_3676;
wire net_4185;
wire net_6143;
wire net_4646;
wire net_4204;
wire net_5630;
wire net_2748;
wire net_9991;
wire net_11561;
wire net_9611;
wire net_7591;
wire net_6072;
wire net_9135;
wire net_8060;
wire net_251;
wire net_6682;
wire net_2054;
wire net_9880;
wire net_128;
wire net_6295;
wire net_840;
wire net_9206;
wire net_10632;
wire net_9133;
wire net_8086;
wire net_14057;
wire net_10901;
wire net_6933;
wire net_15429;
wire net_5789;
wire net_13281;
wire net_15160;
wire net_14133;
wire net_12928;
wire net_11229;
wire net_2793;
wire net_9914;
wire net_411;
wire net_2137;
wire net_1836;
wire net_14971;
wire net_10570;
wire net_8783;
wire net_4310;
wire net_11689;
wire net_15075;
wire net_12220;
wire net_11256;
wire net_12688;
wire net_5922;
wire net_14571;
wire net_13158;
wire net_7874;
wire net_7293;
wire net_11557;
wire net_8975;
wire net_3430;
wire net_8266;
wire net_1862;
wire net_13889;
wire net_10052;
wire net_2317;
wire net_15016;
wire net_6795;
wire net_6248;
wire net_8135;
wire net_14882;
wire net_4244;
wire net_10584;
wire net_7887;
wire net_6035;
wire net_6930;
wire net_6492;
wire net_3583;
wire net_112;
wire net_8183;
wire net_4396;
wire net_6158;
wire net_10536;
wire net_8219;
wire net_2373;
wire net_11694;
wire net_14109;
wire net_9273;
wire net_2398;
wire net_4581;
wire net_12140;
wire net_7811;
wire net_4431;
wire net_15374;
wire net_10943;
wire net_7821;
wire net_7746;
wire net_9282;
wire net_3315;
wire net_2455;
wire net_15137;
wire net_1609;
wire net_402;
wire net_7847;
wire net_4047;
wire net_3448;
wire net_12732;
wire net_7108;
wire net_3248;
wire net_10753;
wire net_12450;
wire net_2274;
wire net_11597;
wire net_8493;
wire net_8744;
wire net_12681;
wire net_1386;
wire net_11488;
wire net_7841;
wire net_13859;
wire net_10950;
wire net_9431;
wire net_12345;
wire net_2359;
wire net_8949;
wire net_6546;
wire net_6115;
wire net_12805;
wire net_10550;
wire net_15038;
wire net_13101;
wire net_12574;
wire net_5991;
wire net_10252;
wire net_5101;
wire net_15432;
wire net_14968;
wire net_11585;
wire net_14989;
wire net_10127;
wire net_4102;
wire net_2186;
wire net_3696;
wire net_13551;
wire net_3473;
wire net_6908;
wire net_1430;
wire net_9964;
wire net_12062;
wire net_6892;
wire net_569;
wire net_2478;
wire net_6429;
wire net_2563;
wire net_13877;
wire net_12435;
wire net_9484;
wire net_9243;
wire net_8051;
wire net_5679;
wire net_12767;
wire net_3408;
wire net_4870;
wire net_630;
wire net_12514;
wire net_8857;
wire net_2202;
wire net_2490;
wire net_8841;
wire x5225;
wire net_4018;
wire net_14861;
wire net_4428;
wire net_1791;
wire net_6826;
wire net_4339;
wire net_1471;
wire net_9975;
wire net_15249;
wire net_8997;
wire net_7667;
wire net_3608;
wire net_13696;
wire net_3124;
wire net_1903;
wire net_2407;
wire net_13467;
wire net_14892;
wire net_10600;
wire net_912;
wire net_13162;
wire net_7412;
wire net_13414;
wire net_13562;
wire net_7018;
wire net_4517;
wire net_15315;
wire net_2078;
wire net_779;
wire net_1928;
wire net_3841;
wire net_12473;
wire net_14438;
wire net_1328;
wire net_9871;
wire net_234;
wire net_2859;
wire net_12634;
wire net_4151;
wire net_2884;
wire net_3848;
wire net_13258;
wire net_5372;
wire net_5142;
wire net_4942;
wire net_13616;
wire net_3205;
wire net_15309;
wire net_1094;
wire net_3487;
wire net_2749;
wire net_7390;
wire net_5764;
wire net_855;
wire net_11469;
wire net_674;
wire net_7732;
wire net_11032;
wire net_9506;
wire net_303;
wire net_10041;
wire net_6583;
wire net_9128;
wire net_9982;
wire net_491;
wire net_2475;
wire net_11460;
wire net_9925;
wire net_1299;
wire net_6679;
wire net_948;
wire net_2937;
wire net_7792;
wire net_7657;
wire net_7400;
wire net_6191;
wire net_11573;
wire net_14744;
wire net_12249;
wire net_12993;
wire net_7865;
wire net_4743;
wire net_13767;
wire net_876;
wire net_2593;
wire net_6479;
wire net_2162;
wire net_10833;
wire net_9478;
wire net_2439;
wire net_15424;
wire net_13297;
wire net_11048;
wire net_7154;
wire net_172;
wire net_9646;
wire net_4341;
wire net_13460;
wire net_8601;
wire net_15300;
wire x4781;
wire net_11960;
wire net_1458;
wire net_4048;
wire net_5587;
wire net_10749;
wire net_4570;
wire net_10184;
wire net_10244;
wire net_5933;
wire net_6689;
wire net_10591;
wire net_905;
wire net_14122;
wire net_12233;
wire net_13934;
wire net_142;
wire net_7034;
wire net_6446;
wire net_8029;
wire net_11939;
wire net_9050;
wire net_6198;
wire net_2229;
wire net_13842;
wire net_10613;
wire net_5774;
wire net_158;
wire net_7370;
wire net_3200;
wire net_14848;
wire net_3733;
wire net_3881;
wire net_12263;
wire net_15457;
wire net_8598;
wire net_5624;
wire net_11944;
wire net_2504;
wire net_11571;
wire net_5650;
wire net_2175;
wire net_3784;
wire net_10519;
wire net_14136;
wire net_15637;
wire net_15481;
wire net_10214;
wire net_8091;
wire net_8057;
wire net_6258;
wire net_8361;
wire net_2116;
wire net_1758;
wire net_4327;
wire net_14701;
wire net_13840;
wire net_11334;
wire net_8813;
wire net_8035;
wire net_14868;
wire net_11802;
wire net_9572;
wire net_8090;
wire net_1769;
wire net_9115;
wire net_6694;
wire net_1967;
wire net_15504;
wire net_11565;
wire net_9333;
wire net_5171;
wire net_1567;
wire net_8020;
wire net_6860;
wire net_6322;
wire x5289;
wire net_12087;
wire net_8754;
wire net_15286;
wire net_465;
wire net_11186;
wire net_8152;
wire net_14676;
wire net_9520;
wire net_1883;
wire net_14930;
wire net_11233;
wire net_476;
wire net_2783;
wire net_14461;
wire net_6055;
wire net_7079;
wire net_382;
wire net_3058;
wire net_11412;
wire net_8484;
wire net_11259;
wire net_5301;
wire net_583;
wire net_1315;
wire net_6994;
wire net_5904;
wire net_7041;
wire net_5358;
wire net_10073;
wire net_9408;
wire net_14173;
wire net_9767;
wire net_5208;
wire net_13144;
wire net_5019;
wire net_9903;
wire net_9376;
wire net_6956;
wire net_13055;
wire net_9695;
wire net_4719;
wire net_10379;
wire net_10138;
wire net_4977;
wire net_15234;
wire net_9005;
wire net_5075;
wire net_4460;
wire net_11646;
wire net_7327;
wire net_220;
wire net_1465;
wire net_293;
wire net_15117;
wire net_11153;
wire net_3666;
wire net_13599;
wire net_11890;
wire net_4982;
wire net_13303;
wire net_1938;
wire net_543;
wire net_15677;
wire net_625;
wire net_3760;
wire net_11411;
wire net_10708;
wire net_14660;
wire net_1823;
wire net_5081;
wire net_15543;
wire net_15516;
wire net_11637;
wire net_14509;
wire net_13790;
wire net_191;
wire net_3576;
wire net_4331;
wire net_2909;
wire net_4953;
wire net_558;
wire net_15021;
wire net_2069;
wire net_15464;
wire net_9607;
wire net_4697;
wire net_5638;
wire x80;
wire net_1618;
wire net_10910;
wire net_14399;
wire net_2497;
wire net_7899;
wire net_15594;
wire net_11594;
wire net_12157;
wire net_10562;
wire net_7006;
wire net_3562;
wire net_15319;
wire net_1694;
wire net_12844;
wire net_15110;
wire net_4991;
wire net_910;
wire net_12356;
wire net_5885;
wire net_15332;
wire net_7112;
wire net_11905;
wire net_5394;
wire net_7944;
wire net_2412;
wire net_4023;
wire net_14720;
wire net_12070;
wire net_4265;
wire net_7755;
wire net_6881;
wire net_4450;
wire net_14563;
wire net_4158;
wire net_15610;
wire net_6942;
wire net_13442;
wire net_1984;
wire net_13959;
wire net_13527;
wire net_315;
wire net_1375;
wire net_4670;
wire net_10734;
wire net_1944;
wire net_4006;
wire net_11545;
wire net_8212;
wire net_1351;
wire net_1775;
wire net_10112;
wire net_10158;
wire net_346;
wire net_297;
wire net_1535;
wire net_2400;
wire net_5543;
wire net_10693;
wire net_13725;
wire net_8661;
wire net_10959;
wire net_2034;
wire net_229;
wire net_15189;
wire net_14835;
wire net_4360;
wire net_14963;
wire net_8921;
wire net_4962;
wire net_1808;
wire net_3256;
wire net_687;
wire net_15073;
wire net_3266;
wire net_13122;
wire net_4160;
wire net_14702;
wire net_13339;
wire net_15003;
wire net_3888;
wire net_14916;
wire net_7072;
wire net_13949;
wire net_13438;
wire net_14303;
wire net_10567;
wire net_3322;
wire net_2533;
wire net_10267;
wire net_3566;
wire net_15263;
wire net_14945;
wire net_1913;
wire net_12297;
wire net_3596;
wire net_13243;
wire net_11526;
wire net_7830;
wire net_9673;
wire net_9016;
wire net_7642;
wire net_10143;
wire net_11904;
wire net_5021;
wire net_9732;
wire net_9264;
wire net_15244;
wire net_6615;
wire net_12279;
wire net_7409;
wire net_13741;
wire net_7671;
wire net_1760;
wire net_9345;
wire net_9296;
wire net_5415;
wire net_13492;
wire net_1184;
wire net_7714;
wire net_4055;
wire net_5339;
wire net_3926;
wire net_6482;
wire net_6961;
wire net_14444;
wire net_4849;
wire net_15363;
wire net_7383;
wire net_10722;
wire net_5758;
wire net_5425;
wire net_3403;
wire net_10002;
wire net_1960;
wire net_6977;
wire net_10718;
wire net_9660;
wire net_3093;
wire net_7935;
wire net_12820;
wire net_6886;
wire net_647;
wire net_3247;
wire net_15622;
wire net_15745;
wire net_12548;
wire net_7435;
wire net_15194;
wire net_6452;
wire net_8684;
wire net_2464;
wire net_12272;
wire net_9492;
wire net_9145;
wire net_4256;
wire net_828;
wire net_6222;
wire net_3839;
wire net_6513;
wire net_4490;
wire net_1603;
wire net_14349;
wire net_12222;
wire x57;
wire net_13031;
wire net_2732;
wire net_10009;
wire net_7446;
wire net_10108;
wire net_13483;
wire net_11809;
wire net_11017;
wire net_8368;
wire net_8385;
wire net_7345;
wire net_3521;
wire net_14877;
wire net_1096;
wire net_795;
wire net_982;
wire net_14874;
wire net_8153;
wire net_11403;
wire net_9610;
wire net_1580;
wire net_1406;
wire net_9093;
wire net_5287;
wire net_3896;
wire net_4384;
wire net_6462;
wire net_9189;
wire net_8490;
wire net_10463;
wire net_9314;
wire net_1434;
wire net_6996;
wire net_3668;
wire net_14728;
wire net_6096;
wire net_9576;
wire x4851;
wire net_9823;
wire net_4912;
wire net_10012;
wire net_5130;
wire net_11870;
wire net_5617;
wire net_4946;
wire net_6002;
wire net_774;
wire net_15101;
wire net_14501;
wire net_10071;
wire net_5748;
wire net_15531;
wire net_12076;
wire net_8180;
wire net_6958;
wire net_11393;
wire net_10869;
wire net_5049;
wire net_8892;
wire net_13235;
wire net_7221;
wire net_11058;
wire net_501;
wire net_8899;
wire net_3679;
wire net_14927;
wire net_225;
wire net_4489;
wire net_12344;
wire net_5818;
wire net_3128;
wire net_4733;
wire net_12937;
wire net_6524;
wire net_6213;
wire net_4692;
wire net_9769;
wire net_6644;
wire net_7481;
wire net_9170;
wire net_15334;
wire net_13327;
wire net_5313;
wire net_447;
wire net_9180;
wire net_871;
wire net_2611;
wire net_14974;
wire net_11804;
wire net_15126;
wire net_390;
wire net_13279;
wire net_5772;
wire net_1154;
wire net_6318;
wire net_11789;
wire net_11219;
wire net_6983;
wire net_6593;
wire net_14031;
wire net_10755;
wire net_13371;
wire net_11782;
wire net_9703;
wire net_12368;
wire net_8952;
wire net_13944;
wire net_4294;
wire net_5128;
wire net_10923;
wire net_6062;
wire net_15723;
wire net_12735;
wire net_7900;
wire net_7494;
wire net_14038;
wire net_4106;
wire net_12798;
wire net_2951;
wire net_8621;
wire net_3631;
wire net_12854;
wire net_2293;
wire net_12132;
wire net_280;
wire net_12027;
wire net_12715;
wire net_495;
wire net_13022;
wire net_10105;
wire net_1802;
wire net_15100;
wire net_10569;
wire net_7694;
wire net_13180;
wire net_2140;
wire net_5482;
wire net_13975;
wire net_6345;
wire net_10456;
wire net_13211;
wire net_7637;
wire net_2517;
wire net_11318;
wire net_8798;
wire net_2316;
wire net_12105;
wire net_8644;
wire net_14525;
wire net_6457;
wire net_2755;
wire net_6100;
wire net_12172;
wire net_6356;
wire net_13850;
wire net_1678;
wire net_2703;
wire net_14997;
wire net_11273;
wire net_13524;
wire net_6638;
wire net_3366;
wire net_14214;
wire net_1441;
wire net_10210;
wire net_15338;
wire net_969;
wire net_9154;
wire net_8271;
wire net_1525;
wire net_7097;
wire net_12710;
wire net_11458;
wire net_7737;
wire net_7206;
wire net_4003;
wire net_821;
wire net_13444;
wire net_6757;
wire net_4177;
wire net_9350;
wire net_8511;
wire net_7757;
wire net_11726;
wire net_15442;
wire net_8936;
wire x3949;
wire net_10934;
wire net_3436;
wire net_8345;
wire net_2335;
wire net_14159;
wire net_11210;
wire net_15500;
wire net_14603;
wire net_3940;
wire net_10812;
wire net_8708;
wire net_7725;
wire net_3911;
wire net_11533;
wire net_13913;
wire net_11161;
wire net_12866;
wire net_5337;
wire net_15557;
wire net_14153;
wire net_2618;
wire net_8638;
wire net_4316;
wire net_3365;
wire net_10711;
wire net_6045;
wire net_14372;
wire net_14099;
wire net_6540;
wire net_14688;
wire net_12698;
wire net_8587;
wire net_7952;
wire net_1114;
wire net_12786;
wire net_10619;
wire net_8670;
wire net_13431;
wire net_7090;
wire net_3388;
wire net_5411;
wire net_12691;
wire net_1748;
wire net_10664;
wire net_4116;
wire net_3078;
wire net_3218;
wire x3683;
wire net_13005;
wire net_11882;
wire net_4632;
wire net_2964;
wire net_12283;
wire net_9946;
wire net_8171;
wire net_7266;
wire net_6738;
wire x1187;
wire net_2232;
wire net_2343;
wire net_726;
wire net_13241;
wire net_6690;
wire net_6565;
wire net_15349;
wire net_3811;
wire net_1028;
wire net_14287;
wire net_1529;
wire net_600;
wire net_14021;
wire net_3237;
wire net_701;
wire net_397;
wire net_808;
wire net_5553;
wire net_11126;
wire net_7602;
wire net_5595;
wire net_10968;
wire net_9121;
wire net_9894;
wire net_1704;
wire net_12373;
wire net_5026;
wire net_4821;
wire net_1384;
wire net_2738;
wire net_8712;
wire net_3918;
wire net_9107;
wire net_5280;
wire net_320;
wire net_6844;
wire net_4916;
wire net_6902;
wire net_15211;
wire net_9251;
wire net_2944;
wire net_9103;
wire net_12530;
wire net_7063;
wire net_986;
wire net_12079;
wire net_1242;
wire net_6556;
wire net_14384;
wire net_4346;
wire net_1241;
wire net_15571;
wire net_13153;
wire net_11953;
wire net_6662;
wire net_3690;
wire net_11176;
wire net_15584;
wire net_13058;
wire net_9451;
wire net_7927;
wire net_7524;
wire net_11833;
wire net_11019;
wire net_13998;
wire net_13197;
wire net_5654;
wire net_13034;
wire net_8827;
wire net_935;
wire net_3001;
wire net_1511;
wire net_3116;
wire net_645;
wire net_14649;
wire net_11436;
wire net_3121;
wire net_10368;
wire net_4841;
wire net_4621;
wire net_10289;
wire net_10217;
wire net_4071;
wire net_1634;
wire net_10305;
wire net_6271;
wire net_609;
wire net_12034;
wire net_13343;
wire net_14242;
wire net_8825;
wire net_10862;
wire net_6155;
wire net_3083;
wire net_5693;
wire net_4533;
wire net_1816;
wire net_9782;
wire net_8076;
wire net_1221;
wire net_15419;
wire net_7909;
wire net_7158;
wire net_4195;
wire net_14085;
wire net_6911;
wire net_4895;
wire net_9851;
wire net_331;
wire net_14943;
wire net_12597;
wire net_816;
wire net_9100;
wire net_4644;
wire net_3264;
wire net_7363;
wire net_2092;
wire net_13209;
wire net_8633;
wire net_7134;
wire net_12745;
wire net_8669;
wire net_2220;
wire net_4762;
wire net_2823;
wire net_1217;
wire net_13879;
wire net_7028;
wire net_9719;
wire net_2933;
wire net_3728;
wire net_8141;
wire net_3381;
wire x4520;
wire net_10818;
wire net_14156;
wire net_8848;
wire net_5724;
wire net_7138;
wire net_4118;
wire net_4577;
wire net_4970;
wire net_1575;
wire net_4884;
wire net_3279;
wire net_12981;
wire net_657;
wire net_8000;
wire net_15537;
wire net_8495;
wire net_5042;
wire net_1727;
wire net_12541;
wire net_13808;
wire net_14333;
wire net_12841;
wire net_12199;
wire x507;
wire net_329;
wire net_5809;
wire net_4600;
wire x6327;
wire net_4753;
wire net_1259;
wire net_14633;
wire net_12848;
wire net_11207;
wire net_1924;
wire net_4225;
wire net_2143;
wire net_2839;
wire net_4287;
wire net_1825;
wire net_2196;
wire net_3791;
wire net_7676;
wire net_3168;
wire net_8059;
wire net_10478;
wire net_10078;
wire net_14714;
wire net_10558;
wire net_11611;
wire net_5275;
wire net_962;
wire net_7914;
wire net_478;
wire net_8695;
wire net_13731;
wire net_7817;
wire net_596;
wire net_11429;
wire net_6608;
wire net_11840;
wire net_1261;
wire net_8733;
wire net_5781;
wire net_4959;
wire net_2120;
wire net_1975;
wire net_15081;
wire net_4705;
wire net_10430;
wire net_14167;
wire net_8958;
wire net_8375;
wire net_7566;
wire net_14735;
wire net_13512;
wire net_13067;
wire net_11948;
wire net_13991;
wire net_12893;
wire net_565;
wire net_2569;
wire net_5600;
wire net_7406;
wire net_2832;
wire net_7530;
wire net_4478;
wire net_7253;
wire net_2149;
wire net_3028;
wire net_11281;
wire net_7087;
wire net_1692;
wire net_13174;
wire net_9736;
wire net_15654;
wire net_12675;
wire net_5079;
wire net_2528;
wire net_2655;
wire net_10611;
wire net_10363;
wire net_5062;
wire net_10854;
wire net_9682;
wire net_6518;
wire net_4236;
wire net_11618;
wire net_1361;
wire net_2450;
wire net_4813;
wire net_9260;
wire net_14118;
wire net_1208;
wire net_14679;
wire net_10986;
wire net_7948;
wire net_232;
wire net_8920;
wire net_6538;
wire net_14273;
wire net_13201;
wire net_12162;
wire net_13769;
wire net_8560;
wire net_9279;
wire net_12954;
wire net_12778;
wire net_2167;
wire net_2880;
wire net_15408;
wire net_7923;
wire net_11062;
wire net_13378;
wire net_4710;
wire net_13810;
wire net_4808;
wire net_2996;
wire net_5506;
wire net_2889;
wire net_9537;
wire net_4544;
wire net_7340;
wire net_13901;
wire net_12187;
wire net_137;
wire net_6398;
wire net_3154;
wire net_6386;
wire net_4828;
wire net_15147;
wire net_4465;
wire net_15568;
wire net_532;
wire net_2501;
wire net_3530;
wire net_13179;
wire net_9862;
wire net_13190;
wire net_3622;
wire net_10398;
wire net_9800;
wire net_10389;
wire net_2729;
wire net_14751;
wire net_4422;
wire net_14817;
wire net_10116;
wire net_302;
wire net_8223;
wire net_1131;
wire net_889;
wire net_12609;
wire net_1116;
wire net_13018;
wire net_753;
wire net_15668;
wire net_9034;
wire net_5253;
wire net_5575;
wire net_4373;
wire net_13135;
wire net_9289;
wire net_9710;
wire net_11521;
wire net_2814;
wire net_13609;
wire net_12464;
wire net_689;
wire net_751;
wire net_8084;
wire net_4155;
wire net_15172;
wire net_13864;
wire net_11297;
wire net_6353;
wire net_15222;
wire net_6722;
wire net_14670;
wire net_8288;
wire net_2363;
wire net_14346;
wire net_6283;
wire net_12861;
wire net_3659;
wire net_6578;
wire net_5232;
wire net_5192;
wire net_13708;
wire net_10512;
wire net_3724;
wire net_13129;
wire net_12301;
wire net_13268;
wire net_1228;
wire net_10146;
wire net_7148;
wire net_4593;
wire net_15615;
wire net_7807;
wire net_15561;
wire net_13092;
wire net_2722;
wire net_9891;
wire net_12139;
wire net_1426;
wire net_12649;
wire net_9399;
wire net_6504;
wire net_11111;
wire net_12013;
wire net_8531;
wire net_13113;
wire net_9813;
wire net_15190;
wire net_1407;
wire net_3147;
wire net_4903;
wire net_15343;
wire net_11548;
wire net_8536;
wire net_11380;
wire net_5409;
wire net_12949;
wire net_13602;
wire net_11795;
wire net_3263;
wire net_10093;
wire net_1057;
wire net_2915;
wire net_14610;
wire net_14129;
wire net_15673;
wire net_7235;
wire net_10895;
wire net_5225;
wire net_4931;
wire net_6161;
wire net_6953;
wire net_10647;
wire net_2987;
wire net_15199;
wire net_10509;
wire net_7261;
wire net_8613;
wire net_8233;
wire net_2253;
wire net_6189;
wire net_1699;
wire net_5114;
wire net_4398;
wire net_9534;
wire net_1042;
wire net_4783;
wire net_4076;
wire net_4792;
wire net_15703;
wire net_12944;
wire net_7788;
wire net_13267;
wire net_15589;
wire net_1000;
wire net_11309;
wire net_11133;
wire net_1995;
wire net_2521;
wire net_12915;
wire net_6246;
wire net_11296;
wire net_2545;
wire net_1016;
wire net_6437;
wire net_15256;
wire net_9035;
wire net_5158;
wire net_11315;
wire net_10017;
wire x3588;
wire net_10323;
wire net_3977;
wire net_4567;
wire net_10417;
wire net_10201;
wire net_1744;
wire net_516;
wire net_2870;
wire net_14769;
wire net_3176;
wire net_3585;
wire net_12655;
wire net_11776;
wire net_12614;
wire net_6182;
wire net_956;
wire net_4320;
wire net_3963;
wire net_11847;
wire net_5799;
wire net_14383;
wire net_2596;
wire net_5496;
wire net_10835;
wire net_2970;
wire net_14388;
wire net_12369;
wire net_438;
wire net_8181;
wire net_8178;
wire net_14001;
wire net_9001;
wire net_2584;
wire net_14052;
wire net_12334;
wire net_2250;
wire net_5278;
wire net_3013;
wire net_5438;
wire net_13826;
wire net_7546;
wire net_11963;
wire net_952;
wire net_3110;
wire net_2967;
wire net_14305;
wire net_4097;
wire net_11743;
wire net_5170;
wire net_3185;
wire net_13821;
wire net_10916;
wire net_8214;
wire net_14290;
wire net_13337;
wire net_9048;
wire net_7598;
wire net_3300;
wire net_6808;
wire net_6438;
wire net_2245;
wire net_10645;
wire net_13185;
wire net_7268;
wire net_12963;
wire net_15471;
wire net_8187;
wire net_7570;
wire net_13773;
wire net_4231;
wire net_383;
wire net_15283;
wire net_4068;
wire net_3570;
wire net_15663;
wire net_14055;
wire net_3140;
wire net_15678;
wire net_15625;
wire net_5916;
wire net_6765;
wire net_9773;
wire net_427;
wire net_7823;
wire net_135;
wire net_2785;
wire net_9693;
wire net_10840;
wire net_1121;
wire net_8575;
wire net_13169;
wire net_8274;
wire net_473;
wire net_13687;
wire net_7288;
wire net_14426;
wire net_13897;
wire net_7559;
wire net_3599;
wire net_7381;
wire net_5099;
wire net_9512;
wire net_8350;
wire net_4329;
wire net_11094;
wire net_6409;
wire net_2777;
wire net_1049;
wire net_13531;
wire net_9440;
wire net_3901;
wire net_454;
wire net_6251;
wire net_5349;
wire net_15518;
wire net_10674;
wire x784;
wire net_14674;
wire net_9364;
wire net_6707;
wire net_709;
wire net_2484;
wire net_8437;
wire net_13535;
wire net_9278;
wire net_7582;
wire net_11342;
wire net_6229;
wire net_8608;
wire net_10791;
wire net_5199;
wire net_12905;
wire net_1066;
wire net_5514;
wire net_12388;
wire net_9293;
wire net_9956;
wire net_15095;
wire net_2591;
wire net_14534;
wire net_4304;
wire net_10552;
wire net_8985;
wire net_10880;
wire net_5847;
wire net_5189;
wire net_11896;
wire net_4560;
wire net_1344;
wire net_5791;
wire net_3968;
wire net_1283;
wire net_1084;
wire net_12875;
wire net_4554;
wire net_1500;
wire net_354;
wire net_9778;
wire net_14607;
wire net_11376;
wire net_1136;
wire net_14010;
wire net_12428;
wire net_5418;
wire net_15001;
wire net_3008;
wire net_11707;
wire net_2763;
wire net_573;
wire net_12099;
wire net_9065;
wire net_3356;
wire net_12412;
wire net_11423;
wire net_7175;
wire net_5465;
wire net_6855;
wire net_13314;
wire net_12640;
wire net_11606;
wire net_3616;
wire net_9494;
wire net_3886;
wire net_7281;
wire net_1592;
wire net_13650;
wire net_2085;
wire net_13352;
wire net_8570;
wire net_5521;
wire net_5037;
wire net_3672;
wire net_11101;
wire net_6089;
wire net_4406;
wire x3698;
wire net_9249;
wire net_14371;
wire net_12557;
wire net_5621;
wire net_15425;
wire net_8764;
wire x3360;
wire net_11879;
wire net_10297;
wire net_1637;
wire net_3702;
wire net_9374;
wire net_6480;
wire net_6425;
wire net_5971;
wire net_5811;
wire net_6220;
wire net_8915;
wire net_941;
wire net_7560;
wire net_7629;
wire net_6038;
wire net_11324;
wire net_5854;
wire net_13292;
wire net_14582;
wire net_14351;
wire net_8129;
wire net_14519;
wire net_4555;
wire net_2070;
wire net_2311;
wire net_9444;
wire net_11661;
wire net_4611;
wire net_7500;
wire net_10605;
wire net_4124;
wire net_1599;
wire net_6587;
wire net_15151;
wire net_10575;
wire net_11087;
wire net_12372;
wire net_3981;
wire net_3828;
wire net_13659;
wire net_11504;
wire net_3132;
wire net_3161;
wire net_9973;
wire net_6107;
wire net_4303;
wire net_1290;
wire net_12924;
wire net_4147;
wire net_12240;
wire net_3053;
wire net_9802;
wire net_15209;
wire net_9579;
wire net_4056;
wire net_7187;
wire net_12589;
wire net_7460;
wire net_3297;
wire net_6601;
wire net_8518;
wire net_2023;
wire net_15041;
wire net_14028;
wire net_13923;
wire net_4523;
wire net_123;
wire net_11766;
wire net_5249;
wire net_1668;
wire net_527;
wire net_262;
wire net_13474;
wire net_12205;
wire net_3424;
wire net_15371;
wire net_12151;
wire net_7552;
wire net_6364;
wire net_10169;
wire net_3139;
wire net_5388;
wire net_4063;
wire net_6399;
wire net_5087;
wire net_13218;
wire net_11983;
wire net_1793;
wire net_15397;
wire net_11714;
wire net_3104;
wire net_3786;
wire net_5508;
wire net_15066;
wire net_2278;
wire net_8261;
wire net_7161;
wire net_3072;
wire net_15409;
wire net_6215;
wire net_7286;
wire net_1021;
wire net_10498;
wire net_5269;
wire net_10488;
wire net_1737;
wire net_9979;
wire net_10657;
wire net_5706;
wire net_6801;
wire net_1859;
wire net_12550;
wire net_145;
wire net_3607;
wire net_4654;
wire net_15299;
wire net_8541;
wire net_4917;
wire net_10699;
wire net_8193;
wire net_1145;
wire net_10431;
wire net_8424;
wire net_4637;
wire x6531;
wire net_2804;
wire net_11134;
wire net_9306;
wire net_2261;
wire net_9411;
wire net_5535;
wire net_188;
wire net_3753;
wire net_3061;
wire net_3319;
wire net_4353;
wire net_7414;
wire net_10160;
wire x1058;
wire net_7141;
wire net_2958;
wire net_1077;
wire net_14163;
wire net_6520;
wire net_2924;
wire net_15700;
wire net_10050;
wire net_8969;
wire net_11328;
wire net_14131;
wire net_12318;
wire net_11825;
wire net_8022;
wire net_5918;
wire net_2410;
wire net_8281;
wire net_10827;
wire net_9208;
wire net_119;
wire net_3108;
wire net_10975;
wire net_10445;
wire net_2185;
wire net_13103;
wire net_6853;
wire net_1321;
wire net_14263;
wire net_13961;
wire net_13624;
wire net_4441;
wire net_6307;
wire net_4192;
wire net_8741;
wire net_5392;
wire net_4949;
wire net_14484;
wire net_1099;
wire net_11977;
wire net_14586;
wire net_11733;
wire net_11141;
wire net_11568;
wire net_90;
wire net_14901;
wire net_7106;
wire net_4583;
wire net_7103;
wire net_14543;
wire net_9885;
wire net_9227;
wire net_15185;
wire net_12290;
wire net_404;
wire net_11683;
wire net_14941;
wire net_6033;
wire net_4663;
wire net_14330;
wire net_11624;
wire net_5455;
wire net_9276;
wire net_2666;
wire net_5822;
wire net_4084;
wire net_4500;
wire net_10929;
wire net_8045;
wire net_8402;
wire net_1239;
wire net_15351;
wire net_10246;
wire net_8663;
wire net_8591;
wire net_5879;
wire net_1463;
wire net_9743;
wire net_14250;
wire net_8793;
wire net_8562;
wire net_12257;
wire net_2056;
wire net_10081;
wire net_5716;
wire net_9266;
wire net_7884;
wire net_3822;
wire net_15139;
wire net_12217;
wire net_10800;
wire net_9147;
wire net_1628;
wire net_3476;
wire net_15162;
wire net_13957;
wire net_6872;
wire net_7347;
wire net_896;
wire net_484;
wire net_7655;
wire net_4823;
wire net_12519;
wire net_2512;
wire net_3223;
wire net_12997;
wire net_5894;
wire net_1936;
wire net_11363;
wire net_3802;
wire net_14749;
wire net_11599;
wire net_10035;
wire net_14339;
wire net_126;
wire net_15135;
wire net_2708;
wire net_8773;
wire net_8705;
wire net_10088;
wire net_10873;
wire net_9795;
wire net_12971;
wire net_9958;
wire net_2211;
wire net_13106;
wire net_11563;
wire net_7425;
wire x1206;
wire net_5479;
wire net_15031;
wire net_13939;
wire net_11794;
wire net_13001;
wire net_13614;
wire net_11550;
wire net_7917;
wire net_1896;
wire net_14090;
wire net_8388;
wire net_8777;
wire net_9998;
wire net_1732;
wire net_1982;
wire net_14577;
wire net_13283;
wire net_12687;
wire net_5926;
wire net_8089;
wire net_7866;
wire net_6348;
wire net_12084;
wire net_10014;
wire net_9390;
wire net_11719;
wire net_12149;
wire net_6509;
wire net_12507;
wire net_900;
wire net_3253;
wire net_10630;
wire net_6935;
wire net_13176;
wire net_7597;
wire net_5498;
wire net_1882;
wire net_12347;
wire net_12229;
wire net_12755;
wire net_7744;
wire net_5528;
wire net_413;
wire net_2001;
wire net_11072;
wire net_1491;
wire net_10879;
wire net_9613;
wire net_14442;
wire net_14982;
wire net_8306;
wire net_6141;
wire net_10918;
wire net_12666;
wire net_5390;
wire net_7876;
wire net_2419;
wire net_10154;
wire net_1034;
wire net_11559;
wire net_14898;
wire net_5753;
wire x73;
wire net_15634;
wire net_7608;
wire net_12203;
wire net_11510;
wire net_14315;
wire net_253;
wire net_11696;
wire net_276;
wire net_9728;
wire net_14229;
wire net_3439;
wire net_12112;
wire x185142;
wire net_8470;
wire net_13899;
wire net_13332;
wire net_10586;
wire net_6490;
wire x304;
wire net_13395;
wire net_9799;
wire net_11398;
wire net_1959;
wire net_616;
wire net_1847;
wire net_15372;
wire net_11506;
wire net_12320;
wire net_14884;
wire net_2717;
wire net_793;
wire net_9137;
wire net_460;
wire net_7356;
wire net_6797;
wire net_2353;
wire net_6074;
wire net_11919;
wire net_2272;
wire net_9231;
wire net_4206;
wire net_9708;
wire net_15566;
wire net_15365;
wire net_1133;
wire net_14788;
wire net_14222;
wire net_6131;
wire net_4104;
wire net_8133;
wire net_3287;
wire net_11712;
wire net_10724;
wire net_14922;
wire net_166;
wire net_11305;
wire net_14429;
wire net_11027;
wire net_2866;
wire net_5866;
wire net_13954;
wire net_5489;
wire net_3025;
wire net_13164;
wire net_3871;
wire net_5407;
wire net_4455;
wire net_7673;
wire net_10995;
wire net_8788;
wire net_3352;
wire net_7507;
wire net_7309;
wire net_10342;
wire net_6071;
wire net_6894;
wire net_3832;
wire net_5663;
wire net_205;
wire net_11702;
wire net_1286;
wire net_6427;
wire net_15204;
wire net_6017;
wire net_10062;
wire net_15290;
wire net_11872;
wire net_9764;
wire net_7617;
wire net_7533;
wire net_6925;
wire net_334;
wire net_1952;
wire net_9214;
wire net_10930;
wire net_9846;
wire net_2453;
wire net_3062;
wire net_11495;
wire net_9586;
wire net_5738;
wire net_12512;
wire net_12629;
wire net_4620;
wire net_14141;
wire net_5696;
wire net_380;
wire net_2847;
wire net_10952;
wire net_6515;
wire net_13797;
wire net_7932;
wire net_12626;
wire net_14042;
wire net_12885;
wire net_1556;
wire net_6803;
wire net_5911;
wire net_6790;
wire net_4337;
wire net_13548;
wire net_3768;
wire net_7976;
wire net_4745;
wire net_1270;
wire net_4905;
wire net_2286;
wire net_15345;
wire net_14178;
wire net_9717;
wire net_1552;
wire x1029;
wire net_13785;
wire net_9380;
wire net_14833;
wire net_14015;
wire net_14454;
wire net_6094;
wire net_7712;
wire x2826;
wire net_14539;
wire net_4940;
wire net_3878;
wire net_5674;
wire net_14532;
wire net_14591;
wire net_7954;
wire net_8132;
wire net_5585;
wire net_3215;
wire net_298;
wire net_1933;
wire net_3717;
wire x637;
wire net_3241;
wire net_998;
wire net_12620;
wire net_4657;
wire net_2157;
wire net_8945;
wire net_7273;
wire net_15491;
wire net_2555;
wire net_10317;
wire net_4864;
wire net_11154;
wire net_13148;
wire net_12457;
wire net_9328;
wire net_3504;
wire net_13763;
wire net_14194;
wire net_2405;
wire net_14929;
wire net_1687;
wire net_835;
wire net_7459;
wire net_5243;
wire net_1762;
wire net_15381;
wire net_7407;
wire net_13683;
wire net_1181;
wire net_9321;
wire net_10685;
wire net_10466;
wire net_6459;
wire net_14795;
wire net_638;
wire net_12299;
wire x3390;
wire x3300;
wire net_7472;
wire net_932;
wire net_313;
wire net_15577;
wire net_5633;
wire net_6082;
wire net_10028;
wire net_5766;
wire net_11519;
wire net_13403;
wire net_10783;
wire net_12488;
wire net_12801;
wire net_4767;
wire net_1783;
wire net_14257;
wire net_5271;
wire net_12814;
wire net_6771;
wire net_7771;
wire net_1874;
wire net_9554;
wire net_7769;
wire net_972;
wire net_14948;
wire net_14308;
wire net_15043;
wire net_9650;
wire net_14447;
wire net_3499;
wire net_5206;
wire net_4725;
wire net_4777;
wire net_14292;
wire net_13192;
wire net_11669;
wire net_6201;
wire net_14108;
wire net_12808;
wire net_785;
wire net_7047;
wire net_9152;
wire net_1489;
wire net_13665;
wire net_5883;
wire net_4343;
wire net_4215;
wire net_10276;
wire net_9874;
wire net_6677;
wire net_10902;
wire net_13633;
wire net_10409;
wire net_9657;
wire net_7479;
wire net_3746;
wire net_1349;
wire net_7794;
wire net_7194;
wire net_979;
wire net_2392;
wire net_156;
wire net_13251;
wire net_11820;
wire net_10278;
wire net_12563;
wire net_2015;
wire net_8441;
wire net_6658;
wire net_13064;
wire net_10266;
wire net_5947;
wire net_1040;
wire net_9676;
wire net_8978;
wire net_5202;
wire net_4877;
wire x555;
wire net_6781;
wire net_4170;
wire net_3089;
wire net_3101;
wire net_12336;
wire net_6268;
wire net_3037;
wire net_4472;
wire net_12723;
wire net_7331;
wire net_4463;
wire net_3876;
wire net_5982;
wire net_2907;
wire net_3686;
wire net_1887;
wire net_13146;
wire net_7444;
wire net_15607;
wire net_5470;
wire net_14851;
wire net_379;
wire net_2243;
wire net_1569;
wire net_4033;
wire net_4245;
wire net_11868;
wire net_9514;
wire net_7795;
wire net_3133;
wire net_5568;
wire net_3047;
wire net_2559;
wire net_8910;
wire net_14451;
wire net_9532;
wire net_6944;
wire net_6883;
wire net_2657;
wire net_14475;
wire net_1358;
wire net_15119;
wire net_8477;
wire x329;
wire net_14708;
wire net_6815;
wire net_12259;
wire net_11438;
wire net_14696;
wire net_8415;
wire net_7742;
wire net_2629;
wire net_2486;
wire net_11405;
wire net_6888;
wire net_15196;
wire net_8927;
wire net_8421;
wire net_7117;
wire x277;
wire net_1206;
wire net_8381;
wire net_3653;
wire net_960;
wire net_13494;
wire x2531;
wire net_3704;
wire net_1166;
wire net_10706;
wire net_8155;
wire net_14957;
wire net_10765;
wire net_801;
wire net_11051;
wire net_2620;
wire net_14062;
wire net_7450;
wire net_1718;
wire net_2581;
wire net_5093;
wire net_12842;
wire net_13365;
wire net_9417;
wire net_7372;
wire net_13996;
wire net_9445;
wire net_6441;
wire net_4348;
wire net_4526;
wire net_11921;
wire net_10391;
wire net_15612;
wire net_8482;
wire net_2129;
wire net_7832;
wire net_5968;
wire net_6234;
wire net_15112;
wire net_9909;
wire net_8991;
wire net_581;
wire net_10564;
wire net_13967;
wire net_8799;
wire net_2899;
wire net_9833;
wire net_8856;
wire net_12421;
wire net_9609;
wire net_11382;
wire net_658;
wire net_7115;
wire net_5906;
wire net_7978;
wire net_14565;
wire net_11391;
wire net_8462;
wire net_13529;
wire net_2090;
wire net_9540;
wire net_7723;
wire net_12509;
wire net_2325;
wire net_8807;
wire net_13715;
wire net_12758;
wire net_806;
wire net_10259;
wire net_11907;
wire net_5801;
wire net_9901;
wire net_8940;
wire net_4021;
wire net_15270;
wire net_8999;
wire net_7026;
wire net_10960;
wire net_5461;
wire net_946;
wire net_1176;
wire net_2676;
wire net_14853;
wire net_6372;
wire net_7032;
wire net_4989;
wire net_2194;
wire net_11609;
wire net_1751;
wire net_13593;
wire net_5010;
wire net_3559;
wire net_8370;
wire net_4682;
wire net_6733;
wire net_15261;
wire net_10114;
wire net_3508;
wire net_10402;
wire net_12499;
wire net_10732;
wire net_2434;
wire net_3564;
wire net_1448;
wire net_2032;
wire net_392;
wire net_118;
wire net_2467;
wire net_5683;
wire net_14499;
wire net_11524;
wire net_7003;
wire net_2452;
wire net_14415;
wire net_11463;
wire net_9916;
wire net_12008;
wire net_10336;
wire net_3523;
wire net_4162;
wire net_5549;
wire net_3712;
wire net_6680;
wire net_8865;
wire net_7223;
wire net_6613;
wire net_246;
wire net_1186;
wire net_4747;
wire net_14829;
wire net_11269;
wire net_13041;
wire net_7074;
wire net_10607;
wire net_10437;
wire net_14914;
wire net_13436;
wire net_10121;
wire net_2216;
wire net_10410;
wire net_8968;
wire net_6725;
wire net_1378;
wire net_7399;
wire net_1773;
wire net_3773;
wire net_9057;
wire net_1600;
wire net_2531;
wire net_12440;
wire net_15743;
wire net_11971;
wire net_8731;
wire net_676;
wire net_11254;
wire net_12492;
wire net_6626;
wire net_15592;
wire net_4263;
wire net_5073;
wire net_2538;
wire net_4452;
wire net_2447;
wire net_7433;
wire net_5133;
wire net_5542;
wire net_14116;
wire net_5417;
wire net_15237;
wire net_5370;
wire net_4260;
wire net_3492;
wire net_8137;
wire net_14643;
wire net_6010;
wire net_182;
wire net_2462;
wire net_4359;
wire net_12760;
wire net_9635;
wire net_9018;
wire net_14506;
wire net_11260;
wire net_8820;
wire net_3324;
wire net_13485;
wire net_9547;
wire net_14872;
wire net_5426;
wire net_6450;
wire net_6138;
wire net_14237;
wire net_8398;
wire net_6979;
wire net_11442;
wire net_7893;
wire net_1435;
wire net_1370;
wire net_14463;
wire net_9600;
wire net_10429;
wire net_8112;
wire net_11274;
wire net_9462;
wire net_7939;
wire net_3568;
wire net_3207;
wire net_13920;
wire net_7810;
wire net_4482;
wire net_6470;
wire net_2204;
wire net_9668;
wire net_5088;
wire net_15485;
wire net_8459;
wire net_2492;
wire net_11188;
wire net_9088;
wire net_1970;
wire net_1306;
wire net_4045;
wire net_15228;
wire net_3843;
wire net_1858;
wire net_10223;
wire net_14551;
wire net_7635;
wire net_6543;
wire net_11005;
wire net_3038;
wire net_14846;
wire net_13560;
wire net_2690;
wire net_11332;
wire x1418;
wire net_7016;
wire net_3924;
wire net_9825;
wire net_11196;
wire net_5226;
wire net_12242;
wire net_791;
wire net_14207;
wire net_10230;
wire net_9422;
wire net_1419;
wire net_3239;
wire net_8554;
wire net_2188;
wire net_8811;
wire net_10546;
wire net_1051;
wire net_12064;
wire net_13882;
wire net_10386;
wire net_10048;
wire net_14770;
wire net_7644;
wire net_14841;
wire net_11034;
wire net_7858;
wire net_7410;
wire net_12471;
wire net_1515;
wire net_1573;
wire net_10356;
wire net_7669;
wire net_7219;
wire x454;
wire net_13272;
wire net_6869;
wire net_4983;
wire net_6824;
wire net_14651;
wire net_361;
wire net_13932;
wire net_2890;
wire net_11547;
wire net_9984;
wire net_7100;
wire net_305;
wire net_4208;
wire net_4515;
wire net_1905;
wire net_12433;
wire net_2540;
wire net_15434;
wire net_12016;
wire net_12452;
wire net_9166;
wire net_14716;
wire net_1125;
wire net_2230;
wire net_15084;
wire net_10195;
wire net_227;
wire net_144;
wire net_13758;
wire net_4183;
wire net_10667;
wire net_10237;
wire x157;
wire net_14664;
wire net_3592;
wire net_5961;
wire net_13728;
wire net_12405;
wire net_12543;
wire net_6687;
wire net_8818;
wire net_15555;
wire x233;
wire net_13592;
wire net_7156;
wire net_14413;
wire net_12636;
wire net_4969;
wire net_9175;
wire net_1415;
wire net_3485;
wire net_7052;
wire net_8859;
wire net_6379;
wire net_2886;
wire net_3317;
wire net_14408;
wire net_11746;
wire net_8140;
wire net_14934;
wire net_1921;
wire net_11638;
wire net_10945;
wire net_9161;
wire net_3853;
wire net_14781;
wire net_9962;
wire net_10120;
wire net_15462;
wire net_11910;
wire net_9091;
wire net_1230;
wire net_2135;
wire net_667;
wire net_853;
wire net_212;
wire net_12265;
wire net_9508;
wire net_6047;
wire net_914;
wire net_10254;
wire net_15418;
wire net_9923;
wire net_12835;
wire net_15245;
wire net_6862;
wire net_6320;
wire net_6064;
wire net_6448;
wire net_875;
wire x2400;
wire net_15455;
wire net_15317;
wire net_14807;
wire net_5619;
wire net_1092;
wire net_12046;
wire net_7585;
wire net_627;
wire net_10597;
wire net_8759;
wire x316;
wire net_2039;
wire net_15313;
wire net_11579;
wire net_12067;
wire net_1456;
wire net_9198;
wire net_11042;
wire net_15444;
wire net_2227;
wire net_15469;
wire net_5636;
wire net_10280;
wire net_8876;
wire net_12231;
wire net_2473;
wire net_6968;
wire net_399;
wire net_15284;
wire net_8107;
wire net_11041;
wire net_5949;
wire net_5069;
wire net_13509;
wire net_13844;
wire net_10678;
wire net_8752;
wire net_1390;
wire net_11209;
wire net_7180;
wire net_5565;
wire net_218;
wire net_12338;
wire net_10517;
wire net_7110;
wire net_1112;
wire net_9335;
wire net_5173;
wire net_1273;
wire net_3283;
wire net_10747;
wire net_15483;
wire net_9025;
wire net_4433;
wire net_13907;
wire net_11995;
wire net_8146;
wire net_5449;
wire net_2114;
wire net_2506;
wire net_11200;
wire net_12085;
wire net_5012;
wire net_9644;
wire net_3230;
wire net_13295;
wire net_7124;
wire net_14494;
wire x3621;
wire net_11235;
wire net_11990;
wire net_10187;
wire net_14073;
wire net_285;
wire net_8316;
wire net_13585;
wire net_14932;
wire net_11486;
wire net_5677;
wire net_5296;
wire net_14171;
wire net_1310;
wire net_9634;
wire net_2499;
wire net_6057;
wire net_11567;
wire net_1297;
wire net_15687;
wire net_7579;
wire net_1304;
wire net_9471;
wire net_8901;
wire net_4381;
wire net_2177;
wire net_11918;
wire net_11378;
wire net_6674;
wire net_13427;
wire net_7863;
wire net_11450;
wire net_11587;
wire net_6581;
wire net_6916;
wire net_10370;
wire net_6127;
wire net_5030;
wire net_13417;
wire net_6058;
wire net_10919;
wire net_2449;
wire net_6070;
wire net_1317;
wire net_6588;
wire net_215;
wire net_416;
wire net_2394;
wire net_1382;
wire net_5629;
wire net_11593;
wire net_13408;
wire net_15513;
wire net_6896;
wire net_6442;
wire net_15487;
wire net_4508;
wire net_14814;
wire x143;
wire net_6642;
wire net_10760;
wire net_8093;
wire net_3498;
wire net_1377;
wire net_1786;
wire net_12831;
wire net_5620;
wire net_13580;
wire net_12031;
wire net_10253;
wire x2890;
wire net_4513;
wire net_14025;
wire net_10940;
wire net_9658;
wire net_5965;
wire net_14439;
wire net_13428;
wire net_11118;
wire net_5586;
wire net_5430;
wire net_5954;
wire net_1393;
wire net_13724;
wire net_14321;
wire net_2169;
wire net_6119;
wire net_8758;
wire net_1324;
wire net_14020;
wire net_9960;
wire net_7114;
wire net_14949;
wire net_12058;
wire net_10672;
wire net_10476;
wire net_8017;
wire net_2207;
wire net_263;
wire net_6997;
wire net_9336;
wire net_4323;
wire net_8805;
wire net_1138;
wire net_3527;
wire net_8509;
wire net_14139;
wire net_3483;
wire net_6838;
wire net_10167;
wire x401;
wire net_10548;
wire net_1439;
wire net_3292;
wire net_8714;
wire net_12528;
wire net_13489;
wire net_9700;
wire net_508;
wire net_1778;
wire net_4189;
wire net_15428;
wire net_9256;
wire net_1090;
wire net_5098;
wire net_6907;
wire net_15617;
wire net_7438;
wire net_14850;
wire net_3685;
wire net_5355;
wire net_8149;
wire net_7030;
wire net_7012;
wire net_14107;
wire net_11962;
wire net_11453;
wire net_9007;
wire net_4285;
wire net_8643;
wire net_4434;
wire net_5413;
wire net_12068;
wire net_4744;
wire net_10726;
wire net_201;
wire net_5077;
wire net_9496;
wire net_6636;
wire net_3280;
wire net_9666;
wire net_3085;
wire net_4043;
wire net_2896;
wire net_14707;
wire net_8371;
wire net_4258;
wire net_7443;
wire net_12838;
wire net_12631;
wire net_12207;
wire net_12454;
wire net_13833;
wire net_9985;
wire net_1852;
wire net_11236;
wire net_11912;
wire net_9515;
wire net_6129;
wire net_1555;
wire net_7301;
wire net_10594;
wire net_2780;
wire net_9349;
wire net_4480;
wire net_789;
wire net_15454;
wire net_15240;
wire net_10131;
wire net_10769;
wire net_3244;
wire net_12819;
wire net_15153;
wire net_9041;
wire net_2171;
wire net_15282;
wire net_12080;
wire net_10233;
wire net_3833;
wire net_6338;
wire net_9967;
wire net_8664;
wire net_7256;
wire net_4521;
wire net_11245;
wire net_2425;
wire net_6112;
wire net_13691;
wire net_8319;
wire net_14870;
wire net_10573;
wire net_8143;
wire net_2509;
wire net_5137;
wire net_11569;
wire net_1860;
wire net_14587;
wire net_8025;
wire net_2156;
wire net_1432;
wire x2333;
wire net_1312;
wire net_9474;
wire net_9177;
wire net_5463;
wire net_14188;
wire net_8843;
wire net_8488;
wire net_8435;
wire net_4801;
wire net_13246;
wire net_6831;
wire net_5334;
wire net_4314;
wire net_5290;
wire net_14958;
wire net_11640;
wire net_10005;
wire net_3343;
wire net_3546;
wire net_8002;
wire net_3326;
wire net_11877;
wire net_1453;
wire net_14328;
wire net_13802;
wire net_2239;
wire net_13075;
wire net_9603;
wire net_3394;
wire net_3542;
wire net_634;
wire net_5374;
wire net_8516;
wire net_14177;
wire net_12846;
wire net_9630;
wire net_8055;
wire net_4680;
wire net_14066;
wire net_371;
wire net_15474;
wire net_13786;
wire net_3903;
wire net_7752;
wire net_15192;
wire net_2787;
wire net_8879;
wire net_4050;
wire net_1571;
wire net_11467;
wire net_9248;
wire net_2466;
wire net_4904;
wire net_8580;
wire net_4699;
wire net_7710;
wire net_7975;
wire net_5090;
wire net_8872;
wire net_10530;
wire net_7574;
wire net_13921;
wire net_850;
wire net_5217;
wire net_12511;
wire net_679;
wire net_1168;
wire net_2680;
wire net_8116;
wire net_8924;
wire net_308;
wire net_10118;
wire net_11008;
wire net_12218;
wire net_9631;
wire net_5545;
wire net_10744;
wire net_6327;
wire net_3090;
wire net_8747;
wire net_15052;
wire net_8387;
wire x19;
wire net_1009;
wire net_715;
wire net_11444;
wire net_890;
wire net_14503;
wire net_13857;
wire net_15693;
wire net_8454;
wire net_11181;
wire net_2546;
wire net_7228;
wire net_12042;
wire net_7056;
wire net_9019;
wire net_13401;
wire net_9162;
wire net_13646;
wire net_13595;
wire net_2471;
wire net_6702;
wire net_11130;
wire net_312;
wire net_2404;
wire net_2627;
wire net_5386;
wire net_147;
wire net_481;
wire net_12490;
wire net_7182;
wire net_5346;
wire x1290;
wire net_8589;
wire net_12137;
wire net_12335;
wire net_7750;
wire x1865;
wire net_2444;
wire net_6891;
wire net_11482;
wire net_13496;
wire net_1188;
wire net_13855;
wire net_12936;
wire net_8148;
wire net_5297;
wire net_9625;
wire net_1446;
wire net_10122;
wire net_541;
wire net_14965;
wire net_8551;
wire net_13380;
wire net_1251;
wire net_8157;
wire net_14148;
wire net_10759;
wire net_8830;
wire net_1697;
wire net_15748;
wire x871;
wire net_15741;
wire net_4222;
wire net_7431;
wire net_12238;
wire net_1753;
wire net_4163;
wire net_5398;
wire net_14418;
wire net_5548;
wire net_245;
wire net_2435;
wire net_6990;
wire net_2383;
wire net_4858;
wire net_14760;
wire net_14298;
wire net_12177;
wire net_4264;
wire net_11013;
wire net_9749;
wire net_3491;
wire net_10829;
wire x65;
wire net_15205;
wire net_8380;
wire net_9908;
wire net_277;
wire net_1965;
wire net_4251;
wire net_11418;
wire net_7525;
wire net_13886;
wire net_3071;
wire net_8611;
wire net_680;
wire net_14238;
wire net_10925;
wire net_9568;
wire net_13435;
wire net_13230;
wire net_338;
wire net_7149;
wire net_9994;
wire net_4494;
wire net_7619;
wire net_15672;
wire net_8397;
wire net_2998;
wire net_14597;
wire net_15549;
wire net_243;
wire net_9971;
wire net_8905;
wire net_10705;
wire net_4089;
wire net_6882;
wire net_13721;
wire net_2854;
wire net_2009;
wire net_10730;
wire net_8867;
wire net_4026;
wire net_4132;
wire net_8925;
wire net_6697;
wire net_106;
wire net_4990;
wire net_1380;
wire net_7721;
wire net_9292;
wire net_14844;
wire net_11056;
wire net_13588;
wire net_8326;
wire net_14731;
wire net_9340;
wire net_1915;
wire net_5176;
wire net_15289;
wire net_13566;
wire net_10992;
wire net_8280;
wire net_4334;
wire net_14650;
wire net_5936;
wire net_11956;
wire net_8937;
wire net_6987;
wire net_15295;
wire net_14550;
wire net_1997;
wire net_13206;
wire net_12738;
wire net_14657;
wire net_13779;
wire net_138;
wire net_12497;
wire net_7718;
wire net_14452;
wire net_13607;
wire net_8553;
wire net_6728;
wire net_15131;
wire net_13698;
wire net_13364;
wire net_11139;
wire net_9195;
wire net_12714;
wire net_14151;
wire net_7164;
wire net_12313;
wire net_6579;
wire net_14645;
wire net_9670;
wire net_15232;
wire net_14684;
wire net_14792;
wire net_7633;
wire net_1418;
wire net_13955;
wire net_8686;
wire net_13393;
wire net_5938;
wire net_8994;
wire net_3202;
wire net_13422;
wire net_8343;
wire net_4059;
wire net_5931;
wire net_6980;
wire net_6376;
wire net_6736;
wire net_7461;
wire net_15226;
wire net_15032;
wire net_12913;
wire net_1713;
wire net_15389;
wire net_10380;
wire net_5612;
wire net_2668;
wire net_4684;
wire net_13480;
wire net_11383;
wire net_2677;
wire net_15307;
wire net_8988;
wire net_14498;
wire net_15545;
wire net_10415;
wire net_2775;
wire net_14594;
wire net_7001;
wire net_11540;
wire net_12007;
wire net_11741;
wire net_14839;
wire net_3916;
wire net_7654;
wire net_163;
wire net_6852;
wire net_6022;
wire net_8312;
wire net_5802;
wire net_15736;
wire net_13937;
wire net_11037;
wire net_8037;
wire net_14466;
wire net_12590;
wire net_9830;
wire net_8444;
wire net_5900;
wire x3632;
wire net_6206;
wire net_13863;
wire net_11580;
wire net_6135;
wire net_3990;
wire net_12595;
wire net_2193;
wire net_12293;
wire net_12002;
wire net_11159;
wire net_10221;
wire net_3856;
wire net_9210;
wire x5722;
wire net_5345;
wire net_6304;
wire net_8363;
wire net_4885;
wire net_11704;
wire net_5574;
wire net_5258;
wire net_14459;
wire net_1886;
wire net_2604;
wire net_3501;
wire net_13689;
wire net_14115;
wire net_12191;
wire net_7862;
wire net_12775;
wire net_4678;
wire net_14307;
wire net_6678;
wire net_15070;
wire net_7916;
wire net_14256;
wire net_13600;
wire net_4866;
wire net_5652;
wire net_8081;
wire net_101;
wire net_15524;
wire net_13982;
wire net_14013;
wire net_8835;
wire net_1272;
wire net_1770;
wire net_2109;
wire net_10273;
wire net_3505;
wire net_4001;
wire net_5059;
wire net_655;
wire net_9326;
wire net_3536;
wire net_6878;
wire net_4703;
wire net_8534;
wire net_10059;
wire net_14530;
wire net_4770;
wire net_12961;
wire net_14049;
wire net_378;
wire net_7770;
wire net_14262;
wire net_9110;
wire net_3309;
wire net_14403;
wire net_5767;
wire net_423;
wire net_3036;
wire net_10032;
wire net_11628;
wire net_328;
wire net_4202;
wire net_10103;
wire net_10565;
wire net_1958;
wire net_7934;
wire net_7977;
wire net_1931;
wire net_15493;
wire net_9060;
wire net_14041;
wire net_3294;
wire net_1549;
wire net_6244;
wire net_10039;
wire net_3016;
wire net_4477;
wire net_7736;
wire net_2929;
wire net_7192;
wire net_12933;
wire net_9117;
wire net_7213;
wire net_5666;
wire net_11717;
wire net_11227;
wire net_8527;
wire net_818;
wire net_3749;
wire net_15103;
wire net_11275;
wire net_2746;
wire net_12592;
wire net_9403;
wire net_1211;
wire net_5024;
wire net_1183;
wire net_5448;
wire net_14574;
wire net_11863;
wire net_2594;
wire net_15574;
wire net_4248;
wire net_14537;
wire net_12337;
wire net_5944;
wire net_15436;
wire net_811;
wire net_1684;
wire net_7241;
wire net_14549;
wire net_9753;
wire net_1462;
wire net_9551;
wire net_9203;
wire net_4674;
wire net_15495;
wire net_2017;
wire net_6791;
wire net_15019;
wire net_9150;
wire net_4993;
wire net_5154;
wire net_11508;
wire net_1926;
wire net_12145;
wire net_2735;
wire net_3115;
wire net_8780;
wire net_14158;
wire net_14809;
wire net_8377;
wire net_3518;
wire net_13069;
wire net_10261;
wire net_8800;
wire net_1621;
wire net_14432;
wire net_3680;
wire net_6926;
wire net_14319;
wire net_3984;
wire net_13317;
wire net_3615;
wire net_1035;
wire net_12253;
wire net_11331;
wire net_9559;
wire net_14076;
wire net_13172;
wire net_3055;
wire net_9844;
wire net_13035;
wire net_5597;
wire x4117;
wire net_6914;
wire net_4656;
wire net_10264;
wire net_3593;
wire net_2845;
wire net_3095;
wire net_6510;
wire net_12585;
wire net_11358;
wire net_4586;
wire net_14986;
wire net_6748;
wire net_2641;
wire net_7711;
wire net_6688;
wire net_13141;
wire net_9389;
wire net_1763;
wire net_6168;
wire net_7291;
wire net_15476;
wire net_12321;
wire net_11067;
wire net_4035;
wire net_9362;
wire net_7816;
wire net_12999;
wire x374;
wire net_9881;
wire net_8948;
wire net_13464;
wire net_9092;
wire net_7919;
wire net_8131;
wire net_2882;
wire net_14440;
wire x1010;
wire net_3278;
wire net_12277;
wire x911;
wire net_4386;
wire net_8837;
wire net_1513;
wire net_14191;
wire net_15014;
wire net_14253;
wire net_10668;
wire net_3064;
wire net_5731;
wire net_12701;
wire net_2276;
wire net_12748;
wire net_4613;
wire net_6369;
wire net_9302;
wire net_11639;
wire net_7763;
wire net_7748;
wire net_11388;
wire net_9426;
wire net_6745;
wire net_10084;
wire net_13716;
wire net_14149;
wire net_798;
wire net_14820;
wire net_3135;
wire net_5266;
wire net_5165;
wire net_2059;
wire net_8473;
wire net_9740;
wire net_8520;
wire net_8860;
wire net_8209;
wire net_1899;
wire net_6018;
wire net_15715;
wire x2767;
wire net_8890;
wire net_1336;
wire net_4746;
wire net_12198;
wire net_9915;
wire net_10033;
wire net_1843;
wire net_6031;
wire net_11739;
wire net_6946;
wire net_12211;
wire net_7019;
wire net_534;
wire net_14114;
wire net_11534;
wire net_3793;
wire net_9261;
wire net_13523;
wire net_11671;
wire net_8659;
wire net_6823;
wire net_3336;
wire net_15502;
wire net_9561;
wire net_903;
wire net_1551;
wire net_14951;
wire net_10025;
wire net_12069;
wire net_486;
wire net_14753;
wire net_13796;
wire net_12898;
wire net_406;
wire net_11395;
wire net_8407;
wire net_7354;
wire net_5986;
wire net_4190;
wire net_2378;
wire net_5391;
wire net_12448;
wire net_11758;
wire net_10461;
wire net_6261;
wire net_8967;
wire net_10319;
wire net_15186;
wire net_8046;
wire net_15378;
wire net_13746;
wire net_7125;
wire net_3640;
wire x941;
wire net_748;
wire net_9865;
wire net_8605;
wire net_95;
wire net_14445;
wire net_10587;
wire net_10010;
wire net_5566;
wire net_6917;
wire net_13124;
wire net_10778;
wire net_3958;
wire net_5281;
wire net_12270;
wire net_8776;
wire net_5427;
wire net_15259;
wire net_11621;
wire net_11684;
wire net_14902;
wire net_10868;
wire net_8772;
wire net_1003;
wire net_2327;
wire net_514;
wire net_15443;
wire net_11255;
wire net_3645;
wire net_7376;
wire net_10310;
wire net_1604;
wire net_6499;
wire net_5755;
wire net_14093;
wire net_5669;
wire net_6122;
wire net_524;
wire net_6497;
wire net_13387;
wire net_11991;
wire net_6060;
wire net_13816;
wire net_13554;
wire net_11513;
wire net_3742;
wire net_445;
wire net_4368;
wire net_7109;
wire net_13398;
wire net_13002;
wire net_10773;
wire net_6673;
wire net_3748;
wire net_12319;
wire net_15164;
wire net_13637;
wire net_10786;
wire net_9355;
wire net_8307;
wire net_2213;
wire net_14789;
wire net_12083;
wire net_2575;
wire net_5067;
wire net_11986;
wire net_10935;
wire x3565;
wire net_1097;
wire net_11756;
wire net_12227;
wire net_14172;
wire net_9219;
wire net_12142;
wire net_762;
wire net_6921;
wire net_3589;
wire net_8445;
wire net_13517;
wire net_4943;
wire net_10876;
wire net_3713;
wire net_8400;
wire net_556;
wire net_6173;
wire net_893;
wire net_3330;
wire net_11163;
wire net_4121;
wire net_255;
wire net_3826;
wire net_620;
wire net_9641;
wire net_619;
wire x6282;
wire net_13618;
wire net_9085;
wire net_8702;
wire net_4659;
wire net_7321;
wire net_14529;
wire net_3932;
wire net_7233;
wire net_14392;
wire net_11177;
wire net_4779;
wire net_5997;
wire net_11150;
wire net_7689;
wire net_14802;
wire net_8156;
wire net_5129;
wire net_7104;
wire net_14909;
wire net_10444;
wire net_7883;
wire net_3444;
wire net_4922;
wire net_6414;
wire net_3800;
wire net_5393;
wire net_3285;
wire net_6937;
wire net_7278;
wire net_7825;
wire net_4425;
wire net_4933;
wire net_5834;
wire net_4044;
wire net_13613;
wire net_14862;
wire net_8855;
wire net_11300;
wire net_1493;
wire net_9167;
wire x3327;
wire net_13285;
wire net_11699;
wire net_5875;
wire net_4630;
wire net_15636;
wire net_11143;
wire net_976;
wire net_6287;
wire net_8498;
wire net_2709;
wire net_5309;
wire net_10321;
wire net_11630;
wire net_8897;
wire net_611;
wire net_7879;
wire net_2579;
wire net_3514;
wire net_4179;
wire net_5441;
wire net_8235;
wire net_9581;
wire net_10296;
wire net_6013;
wire net_7307;
wire net_5873;
wire net_12990;
wire net_1866;
wire net_6077;
wire net_14852;
wire net_10849;
wire net_4907;
wire net_6567;
wire net_4107;
wire net_6934;
wire net_5761;
wire net_2160;
wire net_3211;
wire net_3692;
wire net_13060;
wire net_10820;
wire net_3477;
wire net_391;
wire net_6361;
wire net_9268;
wire net_9723;
wire net_5927;
wire net_7634;
wire net_5040;
wire net_13894;
wire net_11738;
wire net_12754;
wire net_8625;
wire net_5820;
wire net_6692;
wire net_4172;
wire net_11732;
wire net_8342;
wire x6496;
wire net_2516;
wire net_13892;
wire net_8123;
wire net_2807;
wire net_7553;
wire net_12417;
wire net_10676;
wire net_4687;
wire net_1141;
wire net_6253;
wire net_10621;
wire net_3243;
wire net_4867;
wire net_6321;
wire net_7871;
wire net_7584;
wire net_2104;
wire net_5564;
wire net_1288;
wire net_6190;
wire net_4708;
wire net_12554;
wire net_10511;
wire net_2766;
wire net_10559;
wire net_3771;
wire net_12469;
wire net_8119;
wire net_2300;
wire net_2417;
wire net_6710;
wire net_14406;
wire net_8426;
wire net_741;
wire net_7091;
wire net_13915;
wire net_6383;
wire net_4816;
wire net_5509;
wire net_6434;
wire net_11428;
wire net_15092;
wire net_6472;
wire net_7853;
wire net_13765;
wire net_11604;
wire net_3789;
wire net_15664;
wire net_13288;
wire net_5524;
wire net_9598;
wire net_4937;
wire net_11947;
wire net_4199;
wire net_11897;
wire net_1043;
wire net_12977;
wire net_15086;
wire net_2850;
wire net_770;
wire net_13905;
wire net_12901;
wire net_1005;
wire x1598;
wire net_15711;
wire net_9737;
wire net_11792;
wire net_11198;
wire net_6389;
wire net_7493;
wire net_1059;
wire net_1630;
wire net_3891;
wire net_4918;
wire net_2956;
wire net_1082;
wire net_1796;
wire net_10328;
wire net_15645;
wire net_11170;
wire net_10405;
wire net_5187;
wire net_15407;
wire net_7501;
wire net_11368;
wire net_11291;
wire net_11861;
wire net_1507;
wire net_2310;
wire net_257;
wire net_3296;
wire net_11407;
wire net_10096;
wire net_8543;
wire net_7466;
wire net_9978;
wire net_474;
wire net_5500;
wire net_5770;
wire net_12518;
wire net_6576;
wire net_11421;
wire net_958;
wire net_12646;
wire net_11934;
wire net_11940;
wire net_4556;
wire net_6400;
wire net_7947;
wire net_11855;
wire net_11447;
wire net_12244;
wire net_12407;
wire net_944;
wire net_6199;
wire net_1734;
wire net_10189;
wire net_10008;
wire net_11175;
wire net_4308;
wire net_5534;
wire net_13477;
wire net_12538;
wire net_10987;
wire net_11002;
wire net_7199;
wire x5364;
wire net_14510;
wire net_13450;
wire net_7166;
wire net_12580;
wire net_1728;
wire net_3050;
wire net_12883;
wire net_5963;
wire net_15394;
wire net_3956;
wire net_15709;
wire net_12426;
wire net_10218;
wire net_8761;
wire net_8467;
wire net_13669;
wire net_425;
wire net_12028;
wire net_287;
wire net_189;
wire net_5204;
wire net_10414;
wire net_9893;
wire net_9860;
wire net_2205;
wire net_3755;
wire net_6036;
wire net_13154;
wire net_433;
wire net_11709;
wire net_8108;
wire net_8296;
wire net_4443;
wire net_11344;
wire net_13667;
wire net_8064;
wire net_368;
wire net_224;
wire net_4833;
wire net_1898;
wire net_10670;
wire net_9073;
wire net_608;
wire net_1212;
wire net_3604;
wire net_2000;
wire net_13089;
wire net_4383;
wire net_5331;
wire net_14799;
wire net_6226;
wire net_12502;
wire net_13194;
wire net_3706;
wire net_10603;
wire net_1020;
wire net_2984;
wire net_7062;
wire net_12879;
wire net_3282;
wire net_11997;
wire net_8299;
wire net_3122;
wire net_13989;
wire net_8546;
wire net_12832;
wire net_10164;
wire net_10763;
wire net_12521;
wire net_8594;
wire net_11965;
wire net_2094;
wire net_6416;
wire net_2543;
wire net_7282;
wire net_8275;
wire net_13227;
wire net_760;
wire net_2083;
wire net_12050;
wire net_8318;
wire net_873;
wire net_3851;
wire net_1811;
wire net_2488;
wire net_13884;
wire net_4536;
wire net_12374;
wire net_11080;
wire net_5034;
wire net_2588;
wire net_8192;
wire net_7802;
wire net_1870;
wire net_5200;
wire net_9771;
wire net_704;
wire net_12772;
wire net_12906;
wire net_2063;
wire net_3997;
wire net_192;
wire net_1356;
wire net_1739;
wire net_14542;
wire net_2912;
wire net_8913;
wire net_4140;
wire net_4393;
wire net_6541;
wire net_3816;
wire net_6101;
wire net_13254;
wire net_13457;
wire net_735;
wire net_14269;
wire net_5539;
wire net_9056;
wire net_1711;
wire net_3809;
wire net_14527;
wire net_2084;
wire net_8186;
wire net_11590;
wire net_9442;
wire net_9530;
wire net_1081;
wire net_5085;
wire net_7031;
wire net_2037;
wire net_8163;
wire net_7349;
wire net_1237;
wire net_12478;
wire net_1420;
wire net_4789;
wire net_12653;
wire net_9112;
wire net_8680;
wire net_14921;
wire net_4836;
wire net_9587;
wire net_4064;
wire net_9712;
wire net_4237;
wire net_9602;
wire net_9542;
wire net_4559;
wire net_15265;
wire net_11663;
wire net_699;
wire net_3144;
wire net_7782;
wire net_7270;
wire net_359;
wire net_9283;
wire net_12892;
wire net_5239;
wire net_2526;
wire net_9414;
wire net_9068;
wire net_12862;
wire net_7338;
wire net_11316;
wire net_1644;
wire net_2819;
wire net_5827;
wire net_12126;
wire net_882;
wire net_2800;
wire net_14225;
wire net_7940;
wire net_15614;
wire net_1827;
wire net_6433;
wire net_14867;
wire net_8255;
wire x1153;
wire net_12606;
wire net_1190;
wire net_3225;
wire net_4109;
wire net_8903;
wire net_3858;
wire net_14182;
wire net_10813;
wire net_7838;
wire net_4093;
wire net_6449;
wire net_15535;
wire net_4799;
wire net_13812;
wire net_8721;
wire net_15254;
wire net_12021;
wire net_1207;
wire net_2283;
wire net_10436;
wire net_9829;
wire net_6066;
wire net_15140;
wire net_8228;
wire net_2121;
wire net_2191;
wire net_14698;
wire net_14326;
wire net_13318;
wire net_14671;
wire net_13304;
wire net_2252;
wire net_10690;
wire net_4755;
wire net_15077;
wire net_13168;
wire net_12617;
wire net_7951;
wire net_15639;
wire net_12416;
wire net_12352;
wire net_14249;
wire net_2126;
wire net_5022;
wire net_1577;
wire net_1054;
wire net_4595;
wire net_10449;
wire net_9931;
wire net_7342;
wire net_9524;
wire net_2727;
wire net_12461;
wire net_14616;
wire net_5605;
wire net_2257;
wire net_6952;
wire net_10640;
wire net_14741;
wire net_3418;
wire net_3655;
wire net_2304;
wire net_5491;
wire net_14098;
wire net_13217;
wire net_12044;
wire net_2968;
wire net_7314;
wire net_12942;
wire net_10649;
wire net_5989;
wire net_12339;
wire net_7418;
wire net_1593;
wire net_2643;
wire net_5845;
wire net_8918;
wire net_10397;
wire net_9591;
wire net_3380;
wire net_3722;
wire net_15272;
wire net_12794;
wire net_14758;
wire net_11117;
wire net_11762;
wire net_1517;
wire net_14682;
wire net_5115;
wire net_4502;
wire net_15658;
wire x480;
wire net_12275;
wire net_11218;
wire net_5980;
wire net_13131;
wire net_12567;
wire net_2076;
wire net_2218;
wire net_4378;
wire net_6505;
wire net_6705;
wire net_9192;
wire net_6807;
wire net_15217;
wire net_10147;
wire net_1690;
wire net_15219;
wire net_9811;
wire net_1078;
wire net_12340;
wire net_9853;
wire net_14984;
wire net_11924;
wire net_2093;
wire net_2997;
wire net_6813;
wire net_14831;
wire net_6382;
wire net_15027;
wire net_14896;
wire net_5681;
wire net_13126;
wire net_14186;
wire net_10635;
wire net_9076;
wire net_7239;
wire net_14341;
wire net_12269;
wire net_11787;
wire net_5197;
wire net_15099;
wire net_12703;
wire net_13059;
wire net_12856;
wire net_2355;
wire net_13825;
wire net_9549;
wire net_4357;
wire net_3262;
wire net_139;
wire net_2536;
wire x798;
wire net_5890;
wire net_7968;
wire net_2949;
wire net_3429;
wire net_10954;
wire net_9032;
wire net_4495;
wire net_12587;
wire net_1708;
wire net_12398;
wire net_5519;
wire net_12824;
wire net_7454;
wire net_4196;
wire net_13678;
wire net_3974;
wire net_13112;
wire net_4626;
wire net_12575;
wire net_13050;
wire net_8532;
wire net_8478;
wire net_15007;
wire net_722;
wire net_2976;
wire net_13138;
wire net_5420;
wire net_12094;
wire net_988;
wire net_8221;
wire net_14612;
wire net_13099;
wire net_3621;
wire net_5798;
wire net_11351;
wire net_14313;
wire net_5223;
wire net_12441;
wire net_9820;
wire net_8216;
wire net_435;
wire net_12077;
wire net_1830;
wire net_4091;
wire net_12110;
wire net_132;
wire net_2838;
wire net_5156;
wire net_6481;
wire net_1649;
wire net_6603;
wire net_1837;
wire net_1841;
wire net_5219;
wire net_5614;
wire net_6973;
wire net_1249;
wire net_2427;
wire net_4601;
wire net_8075;
wire net_1071;
wire net_3378;
wire net_7973;
wire net_3163;
wire net_4928;
wire net_5004;
wire net_5817;
wire net_6221;
wire net_9776;
wire net_1701;
wire net_4417;
wire net_5675;
wire net_11156;
wire net_822;
wire net_7145;
wire net_14007;
wire net_8678;
wire net_12175;
wire net_1633;
wire net_7084;
wire net_15369;
wire net_11132;
wire net_15523;
wire net_12150;
wire net_6561;
wire net_13470;
wire net_5251;
wire net_15691;
wire net_6842;
wire net_8694;
wire net_1974;
wire net_7701;
wire net_319;
wire net_8010;
wire net_2670;
wire net_4963;
wire net_1743;
wire net_2597;
wire net_5913;
wire net_11480;
wire net_9996;
wire net_9021;
wire net_1544;
wire net_7640;
wire net_11887;
wire net_7366;
wire net_4400;
wire net_10044;
wire net_4139;
wire net_15572;
wire net_2923;
wire x182;
wire net_10340;
wire net_7545;
wire net_512;
wire net_7929;
wire net_1174;
wire net_15168;
wire net_1109;
wire net_6664;
wire net_6731;
wire net_12326;
wire net_3102;
wire net_4224;
wire net_7510;
wire net_13733;
wire net_13513;
wire net_9683;
wire net_3457;
wire net_5780;
wire net_5721;
wire net_10963;
wire net_7904;
wire net_13119;
wire net_11721;
wire net_5276;
wire net_1102;
wire net_4471;
wire net_13644;
wire net_5487;
wire net_4976;
wire net_5640;
wire net_5245;
wire net_11205;
wire net_3371;
wire net_5317;
wire net_14175;
wire net_13953;
wire net_2692;
wire net_6800;
wire net_9375;
wire net_3777;
wire net_12673;
wire net_11322;
wire net_15212;
wire net_1875;
wire net_14355;
wire net_5862;
wire net_3420;
wire net_13353;
wire net_10285;
wire net_14382;
wire net_3887;
wire net_6279;
wire net_7050;
wire net_7516;
wire net_1487;
wire net_7037;
wire net_4572;
wire net_10020;
wire net_2759;
wire net_7484;
wire net_13373;
wire net_5408;
wire net_8243;
wire net_15045;
wire net_14128;
wire net_12486;
wire net_3634;
wire net_12189;
wire net_8736;
wire net_13348;
wire net_12953;
wire net_5178;
wire net_7678;
wire net_2835;
wire net_4543;
wire net_13705;
wire net_4871;
wire net_6599;
wire net_14215;
wire net_1240;
wire net_9213;
wire net_3000;
wire net_12200;
wire net_10338;
wire net_15002;
wire net_10349;
wire net_2564;
wire net_2821;
wire net_12674;
wire net_1658;
wire net_13048;
wire net_5481;
wire net_5688;
wire net_858;
wire net_7318;
wire net_3007;
wire net_9505;
wire net_9338;
wire net_7554;
wire net_4487;
wire net_15412;
wire net_15583;
wire net_14998;
wire net_8986;
wire net_4766;
wire net_9122;
wire x1170;
wire net_3174;
wire net_6004;
wire net_2876;
wire net_6966;
wire net_8504;
wire net_844;
wire net_13549;
wire net_1496;
wire net_9867;
wire net_14470;
wire net_325;
wire net_7995;
wire net_3735;
wire net_1820;
wire net_10870;
wire net_11422;
wire net_14628;
wire net_8175;
wire net_1427;
wire net_5123;
wire net_3921;
wire net_5690;
wire net_7075;
wire net_13274;
wire net_5899;
wire net_4098;
wire net_5478;
wire net_7251;
wire net_10287;
wire net_5956;
wire net_12106;
wire x46;
wire net_9827;
wire net_5014;
wire net_11029;
wire net_4036;
wire net_7517;
wire net_11266;
wire net_14762;
wire net_1521;
wire net_4182;
wire net_6274;
wire net_10308;
wire net_6020;
wire net_7172;
wire net_1677;
wire net_11813;
wire net_7908;
wire net_11727;
wire net_4734;
wire net_7179;
wire net_2991;
wire net_14919;
wire net_13260;
wire net_10077;
wire net_564;
wire net_4276;
wire net_6154;
wire net_10618;
wire net_2050;
wire net_4086;
wire net_13992;
wire net_9082;
wire net_7089;
wire net_2811;
wire net_6788;
wire net_813;
wire net_14105;
wire net_10661;
wire net_5609;
wire net_15279;
wire net_1027;
wire net_2612;
wire net_8791;
wire net_5230;
wire net_2042;
wire net_12403;
wire net_1408;
wire net_265;
wire net_7189;
wire net_13626;
wire net_11649;
wire net_8110;
wire net_6649;
wire net_11720;
wire net_10949;
wire net_3488;
wire net_8673;
wire net_3023;
wire net_13538;
wire net_11097;
wire net_6774;
wire net_5584;
wire net_10834;
wire net_1202;
wire net_14373;
wire net_9351;
wire net_14606;
wire net_10890;
wire net_9258;
wire net_1155;
wire net_925;
wire net_4932;
wire net_6776;
wire net_7452;
wire net_9787;
wire net_12827;
wire net_5384;
wire net_7374;
wire net_15680;
wire net_12764;
wire net_11317;
wire net_10974;
wire net_12074;
wire net_4661;
wire net_2695;
wire net_10331;
wire net_864;
wire net_10196;
wire net_11054;
wire net_14337;
wire net_13336;
wire net_7691;
wire net_13004;
wire net_12851;
wire net_12611;
wire net_7404;
wire net_12787;
wire net_8564;
wire net_12285;
wire net_7783;
wire net_14477;
wire net_4113;
wire net_14992;
wire net_8850;
wire net_10365;
wire net_6284;
wire net_660;
wire net_2298;
wire net_14060;
wire net_9436;
wire net_7132;
wire net_9707;
wire net_2313;
wire net_11655;
wire net_6580;
wire net_9044;
wire net_1908;
wire net_6172;
wire net_7595;
wire net_7647;
wire net_230;
wire net_4214;
wire net_9309;
wire net_3383;
wire net_13020;
wire net_12958;
wire net_6985;
wire net_7265;
wire net_3349;
wire net_4782;
wire net_6751;
wire net_1222;
wire net_3404;
wire net_14080;
wire net_14291;
wire net_3810;
wire net_14560;
wire net_9172;
wire net_3914;
wire net_7607;
wire net_12018;
wire net_6531;
wire net_15689;
wire net_14104;
wire net_6463;
wire net_11973;
wire net_4739;
wire net_6455;
wire net_4156;
wire net_10610;
wire net_5777;
wire net_8823;
wire net_12685;
wire net_13449;
wire net_7576;
wire net_13693;
wire net_12459;
wire net_3440;
wire net_6904;
wire net_3358;
wire net_1776;
wire net_2145;
wire net_6488;
wire net_11109;
wire net_3368;
wire net_5747;
wire net_3311;
wire net_4014;
wire net_14723;
wire net_15626;
wire net_8874;
wire net_11020;
wire net_14036;
wire net_12729;
wire net_10887;
wire net_7204;
wire net_10454;
wire net_2132;
wire net_2292;
wire net_15310;
wire net_9313;
wire net_12367;
wire net_1880;
wire net_10716;
wire net_3862;
wire net_184;
wire net_5103;
wire net_13943;
wire net_4853;
wire net_14775;
wire net_8699;
wire net_5855;
wire net_10757;
wire net_14087;
wire net_11247;
wire net_10427;
wire net_15359;
wire net_10474;
wire net_7203;
wire net_13080;
wire net_11507;
wire net_3538;
wire net_1867;
wire net_9498;
wire net_8205;
wire net_1949;
wire net_2650;
wire net_13568;
wire net_10455;
wire net_1583;
wire net_15564;
wire net_1804;
wire net_9454;
wire net_2331;
wire net_14520;
wire net_4408;
wire net_6667;
wire net_1563;
wire net_4291;
wire net_3898;
wire net_13969;
wire net_12389;
wire net_4948;
wire net_8637;
wire net_7600;
wire net_14483;
wire net_13073;
wire net_5599;
wire net_3361;
wire net_1135;
wire net_1365;
wire net_13019;
wire net_11674;
wire net_10553;
wire net_1346;
wire net_5047;
wire net_14285;
wire net_8578;
wire net_1942;
wire net_11484;
wire net_11478;
wire net_13865;
wire net_10070;
wire net_13835;
wire net_9220;
wire net_12119;
wire net_9277;
wire net_1801;
wire net_13755;
wire net_7891;
wire net_15650;
wire net_14150;
wire net_1267;
wire net_14364;
wire net_6093;
wire net_12570;
wire net_11846;
wire net_3661;
wire net_3944;
wire net_9188;
wire net_4350;
wire net_6029;
wire net_4893;
wire net_12982;
wire net_8955;
wire net_15724;
wire net_669;
wire net_6526;
wire net_937;
wire net_11252;
wire net_10179;
wire net_5888;
wire net_8452;
wire net_9575;
wire net_8030;
wire net_5131;
wire net_2349;
wire net_479;
wire net_11074;
wire net_8740;
wire net_12769;
wire net_1294;
wire net_10350;
wire net_6086;
wire net_14692;
wire net_14450;
wire net_2030;
wire net_1587;
wire net_3520;
wire net_5006;
wire net_13232;
wire net_1354;
wire net_11025;
wire net_15480;
wire net_1308;
wire net_796;
wire net_2904;
wire net_7631;
wire net_12081;
wire net_4332;
wire net_9992;
wire net_1389;
wire net_648;
wire net_11901;
wire net_12114;
wire net_6884;
wire net_12040;
wire net_8150;
wire net_13818;
wire net_4748;
wire net_14300;
wire net_3250;
wire net_14443;
wire net_7054;
wire net_11950;
wire net_7625;
wire net_5304;
wire net_3658;
wire net_10737;
wire net_548;
wire net_12560;
wire net_2402;
wire net_4985;
wire net_6529;
wire net_14146;
wire net_5902;
wire net_6964;
wire net_9148;
wire net_5082;
wire net_15414;
wire net_636;
wire net_10239;
wire net_4269;
wire net_8237;
wire net_8159;
wire net_8556;
wire net_7649;
wire net_12179;
wire net_10739;
wire net_10232;
wire net_8725;
wire net_8471;
wire net_8218;
wire net_4492;
wire net_6700;
wire net_14655;
wire net_1961;
wire net_10831;
wire net_1260;
wire net_12678;
wire net_10124;
wire net_4165;
wire net_4262;
wire net_9832;
wire net_10228;
wire net_1185;
wire net_4506;
wire net_13868;
wire net_5001;
wire net_15375;
wire net_239;
wire net_13396;
wire net_310;
wire net_14599;
wire net_11216;
wire net_10367;
wire net_2437;
wire net_7942;
wire net_10792;
wire net_9401;
wire net_14772;
wire net_8982;
wire net_9917;
wire net_4826;
wire net_1912;
wire net_13498;
wire net_9566;
wire net_11353;
wire net_11263;
wire net_5886;
wire net_14960;
wire net_11416;
wire net_9118;
wire net_11542;
wire net_13711;
wire net_9906;
wire net_682;
wire net_15746;
wire net_1963;
wire net_7122;
wire net_15721;
wire net_1538;
wire net_108;
wire net_14228;
wire net_13558;
wire net_9501;
wire net_12049;
wire net_11499;
wire net_8989;
wire net_13965;
wire net_3560;
wire net_5804;
wire net_1007;
wire net_15497;
wire net_1579;
wire net_7000;
wire net_14837;
wire net_13440;
wire net_4772;
wire net_7007;
wire net_11415;
wire net_1292;
wire net_7197;
wire net_10703;
wire net_10520;
wire net_6484;
wire net_7861;
wire net_10771;
wire net_12262;
wire net_1999;
wire net_1014;
wire net_6669;
wire net_11039;
wire net_1444;
wire net_2796;
wire net_11400;
wire net_2679;
wire net_5016;
wire net_4024;
wire net_6255;
wire net_4082;
wire net_6699;
wire x4359;
wire net_14666;
wire net_11577;
wire net_9544;
wire net_14864;
wire net_14746;
wire net_9083;
wire net_538;
wire net_12994;
wire net_12443;
wire net_4130;
wire net_6280;
wire net_8043;
wire net_1937;
wire net_15114;
wire net_13306;
wire net_9965;
wire net_7215;
wire net_366;
wire net_1854;
wire net_1956;
wire net_11339;
wire net_1917;
wire net_13433;
wire net_1614;
wire net_1755;
wire net_13491;
wire net_12911;
wire net_1359;
wire x427;
wire net_11958;
wire net_7119;
wire net_2460;
wire x1240;
wire net_13228;
wire net_8929;
wire net_10255;
wire net_3209;
wire net_12791;
wire net_14704;
wire net_11238;
wire net_4891;
wire net_15547;
wire net_8688;
wire net_13424;
wire net_11348;
wire net_10874;
wire net_8412;
wire net_14496;
wire net_12618;
wire net_209;
wire net_9242;
wire net_1282;
wire net_7716;
wire net_294;
wire net_15305;
wire net_8211;
wire net_13291;
wire net_9837;
wire net_4041;
wire net_10797;
wire net_2429;
wire net_9217;
wire net_1265;
wire net_3204;
wire net_10822;
wire net_8996;
wire net_6224;
wire net_14694;
wire net_8697;
wire net_11203;
wire net_12315;
wire net_3471;
wire net_9677;
wire net_12984;
wire net_8039;
wire net_1619;
wire net_5468;
wire net_12727;
wire net_2124;
wire net_5934;
wire net_9692;
wire net_12354;
wire net_12966;
wire net_15247;
wire net_1161;
wire net_3512;
wire net_7070;
wire net_4671;
wire net_15387;
wire net_13606;
wire net_12695;
wire net_8907;
wire net_7663;
wire net_11531;
wire net_9394;
wire net_11385;
wire net_10382;
wire net_10177;
wire net_2430;
wire net_10721;
wire net_8433;
wire net_4461;
wire net_7687;
wire net_13598;
wire net_8500;
wire net_1395;
wire net_11942;
wire net_3481;
wire net_8877;
wire net_9360;
wire net_1589;
wire net_14979;
wire net_15005;
wire net_11875;
wire net_8114;
wire net_14678;
wire net_5353;
wire net_2396;
wire net_9098;
wire net_8756;
wire net_5270;
wire net_9921;
wire net_15489;
wire net_13298;
wire net_12456;
wire net_8354;
wire net_2445;
wire net_5815;
wire net_3396;
wire net_6640;
wire net_2856;
wire net_5324;
wire net_15452;
wire net_10592;
wire net_787;
wire net_10789;
wire net_7777;
wire net_8125;
wire net_3603;
wire net_4511;
wire net_7395;
wire net_13419;
wire net_9656;
wire net_2894;
wire net_15643;
wire net_4187;
wire net_8095;
wire net_13714;
wire net_6999;
wire net_1988;
wire net_7388;
wire net_12071;
wire net_14323;
wire net_3718;
wire net_11001;
wire net_8463;
wire net_4419;
wire net_6195;
wire net_15619;
wire net_10767;
wire x1104;
wire net_3579;
wire net_5284;
wire net_11125;
wire net_3525;
wire net_10696;
wire net_11069;
wire net_6850;
wire net_13508;
wire net_8870;
wire net_15638;
wire net_1608;
wire net_2139;
wire net_506;
wire net_5332;
wire net_3769;
wire net_12802;
wire net_8019;
wire net_10250;
wire net_9330;
wire net_12836;
wire net_1910;
wire net_3775;
wire net_8278;
wire net_8103;
wire net_14891;
wire net_12689;
wire net_5432;
wire net_6586;
wire net_3544;
wire net_9517;
wire net_3034;
wire net_5229;
wire net_9488;
wire net_5096;
wire net_7895;
wire net_7938;
wire net_6285;
wire net_7610;
wire net_12817;
wire net_11030;
wire net_9664;
wire net_2493;
wire net_11914;
wire net_919;
wire net_9009;
wire net_7589;
wire net_12055;
wire net_11574;
wire net_6909;
wire net_290;
wire net_6476;
wire net_7044;
wire net_13676;
wire net_6315;
wire net_6836;
wire net_10913;
wire net_3313;
wire net_4008;
wire net_6444;
wire net_12669;
wire net_15280;
wire net_9987;
wire net_2209;
wire net_1372;
wire net_8803;
wire net_11935;
wire net_1757;
wire net_5769;
wire net_3591;
wire net_15601;
wire net_5729;
wire net_13341;
wire net_8816;
wire net_5215;
wire net_15025;
wire net_13084;
wire net_13015;
wire net_11926;
wire net_14547;
wire net_12430;
wire net_4436;
wire net_2682;
wire net_14936;
wire net_7151;
wire net_8053;
wire net_140;
wire net_14562;
wire net_11949;
wire net_2329;
wire net_6612;
wire net_8911;
wire net_7077;
wire net_2150;
wire net_3790;
wire net_7129;
wire net_9141;
wire net_2065;
wire net_15235;
wire net_10003;
wire net_13244;
wire net_10030;
wire net_15275;
wire net_4267;
wire net_8373;
wire net_2927;
wire net_12482;
wire net_7397;
wire net_7328;
wire net_11831;
wire net_11838;
wire net_194;
wire net_4856;
wire net_2178;
wire net_13941;
wire net_11264;
wire net_9448;
wire net_5292;
wire net_1128;
wire net_10134;
wire net_3073;
wire net_2713;
wire net_13161;
wire net_11582;
wire net_15354;
wire net_12539;
wire net_11320;
wire net_8840;
wire net_13846;
wire net_7949;
wire net_804;
wire net_10541;
wire net_1119;
wire net_9637;
wire net_3548;
wire net_1314;
wire net_9400;
wire net_4312;
wire net_8845;
wire net_6325;
wire net_5376;
wire net_531;
wire net_5299;
wire net_8582;
wire net_499;
wire net_8852;
wire net_3345;
wire net_2752;
wire net_10125;
wire net_7855;
wire net_11642;
wire net_11006;
wire net_9126;
wire net_7127;
wire net_7448;
wire net_10701;
wire net_11900;
wire net_9699;
wire net_9476;
wire net_10742;
wire net_3328;
wire net_13413;
wire net_8027;
wire net_3534;
wire net_4390;
wire net_12155;
wire net_1765;
wire net_14812;
wire net_8965;
wire net_10174;
wire x1142;
wire net_2107;
wire net_10424;
wire net_14878;
wire net_180;
wire net_11231;
wire net_6208;
wire net_13462;
wire x6198;
wire net_6859;
wire net_2420;
wire net_2774;
wire net_6068;
wire net_12437;
wire net_5657;
wire net_13410;
wire net_4367;
wire net_1979;
wire net_5135;
wire net_13927;
wire net_3290;
wire net_3731;
wire net_1475;
wire net_1460;
wire net_10241;
wire net_1451;
wire net_14112;
wire net_13978;
wire net_12246;
wire net_10601;
wire net_5446;
wire net_5008;
wire net_5065;
wire net_8419;
wire net_6619;
wire net_12719;
wire net_4803;
wire net_14667;
wire net_15682;
wire net_203;
wire net_2173;
wire net_9053;
wire net_6865;
wire net_6597;
wire net_7539;
wire net_14589;
wire net_11071;
wire net_1602;
wire net_12213;
wire net_14785;
wire net_6263;
wire net_5590;
wire net_9919;
wire net_613;
wire net_237;
wire net_13239;
wire net_11673;
wire net_14334;
wire net_5476;
wire net_14236;
wire net_3744;
wire net_11851;
wire x3314;
wire net_4635;
wire net_1095;
wire net_14912;
wire net_12193;
wire net_578;
wire net_4729;
wire net_15467;
wire net_12236;
wire net_15460;
wire net_6570;
wire net_14787;
wire net_8309;
wire net_11288;
wire net_15360;
wire net_8514;
wire net_6939;
wire net_12968;
wire net_4485;
wire x3534;
wire net_1558;
wire net_14881;
wire net_2743;
wire net_8603;
wire net_4641;
wire net_10958;
wire net_388;
wire net_2159;
wire x1262;
wire net_10806;
wire net_14360;
wire net_3647;
wire net_14138;
wire net_536;
wire net_455;
wire net_11515;
wire net_1332;
wire net_10294;
wire net_115;
wire net_7498;
wire net_10589;
wire net_3276;
wire net_3339;
wire net_393;
wire net_6303;
wire net_11980;
wire net_9428;
wire net_13525;
wire net_7352;
wire net_7468;
wire net_9130;
wire net_408;
wire net_1832;
wire net_12474;
wire net_12622;
wire net_10904;
wire net_1026;
wire net_15207;
wire net_10582;
wire net_2215;
wire net_3246;
wire net_15376;
wire net_1845;
wire net_6453;
wire net_2573;
wire net_10633;
wire net_12225;
wire net_9369;
wire net_9939;
wire net_10312;
wire net_7378;
wire net_15438;
wire net_3390;
wire net_3993;
wire net_15446;
wire net_13673;
wire net_1401;
wire net_2372;
wire net_12579;
wire net_3909;
wire net_12870;
wire net_868;
wire net_11858;
wire net_11223;
wire net_10979;
wire net_7889;
wire net_14394;
wire net_7248;
wire x987;
wire net_6079;
wire net_13311;
wire net_6821;
wire net_13750;
wire net_443;
wire net_5029;
wire net_13871;
wire net_6367;
wire net_6495;
wire net_8486;
wire net_922;
wire net_522;
wire net_270;
wire net_2638;
wire net_9747;
wire net_13355;
wire net_12364;
wire net_7956;
wire net_5429;
wire net_14034;
wire net_11346;
wire net_1990;
wire net_4992;
wire net_7456;
wire net_10442;
wire net_5757;
wire net_6140;
wire net_2264;
wire net_11632;
wire net_977;
wire net_643;
wire net_4780;
wire net_9951;
wire net_7880;
wire net_11278;
wire net_11988;
wire net_11601;
wire net_622;
wire net_14854;
wire net_6876;
wire x3558;
wire net_15340;
wire net_13564;
wire net_11993;
wire net_11165;
wire net_6175;
wire net_3587;
wire net_3762;
wire net_10580;
wire net_3687;
wire net_11277;
wire net_5909;
wire net_10056;
wire net_11225;
wire net_12015;
wire net_10483;
wire net_5307;
wire net_1338;
wire net_4920;
wire net_7842;
wire net_2045;
wire net_3874;
wire net_2053;
wire net_9357;
wire net_11790;
wire net_6623;
wire net_11829;
wire net_2180;
wire net_2869;
wire x33;
wire net_3332;
wire net_4242;
wire net_1892;
wire net_3446;
wire net_1798;
wire net_2119;
wire net_3220;
wire net_4427;
wire net_4720;
wire net_7401;
wire net_13108;
wire net_13109;
wire net_13287;
wire net_8627;
wire net_837;
wire net_7474;
wire net_10723;
wire net_3469;
wire net_9449;
wire net_5920;
wire net_6124;
wire net_8384;
wire net_6992;
wire net_927;
wire net_13519;
wire net_11686;
wire net_2007;
wire net_5143;
wire net_5763;
wire net_7703;
wire net_713;
wire net_10653;
wire net_1519;
wire net_693;
wire net_12633;
wire net_5711;
wire net_6378;
wire net_13338;
wire net_8700;
wire net_11104;
wire net_729;
wire net_11390;
wire net_9222;
wire net_4197;
wire net_13777;
wire net_3964;
wire net_14893;
wire net_12660;
wire net_13156;
wire net_4219;
wire net_7093;
wire net_7324;
wire net_13948;
wire net_9169;
wire net_8447;
wire net_15166;
wire net_9311;
wire net_5366;
wire net_9898;
wire net_14596;
wire net_11865;
wire net_8711;
wire net_14632;
wire net_13571;
wire net_10847;
wire net_341;
wire net_13611;
wire net_13391;
wire net_14733;
wire net_11651;
wire net_10208;
wire net_12992;
wire net_970;
wire net_13362;
wire net_488;
wire net_13389;
wire net_8653;
wire net_15539;
wire net_12009;
wire net_10460;
wire net_4909;
wire net_6034;
wire net_8088;
wire net_5452;
wire net_8324;
wire net_2319;
wire net_13917;
wire net_13184;
wire net_15717;
wire net_3044;
wire net_5929;
wire net_11785;
wire net_5458;
wire net_7102;
wire net_11145;
wire net_8440;
wire net_1532;
wire net_14745;
wire net_8971;
wire net_13726;
wire net_12308;
wire net_6653;
wire net_14071;
wire net_8207;
wire net_4475;
wire net_14233;
wire net_12038;
wire net_11595;
wire net_10100;
wire net_15478;
wire net_2163;
wire net_3417;
wire net_14639;
wire net_3307;
wire net_7765;
wire net_13301;
wire net_12534;
wire net_553;
wire net_4958;
wire net_15215;
wire net_14719;
wire net_4212;
wire net_5057;
wire net_6133;
wire net_1093;
wire net_14947;
wire net_2592;
wire net_7797;
wire net_6230;
wire net_7680;
wire net_8300;
wire net_9876;
wire net_3580;
wire net_15505;
wire net_3259;
wire net_6239;
wire net_9877;
wire net_5260;
wire net_4701;
wire net_10057;
wire net_10889;
wire net_8833;
wire net_8922;
wire net_710;
wire net_14908;
wire net_462;
wire net_418;
wire net_15415;
wire net_15072;
wire net_14754;
wire net_3097;
wire net_14686;
wire net_5836;
wire net_15105;
wire net_161;
wire net_6478;
wire net_7988;
wire net_14401;
wire net_8660;
wire x1974;
wire net_3970;
wire x6351;
wire net_12516;
wire net_1486;
wire net_173;
wire net_2606;
wire net_3018;
wire net_14317;
wire net_1839;
wire net_2320;
wire net_1665;
wire net_11076;
wire net_9237;
wire net_3006;
wire net_6203;
wire net_14515;
wire net_13744;
wire net_10970;
wire net_8525;
wire net_8349;
wire net_1681;
wire net_7936;
wire net_3550;
wire net_12377;
wire net_11172;
wire net_14468;
wire net_7998;
wire net_15511;
wire net_6893;
wire net_9466;
wire net_2224;
wire net_7066;
wire net_10037;
wire net_4272;
wire net_15404;
wire net_6512;
wire net_5733;
wire net_10532;
wire net_746;
wire net_13406;
wire net_5877;
wire net_6147;
wire net_1274;
wire net_1682;
wire net_2458;
wire net_11302;
wire net_9324;
wire net_10788;
wire net_5743;
wire net_14485;
wire net_7910;
wire net_3435;
wire net_10109;
wire x3320;
wire net_3466;
wire net_2635;
wire x715;
wire net_3374;
wire net_5207;
wire net_15490;
wire net_13540;
wire net_4995;
wire net_5572;
wire net_7834;
wire net_1663;
wire net_629;
wire net_14579;
wire net_15068;
wire net_8283;
wire net_1037;
wire net_8666;
wire net_2019;
wire net_4209;
wire net_15326;
wire net_4676;
wire net_9382;
wire net_8395;
wire net_3019;
wire net_6675;
wire net_13784;
wire net_13033;
wire net_7549;
wire net_15017;
wire net_5579;
wire net_14710;
wire net_2351;
wire net_6793;
wire net_14457;
wire net_9628;
wire net_1350;
wire net_1648;
wire net_6242;
wire net_14433;
wire net_15012;
wire net_12594;
wire net_1623;
wire net_2982;
wire net_6219;
wire net_631;
wire net_6948;
wire net_14201;
wire net_12128;
wire net_4410;
wire net_7230;
wire net_10086;
wire net_5785;
wire net_14047;
wire net_14988;
wire net_13143;
wire net_4007;
wire net_8566;
wire net_4499;
wire net_12100;
wire net_14251;
wire net_13657;
wire net_8650;
wire net_7190;
wire net_10907;
wire net_9910;
wire net_15733;
wire net_8596;
wire x198;
wire net_6928;
wire net_670;
wire net_15159;
wire net_10984;
wire net_103;
wire net_6250;
wire net_12147;
wire net_2687;
wire net_12166;
wire net_6651;
wire net_9889;
wire net_5485;
wire net_7023;
wire net_7243;
wire net_12004;
wire net_10750;
wire net_3554;
wire net_9842;
wire net_9721;
wire net_12853;
wire net_12323;
wire net_1920;
wire net_4101;
wire net_3928;
wire net_13369;
wire net_2010;
wire net_14540;
wire x413;
wire net_3854;
wire net_7038;
wire net_11665;
wire net_8782;
wire net_6717;
wire net_6941;
wire net_9793;
wire net_9857;
wire net_8321;
wire net_9139;
wire net_5493;
wire net_13759;
wire net_4672;
wire net_8862;
wire net_6743;
wire net_755;
wire net_9557;
wire net_1723;
wire x389;
wire net_8465;
wire net_14981;
wire net_9285;
wire net_2900;
wire net_7754;
wire net_14790;
wire net_11015;
wire net_5152;
wire net_12545;
wire net_5718;
wire net_8190;
wire net_4376;
wire net_5892;
wire net_14397;
wire net_13468;
wire net_14953;
wire net_3151;
wire net_6763;
wire net_12890;
wire net_2306;
wire net_3628;
wire net_6053;
wire net_12382;
wire net_12023;
wire net_2873;
wire net_3272;
wire net_14479;
wire net_14618;
wire net_12829;
wire net_2254;
wire net_2861;
wire net_11319;
wire net_1652;
wire net_1429;
wire net_11844;
wire net_11061;
wire net_14343;
wire net_14223;
wire net_14895;
wire net_9570;
wire net_4574;
wire net_7130;
wire net_15223;
wire net_1209;
wire net_2725;
wire net_13166;
wire net_3613;
wire net_8964;
wire net_4615;
wire net_13076;
wire net_4038;
wire net_847;
wire net_727;
wire net_11242;
wire net_10157;
wire net_4787;
wire net_9804;
wire net_11740;
wire net_283;
wire net_12864;
wire net_13505;
wire net_12559;
wire net_5117;
wire net_3190;
wire net_4955;
wire net_4690;
wire net_12796;
wire net_3757;
wire net_11457;
wire net_5020;
wire net_15750;
wire net_14126;
wire net_7316;
wire net_12658;
wire net_9224;
wire net_4445;
wire net_15142;
wire net_5445;
wire net_7428;
wire net_10023;
wire net_11115;
wire net_10990;
wire net_14247;
wire net_7958;
wire net_344;
wire net_14102;
wire net_3951;
wire net_14614;
wire net_4757;
wire net_2269;
wire net_884;
wire net_15054;
wire net_14184;
wire net_712;
wire net_13010;
wire net_11635;
wire net_1422;
wire net_2281;
wire net_12940;
wire net_2259;
wire net_12124;
wire net_4497;
wire net_15079;
wire net_11527;
wire net_15107;
wire net_10651;
wire net_6670;
wire net_15061;
wire net_1106;
wire net_4095;
wire net_13629;
wire net_8483;
wire net_2739;
wire net_2972;
wire net_13330;
wire net_5611;
wire net_11715;
wire net_10113;
wire net_2110;
wire net_11311;
wire net_10836;
wire net_2919;
wire net_15252;
wire net_10642;
wire net_2893;
wire net_11435;
wire net_2241;
wire net_13006;
wire net_2358;
wire net_3227;
wire net_12651;
wire net_9522;
wire net_8615;
wire net_8682;
wire net_3057;
wire net_1547;
wire net_15596;
wire net_9039;
wire net_571;
wire net_13053;
wire net_10692;
wire net_8768;
wire net_10543;
wire net_7569;
wire net_14743;
wire net_5122;
wire net_12495;
wire net_10400;
wire net_4935;
wire net_12168;
wire net_3934;
wire net_10385;
wire net_11146;
wire net_5423;
wire net_13972;
wire net_1877;
wire net_720;
wire net_7971;
wire net_6507;
wire net_9912;
wire net_7653;
wire net_9038;
wire net_12152;
wire net_10395;
wire net_14005;
wire net_5209;
wire net_7344;
wire net_2199;
wire net_5055;
wire net_14886;
wire net_10628;
wire net_7303;
wire net_4794;
wire net_684;
wire net_2625;
wire net_4149;
wire net_2648;
wire x5647;
wire net_5687;
wire net_7299;
wire net_7542;
wire net_3720;
wire net_510;
wire net_12922;
wire net_10909;
wire net_6849;
wire net_10292;
wire net_1595;
wire net_5849;
wire net_15656;
wire net_114;
wire net_8885;
wire net_12919;
wire net_2653;
wire net_3432;
wire net_2960;
wire net_2974;
wire net_9078;
wire net_6519;
wire net_14517;
wire net_3895;
wire net_8339;
wire net_8257;
wire net_13660;
wire net_6703;
wire net_12577;
wire net_11736;
wire net_2734;
wire net_12888;
wire net_15508;
wire net_13133;
wire net_494;
wire net_2782;
wire net_7043;
wire net_10637;
wire net_12569;
wire net_6761;
wire net_14857;
wire net_3146;
wire net_6294;
wire net_7827;
wire net_12877;
wire net_10999;
wire net_6390;
wire net_9347;
wire net_10496;
wire net_5237;
wire net_4283;
wire net_14825;
wire net_15726;
wire net_6592;
wire net_13830;
wire net_11553;
wire net_8953;
wire net_3022;
wire net_6084;
wire net_8226;
wire net_3461;
wire net_12365;
wire net_10989;
wire net_10956;
wire net_10327;
wire net_11747;
wire net_7495;
wire net_14366;
wire net_4610;
wire net_9616;
wire net_5741;
wire net_6391;
wire net_8476;
wire net_457;
wire net_4459;
wire net_12096;
wire net_8821;
wire net_2246;
wire net_772;
wire net_6308;
wire net_10180;
wire net_14375;
wire net_4371;
wire net_5700;
wire net_10190;
wire x1547;
wire net_12773;
wire net_7441;
wire net_9671;
wire net_7966;
wire net_11807;
wire net_15405;
wire net_9159;
wire net_1277;
wire net_14567;
wire net_11899;
wire net_2661;
wire net_3893;
wire net_6113;
wire net_14260;
wire net_13459;
wire net_4706;
wire net_12467;
wire net_594;
wire net_5532;
wire net_11336;
wire net_9818;
wire net_4075;
wire net_6421;
wire net_7385;
wire net_14310;
wire net_6051;
wire net_11892;
wire net_8512;
wire net_11690;
wire net_1721;
wire net_2852;
wire net_6188;
wire net_7851;
wire net_12975;
wire net_4633;
wire net_4402;
wire net_6328;
wire net_6605;
wire net_6249;
wire net_5843;
wire net_2074;
wire net_8428;
wire net_5256;
wire net_5274;
wire net_10626;
wire net_10183;
wire net_2577;
wire net_11091;
wire net_8286;
wire net_2954;
wire net_8073;
wire net_1073;
wire net_11932;
wire net_1947;
wire net_3274;
wire net_2953;
wire net_141;
wire net_15731;
wire net_6380;
wire net_467;
wire net_879;
wire net_2910;
wire net_7227;
wire x4041;
wire net_2415;
wire net_8728;
wire net_4851;
wire net_2081;
wire net_15034;
wire net_9245;
wire net_8738;
wire net_10522;
wire net_5195;
wire net_7312;
wire net_11426;
wire net_13225;
wire net_14555;
wire net_3165;
wire net_12644;
wire net_10740;
wire net_1348;
wire net_3197;
wire net_15707;
wire net_9774;
wire net_7276;
wire net_4965;
wire net_7201;
wire net_12295;
wire net_8648;
wire net_2302;
wire net_3422;
wire net_10151;
wire net_199;
wire net_12523;
wire net_2789;
wire net_14601;
wire net_7844;
wire net_12903;
wire net_431;
wire net_3835;
wire net_8545;
wire net_5783;
wire net_13649;
wire net_8250;
wire net_5502;
wire net_6805;
wire net_10898;
wire net_9373;
wire net_6387;
wire net_6403;
wire net_7734;
wire net_13873;
wire net_12409;
wire net_15294;
wire net_2368;
wire net_5186;
wire net_222;
wire net_4362;
wire net_13215;
wire net_15727;
wire net_12908;
wire net_4520;
wire net_3966;
wire net_3999;
wire net_7060;
wire net_7804;
wire net_1788;
wire net_6330;
wire x3022;
wire net_12476;
wire net_607;
wire net_4301;
wire net_12392;
wire net_8106;
wire x3338;
wire net_9739;
wire net_2935;
wire net_4142;
wire net_1045;
wire net_6166;
wire net_3497;
wire net_3905;
wire net_13087;
wire net_4345;
wire net_15392;
wire net_10507;
wire net_9318;
wire net_13249;
wire net_3516;
wire net_4939;
wire net_11799;
wire net_6547;
wire net_3601;
wire net_9933;
wire net_4588;
wire net_1438;
wire net_10374;
wire net_4395;
wire net_4538;
wire net_8502;
wire net_14648;
wire net_13044;
wire net_12052;
wire net_15550;
wire net_1143;
wire net_14580;
wire net_11167;
wire net_12662;
wire net_1088;
wire net_4527;
wire net_9434;
wire net_6410;
wire net_6419;
wire net_8548;
wire net_13262;
wire net_4144;
wire net_4716;
wire net_7586;
wire net_2079;
wire net_3885;
wire net_1731;
wire net_706;
wire net_2052;
wire net_6373;
wire net_9298;
wire net_9089;
wire net_14376;
wire net_9648;
wire net_9463;
wire net_2768;
wire net_6912;
wire net_12813;
wire net_5125;
wire net_13276;
wire net_13479;
wire net_12536;
wire net_551;
wire net_5952;
wire net_5368;
wire net_7873;
wire net_11769;
wire net_15422;
wire net_3636;
wire net_4617;
wire net_7184;
wire net_14095;
wire x223;
wire net_13182;
wire net_4727;
wire net_15000;
wire net_5032;
wire net_11046;
wire net_1536;
wire net_5852;
wire net_6232;
wire net_11033;
wire net_12504;
wire net_12419;
wire net_3478;
wire net_4168;
wire net_12376;
wire net_1498;
wire net_8117;
wire net_11371;
wire net_1199;
wire net_7986;
wire net_15675;
wire net_10815;
wire net_8930;
wire net_14764;
wire net_3627;
wire net_5561;
wire net_15087;
wire net_15296;
wire net_5530;
wire net_5626;
wire net_949;
wire net_4869;
wire net_289;
wire net_450;
wire net_14000;
wire net_12401;
wire net_10936;
wire net_8041;
wire net_7813;
wire net_9046;
wire net_4111;
wire net_14204;
wire net_9392;
wire net_10972;
wire net_1642;
wire net_2614;
wire net_14267;
wire net_12158;
wire net_10616;
wire net_5322;
wire net_12947;
wire net_12287;
wire net_12722;
wire net_14283;
wire net_2524;
wire net_11490;
wire net_8262;
wire net_1224;
wire net_9028;
wire net_2296;
wire net_6786;
wire net_9438;
wire net_13804;
wire net_13994;
wire net_768;
wire net_3385;
wire net_11084;
wire net_357;
wire net_14423;
wire net_14068;
wire net_6954;
wire net_908;
wire net_9179;
wire net_12934;
wire net_13189;
wire net_7849;
wire net_519;
wire net_3451;
wire net_9697;
wire net_7085;
wire net_11773;
wire net_8790;
wire net_2694;
wire net_12280;
wire net_11052;
wire net_5607;
wire net_2096;
wire net_3118;
wire net_5555;
wire net_2697;
wire net_9184;
wire net_15330;
wire net_11501;
wire net_10808;
wire net_1829;
wire net_14240;
wire net_13904;
wire net_14082;
wire net_9190;
wire net_1204;
wire net_6282;
wire net_14089;
wire net_9780;
wire net_2342;
wire net_8331;
wire net_7336;
wire net_6628;
wire net_9969;
wire net_6778;
wire net_662;
wire net_862;
wire net_1986;
wire net_3214;
wire net_14972;
wire net_2307;
wire x285;
wire net_11472;
wire net_7168;
wire net_14822;
wire net_8127;
wire net_4174;
wire net_5396;
wire net_10864;
wire net_738;
wire net_4080;
wire net_4325;
wire net_12881;
wire net_1150;
wire net_504;
wire net_10333;
wire net_9789;
wire net_15321;
wire net_6634;
wire net_8203;
wire net_6467;
wire net_7527;
wire net_12613;
wire net_11537;
wire net_7698;
wire net_9164;
wire net_9012;
wire net_3406;
wire net_11657;
wire net_13110;
wire net_4229;
wire net_15624;
wire net_2130;
wire net_6474;
wire net_10198;
wire net_1148;
wire net_3362;
wire net_3120;
wire net_14324;
wire net_2382;
wire net_13620;
wire net_4504;
wire net_1561;
wire net_10698;
wire net_3442;
wire net_3864;
wire net_5942;
wire net_9271;
wire net_15357;
wire net_12161;
wire net_3269;
wire net_11455;
wire net_10472;
wire net_5796;
wire net_9730;
wire net_4421;
wire net_6666;
wire net_14725;
wire net_9416;
wire x948;
wire net_6975;
wire net_13329;
wire net_9855;
wire net_1940;
wire net_4389;
wire net_13323;
wire net_11449;
wire net_13935;
wire net_11798;
wire net_10452;
wire x921;
wire net_10728;
wire net_8635;
wire net_11516;
wire net_12781;
wire net_10425;
wire net_14621;
wire net_4561;
wire net_11528;
wire net_991;
wire net_3912;
wire net_6528;
wire net_13204;
wire net_11676;
wire net_6753;
wire net_14800;
wire net_3088;
wire net_1473;
wire net_11107;
wire net_4607;
wire net_12484;
wire net_2979;
wire net_10714;
wire net_2772;
wire net_9564;
wire net_8491;
wire net_5775;
wire net_1674;
wire net_4180;
wire net_5582;
wire net_1651;
wire net_15562;
wire net_2375;
wire net_13582;
wire net_5109;
wire net_13839;
wire net_12116;
wire net_1806;
wire net_6422;
wire net_3234;
wire net_12180;
wire net_15666;
wire net_2347;
wire net_8746;
wire net_1363;
wire net_11710;
wire net_1869;
wire net_14777;
wire net_2684;
wire net_3806;
wire net_4053;
wire net_10795;
wire net_10352;
wire net_10526;
wire net_521;
wire net_3972;
wire net_14275;
wire net_13029;
wire net_9003;
wire net_14738;
wire net_2754;
wire net_15713;
wire net_267;
wire net_1585;
wire x5427;
wire net_13748;
wire net_11613;
wire net_9143;
wire net_11099;
wire net_4012;
wire net_6898;
wire net_7421;
wire net_6169;
wire net_3663;
wire net_10885;
wire net_3260;
wire net_5110;
wire net_6647;
wire net_13017;
wire net_9186;
wire net_6465;
wire net_6486;
wire net_3681;
wire net_6048;
wire net_13177;
wire net_6621;
wire net_2716;
wire net_7902;
wire net_13097;
wire net_7503;
wire net_12717;
wire net_7857;
wire net_15180;
wire net_14522;
wire net_11815;
wire net_10015;
wire net_5246;
wire net_351;
wire net_8558;
wire net_6551;
wire net_4750;
wire net_7761;
wire net_13346;
wire net_4558;
wire net_12858;
wire net_12601;
wire x3606;
wire net_10856;
wire net_6006;
wire net_4240;
wire net_7964;
wire net_15581;
wire net_2842;
wire net_8394;
wire net_15521;
wire net_1257;
wire net_2828;
wire net_3158;
wire net_939;
wire net_12749;
wire net_8365;
wire net_824;
wire net_3458;
wire x420;
wire net_1822;
wire net_13781;
wire net_7984;
wire net_9755;
wire net_14411;
wire net_13038;
wire net_10479;
wire net_1972;
wire net_2791;
wire net_15559;
wire net_10111;
wire net_11023;
wire net_12267;
wire net_3126;
wire net_993;
wire net_15047;
wire net_10555;
wire net_8795;
wire net_4271;
wire net_11817;
wire net_9895;
wire net_317;
wire net_856;
wire net_5974;
wire net_11853;
wire net_9456;
wire net_1100;
wire net_7035;
wire net_15121;
wire net_9944;
wire net_14995;
wire net_7920;
wire net_3845;
wire net_2817;
wire net_6686;
wire net_2026;
wire net_10046;
wire net_11822;
wire net_5727;
wire net_15128;
wire net_12195;
wire net_5673;
wire net_5996;
wire net_6730;
wire net_13823;
wire net_1326;
wire net_3033;
wire net_7488;
wire net_134;
wire net_546;
wire net_14059;
wire net_4648;
wire net_14638;
wire net_3373;
wire net_5382;
wire net_11471;
wire net_2672;
wire net_4546;
wire net_5351;
wire net_588;
wire net_10065;
wire net_13735;
wire net_13320;
wire net_2200;
wire net_8641;
wire net_8062;
wire net_1157;
wire net_12424;
wire net_3701;
wire net_14296;
wire net_4736;
wire net_7486;
wire net_7592;
wire net_7785;
wire net_5592;
wire net_5642;
wire net_8012;
wire net_4974;
wire net_7906;
wire net_3883;
wire net_6001;
wire net_9378;
wire net_1542;
wire net_1172;
wire net_14198;
wire net_9124;
wire net_13703;
wire net_8431;
wire net_4230;
wire net_6350;
wire net_14626;
wire net_7993;
wire net_9840;
wire net_14270;
wire net_10560;
wire net_11800;
wire net_13604;
wire net_5603;
wire net_9503;
wire net_1065;
wire net_13117;
wire net_4860;
wire x6303;
wire net_2237;
wire net_2566;
wire net_8352;
wire net_3795;
wire net_3953;
wire net_13046;
wire net_15696;
wire net_3100;
wire net_13375;
wire net_917;
wire net_241;
wire net_9353;
wire net_3730;
wire net_13196;
wire net_13640;
wire net_13515;
wire net_12010;
wire net_2874;
wire net_10965;
wire net_8942;
wire net_13350;
wire x1121;
wire net_14535;
wire net_4597;
wire net_13814;
wire net_599;
wire net_9685;
wire net_4589;
wire net_2993;
wire net_10921;
wire net_3067;
wire net_13950;
wire net_10075;
wire net_4844;
wire net_4288;
wire net_5860;
wire net_3111;
wire net_323;
wire net_5402;
wire net_963;
wire net_10301;
wire net_10346;
wire net_11880;
wire net_13543;
wire x3867;
wire net_9653;
wire net_13575;
wire net_9482;
wire net_8692;
wire net_8356;
wire net_7368;
wire net_3737;
wire net_4689;
wire net_10216;
wire net_153;
wire net_2389;
wire net_12328;
wire net_6276;
wire net_7556;
wire net_15384;
wire net_375;
wire net_562;
wire net_6103;
wire net_364;
wire net_8675;
wire net_12260;
wire net_14380;
wire net_12770;
wire net_11723;
wire net_3172;
wire net_10485;
wire net_9686;
wire net_13772;
wire net_11706;
wire net_4239;
wire net_2849;
wire net_14011;
wire net_12671;
wire net_5516;
wire net_7177;
wire net_10799;
wire net_15641;
wire net_6313;
wire net_15267;
wire net_12693;
wire net_6341;
wire net_5589;
wire net_8161;
wire net_6840;
wire net_12810;
wire net_4873;
wire net_10851;
wire net_3171;
wire net_4298;
wire net_7514;
wire net_15175;
wire net_11286;
wire net_14217;
wire net_12742;
wire net_14472;
wire net_11250;
wire net_8004;
wire net_7170;
wire x4449;
wire net_10091;
wire net_8173;
wire net_1247;
wire net_3673;
wire net_4137;
wire net_11149;
wire net_8528;
wire net_2388;
wire net_5162;
wire net_9870;
wire net_15383;
wire net_14006;
wire net_7561;
wire net_5765;
wire net_3496;
wire net_1215;
wire net_5169;
wire net_15010;
wire net_5248;
wire net_15578;
wire net_13361;
wire net_4216;
wire net_129;
wire net_98;
wire net_4889;
wire net_10371;
wire net_151;
wire net_13638;
wire net_1625;
wire net_8784;
wire net_284;
wire net_6655;
wire net_9930;
wire net_12743;
wire net_439;
wire net_2513;
wire net_259;
wire net_3582;
wire net_3351;
wire net_4094;
wire net_8662;
wire net_7360;
wire net_7142;
wire net_10291;
wire net_10153;
wire net_3119;
wire net_1231;
wire net_187;
wire net_5841;
wire net_14072;
wire net_3305;
wire x957;
wire net_14045;
wire net_160;
wire net_6205;
wire net_832;
wire net_12304;
wire net_815;
wire net_7875;
wire net_11304;
wire net_15049;
wire net_6514;
wire net_6749;
wire net_7728;
wire net_5578;
wire net_13742;
wire net_7670;
wire net_7897;
wire net_5632;
wire net_6501;
wire net_10279;
wire net_586;
wire net_9580;
wire net_10845;
wire net_1347;
wire net_5272;
wire net_1091;
wire net_6240;
wire net_13145;
wire net_3838;
wire net_7812;
wire net_7768;
wire net_11518;
wire net_3745;
wire net_120;
wire net_6260;
wire net_15116;
wire net_12489;
wire net_292;
wire net_5529;
wire net_11713;
wire net_9879;
wire net_3708;
wire net_12141;
wire net_9384;
wire net_96;
wire net_167;
wire net_12371;
wire net_5830;
wire net_5227;
wire net_7536;
wire net_14259;
wire net_7042;
wire net_6073;
wire net_6170;
wire net_7308;
wire net_8864;
wire net_7478;
wire net_15325;
wire net_9847;
wire net_2556;
wire net_8599;
wire net_3519;
wire net_5735;
wire net_2740;
wire net_14756;
wire net_2806;
wire net_7294;
wire net_9679;
wire net_672;
wire net_14624;
wire net_13163;
wire net_4924;
wire net_15015;
wire net_8834;
wire net_4483;
wire net_8391;
wire net_5212;
wire net_2027;
wire net_9367;
wire net_5045;
wire net_13761;
wire net_14441;
wire net_11680;
wire x3249;
wire net_7021;
wire net_11335;
wire net_6237;
wire net_2456;
wire net_3610;
wire net_2753;
wire net_8963;
wire net_14635;
wire net_10036;
wire net_1232;
wire net_9585;
wire net_4540;
wire net_5662;
wire net_5784;
wire net_1953;
wire net_3059;
wire net_15177;
wire net_11625;
wire net_13506;
wire net_10684;
wire net_12540;
wire net_14295;
wire net_3925;
wire net_5444;
wire net_13039;
wire net_464;
wire net_12003;
wire net_3847;
wire net_4473;
wire net_8230;
wire net_4582;
wire net_5699;
wire net_5089;
wire net_4200;
wire net_4547;
wire net_14205;
wire net_5867;
wire net_6300;
wire net_5362;
wire net_7819;
wire net_14455;
wire net_8954;
wire net_15154;
wire net_10136;
wire net_4640;
wire net_10926;
wire net_11602;
wire net_4658;
wire net_14195;
wire net_12625;
wire net_14602;
wire net_1256;
wire net_7071;
wire net_7982;
wire net_13264;
wire net_1413;
wire net_802;
wire net_12194;
wire net_14252;
wire net_15262;
wire net_3556;
wire net_13872;
wire net_3041;
wire net_1840;
wire net_12930;
wire net_12602;
wire net_4997;
wire net_14359;
wire net_9230;
wire net_6620;
wire net_8015;
wire net_5637;
wire net_3427;
wire net_7167;
wire net_1031;
wire net_4824;
wire net_13170;
wire net_15181;
wire net_7049;
wire net_14189;
wire net_13404;
wire net_1636;
wire net_7568;
wire net_9714;
wire net_3257;
wire net_10265;
wire net_13394;
wire net_4458;
wire net_7245;
wire net_10899;
wire net_9744;
wire net_7458;
wire net_10467;
wire net_10344;
wire net_10270;
wire net_10991;
wire net_1334;
wire net_10782;
wire net_757;
wire net_206;
wire x1179;
wire net_8523;
wire net_2020;
wire net_1688;
wire net_10087;
wire net_13522;
wire net_10794;
wire net_13383;
wire net_10894;
wire net_7665;
wire net_15430;
wire net_14134;
wire net_235;
wire net_6126;
wire net_14056;
wire net_15076;
wire net_13121;
wire net_14970;
wire net_11695;
wire net_12223;
wire net_2961;
wire net_4159;
wire net_4324;
wire net_5108;
wire net_2374;
wire net_7322;
wire net_9911;
wire net_4203;
wire net_7652;
wire net_5631;
wire net_3644;
wire net_10571;
wire net_12273;
wire net_250;
wire net_3600;
wire net_8655;
wire net_7260;
wire net_3081;
wire net_5882;
wire net_12927;
wire net_11279;
wire net_2055;
wire net_10283;
wire net_4879;
wire net_6144;
wire net_14570;
wire net_12929;
wire net_2630;
wire net_7420;
wire net_10027;
wire net_1985;
wire net_403;
wire net_3524;
wire net_2340;
wire net_6265;
wire net_13680;
wire net_14421;
wire net_14883;
wire net_12219;
wire net_2275;
wire net_15560;
wire net_14302;
wire net_10752;
wire net_3976;
wire net_9619;
wire net_9899;
wire net_10939;
wire net_12562;
wire net_12202;
wire net_8602;
wire net_13128;
wire net_841;
wire net_10803;
wire net_1750;
wire net_14910;
wire net_6411;
wire net_794;
wire net_2397;
wire net_3346;
wire net_13277;
wire net_8136;
wire net_8269;
wire net_528;
wire net_10537;
wire net_3433;
wire net_335;
wire net_4878;
wire net_3464;
wire net_1468;
wire net_9132;
wire net_181;
wire net_9661;
wire net_4774;
wire net_6784;
wire net_11767;
wire net_12214;
wire net_3333;
wire net_11556;
wire net_6011;
wire net_10631;
wire net_9014;
wire net_8494;
wire net_7350;
wire net_13530;
wire net_6177;
wire net_6796;
wire net_3649;
wire net_2539;
wire net_1130;
wire net_14826;
wire net_5921;
wire net_6216;
wire net_8111;
wire net_386;
wire net_12680;
wire net_9421;
wire net_8239;
wire net_6150;
wire net_10051;
wire net_1790;
wire net_6451;
wire net_7918;
wire net_8166;
wire net_4103;
wire net_6493;
wire net_9281;
wire net_11221;
wire net_6130;
wire net_6309;
wire net_7745;
wire net_2318;
wire net_8787;
wire net_9207;
wire net_5562;
wire net_3449;
wire net_15719;
wire net_10583;
wire net_9134;
wire net_9004;
wire net_12718;
wire net_1039;
wire net_7573;
wire net_1709;
wire net_11972;
wire net_7822;
wire net_10981;
wire net_15499;
wire net_8629;
wire net_400;
wire net_4651;
wire net_14546;
wire net_10080;
wire net_9698;
wire net_1935;
wire net_5707;
wire net_11608;
wire net_13622;
wire net_175;
wire net_13102;
wire net_12650;
wire net_2925;
wire net_1850;
wire net_11873;
wire net_9142;
wire net_4429;
wire net_14956;
wire net_1855;
wire net_4882;
wire net_6365;
wire net_1992;
wire net_1177;
wire net_1163;
wire net_15606;
wire net_12346;
wire net_897;
wire net_7384;
wire net_13890;
wire net_11362;
wire net_10206;
wire net_5466;
wire net_9521;
wire net_2853;
wire net_10578;
wire net_2705;
wire net_7840;
wire net_5164;
wire net_9215;
wire net_615;
wire net_6712;
wire net_11494;
wire net_3273;
wire net_1559;
wire net_441;
wire net_8706;
wire net_5665;
wire net_1620;
wire net_13966;
wire net_2608;
wire net_14266;
wire net_14224;
wire net_6032;
wire net_14856;
wire net_9763;
wire net_2813;
wire net_2663;
wire net_728;
wire net_14559;
wire net_1276;
wire net_5473;
wire net_719;
wire net_7774;
wire net_14905;
wire net_10878;
wire net_170;
wire net_15138;
wire net_8068;
wire net_6873;
wire net_14032;
wire net_2571;
wire net_9888;
wire net_5305;
wire net_10741;
wire net_5703;
wire net_12264;
wire net_9418;
wire net_14325;
wire net_3479;
wire net_8609;
wire net_13617;
wire net_3222;
wire net_14661;
wire net_3321;
wire net_15342;
wire net_6393;
wire net_15631;
wire net_13764;
wire net_8410;
wire net_708;
wire net_15314;
wire net_3552;
wire net_696;
wire net_7685;
wire net_14079;
wire net_10824;
wire net_10777;
wire net_3216;
wire net_5713;
wire net_7427;
wire net_13175;
wire net_13947;
wire net_10401;
wire net_12972;
wire net_12256;
wire net_171;
wire net_15599;
wire net_10448;
wire net_9953;
wire net_15492;
wire net_9796;
wire net_15134;
wire net_10013;
wire net_6563;
wire net_3821;
wire net_9228;
wire net_10528;
wire net_604;
wire net_14101;
wire net_8403;
wire net_14578;
wire net_4503;
wire net_10872;
wire net_15465;
wire net_12385;
wire net_6938;
wire net_3486;
wire net_483;
wire net_15439;
wire net_15241;
wire net_7359;
wire net_1149;
wire net_9937;
wire net_8097;
wire net_5839;
wire net_7955;
wire net_11199;
wire net_8590;
wire net_15507;
wire net_8919;
wire net_9981;
wire net_8302;
wire net_1298;
wire net_15318;
wire net_296;
wire net_2131;
wire net_6681;
wire net_9733;
wire net_5651;
wire net_13461;
wire net_12845;
wire net_12053;
wire net_7004;
wire net_7153;
wire net_13632;
wire net_8941;
wire net_5435;
wire net_11369;
wire net_11461;
wire net_2228;
wire net_12357;
wire net_3020;
wire net_13720;
wire net_786;
wire net_5141;
wire net_11801;
wire net_11564;
wire net_8998;
wire net_9470;
wire net_127;
wire net_10518;
wire net_1339;
wire net_10608;
wire net_3781;
wire net_5685;
wire net_906;
wire net_15450;
wire net_9892;
wire net_9080;
wire net_8461;
wire net_2422;
wire net_5205;
wire net_3577;
wire net_13951;
wire net_10185;
wire net_652;
wire net_12955;
wire net_13958;
wire net_10137;
wire net_13707;
wire net_3840;
wire net_1815;
wire net_4361;
wire net_10590;
wire net_15458;
wire net_10211;
wire net_6145;
wire net_3782;
wire net_14840;
wire net_14513;
wire net_13250;
wire net_2505;
wire net_11185;
wire net_877;
wire net_14680;
wire net_2799;
wire net_10748;
wire net_6139;
wire net_6868;
wire net_6834;
wire net_8092;
wire net_3734;
wire net_14135;
wire net_2683;
wire net_14524;
wire net_8021;
wire net_4812;
wire net_15714;
wire net_9654;
wire net_2165;
wire net_4253;
wire net_11943;
wire net_11570;
wire net_11232;
wire net_8315;
wire net_4066;
wire net_13296;
wire net_6257;
wire net_14869;
wire net_8026;
wire net_3284;
wire net_1474;
wire net_4297;
wire net_15482;
wire net_12088;
wire net_2784;
wire net_6861;
wire net_11049;
wire net_15642;
wire net_13843;
wire net_8753;
wire net_675;
wire net_2562;
wire net_15417;
wire net_8355;
wire net_2867;
wire net_5134;
wire net_14931;
wire net_9129;
wire net_5293;
wire net_7195;
wire net_13841;
wire net_3472;
wire net_9120;
wire x2589;
wire net_10700;
wire net_7578;
wire net_8151;
wire net_5172;
wire net_10092;
wire net_8145;
wire net_2182;
wire net_1768;
wire net_9928;
wire net_8032;
wire net_4718;
wire net_9295;
wire net_150;
wire net_12950;
wire net_6589;
wire net_7677;
wire net_11915;
wire net_304;
wire net_4351;
wire net_6993;
wire net_10951;
wire net_12436;
wire net_9791;
wire net_7326;
wire net_14967;
wire net_4347;
wire net_7666;
wire net_12768;
wire net_10551;
wire net_1703;
wire net_11004;
wire net_7848;
wire net_9420;
wire net_7731;
wire net_15431;
wire net_9690;
wire net_3693;
wire net_12731;
wire net_15517;
wire net_9027;
wire net_5100;
wire net_1316;
wire net_6845;
wire net_6545;
wire net_14849;
wire net_4319;
wire net_792;
wire net_15744;
wire net_13848;
wire net_13695;
wire net_3070;
wire net_6223;
wire net_13782;
wire net_8842;
wire net_3409;
wire net_9481;
wire net_2203;
wire net_4430;
wire net_13415;
wire net_5373;
wire net_4525;
wire net_1904;
wire net_9446;
wire net_3907;
wire net_5678;
wire net_6332;
wire net_219;
wire net_3609;
wire net_10001;
wire net_6584;
wire net_8617;
wire net_9976;
wire net_2187;
wire net_2476;
wire net_13798;
wire net_913;
wire net_10764;
wire net_4518;
wire net_5378;
wire net_5338;
wire net_13242;
wire net_3387;
wire net_14938;
wire net_13591;
wire net_1479;
wire net_7157;
wire net_15423;
wire net_4330;
wire net_7756;
wire net_15611;
wire net_10268;
wire net_4019;
wire net_15037;
wire net_4152;
wire net_6895;
wire net_10066;
wire net_10832;
wire net_3094;
wire net_360;
wire net_13561;
wire net_1927;
wire net_7017;
wire net_14832;
wire net_10243;
wire net_213;
wire net_6910;
wire net_2324;
wire net_11688;
wire net_9244;
wire net_947;
wire net_4805;
wire net_5359;
wire net_7970;
wire net_14715;
wire net_1126;
wire net_11538;
wire net_2004;
wire net_13259;
wire net_1325;
wire net_6943;
wire net_3316;
wire net_10162;
wire net_3032;
wire net_9507;
wire net_5094;
wire net_6298;
wire net_1373;
wire net_1352;
wire net_2885;
wire net_2567;
wire net_10735;
wire net_10258;
wire net_4696;
wire net_8814;
wire net_14029;
wire net_10944;
wire net_1187;
wire net_7643;
wire net_7408;
wire net_7411;
wire net_4988;
wire net_3206;
wire net_1303;
wire net_8050;
wire net_2858;
wire net_6334;
wire net_15470;
wire net_14806;
wire net_14703;
wire net_2102;
wire net_15004;
wire net_4451;
wire net_5569;
wire net_12234;
wire net_12047;
wire net_1442;
wire net_11903;
wire net_1807;
wire net_10042;
wire net_1943;
wire net_1930;
wire x2214;
wire net_11544;
wire net_15188;
wire net_12298;
wire net_1894;
wire net_12113;
wire net_9645;
wire net_10694;
wire net_2431;
wire net_11555;
wire net_4054;
wire net_5544;
wire net_8213;
wire net_633;
wire net_113;
wire net_5054;
wire net_5750;
wire net_10115;
wire net_9674;
wire net_4848;
wire net_1914;
wire net_7791;
wire net_14944;
wire net_2408;
wire x682;
wire net_3889;
wire net_14899;
wire net_9904;
wire net_6627;
wire net_5943;
wire net_14039;
wire net_6974;
wire net_3567;
wire net_15022;
wire net_14669;
wire net_13717;
wire net_15540;
wire net_7831;
wire net_1457;
wire net_11525;
wire net_2741;
wire net_7010;
wire net_5414;
wire net_14876;
wire net_6483;
wire net_4011;
wire net_6616;
wire net_2448;
wire net_1436;
wire net_15285;
wire net_5424;
wire net_5541;
wire net_9199;
wire net_4338;
wire net_13234;
wire net_10719;
wire net_10054;
wire net_3400;
wire net_10725;
wire net_3392;
wire net_9571;
wire net_2551;
wire net_11572;
wire net_14925;
wire net_646;
wire net_12547;
wire net_2731;
wire net_5823;
wire net_14348;
wire net_11016;
wire net_2601;
wire net_6323;
wire net_8902;
wire net_2891;
wire net_8499;
wire net_520;
wire net_14314;
wire net_13482;
wire net_10159;
wire net_11201;
wire net_8928;
wire net_7237;
wire net_11261;
wire net_4722;
wire net_15269;
wire net_14110;
wire net_3231;
wire net_981;
wire net_2401;
wire net_14502;
wire net_9636;
wire net_8895;
wire net_1566;
wire net_15530;
wire net_1305;
wire net_11584;
wire net_2354;
wire net_12156;
wire net_14493;
wire net_9393;
wire net_1387;
wire net_1581;
wire net_10709;
wire net_10378;
wire net_10440;
wire net_15676;
wire net_8858;
wire net_5018;
wire net_7369;
wire net_11808;
wire net_4468;
wire net_2413;
wire net_5013;
wire net_7786;
wire net_11413;
wire net_559;
wire net_14462;
wire net_3042;
wire net_2792;
wire net_345;
wire net_2965;
wire net_2128;
wire net_12804;
wire net_1717;
wire net_7476;
wire net_9990;
wire net_11891;
wire net_6553;
wire net_398;
wire net_5302;
wire net_3399;
wire net_6976;
wire net_11489;
wire net_9344;
wire net_5080;
wire net_6693;
wire net_11140;
wire net_13584;
wire net_12834;
wire net_2117;
wire net_2461;
wire net_14654;
wire net_4085;
wire net_1766;
wire net_13493;
wire net_7393;
wire net_2582;
wire net_10099;
wire net_8974;
wire net_12472;
wire net_7898;
wire net_5905;
wire net_15233;
wire net_9788;
wire net_6724;
wire net_10419;
wire net_3872;
wire net_4956;
wire net_6054;
wire net_11867;
wire net_1572;
wire net_9407;
wire net_4447;
wire net_10357;
wire net_11647;
wire net_10226;
wire net_9265;
wire net_13933;
wire net_9235;
wire net_8990;
wire net_2134;
wire x341;
wire net_5179;
wire net_14166;
wire net_8794;
wire net_15595;
wire net_9834;
wire net_316;
wire net_5011;
wire net_13439;
wire net_4250;
wire net_4961;
wire net_15303;
wire net_4184;
wire net_11462;
wire net_14736;
wire net_12667;
wire net_14398;
wire net_13536;
wire net_13443;
wire net_10387;
wire net_1759;
wire net_14962;
wire net_12996;
wire net_7033;
wire net_15308;
wire net_12752;
wire net_3764;
wire net_4647;
wire net_15649;
wire net_12964;
wire net_4022;
wire net_11636;
wire net_2541;
wire net_12310;
wire net_9618;
wire net_3689;
wire net_12635;
wire net_533;
wire net_7436;
wire net_13282;
wire net_8347;
wire net_10040;
wire net_1695;
wire net_5932;
wire net_911;
wire net_1617;
wire net_7775;
wire net_12017;
wire x1129;
wire net_7005;
wire net_10047;
wire net_9608;
wire net_6637;
wire net_9015;
wire net_7053;
wire x6241;
wire net_5969;
wire net_5570;
wire net_9332;
wire net_15463;
wire net_11745;
wire net_9457;
wire net_568;
wire net_4579;
wire net_13709;
wire net_13809;
wire net_7962;
wire net_4807;
wire net_1227;
wire net_6046;
wire net_6485;
wire net_1008;
wire net_5312;
wire x3613;
wire net_5340;
wire net_5861;
wire net_1443;
wire net_12178;
wire net_11888;
wire net_3069;
wire net_4862;
wire net_8691;
wire net_3170;
wire net_12239;
wire net_2840;
wire net_14721;
wire net_3463;
wire net_4005;
wire net_6008;
wire net_4819;
wire net_11883;
wire net_3199;
wire net_8001;
wire net_3597;
wire net_5671;
wire net_15602;
wire net_14773;
wire net_14533;
wire net_269;
wire net_5043;
wire net_3193;
wire net_3131;
wire net_469;
wire net_10107;
wire net_12171;
wire net_3179;
wire net_1978;
wire net_1945;
wire net_10064;
wire net_7207;
wire net_10858;
wire net_3167;
wire net_4073;
wire net_5159;
wire net_1170;
wire net_1833;
wire net_5656;
wire net_10144;
wire net_8496;
wire net_13202;
wire net_2280;
wire net_2831;
wire net_9174;
wire net_3029;
wire net_9622;
wire net_2366;
wire net_778;
wire net_7818;
wire net_5725;
wire net_12779;
wire net_2930;
wire net_1455;
wire net_9816;
wire net_8252;
wire net_6523;
wire net_14277;
wire net_15651;
wire net_5064;
wire net_5323;
wire net_6024;
wire net_12167;
wire net_6225;
wire net_11780;
wire net_6832;
wire net_5261;
wire net_4730;
wire net_12154;
wire net_6643;
wire net_11123;
wire net_8172;
wire net_15292;
wire net_7912;
wire net_5380;
wire net_10173;
wire net_8519;
wire net_4119;
wire net_5648;
wire net_14246;
wire net_11152;
wire net_13445;
wire net_11251;
wire net_9450;
wire net_9216;
wire net_10644;
wire net_3980;
wire net_10566;
wire net_10335;
wire net_1481;
wire net_10392;
wire net_995;
wire net_5645;
wire net_7922;
wire net_8328;
wire net_7088;
wire net_700;
wire net_5000;
wire net_12232;
wire net_7334;
wire net_11433;
wire net_9947;
wire net_8957;
wire net_1246;
wire net_13325;
wire net_11043;
wire net_6043;
wire net_7705;
wire net_5216;
wire net_15195;
wire net_1774;
wire net_4228;
wire net_11402;
wire net_11819;
wire net_1673;
wire net_3060;
wire net_10712;
wire net_2568;
wire net_11103;
wire net_11941;
wire net_3480;
wire net_321;
wire net_6715;
wire net_9465;
wire net_8933;
wire net_5518;
wire net_4135;
wire net_2995;
wire net_6982;
wire net_15532;
wire net_3526;
wire net_2945;
wire net_934;
wire net_3103;
wire net_12855;
wire net_5941;
wire net_3665;
wire net_544;
wire net_717;
wire net_4896;
wire net_15587;
wire net_12305;
wire net_10505;
wire net_15328;
wire net_8201;
wire net_11952;
wire net_3630;
wire net_1824;
wire net_12037;
wire net_9659;
wire net_3402;
wire net_2223;
wire net_7603;
wire net_4763;
wire net_5074;
wire net_6957;
wire net_8008;
wire net_2673;
wire net_5694;
wire net_3500;
wire net_6164;
wire net_3166;
wire net_9104;
wire net_7065;
wire net_10861;
wire net_9831;
wire net_9358;
wire net_8079;
wire net_5903;
wire net_7513;
wire net_10665;
wire net_9652;
wire net_1245;
wire net_5552;
wire net_3660;
wire net_860;
wire net_5806;
wire net_870;
wire net_9254;
wire net_7135;
wire net_14474;
wire net_2046;
wire net_7176;
wire net_11708;
wire net_7521;
wire net_7926;
wire net_10819;
wire net_7941;
wire net_2878;
wire net_2871;
wire net_13642;
wire net_12012;
wire net_9850;
wire net_3267;
wire net_14581;
wire net_2321;
wire net_6286;
wire net_9108;
wire net_12874;
wire net_12668;
wire net_11645;
wire net_817;
wire net_11667;
wire net_5127;
wire net_15006;
wire net_3414;
wire net_14804;
wire net_7058;
wire net_14155;
wire net_10922;
wire net_10967;
wire net_7362;
wire net_14084;
wire net_13502;
wire net_9766;
wire net_4576;
wire net_13655;
wire net_2920;
wire net_1591;
wire net_14123;
wire net_13344;
wire net_7695;
wire net_13278;
wire net_1747;
wire net_5483;
wire net_2012;
wire net_650;
wire net_7139;
wire net_15080;
wire net_9761;
wire net_5557;
wire net_597;
wire net_9890;
wire net_15178;
wire net_14065;
wire net_743;
wire net_14387;
wire net_3770;
wire net_15333;
wire net_9062;
wire net_1922;
wire net_5984;
wire net_10482;
wire net_8272;
wire net_15109;
wire net_14281;
wire net_6336;
wire net_12481;
wire net_8889;
wire net_10853;
wire net_14620;
wire net_12384;
wire net_603;
wire net_6639;
wire net_8264;
wire net_4913;
wire net_13499;
wire net_2451;
wire net_14332;
wire net_642;
wire net_9806;
wire net_2699;
wire net_1522;
wire net_4031;
wire net_1158;
wire net_6989;
wire net_11496;
wire net_2926;
wire net_8006;
wire net_11082;
wire net_10775;
wire net_12782;
wire net_11530;
wire net_13964;
wire net_12289;
wire net_8042;
wire net_470;
wire x111;
wire net_13751;
wire net_2702;
wire net_430;
wire net_6991;
wire net_2834;
wire net_11659;
wire net_4551;
wire net_15255;
wire net_5972;
wire net_13557;
wire net_12945;
wire net_3943;
wire net_9370;
wire net_14996;
wire net_15183;
wire net_3129;
wire net_4438;
wire net_7675;
wire net_8568;
wire net_12353;
wire net_10839;
wire net_14154;
wire net_8557;
wire net_11771;
wire net_1063;
wire net_4218;
wire net_968;
wire net_13876;
wire net_14644;
wire net_13572;
wire net_9669;
wire net_12692;
wire net_10421;
wire net_12571;
wire net_9127;
wire net_2534;
wire net_6827;
wire net_7297;
wire net_4133;
wire net_13577;
wire net_15089;
wire net_1504;
wire x2968;
wire net_475;
wire net_6737;
wire net_9432;
wire net_7216;
wire net_14272;
wire net_11137;
wire net_3732;
wire x2707;
wire net_14024;
wire net_13768;
wire net_6903;
wire net_2309;
wire net_502;
wire net_8647;
wire net_2470;
wire net_1564;
wire net_11474;
wire net_1568;
wire net_6632;
wire net_14288;
wire net_12282;
wire net_3804;
wire net_15353;
wire net_10883;
wire net_6756;
wire net_9398;
wire net_1526;
wire net_13271;
wire net_13860;
wire net_8290;
wire net_1884;
wire net_12341;
wire net_12209;
wire net_13858;
wire net_3919;
wire net_7990;
wire net_4112;
wire x91;
wire net_2646;
wire net_3868;
wire net_3936;
wire net_7121;
wire net_4364;
wire net_13198;
wire net_5887;
wire net_6645;
wire net_13233;
wire net_2628;
wire net_4512;
wire net_6535;
wire net_9305;
wire net_11692;
wire net_5145;
wire net_12757;
wire net_11439;
wire net_11160;
wire net_1360;
wire net_6344;
wire net_10494;
wire net_9047;
wire net_3364;
wire net_11078;
wire net_13837;
wire net_13800;
wire net_5316;
wire net_664;
wire net_14420;
wire net_1364;
wire net_6003;
wire net_5050;
wire net_14727;
wire net_6292;
wire net_4622;
wire net_827;
wire net_549;
wire net_4605;
wire net_10192;
wire net_11050;
wire net_10450;
wire net_4295;
wire net_10687;
wire net_4563;
wire net_2337;
wire net_15684;
wire net_14928;
wire net_12533;
wire net_6945;
wire net_1369;
wire net_10614;
wire net_5773;
wire net_6900;
wire net_6405;
wire net_11068;
wire net_4695;
wire net_14779;
wire net_13550;
wire net_7469;
wire net_8622;
wire x1231;
wire net_1013;
wire net_1530;
wire net_6210;
wire net_13869;
wire net_3075;
wire net_2952;
wire net_842;
wire net_11783;
wire net_2336;
wire net_1705;
wire net_14977;
wire net_2035;
wire net_6571;
wire net_9500;
wire net_11215;
wire net_8951;
wire net_5070;
wire net_2826;
wire net_6560;
wire net_10325;
wire net_8199;
wire net_3739;
wire net_10451;
wire net_8455;
wire x898;
wire net_492;
wire net_11392;
wire net_3678;
wire net_6847;
wire net_15123;
wire net_2141;
wire net_7234;
wire net_8797;
wire net_2639;
wire net_14211;
wire net_10830;
wire net_8071;
wire net_11803;
wire net_14818;
wire net_13370;
wire net_11213;
wire net_3695;
wire net_3453;
wire net_12648;
wire net_5450;
wire net_5702;
wire net_1327;
wire net_8632;
wire net_110;
wire net_10598;
wire net_9822;
wire net_4968;
wire net_15447;
wire net_1403;
wire net_6097;
wire net_4532;
wire net_15337;
wire net_12734;
wire net_2248;
wire net_2270;
wire net_1667;
wire net_4971;
wire net_11532;
wire net_7208;
wire net_3866;
wire net_8882;
wire x5143;
wire net_1606;
wire net_6772;
wire net_3710;
wire net_13473;
wire net_7787;
wire net_13223;
wire net_15156;
wire net_14548;
wire net_12024;
wire net_3054;
wire net_12920;
wire net_4300;
wire net_9578;
wire net_7683;
wire net_4776;
wire net_8765;
wire net_3978;
wire net_10477;
wire net_4752;
wire net_15403;
wire net_12708;
wire net_15704;
wire net_15167;
wire net_13820;
wire net_2868;
wire net_2029;
wire net_6083;
wire net_5328;
wire net_3698;
wire net_15074;
wire net_8295;
wire net_11560;
wire net_4629;
wire net_2946;
wire net_2587;
wire net_11373;
wire net_1284;
wire net_4397;
wire net_2959;
wire net_13977;
wire net_13732;
wire net_11836;
wire net_1888;
wire net_13095;
wire net_6671;
wire net_9974;
wire net_4311;
wire net_3929;
wire net_9942;
wire net_12583;
wire net_1792;
wire net_2496;
wire x1357;
wire net_4125;
wire net_13888;
wire net_7567;
wire net_15536;
wire net_10656;
wire net_3109;
wire net_2066;
wire net_13925;
wire net_9310;
wire net_1598;
wire net_7415;
wire net_14192;
wire net_14369;
wire net_8109;
wire net_731;
wire net_1146;
wire net_15063;
wire net_13042;
wire net_11679;
wire net_4612;
wire net_9704;
wire net_7287;
wire net_1733;
wire net_4519;
wire net_10576;
wire net_8584;
wire net_5853;
wire net_5511;
wire net_13881;
wire net_7590;
wire net_13962;
wire net_9897;
wire net_11093;
wire net_6708;
wire net_5495;
wire net_10412;
wire net_13071;
wire net_9511;
wire net_8284;
wire net_2762;
wire net_4146;
wire net_11828;
wire net_1724;
wire net_6106;
wire net_6439;
wire net_3703;
wire net_12551;
wire net_6247;
wire net_14569;
wire net_6424;
wire net_4619;
wire net_6377;
wire net_12682;
wire net_10161;
wire net_2089;
wire net_12506;
wire net_6352;
wire net_10843;
wire net_12429;
wire net_965;
wire net_12378;
wire net_3797;
wire net_15472;
wire net_15391;
wire net_9718;
wire net_3535;
wire net_12248;
wire net_1195;
wire net_2916;
wire net_11976;
wire net_8314;
wire net_8184;
wire x355;
wire net_421;
wire net_5348;
wire net_2502;
wire net_1396;
wire net_1104;
wire net_9783;
wire net_4069;
wire net_764;
wire x257;
wire net_4060;
wire net_7225;
wire net_13009;
wire net_5181;
wire net_2737;
wire net_6397;
wire net_5126;
wire net_14828;
wire net_5038;
wire net_12108;
wire net_2481;
wire net_12465;
wire net_4539;
wire net_15698;
wire net_15094;
wire net_1117;
wire net_7289;
wire net_13534;
wire net_10624;
wire net_15552;
wire x101;
wire net_6866;
wire net_7162;
wire net_13770;
wire net_8104;
wire net_3955;
wire net_14531;
wire net_14210;
wire net_2617;
wire net_1060;
wire net_5950;
wire net_12699;
wire net_11893;
wire net_8246;
wire net_9157;
wire net_4846;
wire x494;
wire net_5503;
wire net_7252;
wire net_8303;
wire net_2235;
wire net_11007;
wire net_12101;
wire net_11329;
wire net_1715;
wire net_5846;
wire net_2080;
wire net_3675;
wire net_9913;
wire net_14842;
wire net_2711;
wire net_6714;
wire net_2097;
wire net_7583;
wire net_9234;
wire net_6194;
wire net_11120;
wire net_15221;
wire net_14557;
wire net_6577;
wire net_3619;
wire net_1216;
wire net_4599;
wire net_14583;
wire net_2815;
wire x3645;
wire net_15040;
wire net_3785;
wire net_11240;
wire net_1271;
wire net_1086;
wire net_15362;
wire net_1782;
wire net_9593;
wire net_10978;
wire net_11191;
wire net_8450;
wire net_13453;
wire net_1197;
wire net_7613;
wire net_1278;
wire net_273;
wire net_4863;
wire net_5744;
wire net_5858;
wire x3675;
wire net_11752;
wire net_4714;
wire net_6430;
wire net_3182;
wire net_576;
wire net_8932;
wire net_1654;
wire net_12643;
wire net_2098;
wire net_3355;
wire net_177;
wire net_4232;
wire net_8438;
wire net_3005;
wire net_4305;
wire net_11183;
wire net_7806;
wire net_12902;
wire net_8739;
wire net_10679;
wire net_2803;
wire net_3301;
wire net_11272;
wire net_725;
wire net_12133;
wire net_6370;
wire net_3931;
wire net_6090;
wire net_953;
wire net_6183;
wire net_11600;
wire net_14766;
wire net_11171;
wire net_894;
wire net_1074;
wire net_13914;
wire net_10545;
wire net_1058;
wire net_7186;
wire net_12728;
wire net_11295;
wire net_9535;
wire net_1423;
wire net_13012;
wire net_2902;
wire net_1871;
wire net_517;
wire net_628;
wire net_14004;
wire net_9064;
wire x1215;
wire net_6159;
wire net_3494;
wire net_2489;
wire net_6962;
wire net_6600;
wire net_12123;
wire net_10377;
wire net_14018;
wire net_10204;
wire net_9555;
wire net_9036;
wire net_13829;
wire net_3160;
wire net_2125;
wire net_7622;
wire net_6406;
wire net_10322;
wire net_8179;
wire net_1289;
wire net_9546;
wire net_13078;
wire net_3138;
wire net_14858;
wire net_11982;
wire net_2623;
wire net_13377;
wire net_8448;
wire net_261;
wire net_10654;
wire net_12867;
wire net_2362;
wire x3733;
wire net_6922;
wire net_12837;
wire net_11162;
wire net_5895;
wire net_8869;
wire net_12446;
wire net_4456;
wire net_5876;
wire net_4354;
wire net_1955;
wire net_5111;
wire net_2723;
wire net_15144;
wire net_5157;
wire net_13504;
wire net_2552;
wire net_8507;
wire net_8196;
wire net_3229;
wire net_1001;
wire net_13778;
wire net_3765;
wire net_781;
wire net_12886;
wire net_8479;
wire net_9729;
wire net_15323;
wire net_13063;
wire net_5241;
wire net_7506;
wire net_3012;
wire net_5967;
wire net_13134;
wire net_6818;
wire x27;
wire net_13188;
wire net_6014;
wire net_5367;
wire net_3754;
wire net_10432;
wire net_185;
wire net_7357;
wire net_6075;
wire net_9935;
wire net_14687;
wire net_11356;
wire net_3989;
wire net_13902;
wire net_10515;
wire x1743;
wire net_7304;
wire net_11312;
wire net_10875;
wire net_4321;
wire net_4631;
wire net_5285;
wire net_1994;
wire net_1015;
wire net_10499;
wire net_2980;
wire net_8574;
wire net_14685;
wire net_4668;
wire net_3897;
wire net_9863;
wire net_9288;
wire net_3960;
wire net_91;
wire net_4374;
wire net_3992;
wire net_6152;
wire net_9772;
wire net_2287;
wire net_14590;
wire net_4211;
wire net_11964;
wire net_5794;
wire net_448;
wire net_14748;
wire net_8224;
wire net_886;
wire net_7766;
wire net_3189;
wire net_11759;
wire net_6856;
wire net_15660;
wire net_2988;
wire net_2146;
wire net_405;
wire net_11927;
wire net_6811;
wire net_1111;
wire net_4592;
wire net_11614;
wire net_2651;
wire net_4281;
wire net_8259;
wire net_5279;
wire net_3651;
wire net_3971;
wire net_12182;
wire net_3155;
wire net_14345;
wire net_9059;
wire net_11440;
wire net_7969;
wire net_1470;
wire net_14053;
wire net_13358;
wire net_4627;
wire net_4423;
wire net_831;
wire net_4728;
wire net_5442;
wire net_15348;
wire net_15373;
wire net_14796;
wire net_451;
wire net_13674;
wire net_4233;
wire net_1234;
wire net_750;
wire net_12558;
wire net_4796;
wire net_7650;
wire net_15057;
wire net_8289;
wire net_7835;
wire net_9746;
wire net_15148;
wire net_13662;
wire net_2778;
wire net_2756;
wire net_12896;
wire net_13027;
wire net_12797;
wire net_7274;
wire net_14641;
wire net_11459;
wire net_9605;
wire net_8571;
wire net_1085;
wire net_5915;
wire net_5184;
wire net_592;
wire net_9528;
wire net_8983;
wire net_5788;
wire net_11920;
wire net_8472;
wire net_773;
wire net_4759;
wire net_7531;
wire net_2266;
wire net_11770;
wire net_281;
wire net_9590;
wire net_12493;
wire net_8337;
wire net_14699;
wire net_5254;
wire net_5193;
wire net_11796;
wire net_11622;
wire net_5235;
wire net_8537;
wire net_12098;
wire net_3727;
wire net_13986;
wire net_5520;
wire net_6766;
wire net_13269;
wire net_6355;
wire net_5052;
wire net_15344;
wire net_14400;
wire net_9997;
wire net_10801;
wire net_13532;
wire net_10281;
wire net_8305;
wire net_14091;
wire net_4205;
wire net_526;
wire net_2718;
wire net_834;
wire net_10298;
wire net_694;
wire net_13123;
wire net_13615;
wire net_13556;
wire net_2747;
wire net_13794;
wire net_5925;
wire net_14365;
wire net_9950;
wire net_7609;
wire net_12271;
wire net_9232;
wire net_8778;
wire net_8946;
wire net_8409;
wire net_974;
wire net_1570;
wire net_12348;
wire net_13385;
wire net_4645;
wire net_11777;
wire net_11100;
wire net_13853;
wire net_923;
wire net_10947;
wire net_1707;
wire net_12204;
wire net_9499;
wire net_2190;
wire net_4566;
wire net_1881;
wire net_11228;
wire net_7014;
wire net_10487;
wire net_111;
wire net_7320;
wire net_10900;
wire net_12925;
wire net_8779;
wire net_124;
wire net_252;
wire net_10497;
wire net_3323;
wire net_11697;
wire net_6347;
wire net_7693;
wire net_14897;
wire net_7867;
wire net_2399;
wire net_14508;
wire net_11073;
wire net_8961;
wire net_901;
wire net_6267;
wire net_7846;
wire net_3425;
wire net_12221;
wire net_410;
wire net_1492;
wire net_8134;
wire x6445;
wire net_14312;
wire net_4243;
wire net_6179;
wire net_14940;
wire net_10585;
wire net_10539;
wire net_6363;
wire net_9275;
wire net_8267;
wire x121;
wire net_9136;
wire net_2537;
wire net_11088;
wire net_6798;
wire net_14904;
wire net_6607;
wire net_3767;
wire net_6919;
wire net_12470;
wire net_6408;
wire net_7886;
wire net_4105;
wire net_11984;
wire x4694;
wire net_11397;
wire net_2603;
wire net_5910;
wire net_7824;
wire net_1132;
wire net_5594;
wire net_14144;
wire net_5880;
wire net_6132;
wire net_10351;
wire net_9553;
wire net_9193;
wire net_2442;
wire net_4569;
wire net_5754;
wire net_3026;
wire net_7743;
wire net_13749;
wire net_12317;
wire net_9410;
wire net_5760;
wire net_5923;
wire net_13000;
wire net_2356;
wire net_3288;
wire net_971;
wire net_6214;
wire net_9798;
wire net_11558;
wire net_8194;
wire net_2273;
wire net_2049;
wire net_617;
wire net_11734;
wire net_11026;
wire net_2184;
wire net_6030;
wire net_13456;
wire net_11824;
wire net_8656;
wire net_554;
wire net_14544;
wire net_13625;
wire net_4176;
wire net_4653;
wire net_14232;
wire net_11187;
wire net_8704;
wire net_3740;
wire net_15278;
wire net_14221;
wire net_8317;
wire net_4032;
wire net_4154;
wire net_9294;
wire net_6306;
wire net_9413;
wire net_584;
wire net_13753;
wire net_10446;
wire net_12656;
wire net_10420;
wire net_9794;
wire net_7877;
wire net_9000;
wire net_5917;
wire net_2411;
wire net_3870;
wire net_5709;
wire net_6254;
wire net_13104;
wire net_11511;
wire net_5456;
wire net_165;
wire net_9226;
wire net_15662;
wire net_7105;
wire net_14794;
wire net_8310;
wire net_3438;
wire net_5946;
wire net_3824;
wire net_11662;
wire net_14481;
wire net_8789;
wire net_8742;
wire net_4440;
wire net_6854;
wire net_14132;
wire net_12216;
wire net_8576;
wire net_13766;
wire net_10082;
wire net_13612;
wire net_10170;
wire net_384;
wire x769;
wire net_12970;
wire net_3823;
wire net_9886;
wire net_4191;
wire net_8600;
wire net_3503;
wire net_5792;
wire net_9365;
wire net_13573;
wire net_13366;
wire net_3859;
wire net_15136;
wire net_8044;
wire net_2599;
wire net_2665;
wire net_9200;
wire net_3642;
wire net_15350;
wire net_7885;
wire net_3803;
wire net_2707;
wire net_8607;
wire net_7426;
wire net_11284;
wire net_485;
wire net_15395;
wire net_14338;
wire net_14592;
wire net_11179;
wire net_8880;
wire net_8592;
wire net_7707;
wire net_3334;
wire net_6789;
wire net_3224;
wire net_7772;
wire net_1719;
wire net_15613;
wire net_15030;
wire net_7348;
wire net_11364;
wire net_5715;
wire net_11562;
wire x3507;
wire net_15739;
wire net_11589;
wire net_11081;
wire net_125;
wire net_11464;
wire net_9329;
wire net_15426;
wire net_13402;
wire net_8786;
wire net_14448;
wire net_8034;
wire net_11598;
wire net_2440;
wire net_1685;
wire net_9386;
wire net_6809;
wire net_14043;
wire net_12800;
wire net_4768;
wire net_1379;
wire net_1322;
wire net_12019;
wire net_14239;
wire net_13147;
wire net_2644;
wire net_6102;
wire net_12815;
wire net_14437;
wire net_9538;
wire net_13093;
wire net_8526;
wire net_12143;
wire net_10373;
wire net_1301;
wire net_12066;
wire net_14258;
wire net_12686;
wire net_286;
wire net_11668;
wire net_12487;
wire net_8749;
wire net_7596;
wire net_3584;
wire net_12756;
wire net_7051;
wire net_7247;
wire net_11591;
wire net_5588;
wire net_6932;
wire net_4999;
wire net_7116;
wire net_426;
wire net_5203;
wire net_10275;
wire net_4340;
wire net_4954;
wire net_6095;
wire net_14511;
wire net_414;
wire net_5878;
wire net_15588;
wire net_10277;
wire net_7793;
wire net_1048;
wire net_3048;
wire net_799;
wire net_5102;
wire net_3475;
wire net_8423;
wire net_5576;
wire net_14142;
wire net_15367;
wire net_5832;
wire net_5737;
wire net_12588;
wire net_2014;
wire net_9070;
wire net_8232;
wire net_12608;
wire net_1951;
wire net_7292;
wire net_12724;
wire net_15608;
wire net_9759;
wire net_8976;
wire net_6747;
wire net_13487;
wire net_5999;
wire net_7661;
wire net_15576;
wire net_12000;
wire net_11869;
wire net_9845;
wire net_5567;
wire net_2558;
wire net_4742;
wire net_2454;
wire net_8917;
wire net_8716;
wire net_2040;
wire x1911;
wire x3194;
wire net_1508;
wire net_3379;
wire net_4761;
wire net_14709;
wire net_931;
wire net_4466;
wire net_5983;
wire net_2242;
wire net_8505;
wire net_7672;
wire net_759;
wire net_6802;
wire net_7616;
wire net_15701;
wire net_6016;
wire net_7852;
wire net_11711;
wire net_11155;
wire net_8832;
wire net_10140;
wire net_12621;
wire x86;
wire net_8083;
wire net_247;
wire net_14630;
wire net_6428;
wire net_6742;
wire net_5242;
wire net_12573;
wire net_3413;
wire net_6516;
wire net_6924;
wire net_14430;
wire net_14585;
wire net_9742;
wire net_8619;
wire net_1341;
wire net_12627;
wire net_4541;
wire net_1934;
wire net_5210;
wire net_14180;
wire net_8138;
wire net_3242;
wire net_1835;
wire net_13740;
wire net_12513;
wire net_6235;
wire net_11327;
wire net_1848;
wire net_333;
wire net_15013;
wire net_639;
wire net_4724;
wire net_14491;
wire net_9583;
wire net_9322;
wire net_9114;
wire net_12309;
wire net_5697;
wire net_1238;
wire net_15203;
wire net_14923;
wire net_15184;
wire net_13697;
wire net_4664;
wire net_14074;
wire net_13547;
wire net_5976;
wire net_7599;
wire net_9483;
wire net_1033;
wire net_10155;
wire net_3923;
wire net_10604;
wire net_8839;
wire net_5560;
wire net_12458;
wire net_11333;
wire net_8333;
wire net_7210;
wire net_13149;
wire net_2554;
wire net_12196;
wire net_4479;
wire x1066;
wire net_15708;
wire net_15163;
wire net_12005;
wire net_7931;
wire net_14453;
wire net_12302;
wire net_3107;
wire net_7069;
wire net_14100;
wire net_9716;
wire net_1686;
wire net_11860;
wire net_11481;
wire net_10686;
wire net_10263;
wire net_367;
wire net_3303;
wire net_6354;
wire net_13630;
wire net_9381;
wire net_10928;
wire net_6296;
wire x3349;
wire net_10316;
wire net_10061;
wire net_1842;
wire net_7980;
wire x3828;
wire net_204;
wire net_14885;
wire net_9849;
wire net_13037;
wire net_8774;
wire net_3957;
wire net_1180;
wire net_8561;
wire net_1627;
wire net_4596;
wire net_13065;
wire net_12932;
wire net_10235;
wire net_5869;
wire net_2002;
wire net_1069;
wire net_2022;
wire net_9932;
wire net_12014;
wire net_14750;
wire net_5406;
wire net_2385;
wire net_7626;
wire net_3431;
wire net_7382;
wire net_5829;
wire net_3565;
wire net_7009;
wire net_15461;
wire net_14942;
wire net_1416;
wire net_7656;
wire net_15239;
wire net_13484;
wire net_12045;
wire net_5416;
wire net_6065;
wire net_2433;
wire x293;
wire net_8142;
wire net_15111;
wire net_6726;
wire net_10784;
wire net_4029;
wire net_93;
wire net_1601;
wire net_1916;
wire net_14808;
wire net_11419;
wire net_2468;
wire net_6614;
wire net_4087;
wire net_4255;
wire net_15306;
wire net_9854;
wire net_13437;
wire net_8866;
wire net_348;
wire net_7073;
wire net_7398;
wire net_14416;
wire net_9667;
wire net_626;
wire net_10796;
wire net_10953;
wire net_15260;
wire net_5068;
wire net_11257;
wire net_100;
wire net_1809;
wire net_2195;
wire net_686;
wire net_1615;
wire net_11546;
wire net_11246;
wire net_3421;
wire net_1691;
wire net_10089;
wire net_14037;
wire net_7859;
wire net_9197;
wire net_4578;
wire net_2112;
wire net_5072;
wire net_595;
wire net_12312;
wire net_14505;
wire net_1320;
wire net_1828;
wire net_9461;
wire net_1466;
wire net_5320;
wire net_10438;
wire net_9573;
wire net_7434;
wire net_11268;
wire net_8960;
wire net_157;
wire net_6960;
wire net_1710;
wire net_10994;
wire net_14274;
wire net_11456;
wire net_9017;
wire net_11922;
wire net_6695;
wire net_9006;
wire net_7759;
wire net_15742;
wire net_11443;
wire net_1205;
wire net_11627;
wire net_10524;
wire net_8154;
wire net_5988;
wire net_6978;
wire net_466;
wire net_6969;
wire net_9612;
wire net_1179;
wire net_4336;
wire net_9601;
wire net_15699;
wire net_13030;
wire net_15231;
wire net_4161;
wire net_3039;
wire net_7833;
wire net_13057;
wire net_6207;
wire net_11021;
wire net_2217;
wire net_938;
wire net_1610;
wire net_1761;
wire net_12163;
wire net_3569;
wire net_5682;
wire net_4683;
wire net_183;
wire net_6814;
wire net_13236;
wire net_4246;
wire net_1440;
wire net_7330;
wire net_8893;
wire net_4020;
wire net_6539;
wire net_8389;
wire net_4453;
wire net_15593;
wire net_11018;
wire net_1011;
wire net_8792;
wire net_7118;
wire net_9902;
wire net_1355;
wire net_7040;
wire net_8420;
wire net_800;
wire net_9221;
wire net_644;
wire net_13495;
wire net_12111;
wire net_8847;
wire net_13586;
wire net_12063;
wire net_12750;
wire net_852;
wire net_5992;
wire net_11917;
wire net_11035;
wire net_15118;
wire net_11648;
wire net_9405;
wire net_4046;
wire net_2580;
wire net_14771;
wire net_13834;
wire net_7391;
wire net_13997;
wire net_9696;
wire net_8904;
wire net_13302;
wire net_9961;
wire net_8416;
wire net_8382;
wire net_1385;
wire net_1643;
wire net_1919;
wire net_1534;
wire net_11404;
wire net_15029;
wire net_9836;
wire net_14690;
wire net_14284;
wire net_12843;
wire net_10128;
wire net_8992;
wire net_14162;
wire net_8685;
wire net_11492;
wire net_9491;
wire net_8555;
wire net_4876;
wire net_11410;
wire net_14860;
wire net_9087;
wire net_659;
wire net_8993;
wire net_5871;
wire net_14652;
wire net_14061;
wire net_899;
wire net_1010;
wire net_15243;
wire net_1693;
wire net_10224;
wire net_13883;
wire net_10707;
wire net_3654;
wire net_8853;
wire net_10139;
wire net_3779;
wire net_15542;
wire net_15082;
wire net_4252;
wire net_2908;
wire net_14830;
wire net_2068;
wire net_4981;
wire net_14659;
wire net_3705;
wire net_5907;
wire net_14566;
wire net_11821;
wire net_15020;
wire net_5930;
wire net_6371;
wire net_14576;
wire net_13780;
wire net_13594;
wire net_13813;
wire net_4449;
wire net_11929;
wire net_8939;
wire net_6458;
wire net_7339;
wire net_2675;
wire net_13528;
wire net_2794;
wire net_13567;
wire net_6986;
wire net_15692;
wire net_314;
wire net_1752;
wire net_5395;
wire net_2527;
wire net_15301;
wire net_11906;
wire net_11381;
wire net_9765;
wire net_14478;
wire net_2091;
wire net_2406;
wire net_6289;
wire net_8722;
wire net_12033;
wire net_14964;
wire net_8442;
wire net_4669;
wire net_807;
wire net_3405;
wire net_15456;
wire net_13791;
wire net_12422;
wire net_3270;
wire net_12665;
wire net_5460;
wire net_12479;
wire net_4286;
wire net_6880;
wire net_10238;
wire net_9872;
wire net_3484;
wire net_2474;
wire net_13931;
wire net_945;
wire net_6532;
wire net_2530;
wire net_4380;
wire net_6971;
wire net_12266;
wire net_11578;
wire net_2101;
wire net_7738;
wire net_9472;
wire net_6192;
wire net_6863;
wire net_11451;
wire net_8875;
wire net_8376;
wire net_217;
wire net_7679;
wire net_15246;
wire net_14935;
wire net_6582;
wire net_5800;
wire net_5601;
wire net_5336;
wire net_12086;
wire net_15312;
wire net_13426;
wire net_8844;
wire net_915;
wire net_2226;
wire net_5634;
wire net_3849;
wire net_8099;
wire net_12251;
wire net_8909;
wire net_8808;
wire net_6340;
wire net_8028;
wire net_13256;
wire net_10516;
wire net_9099;
wire net_5174;
wire net_11343;
wire net_8943;
wire net_1784;
wire net_15479;
wire net_14700;
wire net_1296;
wire net_8369;
wire net_15738;
wire net_13081;
wire net_4326;
wire net_2863;
wire net_3507;
wire net_1165;
wire net_5167;
wire net_10245;
wire net_677;
wire net_7159;
wire net_10762;
wire net_1472;
wire net_9735;
wire net_2939;
wire net_13294;
wire net_2424;
wire net_1113;
wire net_1968;
wire net_9945;
wire x4587;
wire net_15364;
wire net_10746;
wire net_10407;
wire net_12291;
wire net_11208;
wire net_4488;
wire net_11619;
wire net_5092;
wire net_5295;
wire net_15316;
wire net_7464;
wire net_8362;
wire net_11040;
wire net_7713;
wire net_2507;
wire net_5120;
wire net_15197;
wire net_14969;
wire net_9633;
wire net_5948;
wire net_15484;
wire net_13908;
wire net_2685;
wire net_5676;
wire net_8357;
wire net_8340;
wire net_14264;
wire net_2898;
wire net_2658;
wire net_6197;
wire net_2174;
wire net_1391;
wire net_9334;
wire net_14875;
wire net_14933;
wire net_9926;
wire net_5132;
wire net_10304;
wire net_784;
wire net_14847;
wire net_1772;
wire net_14552;
wire net_3529;
wire net_6128;
wire net_5437;
wire net_8481;
wire net_8751;
wire net_2498;
wire net_381;
wire net_6021;
wire net_9144;
wire net_6574;
wire net_6889;
wire net_2326;
wire net_11566;
wire net_10710;
wire net_8094;
wire net_3540;
wire net_3783;
wire net_11234;
wire net_1857;
wire net_7445;
wire net_5375;
wire net_11586;
wire net_11010;
wire net_9489;
wire net_12078;
wire net_12059;
wire net_6109;
wire net_15554;
wire net_14414;
wire net_9883;
wire net_3238;
wire net_1318;
wire net_10677;
wire net_15486;
wire net_15227;
wire net_1557;
wire net_6843;
wire net_3852;
wire net_1514;
wire net_7668;
wire net_13072;
wire net_6825;
wire net_13874;
wire net_7155;
wire net_3092;
wire net_14407;
wire net_3575;
wire net_4349;
wire net_9209;
wire net_11195;
wire net_8802;
wire net_6995;
wire net_8023;
wire net_15039;
wire net_6440;
wire net_306;
wire net_4984;
wire net_4516;
wire net_13240;
wire net_9026;
wire net_5371;
wire net_12241;
wire net_500;
wire net_5061;
wire net_5357;
wire net_1906;
wire net_6471;
wire net_9094;
wire net_2610;
wire net_8056;
wire net_5660;
wire net_15410;
wire net_4432;
wire net_14391;
wire net_1329;
wire net_4584;
wire net_362;
wire net_11967;
wire net_3127;
wire net_9959;
wire net_1052;
wire net_14197;
wire net_10911;
wire net_3831;
wire net_14120;
wire net_13974;
wire net_11180;
wire net_14717;
wire net_10130;
wire net_11974;
wire net_9477;
wire net_4401;
wire net_15271;
wire net_3632;
wire net_2189;
wire net_15083;
wire net_2057;
wire net_4859;
wire net_226;
wire net_1124;
wire net_6413;
wire net_13945;
wire net_7645;
wire net_13737;
wire net_5960;
wire net_5615;
wire net_143;
wire net_12434;
wire net_9160;
wire net_190;
wire net_4964;
wire net_7015;
wire net_2887;
wire net_1447;
wire net_15515;
wire net_4207;
wire net_1929;
wire net_7741;
wire net_1983;
wire net_10129;
wire net_8735;
wire net_10248;
wire net_9423;
wire net_3493;
wire net_3030;
wire net_2061;
wire net_13466;
wire net_5288;
wire net_13956;
wire net_10251;
wire net_14030;
wire net_13910;
wire net_13727;
wire net_3842;
wire net_15433;
wire net_14780;
wire net_13710;
wire net_4266;
wire net_1553;
wire net_1895;
wire net_5360;
wire net_509;
wire net_14983;
wire net_4975;
wire net_13421;
wire net_10563;
wire net_9983;
wire net_8819;
wire net_2491;
wire net_211;
wire net_3208;
wire net_2704;
wire net_13430;
wire net_10079;
wire net_6752;
wire net_14564;
wire net_10933;
wire net_15591;
wire net_14663;
wire net_5771;
wire net_5819;
wire net_13541;
wire net_3910;
wire net_1851;
wire net_3941;
wire net_6630;
wire net_13684;
wire net_12604;
wire net_8645;
wire net_10976;
wire net_3445;
wire net_2233;
wire net_8709;
wire net_2941;
wire net_2033;
wire net_12726;
wire net_12091;
wire net_8487;
wire net_3348;
wire net_477;
wire net_15710;
wire net_2123;
wire net_10811;
wire net_12784;
wire net_2943;
wire net_12360;
wire net_9377;
wire net_9049;
wire net_3861;
wire net_5970;
wire net_10892;
wire net_2532;
wire net_6758;
wire net_6905;
wire net_2315;
wire net_8325;
wire net_12785;
wire net_15501;
wire net_13851;
wire net_2231;
wire net_11112;
wire net_1864;
wire net_14646;
wire net_15441;
wire net_14917;
wire net_11725;
wire net_3812;
wire net_1200;
wire net_6156;
wire net_12840;
wire net_9595;
wire net_2518;
wire net_14604;
wire net_9509;
wire net_6950;
wire net_10663;
wire net_12329;
wire net_4062;
wire net_7558;
wire x926;
wire net_12284;
wire net_14353;
wire net_7953;
wire net_1646;
wire net_4115;
wire net_11437;
wire net_11135;
wire net_2776;
wire net_13980;
wire net_11487;
wire net_3389;
wire net_3437;
wire net_12938;
wire net_1562;
wire net_15225;
wire net_2522;
wire net_472;
wire net_14286;
wire net_1510;
wire net_4178;
wire net_14022;
wire net_3077;
wire net_7267;
wire net_8671;
wire net_8639;
wire net_13608;
wire net_4829;
wire net_13878;
wire net_136;
wire net_12987;
wire net_9430;
wire net_1524;
wire net_4171;
wire net_1528;
wire net_10022;
wire net_13579;
wire net_12676;
wire net_15628;
wire net_9396;
wire net_1749;
wire net_15686;
wire net_3367;
wire net_4915;
wire net_8386;
wire net_4784;
wire net_12355;
wire net_601;
wire net_12531;
wire net_9785;
wire net_1362;
wire net_11670;
wire net_2346;
wire net_4385;
wire net_6461;
wire net_9315;
wire net_2511;
wire net_829;
wire net_13025;
wire net_2626;
wire net_12396;
wire net_11856;
wire net_2294;
wire net_2115;
wire net_4110;
wire net_4317;
wire net_13867;
wire net_2299;
wire net_14174;
wire net_4978;
wire net_9307;
wire net_10612;
wire net_2393;
wire net_7123;
wire net_15171;
wire net_3917;
wire net_8812;
wire net_8539;
wire net_13671;
wire net_3376;
wire net_7979;
wire net_1405;
wire net_13845;
wire net_7726;
wire net_14926;
wire net_10072;
wire net_15090;
wire net_13518;
wire net_7218;
wire net_10881;
wire net_6555;
wire net_5319;
wire net_15102;
wire net_716;
wire net_5147;
wire net_13273;
wire net_13200;
wire net_10489;
wire net_11445;
wire net_11045;
wire net_1269;
wire net_6357;
wire net_13757;
wire net_8630;
wire net_3750;
wire net_12637;
wire net_5314;
wire net_3715;
wire net_3533;
wire net_5400;
wire net_5749;
wire net_12736;
wire net_11805;
wire net_10464;
wire net_9687;
wire net_2696;
wire net_14168;
wire net_6026;
wire net_8457;
wire net_10457;
wire net_12406;
wire net_1449;
wire net_4293;
wire net_9176;
wire net_6984;
wire net_5618;
wire net_15740;
wire net_666;
wire net_5310;
wire net_9725;
wire net_8620;
wire net_13114;
wire net_13776;
wire net_4809;
wire net_11308;
wire net_14729;
wire net_12989;
wire net_12706;
wire net_12184;
wire net_1220;
wire net_6212;
wire net_12343;
wire net_11394;
wire net_9702;
wire net_4017;
wire net_4693;
wire net_15125;
wire net_3946;
wire net_10596;
wire net_10194;
wire net_6346;
wire net_5522;
wire net_6319;
wire net_7636;
wire net_12716;
wire net_9024;
wire net_9824;
wire net_1657;
wire net_6063;
wire net_11781;
wire net_3084;
wire x106;
wire net_4945;
wire net_10689;
wire net_10863;
wire net_15097;
wire net_14208;
wire net_9859;
wire net_2334;
wire net_1367;
wire net_3994;
wire net_11764;
wire net_7943;
wire net_14213;
wire net_13645;
wire net_1976;
wire net_7960;
wire net_8510;
wire net_3169;
wire net_14734;
wire net_5647;
wire net_4079;
wire net_3792;
wire net_12104;
wire net_1371;
wire net_13511;
wire net_12542;
wire net_2758;
wire net_9972;
wire net_117;
wire net_8054;
wire net_1826;
wire net_5002;
wire net_6609;
wire net_7837;
wire net_14634;
wire x3889;
wire net_4609;
wire net_10337;
wire net_6517;
wire net_15526;
wire net_2142;
wire net_4704;
wire net_5782;
wire net_11841;
wire net_9843;
wire net_15335;
wire net_7864;
wire net_11885;
wire net_7332;
wire net_920;
wire net_10359;
wire net_11826;
wire net_1461;
wire net_3009;
wire net_12980;
wire net_12799;
wire net_5596;
wire net_7512;
wire net_15653;
wire net_4226;
wire net_3177;
wire net_820;
wire net_7137;
wire net_11249;
wire net_11325;
wire net_8270;
wire net_14526;
wire net_12556;
wire net_10011;
wire net_9459;
wire net_7222;
wire net_13447;
wire net_8891;
wire net_10360;
wire net_6137;
wire net_13465;
wire net_10475;
wire net_10568;
wire net_437;
wire net_3573;
wire net_13208;
wire net_5959;
wire net_9681;
wire net_566;
wire net_10390;
wire net_9861;
wire net_11477;
wire net_5063;
wire net_7519;
wire net_9071;
wire net_7371;
wire net_12498;
wire net_10855;
wire net_7140;
wire net_9768;
wire net_624;
wire net_2148;
wire net_15669;
wire net_13173;
wire net_13811;
wire x3772;
wire net_14427;
wire net_11616;
wire net_4735;
wire net_8517;
wire net_2108;
wire net_14063;
wire net_2529;
wire net_688;
wire net_6005;
wire net_6044;
wire net_4685;
wire net_4732;
wire net_9751;
wire net_8732;
wire net_5808;
wire net_8390;
wire net_5979;
wire net_7551;
wire net_11810;
wire net_8170;
wire net_3027;
wire net_12777;
wire net_14464;
wire net_5343;
wire net_14279;
wire net_15659;
wire net_6625;
wire net_4235;
wire net_15570;
wire net_14117;
wire net_11871;
wire net_14990;
wire net_9940;
wire net_13379;
wire net_4096;
wire net_5497;
wire net_7924;
wire net_9452;
wire x437;
wire net_4117;
wire net_1357;
wire net_5214;
wire net_13990;
wire net_3986;
wire net_4822;
wire net_3637;
wire net_11754;
wire net_5554;
wire net_1243;
wire net_7482;
wire net_12035;
wire net_1660;
wire net_6839;
wire net_1484;
wire net_5864;
wire net_14476;
wire net_8668;
wire net_4604;
wire net_7489;
wire net_6558;
wire net_12598;
wire net_3667;
wire net_419;
wire net_9949;
wire net_6566;
wire net_6041;
wire net_1635;
wire net_12463;
wire x3599;
wire net_5027;
wire net_6779;
wire net_4840;
wire net_5658;
wire net_936;
wire net_12697;
wire net_15400;
wire net_9259;
wire net_8066;
wire net_7808;
wire net_819;
wire net_7133;
wire net_10969;
wire net_11954;
wire net_8241;
wire net_14121;
wire net_9106;
wire net_8828;
wire net_7523;
wire net_13653;
wire net_10306;
wire net_6871;
wire net_7174;
wire net_7020;
wire net_4070;
wire net_9327;
wire net_3002;
wire net_854;
wire net_11173;
wire net_8713;
wire net_2619;
wire net_6272;
wire net_3141;
wire net_5559;
wire net_1670;
wire net_15585;
wire net_2221;
wire net_11424;
wire net_4274;
wire net_3265;
wire net_2801;
wire net_10369;
wire net_5264;
wire net_6959;
wire net_2932;
wire net_4951;
wire net_6447;
wire net_7789;
wire net_13342;
wire net_12420;
wire net_7928;
wire net_8277;
wire net_9181;
wire net_5812;
wire net_1264;
wire net_8077;
wire net_5746;
wire net_4643;
wire net_13601;
wire net_9852;
wire net_332;
wire net_1745;
wire net_1679;
wire net_7364;
wire net_9058;
wire net_4883;
wire net_9300;
wire net_3148;
wire net_1229;
wire net_6316;
wire net_13739;
wire net_12746;
wire net_656;
wire net_5723;
wire net_14385;
wire net_4800;
wire net_6277;
wire net_8489;
wire net_766;
wire net_1153;
wire net_8935;
wire net_3014;
wire net_8469;
wire net_10961;
wire net_9102;
wire net_4284;
wire net_9252;
wire net_6734;
wire net_5692;
wire net_14241;
wire net_7027;
wire net_3113;
wire net_14157;
wire net_10924;
wire net_3454;
wire net_8826;
wire net_6816;
wire net_8614;
wire net_5113;
wire net_3969;
wire net_9533;
wire net_13682;
wire net_12333;
wire net_14768;
wire net_13266;
wire net_7232;
wire net_3729;
wire net_6602;
wire net_9873;
wire net_11164;
wire net_12615;
wire net_7688;
wire net_15198;
wire net_10465;
wire net_6162;
wire net_14347;
wire net_9589;
wire net_2251;
wire net_12914;
wire net_8898;
wire net_1698;
wire net_9623;
wire net_5897;
wire net_7439;
wire net_10418;
wire net_9727;
wire net_12391;
wire net_955;
wire net_1017;
wire net_2585;
wire net_14379;
wire net_14309;
wire net_15670;
wire net_1996;
wire net_7046;
wire net_13635;
wire net_1029;
wire net_15702;
wire net_14293;
wire net_13664;
wire net_13334;
wire net_9812;
wire net_9066;
wire net_412;
wire net_12566;
wire net_8887;
wire net_4798;
wire net_12762;
wire net_9869;
wire net_2986;
wire net_3162;
wire net_4034;
wire net_4791;
wire net_1873;
wire net_3801;
wire x297;
wire net_13082;
wire net_453;
wire net_7547;
wire net_11937;
wire net_10209;
wire net_3510;
wire net_11848;
wire net_10492;
wire net_5835;
wire net_3180;
wire net_3249;
wire net_15277;
wire net_14002;
wire net_10439;
wire net_2263;
wire net_6157;
wire net_6181;
wire net_3624;
wire net_734;
wire net_14152;
wire net_12564;
wire net_7967;
wire net_2544;
wire net_9391;
wire net_11596;
wire net_2086;
wire net_951;
wire net_4930;
wire net_3186;
wire net_11314;
wire net_12869;
wire net_12278;
wire net_7272;
wire net_7096;
wire net_12654;
wire net_8977;
wire net_8177;
wire net_13895;
wire net_14389;
wire net_10222;
wire net_10648;
wire net_12350;
wire net_12121;
wire net_5277;
wire net_14730;
wire net_7269;
wire net_2966;
wire net_15146;
wire net_4372;
wire net_13186;
wire net_1253;
wire net_2500;
wire net_10508;
wire net_9808;
wire net_15398;
wire net_13971;
wire net_1076;
wire net_3900;
wire net_14051;
wire net_10168;
wire net_8234;
wire net_13315;
wire net_10399;
wire net_9711;
wire net_4352;
wire net_15647;
wire net_3153;
wire net_681;
wire net_6721;
wire net_5155;
wire net_5471;
wire net_7346;
wire net_13136;
wire net_6533;
wire net_3598;
wire net_5252;
wire net_146;
wire net_9562;
wire net_8676;
wire net_3938;
wire net_7534;
wire net_11289;
wire net_5752;
wire net_4594;
wire net_9592;
wire net_1502;
wire net_15009;
wire net_4454;
wire net_6290;
wire net_4624;
wire net_11522;
wire net_11282;
wire net_6596;
wire net_7621;
wire net_428;
wire net_9675;
wire net_11065;
wire net_10557;
wire net_11306;
wire net_10329;
wire net_14816;
wire net_12138;
wire net_10117;
wire net_640;
wire net_7780;
wire net_4666;
wire net_2888;
wire net_7508;
wire net_12884;
wire net_775;
wire net_10903;
wire net_752;
wire net_14362;
wire net_3716;
wire net_535;
wire net_498;
wire net_888;
wire net_13066;
wire net_10772;
wire net_13212;
wire net_11298;
wire net_11095;
wire net_9526;
wire net_5191;
wire net_2721;
wire net_8480;
wire net_8900;
wire net_10513;
wire net_2637;
wire net_15380;
wire net_1023;
wire net_4814;
wire net_5233;
wire net_7499;
wire net_3623;
wire net_301;
wire net_4902;
wire net_6768;
wire net_2360;
wire net_5419;
wire net_3617;
wire net_12228;
wire net_299;
wire net_7432;
wire net_1343;
wire net_7147;
wire net_2285;
wire net_12894;
wire net_12690;
wire net_7355;
wire net_7413;
wire net_12387;
wire net_590;
wire net_3879;
wire net_11755;
wire net_2024;
wire net_3240;
wire net_15150;
wire net_8229;
wire net_11549;
wire net_3254;
wire net_9569;
wire net_9779;
wire net_9342;
wire net_9040;
wire net_3725;
wire net_15569;
wire net_12135;
wire net_10094;
wire net_4194;
wire net_12361;
wire net_5464;
wire net_9111;
wire net_8335;
wire net_6088;
wire net_8530;
wire net_5041;
wire net_5857;
wire net_15161;
wire net_15059;
wire net_407;
wire net_10145;
wire net_1736;
wire net_12807;
wire net_4405;
wire net_12258;
wire net_11793;
wire net_9814;
wire net_11660;
wire net_6947;
wire net_8723;
wire net_9801;
wire net_10314;
wire net_2312;
wire net_10574;
wire net_4148;
wire net_9155;
wire net_5048;
wire net_8586;
wire net_1669;
wire net_7869;
wire net_11505;
wire net_12408;
wire net_14096;
wire net_8189;
wire net_2073;
wire net_1041;
wire net_7628;
wire net_9146;
wire x348;
wire net_6385;
wire net_14027;
wire net_2950;
wire net_6056;
wire net_4057;
wire net_6108;
wire net_5851;
wire net_14350;
wire net_5105;
wire net_4778;
wire net_14244;
wire net_11211;
wire net_6081;
wire net_13159;
wire net_14975;
wire net_14863;
wire net_2364;
wire net_5507;
wire net_12173;
wire net_12526;
wire net_942;
wire net_12822;
wire net_8763;
wire net_15339;
wire net_7565;
wire net_1981;
wire x1274;
wire x906;
wire net_4302;
wire net_1218;
wire net_6245;
wire net_15042;
wire net_10606;
wire net_13658;
wire net_10917;
wire net_6436;
wire net_15201;
wire net_1494;
wire net_3286;
wire net_4415;
wire x589;
wire net_2154;
wire net_1726;
wire net_5527;
wire net_4123;
wire net_7082;
wire net_11430;
wire net_5705;
wire net_15604;
wire net_12165;
wire net_3298;
wire net_3099;
wire net_1398;
wire net_12432;
wire net_10658;
wire net_15065;
wire net_13219;
wire net_10503;
wire net_6339;
wire net_4399;
wire net_7380;
wire net_8197;
wire net_1144;
wire net_6117;
wire net_1794;
wire net_9363;
wire net_8297;
wire net_12508;
wire net_6503;
wire net_10646;
wire net_5536;
wire net_1022;
wire net_4638;
wire net_11129;
wire net_2865;
wire net_2260;
wire net_6110;
wire net_8182;
wire net_9770;
wire net_3606;
wire net_702;
wire net_4328;
wire net_3195;
wire net_1477;
wire net_3210;
wire net_13960;
wire net_13221;
wire net_3318;
wire x931;
wire net_9270;
wire net_15401;
wire net_7800;
wire net_8188;
wire net_8122;
wire net_7571;
wire net_11682;
wire net_13152;
wire net_12948;
wire net_12904;
wire net_15214;
wire net_12439;
wire net_12979;
wire net_1193;
wire net_9412;
wire net_1425;
wire net_14673;
wire net_1122;
wire net_4911;
wire net_8436;
wire net_15679;
wire net_10790;
wire net_6228;
wire net_5505;
wire net_10622;
wire net_1813;
wire net_8540;
wire net_4534;
wire net_6252;
wire net_10673;
wire net_7945;
wire net_12411;
wire net_6491;
wire net_983;
wire net_355;
wire net_13898;
wire net_13702;
wire net_4713;
wire net_7258;
wire net_9709;
wire net_9513;
wire net_8102;
wire net_15534;
wire net_12427;
wire net_9002;
wire net_723;
wire net_4307;
wire net_7311;
wire net_11341;
wire net_8292;
wire net_7614;
wire net_2483;
wire net_5513;
wire x3638;
wire net_8248;
wire net_3962;
wire net_14608;
wire net_12026;
wire net_11834;
wire net_4553;
wire net_275;
wire net_10501;
wire net_10202;
wire net_12641;
wire net_15096;
wire net_9486;
wire net_4831;
wire net_2914;
wire net_15050;
wire net_10547;
wire net_11366;
wire net_2590;
wire net_10841;
wire net_7280;
wire net_13293;
wire net_13351;
wire net_1137;
wire net_7424;
wire net_3948;
wire net_4830;
wire net_6142;
wire net_13475;
wire net_13455;
wire net_5036;
wire net_12414;
wire net_12872;
wire net_12860;
wire net_13909;
wire net_9493;
wire net_4865;
wire net_11765;
wire net_8254;
wire net_11945;
wire net_9955;
wire net_14370;
wire net_3819;
wire net_15640;
wire x366;
wire net_11978;
wire net_254;
wire net_11193;
wire net_12581;
wire net_11895;
wire net_1501;
wire net_3003;
wire net_5622;
wire net_12103;
wire net_574;
wire net_3357;
wire net_11375;
wire net_9467;
wire net_14054;
wire net_9694;
wire net_8425;

// Start cells
CLKBUF_X2 inst_12147 ( .A(net_12065), .Z(net_12066) );
OAI21_X2 inst_1783 ( .ZN(net_7674), .B2(net_7589), .A(net_7582), .B1(net_7442) );
CLKBUF_X2 inst_10910 ( .A(net_10828), .Z(net_10829) );
CLKBUF_X2 inst_13999 ( .A(net_12398), .Z(net_13918) );
INV_X2 inst_6916 ( .ZN(net_2857), .A(net_2173) );
NOR2_X2 inst_2685 ( .A2(net_10376), .A1(net_10375), .ZN(net_5213) );
AOI221_X2 inst_9876 ( .B1(net_9783), .B2(net_9098), .A(net_6940), .C2(net_6939), .ZN(net_6825), .C1(net_253) );
NAND2_X2 inst_4123 ( .A1(net_2405), .ZN(net_2329), .A2(net_1605) );
DFF_X2 inst_7766 ( .Q(net_9715), .D(net_6539), .CK(net_13431) );
INV_X2 inst_6919 ( .A(net_2534), .ZN(net_2121) );
OAI21_X2 inst_1751 ( .ZN(net_8649), .A(net_8648), .B1(net_8647), .B2(net_8615) );
CLKBUF_X2 inst_14490 ( .A(net_14408), .Z(net_14409) );
DFF_X2 inst_8140 ( .Q(net_9939), .D(net_5117), .CK(net_13187) );
INV_X4 inst_5359 ( .ZN(net_3744), .A(net_1223) );
OAI211_X2 inst_2235 ( .C1(net_7226), .C2(net_6480), .ZN(net_6469), .B(net_5552), .A(net_3679) );
OR2_X4 inst_779 ( .A1(net_2963), .A2(net_2955), .ZN(net_2953) );
CLKBUF_X2 inst_13828 ( .A(net_13746), .Z(net_13747) );
CLKBUF_X2 inst_11465 ( .A(net_11383), .Z(net_11384) );
INV_X4 inst_6439 ( .A(net_9851), .ZN(net_619) );
INV_X4 inst_5306 ( .A(net_1819), .ZN(net_1294) );
OAI211_X2 inst_2205 ( .C1(net_7186), .C2(net_6501), .ZN(net_6500), .B(net_5678), .A(net_3679) );
NOR2_X2 inst_2858 ( .ZN(net_2536), .A2(net_1182), .A1(x6351) );
AND2_X2 inst_10503 ( .ZN(net_6617), .A1(net_5960), .A2(net_5781) );
CLKBUF_X1 inst_8981 ( .A(x185142), .Z(x906) );
INV_X4 inst_5488 ( .ZN(net_6633), .A(net_1374) );
NAND2_X2 inst_4131 ( .ZN(net_2690), .A1(net_1811), .A2(net_966) );
CLKBUF_X2 inst_13591 ( .A(net_13509), .Z(net_13510) );
AOI221_X2 inst_9805 ( .B1(net_9984), .A(net_7090), .B2(net_7089), .C2(net_7088), .ZN(net_6997), .C1(net_256) );
CLKBUF_X2 inst_13926 ( .A(net_13844), .Z(net_13845) );
CLKBUF_X2 inst_15089 ( .A(net_11452), .Z(net_15008) );
XNOR2_X2 inst_214 ( .ZN(net_4685), .A(net_4271), .B(net_2653) );
CLKBUF_X2 inst_13990 ( .A(net_10589), .Z(net_13909) );
AOI22_X2 inst_9115 ( .A1(net_9669), .A2(net_6402), .ZN(net_6374), .B2(net_5263), .B1(net_107) );
NAND2_X2 inst_4228 ( .ZN(net_1639), .A2(net_1638), .A1(net_1535) );
SDFF_X2 inst_548 ( .D(net_9141), .SE(net_933), .CK(net_10652), .SI(x1911), .Q(x1170) );
CLKBUF_X2 inst_10808 ( .A(net_10559), .Z(net_10727) );
CLKBUF_X2 inst_12017 ( .A(net_11022), .Z(net_11936) );
INV_X4 inst_4647 ( .ZN(net_8659), .A(net_7038) );
NAND2_X2 inst_4372 ( .A2(net_10430), .ZN(net_1765), .A1(net_879) );
DFF_X2 inst_7408 ( .QN(net_9400), .D(net_8365), .CK(net_14030) );
INV_X2 inst_7191 ( .ZN(net_809), .A(x6577) );
CLKBUF_X2 inst_12796 ( .A(net_12714), .Z(net_12715) );
CLKBUF_X2 inst_14747 ( .A(net_14665), .Z(net_14666) );
INV_X4 inst_4709 ( .ZN(net_4738), .A(net_4620) );
AND2_X4 inst_10461 ( .A1(net_10474), .A2(net_2205), .ZN(net_1645) );
CLKBUF_X2 inst_15436 ( .A(net_15354), .Z(net_15355) );
DFF_X1 inst_8488 ( .Q(net_9956), .D(net_7886), .CK(net_14427) );
CLKBUF_X2 inst_14178 ( .A(net_14096), .Z(net_14097) );
CLKBUF_X2 inst_10820 ( .A(net_10738), .Z(net_10739) );
INV_X2 inst_7060 ( .ZN(net_1274), .A(net_1273) );
CLKBUF_X2 inst_14148 ( .A(net_12387), .Z(net_14067) );
CLKBUF_X2 inst_13127 ( .A(net_13045), .Z(net_13046) );
NAND2_X4 inst_3347 ( .A2(net_9018), .A1(net_9017), .ZN(net_8518) );
NAND4_X2 inst_3130 ( .ZN(net_2932), .A1(net_1999), .A2(net_1133), .A3(net_1047), .A4(net_918) );
CLKBUF_X2 inst_11446 ( .A(net_11364), .Z(net_11365) );
AOI22_X2 inst_9568 ( .B1(net_10300), .A1(net_9700), .B2(net_4774), .ZN(net_3751), .A2(net_3039) );
INV_X4 inst_6406 ( .A(net_9644), .ZN(net_613) );
INV_X4 inst_5341 ( .A(net_2005), .ZN(net_1248) );
NAND2_X2 inst_4136 ( .ZN(net_2220), .A1(net_2219), .A2(net_2218) );
CLKBUF_X2 inst_12400 ( .A(net_12246), .Z(net_12319) );
CLKBUF_X2 inst_12585 ( .A(net_12503), .Z(net_12504) );
AOI22_X2 inst_9372 ( .B1(net_9895), .A1(net_6808), .A2(net_5759), .B2(net_5758), .ZN(net_5533) );
OAI22_X2 inst_1228 ( .B1(net_7226), .ZN(net_4891), .A2(net_4890), .B2(net_4889), .A1(net_349) );
CLKBUF_X2 inst_13185 ( .A(net_13103), .Z(net_13104) );
AOI22_X2 inst_9653 ( .A1(net_2357), .ZN(net_2234), .A2(net_2233), .B1(net_2232), .B2(net_2231) );
INV_X4 inst_4985 ( .ZN(net_2887), .A(net_2239) );
NAND2_X2 inst_4221 ( .A2(net_4017), .ZN(net_1663), .A1(net_846) );
SDFF_X2 inst_521 ( .Q(net_9337), .D(net_9337), .SI(net_9329), .SE(net_7588), .CK(net_14690) );
INV_X4 inst_5164 ( .A(net_3746), .ZN(net_1767) );
AOI22_X2 inst_9461 ( .B1(net_10036), .A1(net_9873), .B2(net_5174), .ZN(net_3866), .A2(net_2973) );
INV_X4 inst_6534 ( .A(net_10049), .ZN(net_339) );
AOI222_X1 inst_9736 ( .B2(net_10192), .C2(net_10190), .A2(net_10189), .B1(net_10185), .C1(net_10183), .A1(net_10182), .ZN(net_1343) );
INV_X4 inst_5947 ( .ZN(net_562), .A(net_561) );
MUX2_X1 inst_4473 ( .S(net_6041), .A(net_4304), .B(x6327), .Z(x381) );
OAI221_X2 inst_1685 ( .C1(net_7226), .B2(net_5642), .ZN(net_5477), .C2(net_4905), .A(net_3507), .B1(net_986) );
NOR2_X2 inst_2511 ( .ZN(net_8454), .A2(net_8377), .A1(net_3298) );
OAI221_X2 inst_1655 ( .B1(net_7209), .C2(net_5591), .ZN(net_5519), .C1(net_5518), .B2(net_4902), .A(net_3507) );
CLKBUF_X2 inst_12320 ( .A(net_12238), .Z(net_12239) );
CLKBUF_X2 inst_10720 ( .A(net_10616), .Z(net_10639) );
AOI22_X2 inst_9038 ( .ZN(net_7428), .A2(net_6957), .B1(net_6956), .B2(net_4595), .A1(net_4594) );
INV_X2 inst_6910 ( .ZN(net_2241), .A(net_2240) );
NAND2_X2 inst_3578 ( .A2(net_7560), .ZN(net_7526), .A1(net_7525) );
CLKBUF_X2 inst_15174 ( .A(net_15092), .Z(net_15093) );
AOI22_X2 inst_9257 ( .A2(net_8042), .B2(net_8041), .A1(net_6628), .B1(net_6414), .ZN(net_6049) );
CLKBUF_X2 inst_15477 ( .A(net_10610), .Z(net_15396) );
CLKBUF_X2 inst_14731 ( .A(net_14649), .Z(net_14650) );
AOI221_X2 inst_9938 ( .B2(net_5867), .A(net_5862), .C2(net_5853), .ZN(net_5828), .C1(net_5827), .B1(x5601) );
CLKBUF_X2 inst_14165 ( .A(net_14083), .Z(net_14084) );
DFF_X2 inst_7415 ( .QN(net_9414), .D(net_8350), .CK(net_13947) );
DFF_X1 inst_8731 ( .QN(net_10136), .D(net_5883), .CK(net_10787) );
CLKBUF_X2 inst_12238 ( .A(net_11439), .Z(net_12157) );
INV_X4 inst_4847 ( .ZN(net_3295), .A(net_3294) );
INV_X4 inst_6010 ( .A(net_9229), .ZN(net_527) );
INV_X4 inst_5940 ( .A(net_586), .ZN(net_570) );
CLKBUF_X2 inst_15733 ( .A(net_15651), .Z(net_15652) );
CLKBUF_X2 inst_14010 ( .A(net_13928), .Z(net_13929) );
CLKBUF_X2 inst_13236 ( .A(net_13154), .Z(net_13155) );
OAI22_X2 inst_1066 ( .A2(net_7036), .B2(net_7035), .ZN(net_6963), .A1(net_2519), .B1(net_1698) );
CLKBUF_X2 inst_10825 ( .A(net_10553), .Z(net_10744) );
AOI221_X2 inst_9978 ( .B1(net_9945), .C1(net_9747), .B2(net_6443), .C2(net_6442), .ZN(net_4235), .A(net_3580) );
DFF_X2 inst_7977 ( .QN(net_10312), .D(net_5571), .CK(net_13323) );
NAND2_X2 inst_3392 ( .ZN(net_9004), .A1(net_8702), .A2(net_8700) );
CLKBUF_X2 inst_12122 ( .A(net_12040), .Z(net_12041) );
AND3_X2 inst_10377 ( .A3(net_10329), .A1(net_3129), .ZN(net_3124), .A2(net_1220) );
INV_X4 inst_5063 ( .A(net_2821), .ZN(net_1870) );
CLKBUF_X2 inst_15707 ( .A(net_12781), .Z(net_15626) );
INV_X4 inst_6232 ( .A(net_9981), .ZN(net_461) );
NOR4_X2 inst_2342 ( .ZN(net_3063), .A2(net_3062), .A1(net_2582), .A4(net_1854), .A3(net_668) );
INV_X4 inst_4608 ( .ZN(net_7638), .A(net_7635) );
OAI211_X2 inst_2294 ( .ZN(net_4510), .C1(net_4509), .C2(net_4508), .A(net_4225), .B(net_3087) );
AOI22_X2 inst_9143 ( .A1(net_9693), .A2(net_6420), .ZN(net_6342), .B2(net_5263), .B1(net_3249) );
CLKBUF_X2 inst_14321 ( .A(net_14239), .Z(net_14240) );
CLKBUF_X2 inst_12495 ( .A(net_12413), .Z(net_12414) );
OAI221_X2 inst_1617 ( .B1(net_10305), .C1(net_7245), .A(net_6546), .ZN(net_5593), .B2(net_5591), .C2(net_4902) );
CLKBUF_X2 inst_12553 ( .A(net_12471), .Z(net_12472) );
XNOR2_X2 inst_151 ( .ZN(net_6647), .A(net_6646), .B(net_2348) );
OAI211_X2 inst_2256 ( .C1(net_7249), .C2(net_6501), .ZN(net_6432), .B(net_5436), .A(net_3679) );
INV_X4 inst_4821 ( .ZN(net_3731), .A(net_3298) );
DFF_X1 inst_8696 ( .D(net_6768), .Q(net_116), .CK(net_15437) );
DFF_X2 inst_7519 ( .Q(net_9538), .D(net_7883), .CK(net_13986) );
NAND2_X2 inst_3931 ( .ZN(net_3730), .A2(net_3378), .A1(net_605) );
INV_X4 inst_4880 ( .ZN(net_2987), .A(net_2784) );
CLKBUF_X2 inst_12409 ( .A(net_12327), .Z(net_12328) );
CLKBUF_X2 inst_11637 ( .A(net_11555), .Z(net_11556) );
CLKBUF_X2 inst_12682 ( .A(net_12600), .Z(net_12601) );
INV_X2 inst_7239 ( .ZN(net_3246), .A(net_165) );
AND3_X2 inst_10370 ( .ZN(net_4965), .A2(net_4964), .A3(net_4689), .A1(net_4688) );
NAND2_X2 inst_3867 ( .ZN(net_4366), .A2(net_4232), .A1(net_4083) );
OAI211_X2 inst_2072 ( .C2(net_6778), .ZN(net_6777), .A(net_6346), .B(net_6094), .C1(net_5103) );
OAI221_X2 inst_1603 ( .B1(net_10218), .C1(net_7182), .B2(net_5642), .ZN(net_5633), .C2(net_4905), .A(net_3731) );
CLKBUF_X2 inst_13237 ( .A(net_12685), .Z(net_13156) );
AOI22_X2 inst_9634 ( .B1(net_10005), .A1(net_9973), .ZN(net_3408), .A2(net_2541), .B2(net_2468) );
XNOR2_X2 inst_340 ( .ZN(net_2872), .A(net_2871), .B(net_1722) );
CLKBUF_X2 inst_11590 ( .A(net_11057), .Z(net_11509) );
CLKBUF_X2 inst_14978 ( .A(net_14896), .Z(net_14897) );
CLKBUF_X2 inst_10785 ( .A(net_10622), .Z(net_10704) );
CLKBUF_X2 inst_13098 ( .A(net_11294), .Z(net_13017) );
DFF_X2 inst_8109 ( .Q(net_9940), .D(net_5116), .CK(net_12030) );
DFF_X1 inst_8864 ( .D(net_10408), .QN(net_10348), .CK(net_11157) );
CLKBUF_X2 inst_11075 ( .A(net_10993), .Z(net_10994) );
NAND2_X2 inst_4280 ( .ZN(net_2952), .A2(net_983), .A1(net_684) );
XNOR2_X2 inst_158 ( .ZN(net_6162), .A(net_5315), .B(net_1399) );
DFF_X2 inst_8171 ( .QN(net_10029), .D(net_5042), .CK(net_13694) );
DFF_X2 inst_7493 ( .Q(net_10299), .D(net_8008), .CK(net_14573) );
INV_X4 inst_5411 ( .ZN(net_1601), .A(net_1154) );
CLKBUF_X2 inst_14279 ( .A(net_14197), .Z(net_14198) );
CLKBUF_X2 inst_13529 ( .A(net_13447), .Z(net_13448) );
NAND2_X2 inst_4244 ( .A2(net_9196), .A1(net_9195), .ZN(net_1509) );
OAI221_X2 inst_1490 ( .C1(net_10418), .B2(net_9063), .C2(net_9056), .ZN(net_7373), .B1(net_7249), .A(net_7034) );
SDFF_X2 inst_507 ( .SI(net_8010), .D(net_7922), .SE(net_197), .Q(net_197), .CK(net_12840) );
CLKBUF_X2 inst_15421 ( .A(net_15339), .Z(net_15340) );
INV_X4 inst_4559 ( .ZN(net_8473), .A(net_8418) );
NAND2_X2 inst_4289 ( .ZN(net_2023), .A2(net_1334), .A1(net_1016) );
NAND2_X2 inst_3709 ( .ZN(net_5916), .A1(net_5915), .A2(net_5914) );
CLKBUF_X2 inst_14365 ( .A(net_14283), .Z(net_14284) );
AND2_X2 inst_10566 ( .ZN(net_3491), .A1(net_3024), .A2(net_3023) );
CLKBUF_X2 inst_10934 ( .A(net_10558), .Z(net_10853) );
INV_X4 inst_6319 ( .A(net_9961), .ZN(net_421) );
CLKBUF_X2 inst_12311 ( .A(net_12229), .Z(net_12230) );
OR2_X2 inst_884 ( .A2(net_7038), .ZN(net_6252), .A1(net_6251) );
OR3_X2 inst_711 ( .ZN(net_5748), .A2(net_5747), .A3(net_5365), .A1(net_5364) );
OR2_X4 inst_827 ( .A1(net_10356), .ZN(net_2716), .A2(net_885) );
INV_X4 inst_6542 ( .A(net_9959), .ZN(net_335) );
CLKBUF_X2 inst_15309 ( .A(net_14112), .Z(net_15228) );
CLKBUF_X2 inst_11477 ( .A(net_11395), .Z(net_11396) );
CLKBUF_X2 inst_14452 ( .A(net_10981), .Z(net_14371) );
AOI22_X2 inst_9573 ( .A2(net_6892), .B2(net_6625), .ZN(net_6316), .B1(net_3733), .A1(net_1144) );
CLKBUF_X2 inst_15231 ( .A(net_15149), .Z(net_15150) );
CLKBUF_X2 inst_10730 ( .A(net_10648), .Z(net_10649) );
CLKBUF_X2 inst_14845 ( .A(net_14763), .Z(net_14764) );
AND2_X2 inst_10574 ( .ZN(net_2962), .A1(net_2961), .A2(net_2960) );
INV_X2 inst_7140 ( .A(net_10356), .ZN(net_1303) );
CLKBUF_X2 inst_11213 ( .A(net_11131), .Z(net_11132) );
DFF_X1 inst_8465 ( .QN(net_9589), .D(net_7962), .CK(net_11527) );
NAND4_X2 inst_3040 ( .ZN(net_7831), .A4(net_7792), .A2(net_2868), .A3(net_1039), .A1(net_926) );
CLKBUF_X2 inst_12937 ( .A(net_12855), .Z(net_12856) );
NAND2_X2 inst_4191 ( .A1(net_4026), .ZN(net_2911), .A2(net_1850) );
NAND2_X2 inst_3870 ( .ZN(net_4630), .A2(net_4229), .A1(net_4080) );
CLKBUF_X2 inst_14171 ( .A(net_14089), .Z(net_14090) );
INV_X4 inst_5675 ( .A(net_10356), .ZN(net_810) );
NAND2_X2 inst_4269 ( .A2(net_10220), .ZN(net_2047), .A1(net_1021) );
DFF_X1 inst_8559 ( .Q(net_9869), .D(net_7120), .CK(net_15643) );
INV_X4 inst_4640 ( .A(net_7036), .ZN(net_6154) );
XOR2_X2 inst_18 ( .Z(net_2771), .B(net_2459), .A(net_1110) );
INV_X4 inst_6047 ( .A(net_9559), .ZN(net_8714) );
CLKBUF_X2 inst_15616 ( .A(net_15534), .Z(net_15535) );
NAND2_X2 inst_4128 ( .ZN(net_2924), .A2(net_2846), .A1(net_2320) );
CLKBUF_X2 inst_14534 ( .A(net_11372), .Z(net_14453) );
AOI22_X2 inst_9040 ( .A1(net_7642), .B2(net_7641), .ZN(net_7135), .A2(net_6561), .B1(net_6167) );
AOI21_X2 inst_10154 ( .ZN(net_4131), .A(net_3658), .B2(net_3229), .B1(net_2621) );
OAI211_X2 inst_2263 ( .C1(net_7129), .C2(net_6548), .ZN(net_6284), .B(net_5711), .A(net_3527) );
INV_X4 inst_5608 ( .ZN(net_1150), .A(net_875) );
INV_X4 inst_4861 ( .ZN(net_4969), .A(net_2965) );
INV_X4 inst_4796 ( .ZN(net_3665), .A(net_3664) );
INV_X4 inst_5183 ( .A(net_3744), .ZN(net_1928) );
NAND2_X2 inst_3549 ( .A2(net_9268), .ZN(net_8018), .A1(net_7875) );
CLKBUF_X2 inst_12602 ( .A(net_12520), .Z(net_12521) );
NAND2_X2 inst_3501 ( .ZN(net_8368), .A1(net_8182), .A2(net_8181) );
AOI21_X2 inst_10035 ( .B1(net_10385), .ZN(net_7863), .A(net_6677), .B2(net_263) );
NAND2_X2 inst_3936 ( .A2(net_10280), .A1(net_4015), .ZN(net_3892) );
CLKBUF_X2 inst_13029 ( .A(net_11667), .Z(net_12948) );
CLKBUF_X2 inst_13738 ( .A(net_11735), .Z(net_13657) );
NAND2_X2 inst_4175 ( .ZN(net_3050), .A1(net_1959), .A2(net_1958) );
INV_X4 inst_6069 ( .A(net_9240), .ZN(net_911) );
INV_X2 inst_6675 ( .ZN(net_8353), .A(net_8290) );
AOI221_X2 inst_9783 ( .B1(net_9973), .ZN(net_7092), .A(net_7090), .B2(net_7089), .C1(net_7088), .C2(net_245) );
DFF_X1 inst_8535 ( .Q(net_9990), .D(net_7369), .CK(net_13298) );
INV_X2 inst_7076 ( .A(net_2393), .ZN(net_1205) );
INV_X4 inst_6020 ( .A(net_10498), .ZN(net_523) );
CLKBUF_X2 inst_14217 ( .A(net_14135), .Z(net_14136) );
CLKBUF_X2 inst_12739 ( .A(net_12657), .Z(net_12658) );
INV_X2 inst_6954 ( .A(net_3710), .ZN(net_1882) );
CLKBUF_X2 inst_14663 ( .A(net_14581), .Z(net_14582) );
AOI22_X2 inst_9416 ( .A1(net_10178), .A2(net_4656), .B2(net_4655), .ZN(net_4653), .B1(x4285) );
DFF_X2 inst_7378 ( .QN(net_9371), .D(net_8665), .CK(net_14182) );
AOI22_X2 inst_9217 ( .A1(net_9935), .B1(net_9836), .B2(net_6140), .A2(net_6111), .ZN(net_6094) );
INV_X4 inst_6475 ( .A(net_10196), .ZN(net_3683) );
NAND2_X2 inst_4397 ( .A2(net_10333), .A1(net_10332), .ZN(net_1432) );
CLKBUF_X2 inst_10818 ( .A(net_10736), .Z(net_10737) );
DFF_X2 inst_7392 ( .Q(net_10065), .D(net_8573), .CK(net_11190) );
NAND4_X2 inst_3102 ( .ZN(net_4341), .A2(net_3829), .A3(net_3828), .A4(net_3680), .A1(net_3573) );
CLKBUF_X2 inst_12847 ( .A(net_12765), .Z(net_12766) );
HA_X1 inst_7364 ( .B(net_9324), .A(net_9323), .S(net_2472), .CO(net_1068) );
INV_X4 inst_5816 ( .ZN(net_1093), .A(net_676) );
NOR2_X2 inst_2695 ( .ZN(net_4599), .A2(net_4415), .A1(net_614) );
CLKBUF_X2 inst_13801 ( .A(net_13719), .Z(net_13720) );
CLKBUF_X2 inst_12748 ( .A(net_12666), .Z(net_12667) );
NAND2_X2 inst_3860 ( .ZN(net_4159), .A2(net_4158), .A1(net_1706) );
CLKBUF_X2 inst_14833 ( .A(net_14751), .Z(net_14752) );
CLKBUF_X2 inst_12515 ( .A(net_12433), .Z(net_12434) );
OAI211_X2 inst_2063 ( .B(net_7783), .C2(net_7782), .ZN(net_7739), .A(net_7676), .C1(net_2474) );
CLKBUF_X2 inst_14659 ( .A(net_12273), .Z(net_14578) );
CLKBUF_X2 inst_13635 ( .A(net_13553), .Z(net_13554) );
CLKBUF_X2 inst_14980 ( .A(net_14898), .Z(net_14899) );
CLKBUF_X2 inst_10692 ( .A(net_10598), .Z(net_10611) );
CLKBUF_X2 inst_14917 ( .A(net_14099), .Z(net_14836) );
INV_X4 inst_4801 ( .A(net_3705), .ZN(net_3658) );
CLKBUF_X2 inst_14150 ( .A(net_14068), .Z(net_14069) );
NAND2_X2 inst_3723 ( .A1(net_10504), .ZN(net_5780), .A2(net_5768) );
CLKBUF_X2 inst_13228 ( .A(net_10728), .Z(net_13147) );
NAND2_X2 inst_3521 ( .A2(net_9597), .ZN(net_8185), .A1(net_8117) );
AOI22_X2 inst_9346 ( .B1(net_9822), .A2(net_5766), .B2(net_5765), .ZN(net_5606), .A1(net_260) );
NAND2_X2 inst_3440 ( .A1(net_9446), .ZN(net_8891), .A2(net_8479) );
CLKBUF_X2 inst_15282 ( .A(net_15200), .Z(net_15201) );
CLKBUF_X2 inst_12286 ( .A(net_11764), .Z(net_12205) );
CLKBUF_X2 inst_14350 ( .A(net_12880), .Z(net_14269) );
INV_X4 inst_5386 ( .A(net_4603), .ZN(net_1483) );
NAND2_X2 inst_3985 ( .ZN(net_3237), .A2(net_3236), .A1(net_3115) );
OAI211_X2 inst_2036 ( .C2(net_8102), .B(net_8098), .ZN(net_8097), .A(net_7996), .C1(net_4191) );
INV_X4 inst_5802 ( .A(net_7025), .ZN(net_687) );
NAND2_X2 inst_4001 ( .ZN(net_4095), .A2(net_3390), .A1(net_3170) );
CLKBUF_X2 inst_12249 ( .A(net_12167), .Z(net_12168) );
CLKBUF_X2 inst_11107 ( .A(net_11025), .Z(net_11026) );
AOI221_X2 inst_9853 ( .A(net_6889), .B2(net_6888), .C2(net_6887), .ZN(net_6865), .B1(net_6514), .C1(x3949) );
DFF_X2 inst_7897 ( .QN(net_10104), .D(net_6016), .CK(net_14905) );
OAI211_X2 inst_2049 ( .C2(net_10171), .B(net_8819), .ZN(net_7839), .A(net_7764), .C1(net_6311) );
OR2_X2 inst_868 ( .ZN(net_7711), .A1(net_7548), .A2(net_7415) );
CLKBUF_X2 inst_10747 ( .A(net_10613), .Z(net_10666) );
DFF_X2 inst_8187 ( .QN(net_10258), .D(net_5193), .CK(net_12198) );
AOI22_X2 inst_9188 ( .A1(net_9879), .B1(net_9780), .A2(net_8042), .B2(net_6140), .ZN(net_6126) );
INV_X4 inst_6625 ( .A(net_8966), .ZN(net_8965) );
CLKBUF_X2 inst_11240 ( .A(net_10855), .Z(net_11159) );
INV_X4 inst_6184 ( .ZN(net_1413), .A(net_194) );
XNOR2_X2 inst_201 ( .ZN(net_4957), .A(net_4407), .B(net_2652) );
CLKBUF_X2 inst_10958 ( .A(net_10584), .Z(net_10877) );
NAND2_X2 inst_3627 ( .ZN(net_7098), .A1(net_6873), .A2(net_6676) );
OAI22_X2 inst_1084 ( .A1(net_7157), .ZN(net_6574), .A2(net_5909), .B2(net_5907), .B1(net_371) );
XNOR2_X2 inst_304 ( .ZN(net_3271), .B(net_3270), .A(net_3023) );
CLKBUF_X2 inst_14388 ( .A(net_14306), .Z(net_14307) );
CLKBUF_X2 inst_14922 ( .A(net_14840), .Z(net_14841) );
AOI21_X2 inst_10106 ( .B1(net_9983), .ZN(net_4874), .A(net_4503), .B2(net_2541) );
NAND2_X2 inst_4157 ( .A2(net_2676), .ZN(net_2026), .A1(net_1629) );
OAI22_X2 inst_1027 ( .A2(net_8036), .B2(net_8018), .ZN(net_7985), .A1(net_3975), .B1(net_522) );
DFF_X1 inst_8432 ( .D(net_8639), .QN(net_278), .CK(net_14948) );
INV_X4 inst_5793 ( .ZN(net_2205), .A(net_1107) );
OAI22_X2 inst_1143 ( .A1(net_7226), .A2(net_5134), .B2(net_5133), .ZN(net_5130), .B1(net_476) );
CLKBUF_X2 inst_12823 ( .A(net_12741), .Z(net_12742) );
CLKBUF_X2 inst_11336 ( .A(net_11254), .Z(net_11255) );
CLKBUF_X2 inst_10670 ( .A(net_10587), .Z(net_10589) );
OAI222_X2 inst_1345 ( .A1(net_7665), .B2(net_7664), .C2(net_7663), .ZN(net_7555), .A2(net_7309), .B1(net_4602), .C1(net_1927) );
NOR2_X2 inst_2947 ( .A1(net_9243), .ZN(net_4464), .A2(net_543) );
CLKBUF_X2 inst_12024 ( .A(net_11942), .Z(net_11943) );
AND2_X4 inst_10457 ( .ZN(net_1658), .A2(net_1380), .A1(net_1364) );
INV_X4 inst_5122 ( .A(net_3397), .ZN(net_1607) );
CLKBUF_X2 inst_14225 ( .A(net_11211), .Z(net_14144) );
CLKBUF_X2 inst_12951 ( .A(net_11653), .Z(net_12870) );
CLKBUF_X2 inst_12679 ( .A(net_12597), .Z(net_12598) );
CLKBUF_X2 inst_11824 ( .A(net_11742), .Z(net_11743) );
INV_X4 inst_5638 ( .ZN(net_1265), .A(net_848) );
DFF_X1 inst_8503 ( .QN(net_9272), .D(net_7792), .CK(net_15405) );
NAND2_X2 inst_3608 ( .ZN(net_7258), .A2(net_6860), .A1(net_6597) );
CLKBUF_X2 inst_15235 ( .A(net_15153), .Z(net_15154) );
CLKBUF_X2 inst_10724 ( .A(net_10642), .Z(net_10643) );
INV_X2 inst_7306 ( .A(net_9076), .ZN(net_9075) );
OAI22_X2 inst_1016 ( .A2(net_8247), .B2(net_8246), .ZN(net_8201), .B1(net_8200), .A1(net_4291) );
NAND2_X2 inst_4147 ( .A2(net_2768), .A1(net_2415), .ZN(net_2075) );
OAI221_X2 inst_1538 ( .B2(net_7295), .C2(net_7293), .C1(net_7229), .ZN(net_7228), .A(net_6822), .B1(net_5467) );
CLKBUF_X2 inst_15273 ( .A(net_13101), .Z(net_15192) );
OR2_X2 inst_848 ( .A2(net_9580), .ZN(net_8705), .A1(net_1217) );
CLKBUF_X2 inst_13394 ( .A(net_11610), .Z(net_13313) );
AND4_X2 inst_10349 ( .ZN(net_1048), .A1(net_106), .A2(net_103), .A3(net_102), .A4(net_101) );
CLKBUF_X2 inst_12525 ( .A(net_12443), .Z(net_12444) );
NOR2_X4 inst_2479 ( .A2(net_10529), .ZN(net_3456), .A1(net_2842) );
CLKBUF_X2 inst_14333 ( .A(net_14251), .Z(net_14252) );
INV_X4 inst_6465 ( .A(net_10297), .ZN(net_371) );
INV_X4 inst_6312 ( .A(net_8833), .ZN(net_2707) );
OAI211_X2 inst_2179 ( .C1(net_7192), .C2(net_6548), .ZN(net_6530), .B(net_5658), .A(net_3679) );
NOR2_X2 inst_2578 ( .ZN(net_7087), .A1(net_6674), .A2(net_6249) );
DFF_X2 inst_7514 ( .QN(net_9238), .D(net_7897), .CK(net_11286) );
OAI21_X2 inst_1996 ( .ZN(net_3002), .B1(net_2491), .B2(net_1614), .A(net_1553) );
OAI221_X2 inst_1554 ( .C2(net_7295), .B2(net_7293), .ZN(net_7204), .B1(net_7203), .A(net_6827), .C1(net_1580) );
OAI221_X2 inst_1542 ( .B2(net_9047), .C2(net_7287), .ZN(net_7222), .C1(net_7221), .A(net_6797), .B1(net_5454) );
INV_X8 inst_4511 ( .ZN(net_4021), .A(net_3059) );
DFF_X1 inst_8849 ( .Q(net_10520), .D(net_92), .CK(net_10895) );
DFF_X2 inst_7830 ( .Q(net_10007), .D(net_6481), .CK(net_15426) );
CLKBUF_X2 inst_11580 ( .A(net_11498), .Z(net_11499) );
CLKBUF_X2 inst_12838 ( .A(net_12756), .Z(net_12757) );
NAND2_X4 inst_3340 ( .A2(net_8891), .A1(net_8890), .ZN(net_8526) );
SDFF_X2 inst_644 ( .Q(net_9461), .D(net_9461), .SE(net_3293), .CK(net_12439), .SI(x1865) );
INV_X4 inst_4683 ( .ZN(net_5263), .A(net_4998) );
INV_X4 inst_5015 ( .ZN(net_2810), .A(net_2116) );
OAI222_X2 inst_1380 ( .B2(net_7660), .A2(net_7659), .C2(net_7658), .ZN(net_6005), .B1(net_3952), .A1(net_2531), .C1(net_1903) );
NOR2_X2 inst_2806 ( .ZN(net_3168), .A2(net_2756), .A1(net_2279) );
NAND2_X2 inst_3891 ( .A1(net_4910), .ZN(net_3998), .A2(net_3981) );
CLKBUF_X2 inst_11298 ( .A(net_11015), .Z(net_11217) );
CLKBUF_X2 inst_12484 ( .A(net_12402), .Z(net_12403) );
INV_X2 inst_6736 ( .ZN(net_7415), .A(net_7332) );
NAND2_X2 inst_4008 ( .ZN(net_4697), .A1(net_3134), .A2(net_3133) );
DFF_X2 inst_8318 ( .Q(net_9619), .D(net_3970), .CK(net_14076) );
INV_X4 inst_6449 ( .A(net_10366), .ZN(net_753) );
CLKBUF_X2 inst_10652 ( .A(net_10570), .Z(net_10571) );
INV_X4 inst_4834 ( .ZN(net_3903), .A(net_3372) );
NAND2_X2 inst_3472 ( .A2(net_9441), .A1(net_8952), .ZN(net_8879) );
CLKBUF_X2 inst_12229 ( .A(net_12147), .Z(net_12148) );
INV_X4 inst_4896 ( .A(net_8856), .ZN(net_3133) );
DFF_X1 inst_8736 ( .Q(net_9135), .D(net_5726), .CK(net_10638) );
CLKBUF_X2 inst_14800 ( .A(net_14718), .Z(net_14719) );
AOI221_X2 inst_9933 ( .B2(net_5867), .A(net_5859), .ZN(net_5838), .C1(net_5837), .C2(net_4725), .B1(x5901) );
XNOR2_X2 inst_432 ( .B(net_9360), .ZN(net_1054), .A(net_195) );
XNOR2_X2 inst_282 ( .B(net_9225), .ZN(net_3663), .A(net_3480) );
CLKBUF_X2 inst_15829 ( .A(net_15747), .Z(net_15748) );
CLKBUF_X2 inst_11584 ( .A(net_10885), .Z(net_11503) );
DFF_X1 inst_8428 ( .Q(net_9583), .D(net_8710), .CK(net_11562) );
CLKBUF_X2 inst_12533 ( .A(net_12451), .Z(net_12452) );
AOI22_X2 inst_9605 ( .B1(net_9994), .A2(net_3500), .ZN(net_3462), .B2(net_2468), .A1(net_90) );
NOR4_X2 inst_2322 ( .ZN(net_6450), .A4(net_5444), .A3(net_4072), .A2(net_3927), .A1(net_3349) );
SDFF_X2 inst_513 ( .Q(net_9328), .D(net_9328), .SI(net_9153), .SE(net_7588), .CK(net_13095) );
NAND3_X2 inst_3266 ( .A1(net_6203), .ZN(net_4889), .A2(net_4233), .A3(net_4232) );
NAND3_X2 inst_3171 ( .A2(net_8961), .A1(net_8940), .ZN(net_8592), .A3(net_8591) );
CLKBUF_X2 inst_14340 ( .A(net_13354), .Z(net_14259) );
DFF_X1 inst_8725 ( .QN(net_10137), .D(net_6515), .CK(net_11228) );
DFF_X2 inst_7694 ( .Q(net_9206), .D(net_6653), .CK(net_11330) );
CLKBUF_X2 inst_14910 ( .A(net_14828), .Z(net_14829) );
CLKBUF_X2 inst_14060 ( .A(net_13978), .Z(net_13979) );
OAI221_X2 inst_1630 ( .B1(net_10308), .C1(net_7190), .B2(net_5591), .ZN(net_5577), .C2(net_4902), .A(net_3507) );
CLKBUF_X2 inst_12479 ( .A(net_12293), .Z(net_12398) );
OAI221_X2 inst_1586 ( .C1(net_10210), .C2(net_7295), .B2(net_7293), .B1(net_7127), .ZN(net_7117), .A(net_6925) );
AOI22_X2 inst_9318 ( .B1(net_9723), .A2(net_5755), .B2(net_5754), .ZN(net_5659), .A1(net_260) );
DFF_X2 inst_7887 ( .QN(net_10110), .D(net_6029), .CK(net_14907) );
AOI211_X2 inst_10296 ( .B(net_4009), .ZN(net_3745), .A(net_3744), .C1(net_3340), .C2(net_3323) );
OR2_X4 inst_774 ( .A2(net_7521), .A1(net_5949), .ZN(net_3093) );
OAI211_X2 inst_2292 ( .ZN(net_5072), .B(net_4478), .C2(net_4329), .A(net_4069), .C1(net_3511) );
CLKBUF_X2 inst_13954 ( .A(net_13781), .Z(net_13873) );
INV_X4 inst_6083 ( .A(net_10123), .ZN(net_501) );
NAND2_X2 inst_4256 ( .ZN(net_2919), .A1(net_932), .A2(net_171) );
CLKBUF_X2 inst_14826 ( .A(net_14744), .Z(net_14745) );
CLKBUF_X2 inst_10773 ( .A(net_10642), .Z(net_10692) );
INV_X4 inst_5300 ( .A(net_6828), .ZN(net_1300) );
CLKBUF_X2 inst_12340 ( .A(net_12258), .Z(net_12259) );
NOR2_X2 inst_2766 ( .A2(net_10540), .ZN(net_4324), .A1(net_3298) );
NAND2_X2 inst_4326 ( .A1(net_10439), .A2(net_1691), .ZN(net_1647) );
OAI221_X2 inst_1508 ( .C1(net_10421), .B2(net_9063), .C2(net_9056), .ZN(net_7353), .B1(net_7234), .A(net_7020) );
OAI22_X2 inst_1222 ( .A1(net_7108), .A2(net_5134), .B2(net_5133), .ZN(net_5025), .B1(net_2110) );
AOI22_X2 inst_9151 ( .A1(net_9748), .A2(net_6420), .ZN(net_6333), .B2(net_5263), .B1(net_3123) );
DFF_X2 inst_7938 ( .QN(net_10429), .D(net_5465), .CK(net_11470) );
CLKBUF_X2 inst_13985 ( .A(net_13903), .Z(net_13904) );
CLKBUF_X2 inst_11366 ( .A(net_11284), .Z(net_11285) );
NAND2_X2 inst_3407 ( .ZN(net_8537), .A2(net_8502), .A1(net_8150) );
OAI22_X2 inst_1073 ( .A2(net_6848), .B2(net_6846), .ZN(net_6845), .A1(net_5950), .B1(net_5786) );
NOR4_X2 inst_2323 ( .A1(net_9204), .ZN(net_6441), .A4(net_5695), .A3(net_1997), .A2(net_1815) );
NAND2_X2 inst_3741 ( .A2(net_9598), .ZN(net_8118), .A1(net_7846) );
CLKBUF_X2 inst_14643 ( .A(net_14561), .Z(net_14562) );
OAI221_X2 inst_1449 ( .B2(net_9629), .B1(net_8972), .ZN(net_8176), .A(net_7963), .C2(net_3526), .C1(net_999) );
XNOR2_X2 inst_127 ( .ZN(net_7484), .A(net_7100), .B(net_2270) );
CLKBUF_X2 inst_14754 ( .A(net_14672), .Z(net_14673) );
CLKBUF_X2 inst_11279 ( .A(net_11197), .Z(net_11198) );
CLKBUF_X2 inst_10657 ( .A(net_10561), .Z(net_10576) );
INV_X4 inst_5657 ( .A(net_843), .ZN(net_825) );
CLKBUF_X2 inst_11614 ( .A(net_11532), .Z(net_11533) );
DFF_X2 inst_7872 ( .QN(net_10144), .D(net_6015), .CK(net_13489) );
CLKBUF_X2 inst_14562 ( .A(net_14480), .Z(net_14481) );
XNOR2_X2 inst_187 ( .ZN(net_5208), .A(net_4437), .B(net_2372) );
XNOR2_X2 inst_206 ( .ZN(net_4946), .A(net_4680), .B(net_1742) );
CLKBUF_X2 inst_14270 ( .A(net_14188), .Z(net_14189) );
NAND2_X2 inst_3739 ( .ZN(net_6623), .A2(net_5393), .A1(net_588) );
NOR2_X1 inst_3029 ( .ZN(net_2973), .A1(net_2972), .A2(net_2971) );
OAI22_X2 inst_1268 ( .B1(net_7198), .A2(net_4842), .B2(net_4841), .ZN(net_4805), .A1(net_357) );
XNOR2_X2 inst_122 ( .ZN(net_7552), .A(net_7326), .B(net_7029) );
CLKBUF_X2 inst_15053 ( .A(net_14971), .Z(net_14972) );
XNOR2_X2 inst_405 ( .B(net_9842), .ZN(net_1693), .A(net_193) );
AOI222_X1 inst_9740 ( .B2(net_10192), .C2(net_10190), .A2(net_10189), .B1(net_10179), .C1(net_10177), .A1(net_10176), .ZN(net_1125) );
INV_X4 inst_6436 ( .ZN(net_7249), .A(x5601) );
INV_X4 inst_4788 ( .ZN(net_4182), .A(net_4028) );
AND2_X2 inst_10505 ( .A2(net_10168), .ZN(net_5971), .A1(net_1168) );
INV_X4 inst_6166 ( .A(net_10255), .ZN(net_1115) );
INV_X4 inst_6281 ( .A(net_9980), .ZN(net_439) );
DFF_X2 inst_7540 ( .QN(net_8825), .D(net_7738), .CK(net_13047) );
AOI21_X2 inst_10077 ( .B2(net_10343), .A(net_10342), .ZN(net_5943), .B1(net_1599) );
NAND2_X2 inst_3912 ( .ZN(net_4011), .A1(net_3920), .A2(net_3890) );
CLKBUF_X2 inst_12833 ( .A(net_11349), .Z(net_12752) );
DFF_X1 inst_8499 ( .QN(net_10256), .D(net_7788), .CK(net_11717) );
NOR4_X2 inst_2306 ( .ZN(net_7769), .A4(net_7617), .A1(net_3362), .A2(net_1996), .A3(net_1416) );
INV_X2 inst_6776 ( .ZN(net_6022), .A(net_5838) );
CLKBUF_X2 inst_13087 ( .A(net_13005), .Z(net_13006) );
AOI22_X2 inst_9191 ( .A1(net_9881), .B1(net_9782), .A2(net_8042), .B2(net_6129), .ZN(net_6123) );
INV_X4 inst_5645 ( .A(net_5786), .ZN(net_1114) );
CLKBUF_X2 inst_13046 ( .A(net_12964), .Z(net_12965) );
CLKBUF_X2 inst_14468 ( .A(net_13928), .Z(net_14387) );
CLKBUF_X2 inst_14008 ( .A(net_13926), .Z(net_13927) );
OAI221_X2 inst_1646 ( .B1(net_10441), .C1(net_7237), .A(net_5575), .ZN(net_5542), .B2(net_4477), .C2(net_4455) );
CLKBUF_X2 inst_15361 ( .A(net_15279), .Z(net_15280) );
OAI211_X2 inst_2176 ( .C1(net_7198), .C2(net_6548), .ZN(net_6533), .B(net_5661), .A(net_3527) );
INV_X2 inst_6748 ( .A(net_7281), .ZN(net_6622) );
INV_X4 inst_5773 ( .ZN(net_1332), .A(net_715) );
NOR2_X2 inst_2892 ( .ZN(net_3145), .A1(net_2074), .A2(net_1688) );
DFF_X2 inst_7547 ( .QN(net_9249), .D(net_7706), .CK(net_11273) );
CLKBUF_X2 inst_13664 ( .A(net_13582), .Z(net_13583) );
INV_X2 inst_6741 ( .ZN(net_7162), .A(net_7028) );
INV_X4 inst_6294 ( .A(net_10107), .ZN(net_5858) );
INV_X4 inst_6339 ( .A(net_9736), .ZN(net_1031) );
INV_X4 inst_5550 ( .A(net_10245), .ZN(net_1272) );
OAI22_X2 inst_1102 ( .B2(net_10133), .A1(net_10132), .ZN(net_6210), .A2(net_5960), .B1(net_2096) );
CLKBUF_X2 inst_13024 ( .A(net_11154), .Z(net_12943) );
INV_X4 inst_6368 ( .A(net_9937), .ZN(net_401) );
CLKBUF_X2 inst_14929 ( .A(net_12639), .Z(net_14848) );
CLKBUF_X2 inst_15082 ( .A(net_12846), .Z(net_15001) );
CLKBUF_X2 inst_11663 ( .A(net_11548), .Z(net_11582) );
DFF_X2 inst_7804 ( .Q(net_9921), .D(net_6458), .CK(net_11967) );
CLKBUF_X2 inst_14968 ( .A(net_10871), .Z(net_14887) );
CLKBUF_X2 inst_13329 ( .A(net_10652), .Z(net_13248) );
AOI221_X2 inst_9795 ( .B1(net_9975), .A(net_7090), .B2(net_7089), .C2(net_7088), .ZN(net_7009), .C1(net_247) );
INV_X4 inst_5365 ( .ZN(net_1975), .A(net_1217) );
OR3_X4 inst_702 ( .A3(net_10304), .ZN(net_7665), .A1(net_4169), .A2(net_4160) );
NOR2_X2 inst_2482 ( .ZN(net_8809), .A2(net_8808), .A1(net_8801) );
INV_X4 inst_5860 ( .ZN(net_2565), .A(net_928) );
NOR2_X2 inst_2957 ( .A1(net_10264), .ZN(net_2231), .A2(net_1208) );
CLKBUF_X2 inst_15606 ( .A(net_15524), .Z(net_15525) );
CLKBUF_X2 inst_12448 ( .A(net_12366), .Z(net_12367) );
CLKBUF_X2 inst_15192 ( .A(net_14981), .Z(net_15111) );
CLKBUF_X2 inst_10880 ( .A(net_10798), .Z(net_10799) );
AOI22_X2 inst_9297 ( .B1(net_10000), .A1(net_5743), .B2(net_5742), .ZN(net_5691), .A2(net_240) );
CLKBUF_X2 inst_15551 ( .A(net_12985), .Z(net_15470) );
NOR2_X2 inst_2711 ( .ZN(net_4174), .A2(net_3715), .A1(net_3140) );
CLKBUF_X2 inst_12808 ( .A(net_12726), .Z(net_12727) );
AOI221_X2 inst_9980 ( .C1(net_10184), .B2(net_6442), .ZN(net_4218), .C2(net_4217), .A(net_3587), .B1(net_2000) );
NAND2_X2 inst_3531 ( .A2(net_9625), .A1(net_8975), .ZN(net_8055) );
NOR2_X2 inst_2753 ( .ZN(net_4098), .A2(net_3640), .A1(net_3181) );
NAND2_X2 inst_3672 ( .A1(net_7846), .ZN(net_6904), .A2(net_6238) );
CLKBUF_X2 inst_14329 ( .A(net_11777), .Z(net_14248) );
XNOR2_X2 inst_132 ( .ZN(net_7418), .A(net_7321), .B(net_1861) );
CLKBUF_X2 inst_15484 ( .A(net_15402), .Z(net_15403) );
AND3_X4 inst_10353 ( .ZN(net_8002), .A3(net_7110), .A2(net_7095), .A1(net_6916) );
CLKBUF_X2 inst_13900 ( .A(net_13818), .Z(net_13819) );
CLKBUF_X2 inst_11502 ( .A(net_10888), .Z(net_11421) );
CLKBUF_X2 inst_12233 ( .A(net_12151), .Z(net_12152) );
CLKBUF_X2 inst_12619 ( .A(net_12537), .Z(net_12538) );
CLKBUF_X2 inst_13912 ( .A(net_13830), .Z(net_13831) );
AOI22_X2 inst_9049 ( .B1(net_9672), .A1(net_6684), .B2(net_6683), .ZN(net_6675), .A2(net_241) );
AND3_X2 inst_10369 ( .ZN(net_4967), .A2(net_4966), .A3(net_4698), .A1(net_4697) );
DFF_X2 inst_7935 ( .QN(net_10219), .D(net_5472), .CK(net_14476) );
INV_X4 inst_6149 ( .ZN(net_5964), .A(net_181) );
NAND2_X2 inst_3545 ( .A1(net_8511), .ZN(net_7927), .A2(net_7926) );
CLKBUF_X2 inst_12365 ( .A(net_12283), .Z(net_12284) );
CLKBUF_X2 inst_15681 ( .A(net_15599), .Z(net_15600) );
CLKBUF_X2 inst_13335 ( .A(net_11839), .Z(net_13254) );
NAND2_X2 inst_3611 ( .ZN(net_7255), .A2(net_6875), .A1(net_6591) );
NOR2_X2 inst_2928 ( .A1(net_10368), .ZN(net_2755), .A2(net_1361) );
NAND2_X2 inst_3813 ( .A1(net_10082), .A2(net_4534), .ZN(net_4525) );
XNOR2_X2 inst_400 ( .A(net_3933), .ZN(net_1753), .B(net_1462) );
NOR2_X2 inst_2991 ( .ZN(net_1863), .A2(net_911), .A1(net_728) );
CLKBUF_X2 inst_12612 ( .A(net_12530), .Z(net_12531) );
INV_X4 inst_6309 ( .A(net_10038), .ZN(net_5092) );
NAND2_X2 inst_3513 ( .ZN(net_8249), .A1(net_8141), .A2(net_8140) );
XNOR2_X2 inst_261 ( .B(net_4927), .ZN(net_3993), .A(net_3483) );
CLKBUF_X2 inst_12418 ( .A(net_12336), .Z(net_12337) );
XNOR2_X2 inst_268 ( .ZN(net_3962), .A(net_3647), .B(net_2042) );
OAI221_X2 inst_1518 ( .C1(net_10422), .B2(net_9063), .C2(net_9056), .ZN(net_7314), .B1(net_7139), .A(net_7062) );
CLKBUF_X2 inst_10985 ( .A(net_10903), .Z(net_10904) );
DFF_X2 inst_8198 ( .Q(net_10034), .D(net_5104), .CK(net_14275) );
DFF_X1 inst_8586 ( .Q(net_9867), .D(net_7126), .CK(net_13372) );
CLKBUF_X2 inst_15083 ( .A(net_15001), .Z(net_15002) );
NAND2_X2 inst_3975 ( .A2(net_4723), .A1(net_3591), .ZN(net_3292) );
CLKBUF_X2 inst_11025 ( .A(net_10943), .Z(net_10944) );
CLKBUF_X2 inst_10976 ( .A(net_10784), .Z(net_10895) );
XNOR2_X2 inst_327 ( .ZN(net_3007), .A(net_2803), .B(net_1799) );
AOI22_X2 inst_9199 ( .A1(net_9889), .B1(net_9790), .B2(net_6140), .ZN(net_6114), .A2(net_6111) );
CLKBUF_X2 inst_12264 ( .A(net_11885), .Z(net_12183) );
DFF_X1 inst_8874 ( .Q(net_9505), .D(net_9281), .CK(net_14370) );
DFF_X2 inst_7801 ( .Q(net_9917), .D(net_6490), .CK(net_12791) );
INV_X2 inst_7245 ( .A(net_9417), .ZN(net_8197) );
CLKBUF_X2 inst_14118 ( .A(net_14036), .Z(net_14037) );
NAND2_X2 inst_3509 ( .A1(net_9545), .ZN(net_8371), .A2(net_8113) );
CLKBUF_X2 inst_13936 ( .A(net_13854), .Z(net_13855) );
AOI22_X2 inst_9431 ( .ZN(net_4591), .A1(net_4423), .A2(net_4280), .B2(net_3395), .B1(net_3174) );
CLKBUF_X2 inst_10746 ( .A(net_10664), .Z(net_10665) );
DFF_X2 inst_7971 ( .QN(net_10323), .D(net_5581), .CK(net_14599) );
NAND2_X2 inst_3853 ( .ZN(net_8897), .A1(net_4190), .A2(net_4187) );
DFF_X2 inst_8044 ( .QN(net_9554), .D(net_9260), .CK(net_13759) );
CLKBUF_X2 inst_15132 ( .A(net_15050), .Z(net_15051) );
INV_X2 inst_6702 ( .ZN(net_8266), .A(net_8152) );
CLKBUF_X2 inst_11511 ( .A(net_10664), .Z(net_11430) );
CLKBUF_X2 inst_14304 ( .A(net_14222), .Z(net_14223) );
CLKBUF_X2 inst_12421 ( .A(net_12339), .Z(net_12340) );
DFF_X2 inst_7905 ( .QN(net_10264), .D(net_6001), .CK(net_11664) );
INV_X4 inst_6348 ( .ZN(net_408), .A(x682) );
AOI22_X2 inst_9229 ( .A1(net_9923), .B1(net_9824), .A2(net_8042), .B2(net_6140), .ZN(net_6082) );
DFF_X2 inst_8357 ( .QN(net_9164), .D(net_9163), .CK(net_12997) );
NAND4_X2 inst_3097 ( .ZN(net_4346), .A2(net_3862), .A1(net_3861), .A3(net_3756), .A4(net_3498) );
CLKBUF_X2 inst_10739 ( .A(net_10555), .Z(net_10658) );
AOI22_X2 inst_9625 ( .A1(net_10077), .B1(net_9964), .A2(net_5319), .ZN(net_3422), .B2(net_2541) );
NAND2_X2 inst_3661 ( .ZN(net_8325), .A2(net_7038), .A1(net_3527) );
CLKBUF_X2 inst_13678 ( .A(net_11733), .Z(net_13597) );
SDFF_X2 inst_502 ( .SE(net_9540), .SI(net_8199), .Q(net_287), .D(net_287), .CK(net_12693) );
CLKBUF_X2 inst_14244 ( .A(net_11061), .Z(net_14163) );
CLKBUF_X2 inst_13976 ( .A(net_13894), .Z(net_13895) );
AOI22_X2 inst_9001 ( .A1(net_8961), .ZN(net_8407), .A2(net_8368), .B2(net_8252), .B1(net_8128) );
CLKBUF_X2 inst_11836 ( .A(net_11376), .Z(net_11755) );
DFF_X1 inst_8745 ( .Q(net_9130), .D(net_5690), .CK(net_10580) );
NAND3_X2 inst_3221 ( .A2(net_7420), .ZN(net_5354), .A1(net_5353), .A3(net_5351) );
CLKBUF_X2 inst_14585 ( .A(net_14503), .Z(net_14504) );
CLKBUF_X2 inst_14771 ( .A(net_14689), .Z(net_14690) );
NAND2_X2 inst_3645 ( .A2(net_7278), .ZN(net_6893), .A1(net_6229) );
CLKBUF_X2 inst_15724 ( .A(net_15642), .Z(net_15643) );
OAI221_X2 inst_1598 ( .B1(net_10213), .C1(net_7211), .B2(net_5642), .ZN(net_5639), .C2(net_4905), .A(net_3507) );
CLKBUF_X2 inst_12335 ( .A(net_12253), .Z(net_12254) );
XNOR2_X2 inst_357 ( .ZN(net_2775), .B(net_2631), .A(net_1803) );
CLKBUF_X2 inst_11083 ( .A(net_11001), .Z(net_11002) );
INV_X2 inst_6969 ( .A(net_4675), .ZN(net_1806) );
AOI21_X2 inst_10028 ( .B1(net_9368), .A(net_7916), .B2(net_7915), .ZN(net_7851) );
CLKBUF_X2 inst_15670 ( .A(net_15588), .Z(net_15589) );
AOI21_X2 inst_10167 ( .B2(net_10407), .ZN(net_8447), .A(net_4371), .B1(net_3672) );
INV_X4 inst_6173 ( .ZN(net_6381), .A(net_128) );
NAND2_X2 inst_4092 ( .A1(net_10366), .ZN(net_3101), .A2(net_2528) );
CLKBUF_X2 inst_13865 ( .A(net_10741), .Z(net_13784) );
AOI21_X2 inst_10098 ( .ZN(net_5102), .A(net_5101), .B1(net_5100), .B2(net_3017) );
DFF_X2 inst_7880 ( .Q(net_9748), .D(net_6152), .CK(net_15229) );
NAND2_X2 inst_3980 ( .A2(net_9958), .A1(net_9957), .ZN(net_3258) );
CLKBUF_X2 inst_15073 ( .A(net_14991), .Z(net_14992) );
NAND4_X2 inst_3152 ( .A3(net_9184), .A4(net_4125), .ZN(net_2092), .A1(net_2091), .A2(net_2090) );
CLKBUF_X2 inst_11438 ( .A(net_11356), .Z(net_11357) );
NAND2_X2 inst_4161 ( .A1(net_9513), .ZN(net_6967), .A2(net_797) );
NAND2_X2 inst_3758 ( .A1(net_5388), .ZN(net_5231), .A2(net_4940) );
OR2_X2 inst_912 ( .ZN(net_3887), .A2(net_3612), .A1(net_752) );
CLKBUF_X2 inst_15653 ( .A(net_15571), .Z(net_15572) );
AOI21_X2 inst_10065 ( .ZN(net_6969), .A(net_6968), .B2(net_6967), .B1(net_1894) );
CLKBUF_X2 inst_11678 ( .A(net_11336), .Z(net_11597) );
AOI21_X2 inst_10117 ( .A(net_8859), .ZN(net_4548), .B2(net_4398), .B1(net_4266) );
INV_X4 inst_5869 ( .A(net_3365), .ZN(net_638) );
NAND3_X2 inst_3196 ( .ZN(net_7477), .A3(net_7476), .A2(net_6630), .A1(net_5984) );
CLKBUF_X2 inst_14603 ( .A(net_12170), .Z(net_14522) );
CLKBUF_X2 inst_12724 ( .A(net_12642), .Z(net_12643) );
INV_X4 inst_5872 ( .A(net_637), .ZN(net_636) );
CLKBUF_X2 inst_15452 ( .A(net_15370), .Z(net_15371) );
INV_X4 inst_6525 ( .A(net_10333), .ZN(net_1344) );
NAND2_X2 inst_4025 ( .ZN(net_3357), .A1(net_3067), .A2(net_2225) );
XNOR2_X2 inst_322 ( .ZN(net_3031), .A(net_2832), .B(net_2497) );
AOI21_X2 inst_10070 ( .B1(net_10385), .ZN(net_6970), .A(net_6677), .B2(net_264) );
NAND2_X2 inst_3516 ( .A2(net_9589), .A1(net_9096), .ZN(net_8153) );
INV_X2 inst_6988 ( .A(net_2074), .ZN(net_1651) );
NAND2_X2 inst_4200 ( .A1(net_1796), .ZN(net_1794), .A2(net_1793) );
NAND2_X2 inst_4188 ( .ZN(net_2905), .A2(net_1971), .A1(net_1856) );
CLKBUF_X2 inst_14888 ( .A(net_14806), .Z(net_14807) );
CLKBUF_X2 inst_14405 ( .A(net_13576), .Z(net_14324) );
NAND2_X2 inst_4169 ( .ZN(net_2661), .A2(net_1378), .A1(net_1073) );
NAND2_X2 inst_3902 ( .ZN(net_3904), .A2(net_3903), .A1(net_100) );
CLKBUF_X2 inst_10858 ( .A(net_10572), .Z(net_10777) );
AOI221_X2 inst_9894 ( .B1(net_9861), .B2(net_9101), .A(net_6945), .C2(net_6944), .C1(net_6828), .ZN(net_6800) );
INV_X4 inst_6191 ( .A(net_10365), .ZN(net_773) );
INV_X2 inst_6863 ( .A(net_3425), .ZN(net_3279) );
CLKBUF_X2 inst_10647 ( .A(net_10565), .Z(net_10566) );
INV_X4 inst_6243 ( .A(net_10249), .ZN(net_759) );
DFF_X2 inst_8302 ( .QN(net_10139), .D(net_4438), .CK(net_10856) );
INV_X2 inst_6908 ( .A(net_5331), .ZN(net_2808) );
INV_X4 inst_5346 ( .A(net_8803), .ZN(net_8801) );
INV_X4 inst_6289 ( .A(net_9731), .ZN(net_724) );
NAND2_X2 inst_4181 ( .ZN(net_2548), .A2(net_1521), .A1(net_1252) );
CLKBUF_X2 inst_12662 ( .A(net_11238), .Z(net_12581) );
NOR4_X2 inst_2315 ( .A3(net_10409), .A1(net_10408), .ZN(net_7412), .A4(net_7064), .A2(net_355) );
OAI33_X1 inst_962 ( .ZN(net_4072), .A2(net_4071), .A3(net_4070), .B1(net_3914), .A1(net_3091), .B2(net_1959), .B3(net_648) );
CLKBUF_X2 inst_10865 ( .A(net_10783), .Z(net_10784) );
INV_X4 inst_6350 ( .A(net_9373), .ZN(net_7634) );
OAI21_X2 inst_2008 ( .ZN(net_2314), .B2(net_2302), .A(net_1675), .B1(net_1094) );
SDFF_X2 inst_641 ( .Q(net_9463), .D(net_9463), .SE(net_3293), .CK(net_11888), .SI(x1743) );
SDFF_X2 inst_498 ( .SE(net_9540), .SI(net_8211), .Q(net_284), .D(net_284), .CK(net_12697) );
OAI21_X2 inst_1988 ( .ZN(net_2898), .B2(net_2685), .B1(net_2202), .A(net_2035) );
CLKBUF_X2 inst_11489 ( .A(net_11407), .Z(net_11408) );
AOI222_X2 inst_9673 ( .ZN(net_3119), .A1(net_3118), .C2(net_3117), .B2(net_3117), .A2(net_2261), .C1(net_1756), .B1(net_1151) );
DFF_X2 inst_8374 ( .QN(net_8831), .D(net_1499), .CK(net_12467) );
CLKBUF_X2 inst_12346 ( .A(net_12264), .Z(net_12265) );
DFF_X2 inst_8287 ( .Q(net_10088), .D(net_4847), .CK(net_10717) );
CLKBUF_X2 inst_11971 ( .A(net_11889), .Z(net_11890) );
DFF_X2 inst_7955 ( .QN(net_10216), .D(net_5635), .CK(net_13258) );
INV_X4 inst_5517 ( .ZN(net_4918), .A(net_971) );
OAI21_X2 inst_1912 ( .ZN(net_4633), .B1(net_4378), .B2(net_4210), .A(net_3086) );
CLKBUF_X2 inst_14478 ( .A(net_14396), .Z(net_14397) );
CLKBUF_X2 inst_14044 ( .A(net_13962), .Z(net_13963) );
OAI21_X2 inst_1831 ( .B1(net_7157), .ZN(net_6451), .A(net_5696), .B2(net_5410) );
CLKBUF_X2 inst_13438 ( .A(net_13356), .Z(net_13357) );
AOI22_X2 inst_9308 ( .B1(net_9695), .A1(net_6828), .A2(net_5755), .B2(net_5754), .ZN(net_5670) );
INV_X2 inst_6714 ( .ZN(net_7942), .A(net_7918) );
INV_X2 inst_6683 ( .ZN(net_8345), .A(net_8279) );
CLKBUF_X2 inst_14339 ( .A(net_10974), .Z(net_14258) );
CLKBUF_X2 inst_13671 ( .A(net_13589), .Z(net_13590) );
NAND2_X2 inst_3468 ( .ZN(net_8546), .A2(net_8454), .A1(net_8124) );
CLKBUF_X2 inst_11876 ( .A(net_11794), .Z(net_11795) );
XNOR2_X2 inst_350 ( .B(net_2876), .ZN(net_2816), .A(net_2510) );
CLKBUF_X2 inst_11322 ( .A(net_11240), .Z(net_11241) );
NOR3_X2 inst_2395 ( .ZN(net_7792), .A1(net_7695), .A3(net_7694), .A2(net_5284) );
XNOR2_X2 inst_231 ( .ZN(net_4387), .A(net_3939), .B(net_2020) );
AOI22_X2 inst_9024 ( .B1(net_9524), .A1(net_8002), .B2(net_8001), .ZN(net_7995), .A2(net_7950) );
AND2_X4 inst_10403 ( .ZN(net_5445), .A2(net_4998), .A1(net_4197) );
NAND3_X2 inst_3309 ( .ZN(net_2791), .A1(net_2169), .A2(net_1728), .A3(net_1719) );
CLKBUF_X2 inst_14437 ( .A(net_14355), .Z(net_14356) );
INV_X4 inst_5104 ( .ZN(net_2321), .A(net_1687) );
AOI221_X2 inst_9952 ( .B2(net_7770), .C1(net_7697), .ZN(net_5005), .B1(net_5004), .A(net_4463), .C2(net_2526) );
INV_X4 inst_5676 ( .A(net_10230), .ZN(net_1282) );
CLKBUF_X2 inst_15459 ( .A(net_15377), .Z(net_15378) );
CLKBUF_X2 inst_12851 ( .A(net_12769), .Z(net_12770) );
NOR4_X2 inst_2317 ( .ZN(net_7174), .A1(net_6613), .A3(net_6381), .A4(net_6379), .A2(net_3614) );
CLKBUF_X2 inst_11901 ( .A(net_11330), .Z(net_11820) );
CLKBUF_X2 inst_11365 ( .A(net_11283), .Z(net_11284) );
DFF_X1 inst_8518 ( .Q(net_8822), .D(net_7473), .CK(net_14495) );
CLKBUF_X2 inst_15816 ( .A(net_15193), .Z(net_15735) );
DFF_X2 inst_7506 ( .QN(net_9591), .D(net_7970), .CK(net_11490) );
OAI221_X2 inst_1452 ( .ZN(net_8060), .C2(net_7880), .A(net_7877), .B2(net_7833), .B1(net_7793), .C1(net_6836) );
CLKBUF_X2 inst_13740 ( .A(net_12829), .Z(net_13659) );
CLKBUF_X2 inst_11867 ( .A(net_11482), .Z(net_11786) );
INV_X2 inst_6756 ( .A(net_9561), .ZN(net_9011) );
INV_X4 inst_6549 ( .A(net_8824), .ZN(net_7640) );
CLKBUF_X2 inst_15208 ( .A(net_15126), .Z(net_15127) );
INV_X4 inst_5000 ( .ZN(net_4713), .A(net_2605) );
CLKBUF_X2 inst_12967 ( .A(net_12885), .Z(net_12886) );
NAND2_X2 inst_4077 ( .A1(net_9535), .ZN(net_7341), .A2(net_2200) );
NAND4_X2 inst_3139 ( .ZN(net_3129), .A3(net_2716), .A1(net_2705), .A4(net_2704), .A2(net_1621) );
CLKBUF_X2 inst_12801 ( .A(net_12719), .Z(net_12720) );
NOR2_X2 inst_2558 ( .ZN(net_7767), .A2(net_7766), .A1(net_7274) );
OAI222_X2 inst_1396 ( .A2(net_7732), .C2(net_7731), .B2(net_7730), .ZN(net_5702), .A1(net_2884), .B1(net_1801), .C1(net_1488) );
XNOR2_X2 inst_352 ( .ZN(net_2813), .B(net_2296), .A(net_1853) );
XNOR2_X2 inst_286 ( .ZN(net_8766), .A(net_2996), .B(net_2447) );
CLKBUF_X2 inst_13354 ( .A(net_13272), .Z(net_13273) );
AOI21_X2 inst_10112 ( .A(net_8861), .ZN(net_4579), .B2(net_4400), .B1(net_4267) );
INV_X2 inst_6880 ( .A(net_3917), .ZN(net_2848) );
CLKBUF_X2 inst_15328 ( .A(net_11626), .Z(net_15247) );
CLKBUF_X2 inst_15768 ( .A(net_15216), .Z(net_15687) );
CLKBUF_X2 inst_15663 ( .A(net_13125), .Z(net_15582) );
AND2_X4 inst_10447 ( .ZN(net_1679), .A2(net_1385), .A1(net_1381) );
CLKBUF_X2 inst_14959 ( .A(net_14877), .Z(net_14878) );
CLKBUF_X2 inst_12984 ( .A(net_12533), .Z(net_12903) );
CLKBUF_X2 inst_15524 ( .A(net_14972), .Z(net_15443) );
CLKBUF_X2 inst_13006 ( .A(net_12924), .Z(net_12925) );
DFF_X2 inst_7961 ( .QN(net_10205), .D(net_5627), .CK(net_14217) );
CLKBUF_X2 inst_15311 ( .A(net_12182), .Z(net_15230) );
NOR2_X2 inst_3003 ( .ZN(net_2434), .A2(net_1118), .A1(net_513) );
INV_X2 inst_6792 ( .A(net_8118), .ZN(net_6160) );
CLKBUF_X2 inst_15058 ( .A(net_14466), .Z(net_14977) );
CLKBUF_X2 inst_12169 ( .A(net_12087), .Z(net_12088) );
INV_X4 inst_5579 ( .ZN(net_1448), .A(net_891) );
NAND2_X2 inst_3841 ( .ZN(net_4439), .A2(net_4296), .A1(net_2600) );
CLKBUF_X2 inst_13134 ( .A(net_13052), .Z(net_13053) );
AOI22_X2 inst_9555 ( .A1(net_10395), .B1(net_9879), .A2(net_4062), .ZN(net_3765), .B2(net_2973) );
AOI22_X2 inst_9165 ( .A2(net_6382), .ZN(net_6307), .B2(net_5263), .A1(net_4037), .B1(net_3000) );
DFF_X1 inst_8550 ( .Q(net_9986), .D(net_7355), .CK(net_14775) );
OAI211_X2 inst_2185 ( .C1(net_7186), .C2(net_6542), .ZN(net_6524), .B(net_5619), .A(net_3679) );
NAND2_X2 inst_4050 ( .ZN(net_3013), .A2(net_2810), .A1(net_1576) );
DFF_X2 inst_7737 ( .Q(net_9897), .D(net_6194), .CK(net_11977) );
INV_X2 inst_6972 ( .ZN(net_2442), .A(net_1714) );
CLKBUF_X2 inst_12203 ( .A(net_12121), .Z(net_12122) );
AOI22_X2 inst_9427 ( .A1(net_9753), .B1(net_6813), .ZN(net_4620), .A2(net_4618), .B2(net_4617) );
NOR3_X2 inst_2370 ( .A3(net_8190), .ZN(net_8161), .A2(net_7694), .A1(net_3867) );
CLKBUF_X2 inst_14069 ( .A(net_13987), .Z(net_13988) );
INV_X4 inst_5887 ( .ZN(net_860), .A(net_615) );
NAND2_X2 inst_3882 ( .ZN(net_4023), .A1(net_4022), .A2(net_4021) );
CLKBUF_X2 inst_11598 ( .A(net_10967), .Z(net_11517) );
CLKBUF_X2 inst_13452 ( .A(net_11624), .Z(net_13371) );
NOR2_X2 inst_2811 ( .ZN(net_2650), .A1(net_2649), .A2(net_2648) );
CLKBUF_X2 inst_12001 ( .A(net_11919), .Z(net_11920) );
INV_X4 inst_6120 ( .A(net_10008), .ZN(net_488) );
INV_X4 inst_4615 ( .ZN(net_7337), .A(net_7152) );
XNOR2_X2 inst_137 ( .ZN(net_7399), .A(net_6913), .B(net_1835) );
INV_X2 inst_6889 ( .ZN(net_2695), .A(net_2414) );
XNOR2_X2 inst_425 ( .B(net_9844), .A(net_1417), .ZN(net_1355) );
NOR2_X2 inst_2567 ( .ZN(net_7517), .A2(net_7352), .A1(net_7044) );
CLKBUF_X2 inst_11384 ( .A(net_11302), .Z(net_11303) );
NAND3_X2 inst_3206 ( .ZN(net_6911), .A3(net_5968), .A1(net_3819), .A2(net_3818) );
CLKBUF_X2 inst_11742 ( .A(net_11660), .Z(net_11661) );
DFF_X1 inst_8416 ( .QN(net_9362), .D(net_8788), .CK(net_11930) );
DFF_X1 inst_8591 ( .Q(net_9669), .D(net_7112), .CK(net_11622) );
CLKBUF_X2 inst_15298 ( .A(net_15216), .Z(net_15217) );
NOR2_X2 inst_2572 ( .ZN(net_7431), .A2(net_7318), .A1(net_7046) );
CLKBUF_X2 inst_13764 ( .A(net_13682), .Z(net_13683) );
AOI22_X2 inst_9380 ( .B1(net_10021), .A1(net_6811), .A2(net_5743), .B2(net_5742), .ZN(net_5525) );
INV_X2 inst_6755 ( .A(net_9545), .ZN(net_6247) );
CLKBUF_X2 inst_13111 ( .A(net_12101), .Z(net_13030) );
AOI21_X2 inst_10245 ( .ZN(net_8865), .B1(net_4553), .B2(net_2396), .A(net_2395) );
NAND2_X2 inst_4046 ( .A2(net_8831), .ZN(net_2825), .A1(net_2824) );
NAND2_X4 inst_3365 ( .A2(net_8898), .A1(net_8897), .ZN(net_7277) );
INV_X2 inst_7179 ( .A(net_9402), .ZN(net_8230) );
NAND3_X2 inst_3254 ( .A3(net_8847), .ZN(net_4507), .A1(net_4506), .A2(net_872) );
CLKBUF_X2 inst_11752 ( .A(net_10868), .Z(net_11671) );
OAI22_X2 inst_983 ( .A2(net_8962), .B2(net_8659), .ZN(net_8657), .A1(net_6220), .B1(net_5803) );
INV_X4 inst_4980 ( .A(net_2601), .ZN(net_2587) );
DFF_X2 inst_8026 ( .QN(net_10431), .D(net_5463), .CK(net_11463) );
DFF_X2 inst_8112 ( .Q(net_9749), .D(net_5141), .CK(net_14743) );
DFF_X1 inst_8511 ( .QN(net_10478), .D(net_7581), .CK(net_11418) );
OAI21_X2 inst_1897 ( .B1(net_7249), .B2(net_4862), .ZN(net_4855), .A(net_4527) );
AND2_X2 inst_10615 ( .ZN(net_2510), .A2(net_1741), .A1(net_878) );
DFF_X2 inst_7773 ( .Q(net_9724), .D(net_6529), .CK(net_12053) );
CLKBUF_X2 inst_11810 ( .A(net_11728), .Z(net_11729) );
NAND4_X2 inst_3159 ( .ZN(net_1736), .A2(net_880), .A3(net_144), .A4(net_143), .A1(net_142) );
CLKBUF_X2 inst_15587 ( .A(net_15505), .Z(net_15506) );
CLKBUF_X2 inst_15786 ( .A(net_15704), .Z(net_15705) );
CLKBUF_X2 inst_11291 ( .A(net_10767), .Z(net_11210) );
CLKBUF_X2 inst_11196 ( .A(net_11114), .Z(net_11115) );
INV_X4 inst_4776 ( .ZN(net_4311), .A(net_4182) );
INV_X2 inst_7130 ( .A(net_1096), .ZN(net_869) );
INV_X4 inst_6237 ( .ZN(net_3733), .A(net_266) );
OAI221_X2 inst_1569 ( .C1(net_10321), .C2(net_9047), .B2(net_7287), .B1(net_7186), .ZN(net_7181), .A(net_6804) );
CLKBUF_X2 inst_11722 ( .A(net_11557), .Z(net_11641) );
CLKBUF_X2 inst_12990 ( .A(net_12908), .Z(net_12909) );
NOR2_X2 inst_2633 ( .A2(net_5927), .ZN(net_5922), .A1(net_961) );
CLKBUF_X2 inst_13565 ( .A(net_12604), .Z(net_13484) );
INV_X2 inst_7314 ( .A(net_9095), .ZN(net_9094) );
INV_X2 inst_7080 ( .ZN(net_1182), .A(net_1181) );
OAI21_X2 inst_1772 ( .ZN(net_8007), .A(net_7871), .B2(net_7864), .B1(net_3984) );
INV_X2 inst_6947 ( .ZN(net_1901), .A(net_1900) );
INV_X4 inst_6274 ( .A(net_10007), .ZN(net_444) );
CLKBUF_X2 inst_13725 ( .A(net_13564), .Z(net_13644) );
CLKBUF_X2 inst_14738 ( .A(net_14656), .Z(net_14657) );
OAI211_X2 inst_2143 ( .C2(net_6778), .ZN(net_6705), .A(net_6332), .B(net_6068), .C1(net_5084) );
CLKBUF_X2 inst_14233 ( .A(net_14151), .Z(net_14152) );
OAI22_X2 inst_1291 ( .ZN(net_4261), .B2(net_3238), .A1(net_2987), .A2(net_2986), .B1(net_2783) );
DFF_X2 inst_7671 ( .D(net_6705), .QN(net_185), .CK(net_15353) );
INV_X2 inst_7029 ( .ZN(net_1486), .A(net_1485) );
OAI211_X2 inst_2130 ( .C2(net_6778), .ZN(net_6718), .A(net_6343), .B(net_6082), .C1(net_373) );
XNOR2_X2 inst_359 ( .ZN(net_2772), .B(net_2299), .A(net_2044) );
DFF_X2 inst_8239 ( .Q(net_10502), .D(net_4879), .CK(net_15210) );
NAND2_X2 inst_4388 ( .ZN(net_5166), .A1(net_3123), .A2(net_183) );
OAI22_X2 inst_1055 ( .B2(net_10345), .A1(net_10344), .ZN(net_7458), .A2(net_7457), .B1(net_3214) );
CLKBUF_X2 inst_12382 ( .A(net_12300), .Z(net_12301) );
CLKBUF_X2 inst_13114 ( .A(net_12252), .Z(net_13033) );
OAI211_X2 inst_2100 ( .C2(net_6778), .ZN(net_6748), .A(net_6375), .B(net_6106), .C1(net_434) );
OAI211_X2 inst_2284 ( .C1(net_7108), .C2(net_6542), .ZN(net_6195), .B(net_5721), .A(net_3679) );
OAI21_X2 inst_1962 ( .B1(net_9106), .ZN(net_4332), .B2(net_3703), .A(net_3531) );
INV_X4 inst_4829 ( .A(net_7157), .ZN(net_5637) );
INV_X4 inst_4757 ( .A(net_7663), .ZN(net_4307) );
OR2_X2 inst_923 ( .ZN(net_4688), .A1(net_3136), .A2(net_3135) );
CLKBUF_X2 inst_13037 ( .A(net_12955), .Z(net_12956) );
CLKBUF_X2 inst_12153 ( .A(net_10964), .Z(net_12072) );
CLKBUF_X2 inst_13582 ( .A(net_13500), .Z(net_13501) );
AND2_X2 inst_10492 ( .ZN(net_6987), .A2(net_6986), .A1(net_1411) );
DFF_X1 inst_8671 ( .D(net_6750), .QN(net_131), .CK(net_13277) );
CLKBUF_X2 inst_11551 ( .A(net_11469), .Z(net_11470) );
DFF_X1 inst_8599 ( .Q(net_9687), .D(net_7299), .CK(net_15249) );
CLKBUF_X2 inst_15334 ( .A(net_15252), .Z(net_15253) );
CLKBUF_X2 inst_11604 ( .A(net_11522), .Z(net_11523) );
CLKBUF_X2 inst_12925 ( .A(net_12843), .Z(net_12844) );
INV_X4 inst_5283 ( .A(net_3173), .ZN(net_1325) );
CLKBUF_X2 inst_15635 ( .A(net_15553), .Z(net_15554) );
CLKBUF_X2 inst_13470 ( .A(net_13388), .Z(net_13389) );
INV_X2 inst_6975 ( .ZN(net_1685), .A(net_1684) );
DFF_X2 inst_8168 ( .QN(net_9831), .D(net_5047), .CK(net_14444) );
INV_X4 inst_6174 ( .A(net_10027), .ZN(net_842) );
CLKBUF_X2 inst_11819 ( .A(net_11262), .Z(net_11738) );
DFF_X2 inst_7564 ( .QN(net_9247), .D(net_7613), .CK(net_11263) );
XNOR2_X2 inst_194 ( .B(net_5798), .ZN(net_5199), .A(net_4939) );
DFF_X1 inst_8421 ( .D(net_8753), .Q(net_246), .CK(net_12690) );
INV_X2 inst_7109 ( .A(net_9354), .ZN(net_1012) );
INV_X4 inst_5890 ( .A(net_1211), .ZN(net_611) );
NAND2_X2 inst_3453 ( .A1(net_9496), .A2(net_8473), .ZN(net_8471) );
DFF_X1 inst_8793 ( .Q(net_9133), .D(net_4334), .CK(net_10605) );
DFF_X2 inst_7686 ( .QN(net_9202), .D(net_6557), .CK(net_11334) );
CLKBUF_X2 inst_12946 ( .A(net_10962), .Z(net_12865) );
NAND2_X2 inst_3766 ( .A2(net_9160), .A1(net_9151), .ZN(net_6184) );
CLKBUF_X2 inst_15594 ( .A(net_15258), .Z(net_15513) );
CLKBUF_X2 inst_12480 ( .A(net_12398), .Z(net_12399) );
CLKBUF_X2 inst_14181 ( .A(net_14099), .Z(net_14100) );
INV_X4 inst_5935 ( .A(net_10529), .ZN(net_955) );
DFF_X1 inst_8714 ( .Q(net_9208), .D(net_6640), .CK(net_11357) );
INV_X4 inst_6136 ( .ZN(net_3123), .A(net_184) );
DFF_X2 inst_7704 ( .Q(net_10005), .D(net_6446), .CK(net_12583) );
CLKBUF_X2 inst_11317 ( .A(net_11235), .Z(net_11236) );
NOR2_X2 inst_2536 ( .A2(net_9595), .ZN(net_8146), .A1(net_8116) );
CLKBUF_X2 inst_11730 ( .A(net_10653), .Z(net_11649) );
CLKBUF_X2 inst_13103 ( .A(net_10713), .Z(net_13022) );
AOI22_X2 inst_9389 ( .B1(net_9804), .A1(net_5766), .B2(net_5765), .ZN(net_5434), .A2(net_242) );
INV_X2 inst_7100 ( .A(net_10327), .ZN(net_1061) );
XNOR2_X2 inst_442 ( .B(net_9304), .ZN(net_918), .A(net_212) );
AOI22_X2 inst_9618 ( .A1(net_9849), .B1(net_9786), .A2(net_6413), .ZN(net_3435), .B2(net_2462) );
NOR2_X2 inst_2507 ( .A2(net_8424), .ZN(net_8422), .A1(net_8240) );
AOI22_X2 inst_9337 ( .B1(net_9813), .A2(net_5766), .B2(net_5765), .ZN(net_5615), .A1(net_251) );
DFF_X2 inst_8338 ( .Q(net_9616), .D(net_3244), .CK(net_13545) );
OAI211_X2 inst_2245 ( .C1(net_7237), .C2(net_6542), .ZN(net_6459), .B(net_5603), .A(net_3679) );
CLKBUF_X2 inst_14751 ( .A(net_13831), .Z(net_14670) );
CLKBUF_X2 inst_15467 ( .A(net_15385), .Z(net_15386) );
CLKBUF_X2 inst_14036 ( .A(net_13954), .Z(net_13955) );
CLKBUF_X2 inst_12620 ( .A(net_11291), .Z(net_12539) );
INV_X2 inst_6870 ( .ZN(net_3046), .A(net_3045) );
INV_X4 inst_5237 ( .ZN(net_1926), .A(net_1477) );
CLKBUF_X2 inst_13300 ( .A(net_13218), .Z(net_13219) );
INV_X4 inst_5915 ( .ZN(net_1370), .A(net_1015) );
INV_X4 inst_6097 ( .A(net_10434), .ZN(net_2702) );
CLKBUF_X2 inst_10998 ( .A(net_10916), .Z(net_10917) );
OAI21_X2 inst_1925 ( .B2(net_10279), .ZN(net_4514), .B1(net_3741), .A(x3772) );
NAND2_X2 inst_4298 ( .A2(net_10230), .A1(net_10229), .ZN(net_1684) );
CLKBUF_X2 inst_14593 ( .A(net_12287), .Z(net_14512) );
CLKBUF_X2 inst_11242 ( .A(net_11160), .Z(net_11161) );
XOR2_X2 inst_40 ( .A(net_9230), .Z(net_1713), .B(net_1440) );
MUX2_X1 inst_4437 ( .S(net_6041), .A(net_309), .B(x4117), .Z(x46) );
INV_X2 inst_7212 ( .A(net_9238), .ZN(net_451) );
OAI22_X2 inst_1249 ( .B1(net_7229), .ZN(net_4827), .A2(net_4826), .B2(net_4825), .A1(net_450) );
CLKBUF_X2 inst_15815 ( .A(net_15733), .Z(net_15734) );
NAND2_X2 inst_4099 ( .ZN(net_2842), .A2(net_2463), .A1(net_447) );
DFF_X1 inst_8765 ( .Q(net_10450), .D(net_5008), .CK(net_11078) );
INV_X4 inst_5403 ( .A(net_6314), .ZN(net_1164) );
INV_X4 inst_4740 ( .ZN(net_7142), .A(net_4452) );
OAI222_X2 inst_1416 ( .A2(net_7665), .C2(net_7664), .B2(net_7663), .ZN(net_5194), .A1(net_2632), .B1(net_1888), .C1(net_1547) );
INV_X4 inst_5967 ( .A(net_10032), .ZN(net_1107) );
CLKBUF_X2 inst_12066 ( .A(net_11984), .Z(net_11985) );
OAI22_X2 inst_1318 ( .A2(net_2878), .B2(net_2134), .ZN(net_2130), .B1(net_2129), .A1(net_1308) );
INV_X2 inst_7219 ( .A(net_8825), .ZN(net_438) );
INV_X2 inst_6894 ( .ZN(net_2591), .A(net_2590) );
INV_X2 inst_7280 ( .A(net_8965), .ZN(net_8964) );
XNOR2_X2 inst_439 ( .ZN(net_1039), .A(net_217), .B(net_194) );
CLKBUF_X2 inst_11567 ( .A(net_11485), .Z(net_11486) );
INV_X8 inst_4529 ( .A(net_9061), .ZN(net_9060) );
CLKBUF_X2 inst_15216 ( .A(net_12593), .Z(net_15135) );
INV_X4 inst_4584 ( .ZN(net_8066), .A(net_8024) );
OAI22_X2 inst_1070 ( .B2(net_10378), .ZN(net_6907), .A2(net_6629), .A1(net_6628), .B1(net_6047) );
CLKBUF_X2 inst_12037 ( .A(net_10755), .Z(net_11956) );
NOR3_X2 inst_2454 ( .A1(net_9523), .A2(net_9522), .ZN(net_3625), .A3(net_1026) );
CLKBUF_X2 inst_12255 ( .A(net_12173), .Z(net_12174) );
DFF_X2 inst_8280 ( .QN(net_10248), .D(net_4923), .CK(net_12181) );
NAND2_X2 inst_3601 ( .ZN(net_7265), .A2(net_6858), .A1(net_6604) );
CLKBUF_X2 inst_14612 ( .A(net_14530), .Z(net_14531) );
AOI222_X1 inst_9693 ( .B1(net_9504), .ZN(net_8288), .A2(net_8286), .B2(net_8285), .C2(net_8284), .C1(net_8220), .A1(x1792) );
INV_X4 inst_4536 ( .ZN(net_8731), .A(net_8726) );
CLKBUF_X2 inst_13309 ( .A(net_10667), .Z(net_13228) );
CLKBUF_X2 inst_13475 ( .A(net_13393), .Z(net_13394) );
AOI22_X2 inst_9478 ( .A1(net_10186), .B1(net_9813), .A2(net_4217), .ZN(net_3845), .B2(net_2556) );
CLKBUF_X2 inst_11854 ( .A(net_11772), .Z(net_11773) );
INV_X4 inst_5601 ( .A(net_3739), .ZN(net_1681) );
INV_X2 inst_6763 ( .ZN(net_6187), .A(net_6186) );
SDFF_X2 inst_654 ( .SI(net_9488), .Q(net_9488), .SE(net_3073), .CK(net_12424), .D(x2165) );
OAI221_X2 inst_1673 ( .C1(net_7219), .B2(net_5642), .ZN(net_5496), .C2(net_4905), .A(net_3527), .B1(net_917) );
INV_X4 inst_5745 ( .A(net_7333), .ZN(net_923) );
CLKBUF_X2 inst_13616 ( .A(net_13534), .Z(net_13535) );
CLKBUF_X2 inst_15163 ( .A(net_12524), .Z(net_15082) );
CLKBUF_X2 inst_14373 ( .A(net_14291), .Z(net_14292) );
CLKBUF_X2 inst_13656 ( .A(net_12302), .Z(net_13575) );
OAI221_X2 inst_1708 ( .ZN(net_4102), .B1(net_4101), .C1(net_4100), .A(net_3627), .B2(net_3143), .C2(net_2765) );
CLKBUF_X2 inst_15264 ( .A(net_15182), .Z(net_15183) );
OAI22_X2 inst_1153 ( .A1(net_7139), .A2(net_5139), .B2(net_5138), .ZN(net_5120), .B1(net_431) );
DFF_X2 inst_7959 ( .QN(net_10203), .D(net_5629), .CK(net_13247) );
DFF_X2 inst_7632 ( .D(net_6761), .QN(net_122), .CK(net_13340) );
NAND2_X2 inst_3823 ( .A2(net_9530), .ZN(net_4907), .A1(net_797) );
CLKBUF_X2 inst_15096 ( .A(net_15014), .Z(net_15015) );
CLKBUF_X2 inst_10905 ( .A(net_10823), .Z(net_10824) );
INV_X1 inst_7325 ( .A(net_8847), .ZN(x472) );
XNOR2_X2 inst_391 ( .B(net_9222), .ZN(net_2171), .A(net_1845) );
CLKBUF_X2 inst_11997 ( .A(net_11915), .Z(net_11916) );
NAND2_X2 inst_4107 ( .A2(net_8913), .ZN(net_2370), .A1(net_2369) );
CLKBUF_X2 inst_15020 ( .A(net_11838), .Z(net_14939) );
AND2_X4 inst_10440 ( .ZN(net_3293), .A1(net_1848), .A2(net_782) );
CLKBUF_X2 inst_11004 ( .A(net_10718), .Z(net_10923) );
NOR2_X2 inst_2738 ( .ZN(net_4152), .A2(net_3701), .A1(net_3298) );
SDFF_X2 inst_634 ( .Q(net_9466), .D(net_9466), .SE(net_3293), .CK(net_11893), .SI(x1547) );
NAND4_X2 inst_3122 ( .ZN(net_3345), .A2(net_3344), .A1(net_2855), .A3(net_2736), .A4(net_1731) );
CLKBUF_X2 inst_15229 ( .A(net_14866), .Z(net_15148) );
CLKBUF_X2 inst_14092 ( .A(net_14010), .Z(net_14011) );
AOI22_X2 inst_9090 ( .A1(net_9703), .ZN(net_6403), .A2(net_6402), .B2(net_5263), .B1(net_143) );
CLKBUF_X2 inst_10896 ( .A(net_10814), .Z(net_10815) );
DFF_X2 inst_8035 ( .Q(net_9229), .D(net_5450), .CK(net_11812) );
AOI22_X2 inst_9232 ( .A1(net_9896), .B1(net_9797), .A2(net_8042), .B2(net_6133), .ZN(net_6079) );
AND2_X4 inst_10420 ( .ZN(net_4394), .A2(net_4253), .A1(net_4110) );
INV_X4 inst_6074 ( .ZN(net_7182), .A(x4937) );
OAI221_X2 inst_1477 ( .ZN(net_7673), .B1(net_7672), .C2(net_7671), .A(net_7587), .C1(net_7434), .B2(net_4321) );
CLKBUF_X2 inst_13774 ( .A(net_13692), .Z(net_13693) );
AOI22_X2 inst_9263 ( .B2(net_10341), .A1(net_10340), .ZN(net_5932), .A2(net_5186), .B1(net_4927) );
DFF_X2 inst_8403 ( .Q(net_9154), .CK(net_11296), .D(x3606) );
INV_X2 inst_7043 ( .ZN(net_1360), .A(net_1359) );
OAI21_X2 inst_1799 ( .ZN(net_7375), .A(net_7374), .B2(net_6563), .B1(net_5331) );
AOI221_X2 inst_9813 ( .B1(net_9962), .A(net_7090), .B2(net_7089), .C2(net_7088), .ZN(net_6989), .C1(net_6808) );
SDFF_X2 inst_529 ( .SI(net_9339), .Q(net_9284), .D(net_9284), .SE(net_7588), .CK(net_14669) );
CLKBUF_X2 inst_15129 ( .A(net_15047), .Z(net_15048) );
MUX2_X1 inst_4442 ( .S(net_6041), .A(net_304), .B(x4520), .Z(x86) );
DFF_X2 inst_7385 ( .D(net_8657), .QN(net_269), .CK(net_12640) );
OAI221_X2 inst_1528 ( .B1(net_10200), .B2(net_7295), .C2(net_7293), .ZN(net_7246), .C1(net_7245), .A(net_6835) );
CLKBUF_X2 inst_11192 ( .A(net_11110), .Z(net_11111) );
AOI22_X2 inst_9326 ( .B1(net_9991), .A1(net_6834), .A2(net_5743), .B2(net_5742), .ZN(net_5649) );
CLKBUF_X2 inst_15705 ( .A(net_15623), .Z(net_15624) );
NAND2_X2 inst_3458 ( .A1(net_9465), .A2(net_8475), .ZN(net_8466) );
INV_X4 inst_5788 ( .ZN(net_7504), .A(net_7336) );
CLKBUF_X2 inst_11788 ( .A(net_11706), .Z(net_11707) );
INV_X4 inst_4694 ( .ZN(net_4833), .A(net_4649) );
OAI22_X2 inst_1313 ( .ZN(net_2238), .A1(net_2237), .B2(net_2236), .B1(net_1365), .A2(net_1138) );
CLKBUF_X2 inst_15460 ( .A(net_12773), .Z(net_15379) );
CLKBUF_X2 inst_14267 ( .A(net_14185), .Z(net_14186) );
CLKBUF_X2 inst_11030 ( .A(net_10948), .Z(net_10949) );
CLKBUF_X2 inst_14572 ( .A(net_14490), .Z(net_14491) );
CLKBUF_X2 inst_11104 ( .A(net_11022), .Z(net_11023) );
DFF_X2 inst_8098 ( .QN(net_9834), .D(net_5030), .CK(net_11735) );
SDFF_X2 inst_675 ( .SI(net_9484), .Q(net_9484), .SE(net_3073), .CK(net_14131), .D(x2400) );
DFF_X1 inst_8632 ( .Q(net_9880), .D(net_7197), .CK(net_12164) );
NAND2_X2 inst_4068 ( .A2(net_3695), .A1(net_3692), .ZN(net_3058) );
CLKBUF_X2 inst_11953 ( .A(net_11871), .Z(net_11872) );
CLKBUF_X2 inst_13706 ( .A(net_13624), .Z(net_13625) );
INV_X4 inst_5729 ( .ZN(net_841), .A(net_754) );
NAND2_X2 inst_4116 ( .ZN(net_2350), .A1(net_2349), .A2(net_1633) );
NOR2_X2 inst_2886 ( .ZN(net_2532), .A2(net_1785), .A1(net_1211) );
CLKBUF_X2 inst_15146 ( .A(net_15064), .Z(net_15065) );
NOR2_X2 inst_2705 ( .ZN(net_4752), .A2(net_4325), .A1(net_4323) );
CLKBUF_X2 inst_14851 ( .A(net_14057), .Z(net_14770) );
INV_X4 inst_6523 ( .A(net_9747), .ZN(net_341) );
INV_X4 inst_5150 ( .ZN(net_1904), .A(net_1585) );
CLKBUF_X2 inst_13291 ( .A(net_13209), .Z(net_13210) );
CLKBUF_X2 inst_13747 ( .A(net_13665), .Z(net_13666) );
CLKBUF_X2 inst_12902 ( .A(net_12263), .Z(net_12821) );
AOI22_X2 inst_9613 ( .B1(net_10291), .A2(net_6413), .B2(net_4774), .ZN(net_3440), .A1(net_688) );
CLKBUF_X2 inst_12924 ( .A(net_12842), .Z(net_12843) );
CLKBUF_X2 inst_10978 ( .A(net_10896), .Z(net_10897) );
INV_X4 inst_5737 ( .A(net_1088), .ZN(net_986) );
CLKBUF_X2 inst_13199 ( .A(net_13117), .Z(net_13118) );
INV_X4 inst_5332 ( .ZN(net_5452), .A(net_1453) );
NOR2_X2 inst_2773 ( .ZN(net_3231), .A2(net_3230), .A1(net_2134) );
OAI211_X2 inst_2081 ( .C2(net_6778), .ZN(net_6767), .A(net_6394), .B(net_6127), .C1(net_337) );
NAND3_X2 inst_3261 ( .ZN(net_4698), .A1(net_4412), .A3(net_4411), .A2(net_3134) );
DFF_X1 inst_8717 ( .Q(net_9543), .D(net_6985), .CK(net_12762) );
CLKBUF_X2 inst_13606 ( .A(net_10791), .Z(net_13525) );
CLKBUF_X2 inst_15796 ( .A(net_15714), .Z(net_15715) );
CLKBUF_X2 inst_11144 ( .A(net_11062), .Z(net_11063) );
OAI22_X2 inst_1211 ( .A1(net_7192), .A2(net_5134), .B2(net_5133), .ZN(net_5038), .B1(net_2630) );
AOI22_X2 inst_9078 ( .B1(net_9677), .A1(net_6684), .B2(net_6683), .ZN(net_6558), .A2(net_246) );
NAND2_X2 inst_3751 ( .ZN(net_5299), .A2(net_4777), .A1(net_3773) );
OAI22_X2 inst_1192 ( .A1(net_7127), .A2(net_5107), .B2(net_5105), .ZN(net_5062), .B1(net_5061) );
OR4_X4 inst_682 ( .A4(net_4631), .A2(net_4460), .ZN(net_4454), .A1(net_4333), .A3(net_4332) );
XNOR2_X2 inst_238 ( .ZN(net_4259), .A(net_4258), .B(net_1771) );
CLKBUF_X2 inst_12463 ( .A(net_12381), .Z(net_12382) );
CLKBUF_X2 inst_12394 ( .A(net_11633), .Z(net_12313) );
INV_X2 inst_6735 ( .ZN(net_7416), .A(net_7334) );
INV_X4 inst_6643 ( .ZN(net_9091), .A(net_9088) );
AOI22_X2 inst_9123 ( .A1(net_9707), .A2(net_6420), .ZN(net_6366), .B2(net_5263), .B1(net_147) );
OAI211_X2 inst_2222 ( .C1(net_7241), .C2(net_6501), .ZN(net_6483), .B(net_5558), .A(net_3679) );
INV_X4 inst_4578 ( .ZN(net_8072), .A(net_8032) );
NAND2_X4 inst_3333 ( .A2(net_9021), .A1(net_9020), .ZN(net_8581) );
AOI21_X2 inst_10021 ( .ZN(net_8299), .A(net_8082), .B2(net_7986), .B1(net_1974) );
CLKBUF_X2 inst_12102 ( .A(net_12020), .Z(net_12021) );
NAND2_X2 inst_4059 ( .A2(net_3630), .ZN(net_3187), .A1(net_949) );
NAND4_X2 inst_3109 ( .ZN(net_4334), .A4(net_3863), .A2(net_3778), .A1(net_3408), .A3(net_3407) );
AOI21_X2 inst_10046 ( .B1(net_9531), .B2(net_9503), .ZN(net_7426), .A(net_2228) );
OAI21_X2 inst_1755 ( .A(net_9575), .B2(net_9574), .ZN(net_8533), .B1(net_1533) );
CLKBUF_X2 inst_14995 ( .A(net_14913), .Z(net_14914) );
OAI211_X2 inst_2240 ( .C1(net_7192), .C2(net_6480), .ZN(net_6464), .B(net_5526), .A(net_3679) );
CLKBUF_X2 inst_11680 ( .A(net_11598), .Z(net_11599) );
OAI22_X2 inst_1210 ( .A1(net_7190), .A2(net_5151), .B2(net_5150), .ZN(net_5039), .B1(net_3353) );
INV_X4 inst_6090 ( .A(net_10391), .ZN(net_496) );
CLKBUF_X2 inst_14674 ( .A(net_14592), .Z(net_14593) );
CLKBUF_X2 inst_12759 ( .A(net_12536), .Z(net_12678) );
CLKBUF_X2 inst_15390 ( .A(net_15308), .Z(net_15309) );
CLKBUF_X2 inst_15154 ( .A(net_13888), .Z(net_15073) );
CLKBUF_X2 inst_15027 ( .A(net_14945), .Z(net_14946) );
NOR3_X2 inst_2437 ( .A1(net_9045), .ZN(net_3099), .A2(net_2849), .A3(net_1231) );
CLKBUF_X2 inst_12715 ( .A(net_12633), .Z(net_12634) );
OR2_X4 inst_806 ( .A1(net_10156), .ZN(net_1770), .A2(net_1374) );
INV_X8 inst_4521 ( .A(net_8933), .ZN(net_8932) );
DFF_X2 inst_8324 ( .Q(net_9618), .D(net_3517), .CK(net_14071) );
INV_X2 inst_7119 ( .ZN(net_1283), .A(net_952) );
OAI21_X2 inst_1981 ( .ZN(net_3607), .A(net_2756), .B2(net_1789), .B1(net_313) );
INV_X2 inst_7232 ( .A(net_9386), .ZN(net_657) );
INV_X4 inst_6324 ( .A(net_9840), .ZN(net_417) );
SDFF_X2 inst_491 ( .SE(net_9540), .SI(net_8218), .Q(net_307), .D(net_307), .CK(net_11657) );
INV_X4 inst_5960 ( .ZN(net_7192), .A(x5961) );
AND2_X2 inst_10485 ( .ZN(net_9005), .A1(net_8968), .A2(net_8397) );
INV_X4 inst_6027 ( .A(net_9532), .ZN(net_751) );
INV_X4 inst_4943 ( .ZN(net_7095), .A(net_6165) );
CLKBUF_X2 inst_13219 ( .A(net_13137), .Z(net_13138) );
CLKBUF_X2 inst_13515 ( .A(net_13433), .Z(net_13434) );
CLKBUF_X2 inst_15122 ( .A(net_15040), .Z(net_15041) );
DFF_X2 inst_8309 ( .QN(net_9160), .D(net_4289), .CK(net_11810) );
CLKBUF_X2 inst_10987 ( .A(net_10905), .Z(net_10906) );
NAND2_X2 inst_3775 ( .ZN(net_5879), .A1(net_4784), .A2(net_4783) );
CLKBUF_X2 inst_13762 ( .A(net_13680), .Z(net_13681) );
CLKBUF_X2 inst_14900 ( .A(net_14818), .Z(net_14819) );
CLKBUF_X2 inst_12097 ( .A(net_11765), .Z(net_12016) );
NOR2_X4 inst_2472 ( .ZN(net_9027), .A2(net_8906), .A1(net_8905) );
AOI22_X2 inst_9441 ( .A1(net_6892), .B2(net_6625), .ZN(net_6427), .B1(net_4273), .A2(net_3519) );
NAND4_X2 inst_3086 ( .ZN(net_4501), .A4(net_4059), .A1(net_3282), .A3(net_3190), .A2(net_2742) );
NOR2_X2 inst_2791 ( .ZN(net_3423), .A2(net_3015), .A1(net_557) );
CLKBUF_X2 inst_12090 ( .A(net_12008), .Z(net_12009) );
CLKBUF_X2 inst_11239 ( .A(net_11152), .Z(net_11158) );
INV_X4 inst_5583 ( .A(net_908), .ZN(net_887) );
AOI21_X2 inst_10243 ( .ZN(net_8863), .B1(net_2404), .B2(net_2403), .A(net_2402) );
DFF_X2 inst_8293 ( .QN(net_10092), .D(net_5235), .CK(net_10876) );
OR2_X2 inst_872 ( .A2(net_7557), .ZN(net_6981), .A1(net_6949) );
INV_X4 inst_6641 ( .A(net_9082), .ZN(net_9080) );
CLKBUF_X2 inst_15633 ( .A(net_15551), .Z(net_15552) );
CLKBUF_X2 inst_14814 ( .A(net_11727), .Z(net_14733) );
CLKBUF_X2 inst_14821 ( .A(net_14739), .Z(net_14740) );
CLKBUF_X2 inst_11479 ( .A(net_10762), .Z(net_11398) );
AOI22_X2 inst_9210 ( .A1(net_9892), .B1(net_9793), .B2(net_6133), .A2(net_6111), .ZN(net_6101) );
NAND2_X1 inst_4419 ( .ZN(net_8742), .A2(net_8741), .A1(net_8619) );
INV_X4 inst_5234 ( .ZN(net_1921), .A(net_1483) );
CLKBUF_X2 inst_14907 ( .A(net_10626), .Z(net_14826) );
CLKBUF_X2 inst_12579 ( .A(net_12236), .Z(net_12498) );
INV_X2 inst_6850 ( .ZN(net_3393), .A(net_3392) );
OAI221_X2 inst_1667 ( .C1(net_7224), .C2(net_5520), .ZN(net_5502), .B2(net_4547), .B1(net_4373), .A(net_3731) );
CLKBUF_X2 inst_15375 ( .A(net_12705), .Z(net_15294) );
INV_X2 inst_6698 ( .ZN(net_8240), .A(net_8239) );
OAI222_X2 inst_1349 ( .B1(net_7732), .A2(net_7731), .C2(net_7730), .ZN(net_7432), .B2(net_7042), .A1(net_4681), .C1(net_768) );
CLKBUF_X2 inst_15339 ( .A(net_15257), .Z(net_15258) );
SDFF_X2 inst_462 ( .SE(net_8747), .SI(net_8696), .Q(net_239), .D(net_108), .CK(net_13852) );
INV_X2 inst_7012 ( .A(net_5993), .ZN(net_1593) );
CLKBUF_X2 inst_12744 ( .A(net_11651), .Z(net_12663) );
AOI211_X2 inst_10261 ( .ZN(net_7933), .C2(net_7932), .B(net_7804), .A(net_7520), .C1(net_3977) );
NAND2_X2 inst_3745 ( .ZN(net_5305), .A2(net_4766), .A1(net_4055) );
CLKBUF_X2 inst_15345 ( .A(net_12501), .Z(net_15264) );
AOI22_X2 inst_9398 ( .B2(net_10446), .A1(net_10445), .ZN(net_5385), .A2(net_4678), .B1(net_4554) );
INV_X4 inst_5572 ( .ZN(net_1221), .A(net_907) );
NAND2_X2 inst_4347 ( .A2(net_9833), .ZN(net_2034), .A1(net_962) );
AND2_X2 inst_10579 ( .A1(net_10437), .A2(net_3492), .ZN(net_2762) );
INV_X2 inst_7223 ( .A(net_9419), .ZN(net_8215) );
INV_X4 inst_5962 ( .A(net_10248), .ZN(net_745) );
OAI211_X2 inst_2224 ( .C1(net_7186), .ZN(net_6481), .C2(net_6480), .B(net_5532), .A(net_3527) );
CLKBUF_X2 inst_13381 ( .A(net_13299), .Z(net_13300) );
AOI21_X4 inst_10002 ( .A(net_9046), .ZN(net_3059), .B2(net_2420), .B1(net_2218) );
AOI21_X2 inst_10185 ( .ZN(net_3424), .A(net_3423), .B2(net_3015), .B1(net_1075) );
INV_X2 inst_6661 ( .ZN(net_8367), .A(net_8313) );
INV_X4 inst_5226 ( .A(net_2205), .ZN(net_1935) );
CLKBUF_X2 inst_13012 ( .A(net_12930), .Z(net_12931) );
AND2_X4 inst_10389 ( .ZN(net_7326), .A2(net_7325), .A1(net_1154) );
INV_X4 inst_4909 ( .A(net_3103), .ZN(net_2838) );
INV_X2 inst_7114 ( .A(net_1367), .ZN(net_997) );
INV_X4 inst_5310 ( .ZN(net_1288), .A(net_685) );
INV_X2 inst_6836 ( .ZN(net_3893), .A(net_3892) );
DFF_X1 inst_8412 ( .Q(net_9604), .D(net_8795), .CK(net_15192) );
DFF_X2 inst_7611 ( .QN(net_9346), .D(net_7132), .CK(net_15282) );
OAI21_X2 inst_1914 ( .A(net_4679), .ZN(net_4609), .B2(net_4306), .B1(net_1512) );
CLKBUF_X2 inst_14702 ( .A(net_14620), .Z(net_14621) );
INV_X4 inst_6219 ( .A(net_9295), .ZN(net_3311) );
INV_X4 inst_4996 ( .ZN(net_2578), .A(net_1975) );
OAI21_X2 inst_1975 ( .ZN(net_4671), .A(net_2958), .B1(net_2873), .B2(net_1981) );
OAI21_X2 inst_1890 ( .B1(net_7243), .ZN(net_4863), .B2(net_4862), .A(net_4535) );
NOR4_X2 inst_2308 ( .ZN(net_7601), .A2(net_7438), .A4(net_4086), .A3(net_3915), .A1(net_2191) );
INV_X4 inst_6647 ( .ZN(net_9109), .A(net_577) );
NAND2_X2 inst_4093 ( .ZN(net_2833), .A1(net_2545), .A2(net_2544) );
AOI222_X1 inst_9728 ( .B1(net_10292), .C1(net_9980), .A2(net_6413), .B2(net_4774), .ZN(net_3627), .C2(net_2541), .A1(net_2021) );
INV_X4 inst_4806 ( .ZN(net_4229), .A(net_3617) );
AOI22_X2 inst_9585 ( .A1(net_10068), .B1(net_10016), .A2(net_5320), .ZN(net_3575), .B2(net_2468) );
NOR2_X2 inst_2879 ( .ZN(net_2720), .A2(net_1884), .A1(net_1643) );
DFF_X2 inst_8117 ( .Q(net_9175), .D(net_5083), .CK(net_11242) );
CLKBUF_X2 inst_14676 ( .A(net_14594), .Z(net_14595) );
CLKBUF_X2 inst_12362 ( .A(net_12280), .Z(net_12281) );
DFF_X2 inst_7482 ( .D(net_8064), .Q(net_217), .CK(net_12528) );
NOR4_X2 inst_2338 ( .ZN(net_4974), .A2(net_4499), .A1(net_4356), .A4(net_4355), .A3(net_3317) );
CLKBUF_X2 inst_11893 ( .A(net_11811), .Z(net_11812) );
NAND2_X2 inst_3475 ( .A1(net_9454), .A2(net_8951), .ZN(net_8903) );
NOR2_X2 inst_3017 ( .A2(net_9525), .A1(net_9524), .ZN(net_1025) );
INV_X4 inst_6389 ( .A(net_10154), .ZN(net_631) );
CLKBUF_X2 inst_13170 ( .A(net_13088), .Z(net_13089) );
CLKBUF_X2 inst_15547 ( .A(net_15465), .Z(net_15466) );
DFF_X2 inst_7818 ( .Q(net_9994), .D(net_6462), .CK(net_13196) );
CLKBUF_X2 inst_11431 ( .A(net_10848), .Z(net_11350) );
OR2_X2 inst_845 ( .A1(net_9586), .A2(net_9585), .ZN(net_8776) );
NAND2_X2 inst_3554 ( .ZN(net_7904), .A2(net_7790), .A1(net_7635) );
OAI222_X2 inst_1367 ( .B1(net_7732), .A2(net_7731), .C2(net_7730), .ZN(net_6283), .B2(net_5739), .A1(net_4133), .C1(net_2089) );
INV_X4 inst_6516 ( .A(net_10291), .ZN(net_347) );
DFF_X1 inst_8649 ( .Q(net_8838), .D(net_7302), .CK(net_12312) );
INV_X4 inst_5198 ( .ZN(net_5175), .A(net_1189) );
INV_X4 inst_5909 ( .A(net_1948), .ZN(net_969) );
CLKBUF_X2 inst_10980 ( .A(net_10898), .Z(net_10899) );
AOI22_X2 inst_9175 ( .A1(net_9900), .B1(net_9801), .A2(net_8042), .B2(net_8041), .ZN(net_6143) );
CLKBUF_X2 inst_10898 ( .A(net_10816), .Z(net_10817) );
OAI21_X2 inst_2016 ( .ZN(net_8855), .B1(net_4409), .B2(net_2682), .A(net_2681) );
NAND2_X2 inst_3687 ( .A2(net_9264), .A1(net_8960), .ZN(net_6243) );
CLKBUF_X2 inst_15426 ( .A(net_15344), .Z(net_15345) );
CLKBUF_X2 inst_10837 ( .A(net_10627), .Z(net_10756) );
CLKBUF_X2 inst_15679 ( .A(net_15597), .Z(net_15598) );
CLKBUF_X2 inst_12723 ( .A(net_12641), .Z(net_12642) );
DFF_X1 inst_8434 ( .QN(net_9581), .D(net_8630), .CK(net_11558) );
NAND2_X2 inst_4012 ( .A1(net_9538), .ZN(net_3693), .A2(net_3084) );
AOI21_X2 inst_10103 ( .B1(net_10051), .B2(net_5174), .ZN(net_4898), .A(net_4501) );
NAND4_X2 inst_3053 ( .ZN(net_5871), .A4(net_4981), .A3(net_3792), .A2(net_3788), .A1(net_3759) );
DFF_X2 inst_8385 ( .QN(net_8839), .D(net_5464), .CK(net_11143) );
CLKBUF_X2 inst_15152 ( .A(net_11641), .Z(net_15071) );
AOI22_X2 inst_9289 ( .B1(net_9703), .A1(net_5755), .B2(net_5754), .ZN(net_5711), .A2(net_240) );
DFF_X2 inst_7630 ( .D(net_6765), .QN(net_119), .CK(net_12828) );
AOI221_X2 inst_9920 ( .ZN(net_5868), .B2(net_5867), .C1(net_5866), .A(net_5862), .C2(net_4725), .B1(x6102) );
DFF_X2 inst_7829 ( .Q(net_9818), .D(net_6512), .CK(net_15686) );
XNOR2_X2 inst_393 ( .B(net_9175), .ZN(net_2087), .A(net_1034) );
AND2_X4 inst_10409 ( .ZN(net_5758), .A2(net_4789), .A1(net_4788) );
INV_X4 inst_4810 ( .ZN(net_3562), .A(net_3398) );
AOI221_X2 inst_9962 ( .C1(net_10495), .B1(net_10285), .C2(net_6415), .B2(net_4774), .ZN(net_4769), .A(net_4340) );
INV_X4 inst_5969 ( .A(net_10302), .ZN(net_544) );
OAI21_X2 inst_1813 ( .ZN(net_6926), .B2(net_6660), .A(net_3200), .B1(net_2178) );
XNOR2_X2 inst_92 ( .ZN(net_8558), .A(net_8503), .B(net_8269) );
CLKBUF_X2 inst_15405 ( .A(net_10754), .Z(net_15324) );
CLKBUF_X2 inst_11168 ( .A(net_11086), .Z(net_11087) );
CLKBUF_X2 inst_10708 ( .A(net_10626), .Z(net_10627) );
XNOR2_X2 inst_345 ( .ZN(net_2863), .B(net_2862), .A(net_1577) );
NAND4_X2 inst_3103 ( .ZN(net_4340), .A2(net_3822), .A3(net_3821), .A1(net_3572), .A4(net_3571) );
AOI22_X2 inst_9086 ( .A1(net_9742), .A2(net_6420), .ZN(net_6409), .B1(net_6408), .B2(net_5263) );
CLKBUF_X2 inst_11985 ( .A(net_11903), .Z(net_11904) );
CLKBUF_X2 inst_11856 ( .A(net_11774), .Z(net_11775) );
DFF_X2 inst_7520 ( .QN(net_9237), .D(net_7830), .CK(net_11278) );
NAND3_X2 inst_3304 ( .ZN(net_2137), .A3(net_1446), .A2(net_958), .A1(net_803) );
AOI21_X2 inst_10233 ( .ZN(net_2310), .A(net_1820), .B1(net_1819), .B2(net_570) );
DFF_X2 inst_7762 ( .Q(net_9712), .D(net_6545), .CK(net_14234) );
AOI21_X2 inst_10087 ( .B2(net_9660), .B1(net_9659), .ZN(net_5894), .A(net_5329) );
INV_X4 inst_6362 ( .ZN(net_404), .A(net_280) );
INV_X4 inst_5384 ( .ZN(net_3631), .A(net_2318) );
DFF_X2 inst_8076 ( .QN(net_10470), .D(net_5307), .CK(net_11451) );
CLKBUF_X2 inst_13806 ( .A(net_12903), .Z(net_13725) );
CLKBUF_X2 inst_11009 ( .A(net_10927), .Z(net_10928) );
AND2_X2 inst_10585 ( .ZN(net_3022), .A2(net_2511), .A1(net_491) );
XOR2_X1 inst_57 ( .A(net_9350), .Z(net_1987), .B(net_1986) );
INV_X4 inst_4723 ( .ZN(net_4615), .A(net_4496) );
NAND2_X2 inst_3655 ( .A2(net_8659), .ZN(net_6656), .A1(net_6655) );
DFF_X2 inst_7532 ( .QN(net_9325), .D(net_7777), .CK(net_13049) );
CLKBUF_X2 inst_12145 ( .A(net_12063), .Z(net_12064) );
INV_X2 inst_6692 ( .ZN(net_8332), .A(net_8268) );
AOI22_X2 inst_9312 ( .B1(net_9717), .A1(net_6823), .A2(net_5755), .B2(net_5754), .ZN(net_5665) );
INV_X4 inst_6617 ( .A(net_8939), .ZN(net_8938) );
NOR2_X2 inst_2843 ( .A1(net_2576), .ZN(net_2319), .A2(net_1616) );
OAI21_X2 inst_1888 ( .B1(net_7785), .ZN(net_4900), .A(net_4507), .B2(net_4506) );
NAND2_X4 inst_3379 ( .ZN(net_3531), .A1(net_771), .A2(net_187) );
OAI21_X2 inst_1763 ( .ZN(net_8925), .A(net_8372), .B2(net_8371), .B1(net_8253) );
OAI22_X2 inst_1307 ( .A1(net_10354), .ZN(net_2411), .A2(net_2410), .B2(net_1652), .B1(net_939) );
CLKBUF_X2 inst_13071 ( .A(net_12602), .Z(net_12990) );
DFF_X2 inst_7759 ( .Q(net_9694), .D(net_6550), .CK(net_12061) );
CLKBUF_X2 inst_10878 ( .A(net_10796), .Z(net_10797) );
DFF_X1 inst_8565 ( .Q(net_9774), .D(net_7212), .CK(net_15568) );
INV_X2 inst_6789 ( .ZN(net_5797), .A(net_5796) );
INV_X2 inst_7190 ( .A(net_9413), .ZN(net_8220) );
CLKBUF_X2 inst_13685 ( .A(net_12132), .Z(net_13604) );
CLKBUF_X2 inst_14309 ( .A(net_14227), .Z(net_14228) );
OAI22_X2 inst_1094 ( .A1(net_9187), .ZN(net_6301), .A2(net_6299), .B2(net_6298), .B1(net_2786) );
CLKBUF_X2 inst_12960 ( .A(net_12878), .Z(net_12879) );
NAND2_X2 inst_4145 ( .ZN(net_2082), .A1(net_2081), .A2(net_1377) );
INV_X4 inst_4590 ( .A(net_8036), .ZN(net_7922) );
INV_X2 inst_7124 ( .A(net_1332), .ZN(net_934) );
INV_X4 inst_6376 ( .A(net_9838), .ZN(net_398) );
NAND2_X2 inst_3680 ( .ZN(net_7248), .A2(net_6205), .A1(net_5938) );
INV_X2 inst_7168 ( .A(net_9420), .ZN(net_8198) );
INV_X4 inst_4878 ( .ZN(net_3488), .A(net_3014) );
OAI221_X2 inst_1699 ( .C1(net_7221), .B2(net_5591), .ZN(net_5455), .B1(net_5454), .C2(net_4902), .A(net_3507) );
DFF_X1 inst_8616 ( .Q(net_9678), .D(net_7270), .CK(net_13287) );
OR2_X2 inst_851 ( .A2(net_9432), .ZN(net_8413), .A1(net_8412) );
CLKBUF_X2 inst_12685 ( .A(net_12603), .Z(net_12604) );
OR2_X4 inst_831 ( .A1(net_10530), .ZN(net_1121), .A2(net_561) );
XOR2_X2 inst_50 ( .A(net_9325), .B(net_9324), .Z(net_1772) );
CLKBUF_X2 inst_11762 ( .A(net_11680), .Z(net_11681) );
INV_X4 inst_5824 ( .ZN(net_1020), .A(net_839) );
NAND2_X2 inst_4264 ( .ZN(net_4115), .A2(net_1111), .A1(net_912) );
NOR2_X2 inst_2589 ( .ZN(net_7049), .A1(net_7048), .A2(net_6615) );
CLKBUF_X2 inst_10626 ( .A(net_10544), .Z(net_10545) );
CLKBUF_X2 inst_11448 ( .A(net_10964), .Z(net_11367) );
MUX2_X2 inst_4430 ( .B(net_9159), .S(net_7553), .Z(net_7496), .A(net_7495) );
DFF_X1 inst_8699 ( .D(net_6713), .Q(net_141), .CK(net_12833) );
OAI221_X2 inst_1650 ( .B1(net_10417), .C1(net_7136), .ZN(net_5538), .B2(net_4477), .C2(net_4455), .A(net_3731) );
CLKBUF_X2 inst_15007 ( .A(net_14925), .Z(net_14926) );
CLKBUF_X2 inst_11174 ( .A(net_11092), .Z(net_11093) );
OAI221_X2 inst_1497 ( .C2(net_9063), .B2(net_9056), .ZN(net_7366), .C1(net_7201), .A(net_7001), .B1(net_5462) );
DFF_X2 inst_8250 ( .Q(net_10179), .D(net_4836), .CK(net_12958) );
DFF_X2 inst_7469 ( .QN(net_9518), .D(net_8101), .CK(net_14968) );
MUX2_X1 inst_4439 ( .S(net_6041), .A(net_307), .B(x4285), .Z(x65) );
INV_X4 inst_5706 ( .A(net_1361), .ZN(net_774) );
NOR2_X2 inst_2872 ( .ZN(net_2505), .A2(net_1950), .A1(net_1073) );
DFF_X1 inst_8683 ( .D(net_6732), .Q(net_135), .CK(net_15442) );
OAI22_X2 inst_1002 ( .B2(net_8545), .ZN(net_8544), .A2(net_8456), .B1(net_8455), .A1(net_8203) );
CLKBUF_X2 inst_12076 ( .A(net_11994), .Z(net_11995) );
DFF_X2 inst_8057 ( .QN(net_10116), .D(net_5505), .CK(net_12332) );
CLKBUF_X2 inst_13179 ( .A(net_13097), .Z(net_13098) );
SDFF_X2 inst_478 ( .SE(net_9540), .SI(net_8231), .Q(net_281), .D(net_281), .CK(net_12713) );
DFF_X1 inst_8630 ( .Q(net_9790), .D(net_7214), .CK(net_13351) );
NAND2_X2 inst_3380 ( .A2(net_8912), .A1(net_8911), .ZN(net_8790) );
CLKBUF_X2 inst_15832 ( .A(net_15750), .Z(net_15751) );
INV_X4 inst_5666 ( .ZN(net_1141), .A(net_818) );
OR2_X4 inst_804 ( .ZN(net_2782), .A2(net_1378), .A1(net_1073) );
NAND3_X2 inst_3290 ( .A2(net_4041), .ZN(net_3057), .A3(net_3056), .A1(net_2941) );
CLKBUF_X2 inst_13953 ( .A(net_13871), .Z(net_13872) );
DFF_X1 inst_8824 ( .QN(net_9188), .D(net_2738), .CK(net_13598) );
XOR2_X2 inst_13 ( .Z(net_2870), .B(net_2869), .A(net_1975) );
CLKBUF_X2 inst_12173 ( .A(net_12091), .Z(net_12092) );
CLKBUF_X2 inst_14126 ( .A(net_14044), .Z(net_14045) );
INV_X4 inst_5378 ( .A(net_2938), .ZN(net_1584) );
NOR2_X2 inst_2584 ( .ZN(net_7064), .A2(net_6636), .A1(net_3745) );
INV_X4 inst_5665 ( .ZN(net_2249), .A(net_1370) );
INV_X4 inst_4931 ( .ZN(net_2875), .A(net_2604) );
CLKBUF_X2 inst_11540 ( .A(net_11458), .Z(net_11459) );
CLKBUF_X2 inst_15111 ( .A(net_15029), .Z(net_15030) );
CLKBUF_X2 inst_14527 ( .A(net_14445), .Z(net_14446) );
HA_X1 inst_7334 ( .S(net_7463), .CO(net_7462), .B(net_7308), .A(net_971) );
OR2_X4 inst_799 ( .A1(net_10259), .ZN(net_3112), .A2(net_1370) );
CLKBUF_X2 inst_12906 ( .A(net_12824), .Z(net_12825) );
NAND2_X2 inst_3481 ( .A2(net_9460), .A1(net_8951), .ZN(net_8876) );
OR2_X4 inst_738 ( .A2(net_9101), .ZN(net_9047), .A1(net_4901) );
CLKBUF_X2 inst_13666 ( .A(net_13584), .Z(net_13585) );
INV_X4 inst_6481 ( .ZN(net_572), .A(net_199) );
NOR2_X2 inst_2755 ( .A2(net_9197), .ZN(net_4224), .A1(net_3607) );
AOI22_X2 inst_9393 ( .A2(net_9093), .B2(net_9068), .ZN(net_5418), .B1(net_2938), .A1(net_1733) );
AOI22_X2 inst_9101 ( .A1(net_9663), .A2(net_6402), .ZN(net_6391), .B2(net_5263), .B1(net_101) );
OAI21_X2 inst_1819 ( .ZN(net_6635), .A(net_6634), .B1(net_6633), .B2(net_5971) );
CLKBUF_X2 inst_14718 ( .A(net_14636), .Z(net_14637) );
CLKBUF_X2 inst_14284 ( .A(net_11194), .Z(net_14203) );
XNOR2_X2 inst_255 ( .ZN(net_4105), .A(net_3474), .B(net_2025) );
NOR2_X2 inst_2726 ( .A1(net_9613), .ZN(net_3970), .A2(net_3330) );
XNOR2_X1 inst_453 ( .B(net_9843), .A(net_1413), .ZN(net_1410) );
SDFF_X2 inst_493 ( .SE(net_9540), .SI(net_8216), .Q(net_310), .D(net_310), .CK(net_11650) );
AND2_X2 inst_10555 ( .ZN(net_3655), .A2(net_3309), .A1(net_342) );
NOR2_X2 inst_2674 ( .ZN(net_5292), .A2(net_4785), .A1(net_3298) );
XOR2_X2 inst_23 ( .Z(net_2409), .B(net_2010), .A(net_1387) );
CLKBUF_X2 inst_14471 ( .A(net_14267), .Z(net_14390) );
AND2_X4 inst_10390 ( .ZN(net_7324), .A2(net_7323), .A1(net_1247) );
AOI211_X2 inst_10279 ( .C1(net_9050), .B(net_7110), .ZN(net_7094), .C2(net_6669), .A(net_3690) );
INV_X2 inst_6686 ( .ZN(net_8342), .A(net_8276) );
DFF_X1 inst_8784 ( .QN(net_9192), .D(net_4588), .CK(net_11349) );
OAI22_X2 inst_1113 ( .ZN(net_6261), .A2(net_5227), .B2(net_5226), .B1(net_3706), .A1(net_2641) );
OAI21_X2 inst_1822 ( .ZN(net_6611), .A(net_5941), .B2(net_5940), .B1(net_3984) );
NAND2_X2 inst_3790 ( .ZN(net_6678), .A2(net_5908), .A1(net_4634) );
CLKBUF_X2 inst_12438 ( .A(net_12356), .Z(net_12357) );
NAND2_X2 inst_4206 ( .A2(net_9038), .ZN(net_2723), .A1(net_1774) );
CLKBUF_X2 inst_12551 ( .A(net_11409), .Z(net_12470) );
INV_X4 inst_5415 ( .ZN(net_5993), .A(net_1150) );
CLKBUF_X2 inst_15574 ( .A(net_15492), .Z(net_15493) );
INV_X2 inst_6701 ( .ZN(net_8154), .A(net_8153) );
AND4_X4 inst_10340 ( .A1(net_9646), .A2(net_9645), .A3(net_9644), .A4(net_9643), .ZN(net_1790) );
CLKBUF_X2 inst_14798 ( .A(net_13838), .Z(net_14717) );
AND4_X2 inst_10347 ( .ZN(net_3319), .A4(net_2967), .A3(net_2862), .A1(net_1386), .A2(net_1073) );
OR2_X4 inst_812 ( .ZN(net_3115), .A2(net_1366), .A1(net_1127) );
CLKBUF_X2 inst_15535 ( .A(net_15128), .Z(net_15454) );
XNOR2_X2 inst_179 ( .ZN(net_5252), .A(net_4976), .B(net_207) );
CLKBUF_X2 inst_15603 ( .A(net_13826), .Z(net_15522) );
INV_X4 inst_5698 ( .ZN(net_956), .A(net_783) );
OAI21_X2 inst_1730 ( .A(net_8783), .ZN(net_8782), .B1(net_8772), .B2(net_8763) );
NAND2_X2 inst_3799 ( .ZN(net_5973), .A1(net_4310), .A2(net_4184) );
DFF_X2 inst_8101 ( .QN(net_9729), .D(net_5039), .CK(net_12266) );
NAND2_X2 inst_3734 ( .A1(net_10195), .ZN(net_5432), .A2(net_5431) );
OAI211_X2 inst_2191 ( .C1(net_7201), .C2(net_6542), .ZN(net_6518), .B(net_5614), .A(net_3679) );
XNOR2_X2 inst_76 ( .ZN(net_8663), .B(net_8644), .A(net_8623) );
INV_X4 inst_5296 ( .ZN(net_6839), .A(net_1307) );
OAI22_X2 inst_1127 ( .A1(net_7243), .ZN(net_5153), .A2(net_5151), .B2(net_5150), .B1(net_1828) );
INV_X2 inst_6769 ( .ZN(net_6033), .A(net_5860) );
XNOR2_X2 inst_172 ( .ZN(net_5738), .A(net_4792), .B(net_1480) );
CLKBUF_X2 inst_12184 ( .A(net_12102), .Z(net_12103) );
CLKBUF_X2 inst_11228 ( .A(net_11146), .Z(net_11147) );
XNOR2_X2 inst_362 ( .B(net_7495), .ZN(net_2620), .A(net_216) );
NAND2_X2 inst_4366 ( .A2(net_10143), .ZN(net_1761), .A1(net_724) );
XNOR2_X2 inst_277 ( .ZN(net_8762), .B(net_3932), .A(net_3193) );
DFF_X2 inst_7787 ( .Q(net_9821), .D(net_6509), .CK(net_11969) );
XNOR2_X2 inst_83 ( .ZN(net_8622), .A(net_8584), .B(net_8393) );
XNOR2_X2 inst_306 ( .B(net_4281), .ZN(net_3251), .A(net_3009) );
NAND2_X2 inst_4186 ( .ZN(net_3198), .A2(net_1863), .A1(net_1000) );
INV_X4 inst_5566 ( .A(net_9245), .ZN(net_1129) );
DFF_X1 inst_8662 ( .Q(net_9122), .D(net_6910), .CK(net_10588) );
CLKBUF_X2 inst_13499 ( .A(net_13417), .Z(net_13418) );
AOI22_X2 inst_9460 ( .B1(net_10193), .B2(net_4217), .ZN(net_3912), .A2(net_3500), .A1(net_91) );
DFF_X2 inst_7946 ( .QN(net_10467), .D(net_5704), .CK(net_11468) );
NAND2_X2 inst_3386 ( .A2(net_8765), .ZN(net_8764), .A1(net_8762) );
NAND4_X2 inst_3095 ( .ZN(net_4350), .A2(net_3815), .A3(net_3550), .A1(net_3185), .A4(net_2743) );
AOI221_X2 inst_9884 ( .B1(net_9763), .B2(net_9098), .A(net_6940), .C2(net_6939), .ZN(net_6814), .C1(net_6813) );
OAI221_X2 inst_1715 ( .ZN(net_3622), .A(net_3156), .C2(net_2310), .B1(net_2308), .B2(net_1598), .C1(net_897) );
CLKBUF_X2 inst_13673 ( .A(net_13591), .Z(net_13592) );
INV_X4 inst_6396 ( .A(net_9927), .ZN(net_1212) );
HA_X1 inst_7355 ( .A(net_9179), .S(net_2738), .CO(net_2737), .B(net_2195) );
XNOR2_X2 inst_140 ( .ZN(net_7315), .A(net_6926), .B(net_2640) );
XNOR2_X2 inst_267 ( .B(net_4304), .ZN(net_3971), .A(net_3652) );
DFF_X2 inst_7990 ( .QN(net_10417), .D(net_5538), .CK(net_13317) );
NOR2_X2 inst_2824 ( .ZN(net_3035), .A2(net_2546), .A1(net_576) );
INV_X4 inst_5945 ( .ZN(net_981), .A(net_898) );
OR3_X2 inst_716 ( .ZN(net_3636), .A3(net_3198), .A1(net_2936), .A2(net_834) );
NAND2_X2 inst_3594 ( .ZN(net_7272), .A1(net_6882), .A2(net_6558) );
OAI21_X2 inst_1906 ( .B1(net_7229), .B2(net_4862), .ZN(net_4846), .A(net_4518) );
OR2_X4 inst_792 ( .A1(net_10367), .ZN(net_2417), .A2(net_1379) );
DFF_X2 inst_8155 ( .Q(net_10530), .D(net_5072), .CK(net_14886) );
OAI211_X2 inst_2024 ( .C2(net_9564), .ZN(net_8795), .B(net_8792), .C1(net_4982), .A(net_3554) );
NAND4_X2 inst_3124 ( .A1(net_5813), .ZN(net_3138), .A4(net_3137), .A3(net_2201), .A2(net_1775) );
AOI221_X2 inst_9984 ( .C1(net_10183), .B1(net_9742), .B2(net_6442), .C2(net_4217), .ZN(net_4213), .A(net_3645) );
DFF_X2 inst_7993 ( .QN(net_9171), .D(net_5720), .CK(net_11312) );
NOR2_X2 inst_2952 ( .A1(net_10145), .ZN(net_2395), .A2(net_1213) );
CLKBUF_X2 inst_11896 ( .A(net_11814), .Z(net_11815) );
AOI22_X2 inst_9061 ( .B1(net_9663), .A1(net_6828), .A2(net_6684), .B2(net_6683), .ZN(net_6605) );
AND2_X4 inst_10476 ( .A2(net_10258), .A1(net_10257), .ZN(net_2014) );
CLKBUF_X2 inst_14990 ( .A(net_14908), .Z(net_14909) );
OAI211_X2 inst_2216 ( .C1(net_7224), .C2(net_6501), .ZN(net_6489), .B(net_5555), .A(net_3679) );
CLKBUF_X2 inst_11558 ( .A(net_11476), .Z(net_11477) );
XNOR2_X2 inst_174 ( .ZN(net_5645), .B(net_5314), .A(net_5313) );
NOR2_X2 inst_2988 ( .A1(net_10354), .ZN(net_2393), .A2(net_676) );
CLKBUF_X2 inst_15043 ( .A(net_14961), .Z(net_14962) );
DFF_X1 inst_8658 ( .Q(net_9767), .D(net_7125), .CK(net_11620) );
INV_X8 inst_4494 ( .ZN(net_6683), .A(net_5937) );
CLKBUF_X2 inst_12293 ( .A(net_12211), .Z(net_12212) );
CLKBUF_X2 inst_11186 ( .A(net_11104), .Z(net_11105) );
OAI211_X2 inst_2105 ( .C2(net_6778), .ZN(net_6743), .A(net_6371), .B(net_6101), .C1(net_499) );
OAI22_X2 inst_1199 ( .A1(net_7136), .A2(net_5107), .B2(net_5105), .ZN(net_5054), .B1(net_5053) );
XOR2_X2 inst_5 ( .B(net_9529), .Z(net_5986), .A(net_5800) );
OR2_X4 inst_729 ( .A2(net_9503), .ZN(net_7486), .A1(net_3088) );
INV_X4 inst_6567 ( .A(net_9215), .ZN(net_836) );
CLKBUF_X2 inst_11520 ( .A(net_11438), .Z(net_11439) );
INV_X4 inst_6506 ( .ZN(net_4026), .A(net_124) );
OAI211_X2 inst_2157 ( .C2(net_6778), .ZN(net_6691), .A(net_6307), .B(net_6050), .C1(net_5043) );
OAI221_X2 inst_1662 ( .C1(net_7231), .A(net_5637), .C2(net_5520), .ZN(net_5507), .B2(net_4547), .B1(net_2295) );
CLKBUF_X2 inst_10891 ( .A(net_10809), .Z(net_10810) );
INV_X4 inst_4553 ( .ZN(net_8557), .A(net_8537) );
NOR2_X2 inst_2783 ( .ZN(net_3425), .A2(net_3105), .A1(net_520) );
DFF_X2 inst_7508 ( .QN(net_9375), .D(net_7940), .CK(net_14176) );
INV_X4 inst_5804 ( .ZN(net_1002), .A(net_929) );
SDFF_X2 inst_604 ( .Q(net_10518), .D(net_10518), .SE(net_4560), .CK(net_10555), .SI(x5961) );
AOI22_X2 inst_9004 ( .A1(net_9955), .B1(net_9856), .ZN(net_8043), .A2(net_8042), .B2(net_8041) );
CLKBUF_X2 inst_13240 ( .A(net_13158), .Z(net_13159) );
CLKBUF_X2 inst_11251 ( .A(net_11169), .Z(net_11170) );
CLKBUF_X2 inst_13872 ( .A(net_13790), .Z(net_13791) );
DFF_X2 inst_7539 ( .D(net_7755), .CK(net_15319), .Q(x589) );
INV_X2 inst_7085 ( .A(net_2621), .ZN(net_1149) );
OAI22_X2 inst_1285 ( .A2(net_4092), .ZN(net_4086), .A1(net_4085), .B1(net_3068), .B2(net_1836) );
XNOR2_X2 inst_380 ( .B(net_9303), .ZN(net_2993), .A(net_2448) );
NAND2_X2 inst_4057 ( .A2(net_8859), .ZN(net_4435), .A1(net_2767) );
OAI22_X2 inst_1179 ( .A1(net_7224), .A2(net_5134), .B2(net_5133), .ZN(net_5080), .B1(net_3163) );
XNOR2_X2 inst_292 ( .B(net_9306), .ZN(net_3725), .A(net_2867) );
NAND2_X2 inst_3650 ( .A2(net_9351), .ZN(net_7783), .A1(net_5393) );
CLKBUF_X2 inst_11661 ( .A(net_10804), .Z(net_11580) );
CLKBUF_X2 inst_14711 ( .A(net_14629), .Z(net_14630) );
CLKBUF_X2 inst_13508 ( .A(net_13426), .Z(net_13427) );
OAI21_X2 inst_2012 ( .B2(net_3899), .A(net_3894), .ZN(net_1710), .B1(net_1708) );
CLKBUF_X2 inst_11350 ( .A(net_11268), .Z(net_11269) );
CLKBUF_X2 inst_10900 ( .A(net_10721), .Z(net_10819) );
DFF_X2 inst_7423 ( .QN(net_9394), .D(net_8336), .CK(net_13946) );
INV_X4 inst_4970 ( .A(net_7437), .ZN(net_2941) );
CLKBUF_X2 inst_12583 ( .A(net_12501), .Z(net_12502) );
OR3_X2 inst_706 ( .ZN(net_7923), .A2(net_7813), .A1(net_7346), .A3(net_5890) );
CLKBUF_X2 inst_14692 ( .A(net_13931), .Z(net_14611) );
CLKBUF_X2 inst_10874 ( .A(net_10792), .Z(net_10793) );
INV_X4 inst_6605 ( .A(net_9637), .ZN(net_3385) );
AOI221_X2 inst_9834 ( .A(net_6889), .B2(net_6888), .C2(net_6887), .ZN(net_6884), .B1(net_5856), .C1(x5289) );
OR2_X4 inst_839 ( .A2(net_10147), .A1(net_10146), .ZN(net_2105) );
CLKBUF_X2 inst_13366 ( .A(net_11212), .Z(net_13285) );
DFF_X2 inst_7985 ( .QN(net_10411), .D(net_5595), .CK(net_14589) );
INV_X4 inst_4734 ( .A(net_10058), .ZN(net_8511) );
XNOR2_X2 inst_240 ( .ZN(net_4256), .A(net_4255), .B(net_2079) );
CLKBUF_X2 inst_15033 ( .A(net_14951), .Z(net_14952) );
CLKBUF_X2 inst_13055 ( .A(net_12973), .Z(net_12974) );
INV_X4 inst_5455 ( .A(net_4331), .ZN(net_1557) );
DFF_X2 inst_7501 ( .Q(net_9274), .D(net_8035), .CK(net_11477) );
NAND2_X2 inst_3966 ( .ZN(net_4319), .A2(net_4070), .A1(net_761) );
XNOR2_X2 inst_110 ( .B(net_9601), .A(net_8956), .ZN(net_8096) );
CLKBUF_X2 inst_13681 ( .A(net_13599), .Z(net_13600) );
OAI211_X2 inst_2047 ( .B(net_9288), .A(net_8057), .ZN(net_7841), .C1(net_7597), .C2(net_6320) );
INV_X4 inst_4545 ( .A(net_9578), .ZN(net_8600) );
NAND2_X2 inst_3825 ( .ZN(net_9078), .A2(net_4179), .A1(net_4032) );
INV_X4 inst_6634 ( .A(net_9042), .ZN(net_9041) );
XNOR2_X2 inst_99 ( .B(net_9434), .ZN(net_8410), .A(net_6585) );
AOI21_X4 inst_9997 ( .ZN(net_8720), .B1(net_8708), .A(net_8552), .B2(net_8538) );
CLKBUF_X2 inst_13210 ( .A(net_13128), .Z(net_13129) );
DFF_X2 inst_7876 ( .QN(net_10156), .D(net_6006), .CK(net_13483) );
CLKBUF_X2 inst_13152 ( .A(net_13070), .Z(net_13071) );
CLKBUF_X2 inst_10842 ( .A(net_10760), .Z(net_10761) );
CLKBUF_X2 inst_11927 ( .A(net_11729), .Z(net_11846) );
CLKBUF_X2 inst_11050 ( .A(net_10968), .Z(net_10969) );
NAND2_X2 inst_4384 ( .A2(net_10246), .ZN(net_1337), .A1(net_649) );
DFF_X2 inst_7846 ( .Q(net_9912), .D(net_6495), .CK(net_15661) );
OAI211_X2 inst_2059 ( .A(net_7783), .C2(net_7782), .ZN(net_7774), .B(net_7678), .C1(net_2475) );
CLKBUF_X2 inst_13851 ( .A(net_13769), .Z(net_13770) );
INV_X2 inst_7023 ( .ZN(net_1518), .A(net_908) );
AOI22_X2 inst_9473 ( .B1(net_10394), .A1(net_9878), .B2(net_4062), .ZN(net_3850), .A2(net_2973) );
AOI22_X2 inst_9445 ( .A1(net_10525), .B1(net_9798), .A2(net_4056), .ZN(net_4054), .B2(net_2556) );
NOR2_X2 inst_2949 ( .A2(net_4157), .ZN(net_1627), .A1(net_1244) );
NOR3_X2 inst_2414 ( .ZN(net_5380), .A3(net_4670), .A1(net_3216), .A2(net_2433) );
AOI22_X2 inst_9656 ( .ZN(net_2700), .A1(net_2207), .A2(net_2206), .B1(net_2205), .B2(net_1645) );
XNOR2_X2 inst_311 ( .ZN(net_3225), .B(net_2525), .A(net_2473) );
CLKBUF_X2 inst_12461 ( .A(net_12379), .Z(net_12380) );
AOI221_X2 inst_9914 ( .B1(net_9947), .C1(net_9749), .ZN(net_6444), .B2(net_6443), .C2(net_6442), .A(net_5722) );
CLKBUF_X2 inst_13205 ( .A(net_13123), .Z(net_13124) );
AND2_X4 inst_10429 ( .A1(net_4233), .ZN(net_3928), .A2(net_3452) );
CLKBUF_X2 inst_13180 ( .A(net_13098), .Z(net_13099) );
DFF_X2 inst_8139 ( .Q(net_9948), .D(net_5118), .CK(net_14729) );
OAI211_X2 inst_2203 ( .C1(net_7241), .C2(net_6542), .ZN(net_6504), .B(net_5601), .A(net_3527) );
CLKBUF_X2 inst_11132 ( .A(net_11050), .Z(net_11051) );
DFF_X2 inst_7901 ( .QN(net_10368), .D(net_5958), .CK(net_13656) );
CLKBUF_X2 inst_15189 ( .A(net_15107), .Z(net_15108) );
AND2_X2 inst_10495 ( .A2(net_10240), .ZN(net_6668), .A1(net_1477) );
INV_X2 inst_6981 ( .A(net_2078), .ZN(net_1672) );
CLKBUF_X2 inst_14413 ( .A(net_13818), .Z(net_14332) );
CLKBUF_X2 inst_11695 ( .A(net_11449), .Z(net_11614) );
CLKBUF_X2 inst_14648 ( .A(net_14566), .Z(net_14567) );
INV_X2 inst_7316 ( .A(net_9100), .ZN(net_9099) );
CLKBUF_X2 inst_15002 ( .A(net_14920), .Z(net_14921) );
OAI21_X2 inst_1930 ( .ZN(net_4410), .B1(net_4409), .B2(net_4408), .A(net_3135) );
CLKBUF_X2 inst_14440 ( .A(net_14358), .Z(net_14359) );
OR2_X2 inst_889 ( .A1(net_10377), .ZN(net_6629), .A2(net_5970) );
SDFF_X2 inst_577 ( .D(net_9132), .SE(net_933), .CK(net_10947), .SI(x2477), .Q(x1240) );
INV_X4 inst_5536 ( .A(net_9354), .ZN(net_5405) );
CLKBUF_X2 inst_12305 ( .A(net_12164), .Z(net_12224) );
CLKBUF_X2 inst_13497 ( .A(net_13415), .Z(net_13416) );
DFF_X1 inst_8533 ( .Q(net_9965), .D(net_7335), .CK(net_14268) );
CLKBUF_X2 inst_15269 ( .A(net_15187), .Z(net_15188) );
INV_X4 inst_4975 ( .ZN(net_2311), .A(net_2310) );
INV_X2 inst_6760 ( .ZN(net_6229), .A(net_6228) );
CLKBUF_X2 inst_12457 ( .A(net_12024), .Z(net_12376) );
INV_X4 inst_5188 ( .A(net_1554), .ZN(net_1548) );
NOR3_X2 inst_2379 ( .ZN(net_7898), .A3(net_7773), .A1(net_3984), .A2(x3390) );
NAND2_X2 inst_3938 ( .A1(net_9912), .A2(net_4969), .ZN(net_3552) );
AND3_X4 inst_10358 ( .ZN(net_5759), .A2(net_4788), .A3(net_4629), .A1(net_4462) );
DFF_X1 inst_8774 ( .Q(net_10484), .D(net_4957), .CK(net_11411) );
CLKBUF_X2 inst_11754 ( .A(net_11672), .Z(net_11673) );
CLKBUF_X2 inst_11244 ( .A(net_11162), .Z(net_11163) );
NOR2_X2 inst_2865 ( .A2(net_2425), .ZN(net_2046), .A1(net_2045) );
CLKBUF_X2 inst_15047 ( .A(net_14965), .Z(net_14966) );
CLKBUF_X2 inst_14933 ( .A(net_14851), .Z(net_14852) );
AND3_X2 inst_10382 ( .ZN(net_880), .A1(net_147), .A2(net_146), .A3(net_145) );
INV_X4 inst_5986 ( .A(net_9932), .ZN(net_1347) );
INV_X4 inst_4916 ( .ZN(net_2974), .A(net_2769) );
DFF_X2 inst_8149 ( .QN(net_9751), .D(net_5082), .CK(net_14535) );
INV_X4 inst_4891 ( .ZN(net_3285), .A(net_2925) );
NAND2_X2 inst_3571 ( .ZN(net_7656), .A1(net_7655), .A2(net_7596) );
CLKBUF_X2 inst_15757 ( .A(net_15675), .Z(net_15676) );
INV_X4 inst_6132 ( .A(net_9650), .ZN(net_484) );
OAI22_X2 inst_1190 ( .A1(net_7127), .A2(net_5134), .B2(net_5133), .ZN(net_5064), .B1(net_1313) );
CLKBUF_X2 inst_14520 ( .A(net_12935), .Z(net_14439) );
XNOR2_X2 inst_444 ( .B(net_9304), .ZN(net_862), .A(net_227) );
DFF_X1 inst_8865 ( .D(net_10303), .QN(net_10243), .CK(net_11128) );
DFF_X2 inst_7460 ( .QN(net_8833), .D(net_8125), .CK(net_14764) );
CLKBUF_X2 inst_11092 ( .A(net_11010), .Z(net_11011) );
CLKBUF_X2 inst_11016 ( .A(net_10860), .Z(net_10935) );
DFF_X2 inst_7489 ( .D(net_7984), .Q(net_206), .CK(net_14762) );
DFF_X2 inst_8246 ( .Q(net_10084), .D(net_4851), .CK(net_10723) );
INV_X4 inst_6264 ( .A(net_9994), .ZN(net_449) );
CLKBUF_X2 inst_12816 ( .A(net_12734), .Z(net_12735) );
AOI22_X2 inst_9064 ( .B1(net_9684), .A2(net_6684), .B2(net_6683), .ZN(net_6602), .A1(net_253) );
AOI21_X2 inst_10033 ( .B1(net_10175), .ZN(net_7867), .A(net_6679), .B2(net_263) );
CLKBUF_X2 inst_14196 ( .A(net_13313), .Z(net_14115) );
CLKBUF_X2 inst_14556 ( .A(net_11112), .Z(net_14475) );
DFF_X1 inst_8705 ( .Q(net_9139), .D(net_6780), .CK(net_11013) );
CLKBUF_X2 inst_11720 ( .A(net_11638), .Z(net_11639) );
INV_X2 inst_7040 ( .ZN(net_1377), .A(net_1376) );
INV_X4 inst_4905 ( .A(net_9421), .ZN(net_8082) );
XNOR2_X2 inst_63 ( .ZN(net_8730), .A(net_8709), .B(net_8139) );
INV_X4 inst_5833 ( .ZN(net_1225), .A(net_1213) );
CLKBUF_X2 inst_12047 ( .A(net_11965), .Z(net_11966) );
XNOR2_X2 inst_119 ( .B(net_9424), .ZN(net_7670), .A(net_6287) );
NAND3_X2 inst_3181 ( .ZN(net_8112), .A1(net_8052), .A3(net_7957), .A2(net_3729) );
OR2_X2 inst_939 ( .A2(net_2396), .ZN(net_1813), .A1(net_1812) );
DFF_X2 inst_7968 ( .QN(net_10319), .D(net_5585), .CK(net_14791) );
AOI222_X1 inst_9722 ( .C1(net_10496), .B1(net_10391), .A1(net_9921), .C2(net_6415), .A2(net_4969), .B2(net_4062), .ZN(net_4059) );
CLKBUF_X2 inst_10770 ( .A(net_10688), .Z(net_10689) );
INV_X4 inst_5469 ( .ZN(net_6056), .A(net_1020) );
OAI22_X2 inst_1233 ( .B1(net_7186), .A2(net_4890), .B2(net_4889), .ZN(net_4884), .A1(net_506) );
AND2_X4 inst_10445 ( .ZN(net_1738), .A2(net_1570), .A1(net_222) );
DFF_X2 inst_8205 ( .Q(net_10181), .D(net_4829), .CK(net_12969) );
NOR2_X2 inst_2924 ( .A1(net_10247), .ZN(net_1820), .A2(net_824) );
CLKBUF_X2 inst_15389 ( .A(net_15307), .Z(net_15308) );
CLKBUF_X2 inst_11117 ( .A(net_10630), .Z(net_11036) );
OAI22_X2 inst_1019 ( .ZN(net_8037), .A2(net_8036), .B2(net_8018), .A1(net_4541), .B1(net_365) );
CLKBUF_X2 inst_13490 ( .A(net_12750), .Z(net_13409) );
OAI21_X2 inst_2006 ( .B1(net_5462), .ZN(net_2141), .A(net_1464), .B2(net_1197) );
AND4_X4 inst_10337 ( .ZN(net_3215), .A3(net_2432), .A1(net_2186), .A4(net_2058), .A2(net_1009) );
CLKBUF_X2 inst_15672 ( .A(net_11589), .Z(net_15591) );
OAI21_X2 inst_1827 ( .B2(net_9170), .ZN(net_6566), .A(net_4717), .B1(net_4041) );
CLKBUF_X2 inst_10830 ( .A(net_10748), .Z(net_10749) );
OR2_X4 inst_742 ( .A1(net_9162), .ZN(net_5940), .A2(net_5939) );
CLKBUF_X2 inst_13372 ( .A(net_12574), .Z(net_13291) );
NOR2_X2 inst_2619 ( .ZN(net_7154), .A2(net_6202), .A1(net_6165) );
CLKBUF_X2 inst_15625 ( .A(net_15543), .Z(net_15544) );
INV_X2 inst_7057 ( .ZN(net_1290), .A(net_1289) );
NAND2_X2 inst_3465 ( .A1(net_9500), .A2(net_8473), .ZN(net_8458) );
OAI211_X2 inst_2033 ( .C2(net_8102), .ZN(net_8101), .A(net_8000), .B(net_3507), .C1(net_2140) );
CLKBUF_X2 inst_14131 ( .A(net_14049), .Z(net_14050) );
DFF_X2 inst_7850 ( .Q(net_10021), .D(net_6463), .CK(net_12037) );
MUX2_X1 inst_4481 ( .S(net_9201), .A(net_9064), .Z(net_8853), .B(net_6639) );
DFF_X2 inst_7675 ( .D(net_6721), .QN(net_163), .CK(net_11995) );
NOR2_X2 inst_2559 ( .A2(net_7805), .ZN(net_7760), .A1(net_2850) );
CLKBUF_X2 inst_13898 ( .A(net_13816), .Z(net_13817) );
CLKBUF_X2 inst_13545 ( .A(net_13463), .Z(net_13464) );
CLKBUF_X2 inst_13336 ( .A(net_12018), .Z(net_13255) );
HA_X1 inst_7345 ( .S(net_5237), .CO(net_5236), .B(net_4433), .A(net_1301) );
CLKBUF_X2 inst_12039 ( .A(net_10698), .Z(net_11958) );
INV_X4 inst_5289 ( .A(net_3171), .ZN(net_2488) );
AOI21_X2 inst_10201 ( .ZN(net_2819), .B1(net_2818), .A(net_2170), .B2(net_1525) );
AOI22_X2 inst_9121 ( .A1(net_9706), .A2(net_6404), .ZN(net_6368), .B2(net_5263), .B1(net_146) );
DFF_X2 inst_8386 ( .Q(net_10303), .D(net_904), .CK(net_11422) );
INV_X2 inst_6997 ( .ZN(net_1630), .A(net_1571) );
OAI21_X2 inst_1955 ( .ZN(net_4258), .A(net_3326), .B2(net_3240), .B1(net_3117) );
DFF_X1 inst_8837 ( .Q(net_9859), .D(net_2158), .CK(net_10759) );
INV_X4 inst_6125 ( .ZN(net_6379), .A(net_129) );
CLKBUF_X2 inst_12657 ( .A(net_12575), .Z(net_12576) );
NAND2_X2 inst_3618 ( .ZN(net_7112), .A1(net_6871), .A2(net_6685) );
OAI22_X2 inst_1269 ( .B1(net_7186), .A2(net_4826), .B2(net_4825), .ZN(net_4804), .A1(net_455) );
CLKBUF_X2 inst_13575 ( .A(net_13493), .Z(net_13494) );
CLKBUF_X2 inst_14768 ( .A(net_14686), .Z(net_14687) );
CLKBUF_X2 inst_14807 ( .A(net_13392), .Z(net_14726) );
CLKBUF_X2 inst_14430 ( .A(net_14348), .Z(net_14349) );
CLKBUF_X2 inst_14945 ( .A(net_14863), .Z(net_14864) );
AOI22_X2 inst_9181 ( .A1(net_9860), .B1(net_9761), .B2(net_8041), .A2(net_6141), .ZN(net_6135) );
INV_X2 inst_7202 ( .A(net_10244), .ZN(net_904) );
AOI221_X2 inst_9781 ( .C1(net_9349), .B1(net_9158), .A(net_7157), .B2(net_7155), .C2(net_7154), .ZN(net_7153) );
NAND3_X2 inst_3241 ( .A1(net_7142), .A3(net_4719), .ZN(net_4712), .A2(net_3056) );
NOR2_X2 inst_2704 ( .ZN(net_4746), .A2(net_4325), .A1(net_4324) );
CLKBUF_X2 inst_11842 ( .A(net_11760), .Z(net_11761) );
OAI221_X2 inst_1620 ( .B1(net_10317), .C1(net_7139), .A(net_5637), .B2(net_5591), .ZN(net_5587), .C2(net_4902) );
INV_X4 inst_4958 ( .A(net_4713), .ZN(net_2542) );
CLKBUF_X2 inst_13344 ( .A(net_11280), .Z(net_13263) );
DFF_X2 inst_8349 ( .QN(net_10479), .D(net_2779), .CK(net_11429) );
CLKBUF_X2 inst_11461 ( .A(net_11379), .Z(net_11380) );
AND2_X2 inst_10572 ( .ZN(net_3452), .A2(net_3182), .A1(net_955) );
INV_X4 inst_5924 ( .ZN(net_2202), .A(net_581) );
XNOR2_X2 inst_347 ( .ZN(net_2859), .A(net_1831), .B(net_1578) );
CLKBUF_X2 inst_14551 ( .A(net_14469), .Z(net_14470) );
INV_X4 inst_5438 ( .A(net_4986), .ZN(net_1582) );
CLKBUF_X2 inst_11600 ( .A(net_11188), .Z(net_11519) );
CLKBUF_X2 inst_13327 ( .A(net_13245), .Z(net_13246) );
OR2_X4 inst_755 ( .ZN(net_4401), .A2(net_4400), .A1(net_1668) );
AOI22_X2 inst_9508 ( .B1(net_9891), .A1(net_9855), .A2(net_6413), .ZN(net_3815), .B2(net_2973) );
OAI21_X4 inst_1724 ( .ZN(net_8950), .B2(net_8505), .A(net_8495), .B1(net_8424) );
DFF_X2 inst_7918 ( .QN(net_9552), .D(net_5804), .CK(net_13768) );
AOI222_X1 inst_9701 ( .B1(net_9510), .A2(net_8286), .B2(net_8285), .C2(net_8284), .ZN(net_8277), .C1(net_8215), .A1(x1459) );
INV_X4 inst_5855 ( .ZN(net_932), .A(net_642) );
CLKBUF_X2 inst_13149 ( .A(net_13067), .Z(net_13068) );
INV_X8 inst_4505 ( .ZN(net_6420), .A(net_5295) );
NOR2_X2 inst_2610 ( .ZN(net_6246), .A1(net_5764), .A2(net_4161) );
DFF_X1 inst_8819 ( .Q(net_10059), .D(net_3260), .CK(net_11107) );
INV_X4 inst_5473 ( .A(net_4160), .ZN(net_1165) );
OAI22_X2 inst_1043 ( .A1(net_9075), .A2(net_8921), .B1(net_8920), .ZN(net_7921), .B2(net_2826) );
CLKBUF_X2 inst_12327 ( .A(net_12038), .Z(net_12246) );
NAND2_X2 inst_4030 ( .ZN(net_3471), .A2(net_3003), .A1(net_2036) );
AOI22_X2 inst_9234 ( .A1(net_9898), .B1(net_9799), .A2(net_8042), .B2(net_6129), .ZN(net_6077) );
INV_X2 inst_7230 ( .A(net_9325), .ZN(net_393) );
CLKBUF_X2 inst_15014 ( .A(net_14932), .Z(net_14933) );
INV_X4 inst_4817 ( .ZN(net_4027), .A(net_3059) );
MUX2_X1 inst_4456 ( .S(net_6041), .A(net_290), .B(x5548), .Z(x208) );
INV_X4 inst_4926 ( .ZN(net_4964), .A(net_2229) );
AOI221_X2 inst_9769 ( .B2(net_10380), .ZN(net_7545), .C2(net_7476), .A(net_7289), .C1(net_6907), .B1(net_2163) );
INV_X2 inst_6846 ( .A(net_10479), .ZN(net_3461) );
OAI21_X2 inst_1792 ( .B2(net_10242), .A(net_10241), .ZN(net_7482), .B1(net_7481) );
NAND2_X1 inst_4426 ( .ZN(net_2614), .A1(net_2613), .A2(net_2612) );
CLKBUF_X2 inst_13840 ( .A(net_13758), .Z(net_13759) );
INV_X4 inst_6017 ( .A(net_10330), .ZN(net_1361) );
INV_X4 inst_4571 ( .ZN(net_8241), .A(net_8129) );
AOI21_X2 inst_10231 ( .B2(net_10327), .ZN(net_2312), .A(net_2006), .B1(net_2005) );
INV_X4 inst_5111 ( .ZN(net_3487), .A(net_1652) );
NAND2_X2 inst_3928 ( .A2(net_4319), .ZN(net_3878), .A1(net_2887) );
NAND2_X4 inst_3353 ( .ZN(net_8420), .A2(net_8385), .A1(net_8382) );
NAND2_X2 inst_3634 ( .A1(net_10296), .ZN(net_6980), .A2(net_6972) );
CLKBUF_X2 inst_12877 ( .A(net_12795), .Z(net_12796) );
CLKBUF_X2 inst_12212 ( .A(net_11051), .Z(net_12131) );
CLKBUF_X2 inst_11849 ( .A(net_11524), .Z(net_11768) );
NAND2_X2 inst_4017 ( .A2(net_7095), .ZN(net_3514), .A1(net_1774) );
INV_X2 inst_7121 ( .A(net_1380), .ZN(net_1178) );
INV_X4 inst_4598 ( .ZN(net_8783), .A(net_8691) );
INV_X4 inst_4681 ( .ZN(net_5001), .A(net_4743) );
INV_X4 inst_5135 ( .A(net_2693), .ZN(net_1936) );
CLKBUF_X2 inst_12879 ( .A(net_11002), .Z(net_12798) );
CLKBUF_X2 inst_13050 ( .A(net_11155), .Z(net_12969) );
AOI221_X2 inst_9772 ( .B2(net_10485), .ZN(net_7494), .C2(net_7407), .A(net_7075), .C1(net_6654), .B1(net_2205) );
CLKBUF_X2 inst_11204 ( .A(net_11122), .Z(net_11123) );
INV_X4 inst_5760 ( .ZN(net_801), .A(net_727) );
DFF_X2 inst_7556 ( .QN(net_9320), .D(net_7689), .CK(net_13035) );
CLKBUF_X2 inst_11513 ( .A(net_11431), .Z(net_11432) );
INV_X2 inst_7037 ( .A(net_3748), .ZN(net_1395) );
INV_X2 inst_7294 ( .A(net_9045), .ZN(net_9044) );
INV_X4 inst_5095 ( .ZN(net_2490), .A(net_1624) );
CLKBUF_X2 inst_14591 ( .A(net_13051), .Z(net_14510) );
XNOR2_X2 inst_426 ( .B(net_9357), .ZN(net_1331), .A(net_502) );
NAND4_X2 inst_3145 ( .ZN(net_2162), .A4(net_1251), .A2(net_1052), .A3(net_735), .A1(net_630) );
INV_X4 inst_5144 ( .ZN(net_6305), .A(net_1590) );
SDFF_X2 inst_648 ( .SI(net_9489), .Q(net_9489), .SE(net_3073), .CK(net_12432), .D(x2098) );
AND2_X2 inst_10600 ( .A2(net_4114), .ZN(net_2079), .A1(net_2078) );
INV_X4 inst_6035 ( .A(net_10531), .ZN(net_561) );
DFF_X2 inst_7857 ( .Q(net_9182), .D(net_6272), .CK(net_13569) );
CLKBUF_X2 inst_13718 ( .A(net_13636), .Z(net_13637) );
XNOR2_X2 inst_270 ( .ZN(net_3957), .A(net_3237), .B(net_2894) );
OAI21_X2 inst_1901 ( .B1(net_7231), .B2(net_4862), .ZN(net_4851), .A(net_4523) );
CLKBUF_X2 inst_13856 ( .A(net_13774), .Z(net_13775) );
NAND2_X2 inst_4302 ( .A2(net_9040), .ZN(net_7442), .A1(net_6949) );
CLKBUF_X2 inst_11654 ( .A(net_11414), .Z(net_11573) );
CLKBUF_X2 inst_11068 ( .A(net_10776), .Z(net_10987) );
DFF_X2 inst_8092 ( .QN(net_9932), .D(net_5055), .CK(net_14352) );
INV_X4 inst_6560 ( .A(net_10430), .ZN(net_701) );
DFF_X2 inst_7725 ( .Q(net_9902), .D(net_6277), .CK(net_15062) );
NAND2_X2 inst_4104 ( .ZN(net_2383), .A1(net_2145), .A2(net_1659) );
INV_X4 inst_6341 ( .A(net_9969), .ZN(net_411) );
CLKBUF_X2 inst_11826 ( .A(net_11744), .Z(net_11745) );
DFF_X1 inst_8608 ( .Q(net_9860), .D(net_7240), .CK(net_12094) );
NOR2_X2 inst_2552 ( .A2(net_9272), .ZN(net_8029), .A1(net_6165) );
CLKBUF_X2 inst_11809 ( .A(net_11089), .Z(net_11728) );
SDFF_X2 inst_631 ( .Q(net_9454), .D(net_9454), .SE(net_3293), .CK(net_11898), .SI(x2278) );
CLKBUF_X2 inst_11163 ( .A(net_10553), .Z(net_11082) );
DFF_X1 inst_8544 ( .Q(net_9978), .D(net_7367), .CK(net_14783) );
AOI22_X2 inst_9247 ( .A1(net_9953), .B1(net_9854), .A2(net_6141), .B2(net_6133), .ZN(net_6064) );
INV_X4 inst_6427 ( .A(net_9372), .ZN(net_7632) );
CLKBUF_X2 inst_15070 ( .A(net_14988), .Z(net_14989) );
NAND2_X2 inst_3674 ( .A1(net_9073), .ZN(net_6903), .A2(net_6235) );
AOI221_X2 inst_9904 ( .B1(net_9889), .B2(net_9101), .A(net_6945), .C2(net_6944), .ZN(net_6790), .C1(net_260) );
CLKBUF_X2 inst_12835 ( .A(net_11954), .Z(net_12754) );
CLKBUF_X2 inst_11346 ( .A(net_11264), .Z(net_11265) );
CLKBUF_X2 inst_13505 ( .A(net_13423), .Z(net_13424) );
CLKBUF_X2 inst_15182 ( .A(net_15100), .Z(net_15101) );
CLKBUF_X2 inst_13789 ( .A(net_13707), .Z(net_13708) );
CLKBUF_X2 inst_12558 ( .A(net_12476), .Z(net_12477) );
DFF_X2 inst_8136 ( .Q(net_9924), .D(net_5140), .CK(net_12124) );
CLKBUF_X2 inst_15645 ( .A(net_15563), .Z(net_15564) );
NAND2_X2 inst_3995 ( .ZN(net_3909), .A2(net_3390), .A1(net_1522) );
NAND2_X2 inst_4211 ( .ZN(net_2117), .A2(net_1745), .A1(net_896) );
INV_X4 inst_5074 ( .A(net_3177), .ZN(net_1831) );
OAI21_X2 inst_1745 ( .B1(net_8691), .ZN(net_8683), .B2(net_8663), .A(net_7851) );
NAND2_X2 inst_3831 ( .A1(net_8863), .ZN(net_4407), .A2(net_4406) );
OAI211_X2 inst_2079 ( .C2(net_6778), .ZN(net_6769), .A(net_6396), .B(net_6130), .C1(net_533) );
XNOR2_X2 inst_102 ( .B(net_9430), .ZN(net_8321), .A(net_6182) );
AND2_X2 inst_10534 ( .ZN(net_4171), .A1(net_3853), .A2(net_3852) );
CLKBUF_X2 inst_15506 ( .A(net_15424), .Z(net_15425) );
CLKBUF_X2 inst_14749 ( .A(net_14667), .Z(net_14668) );
NOR2_X2 inst_2527 ( .A2(net_8930), .ZN(net_8330), .A1(net_8164) );
INV_X2 inst_6819 ( .A(net_4968), .ZN(net_4673) );
NAND3_X2 inst_3277 ( .ZN(net_4370), .A1(net_3630), .A3(net_3383), .A2(net_2763) );
CLKBUF_X2 inst_14883 ( .A(net_14801), .Z(net_14802) );
CLKBUF_X2 inst_12042 ( .A(net_11960), .Z(net_11961) );
AOI22_X2 inst_9299 ( .B1(net_10017), .A2(net_5743), .B2(net_5742), .ZN(net_5679), .A1(net_257) );
CLKBUF_X2 inst_14053 ( .A(net_13971), .Z(net_13972) );
INV_X4 inst_5352 ( .ZN(net_1561), .A(net_692) );
NOR2_X2 inst_2786 ( .A2(net_7644), .ZN(net_7424), .A1(net_3088) );
CLKBUF_X2 inst_11045 ( .A(net_10963), .Z(net_10964) );
AOI21_X2 inst_10043 ( .ZN(net_7471), .A(net_7470), .B2(net_7385), .B1(net_1895) );
OAI22_X2 inst_1224 ( .A1(net_7108), .A2(net_5151), .B2(net_5150), .ZN(net_5023), .B1(net_2561) );
NAND2_X2 inst_3905 ( .ZN(net_3900), .A1(net_3899), .A2(net_3059) );
DFF_X2 inst_7666 ( .D(net_6730), .QN(net_155), .CK(net_12809) );
INV_X4 inst_6554 ( .A(net_10039), .ZN(net_5090) );
INV_X4 inst_5615 ( .A(net_10350), .ZN(net_1120) );
CLKBUF_X2 inst_11797 ( .A(net_11715), .Z(net_11716) );
OAI22_X2 inst_1170 ( .A1(net_7186), .A2(net_5107), .B2(net_5105), .ZN(net_5093), .B1(net_5092) );
CLKBUF_X2 inst_14729 ( .A(net_14647), .Z(net_14648) );
CLKBUF_X2 inst_14246 ( .A(net_12386), .Z(net_14165) );
CLKBUF_X2 inst_15219 ( .A(net_15137), .Z(net_15138) );
CLKBUF_X2 inst_12081 ( .A(net_11999), .Z(net_12000) );
NOR2_X2 inst_2596 ( .A2(net_7461), .A1(net_7276), .ZN(net_6896) );
CLKBUF_X2 inst_11659 ( .A(net_11577), .Z(net_11578) );
INV_X4 inst_6599 ( .A(net_9223), .ZN(net_317) );
INV_X4 inst_6242 ( .A(net_10110), .ZN(net_5851) );
DFF_X1 inst_8752 ( .Q(net_9127), .D(net_5282), .CK(net_10970) );
DFF_X1 inst_8579 ( .Q(net_9677), .D(net_7272), .CK(net_13887) );
NOR2_X2 inst_3022 ( .ZN(net_621), .A2(net_274), .A1(net_273) );
CLKBUF_X2 inst_12133 ( .A(net_11618), .Z(net_12052) );
SDFF_X2 inst_680 ( .D(net_9584), .SI(net_2183), .SE(net_758), .Q(net_258), .CK(net_11566) );
INV_X4 inst_6575 ( .ZN(net_7241), .A(x5850) );
OR2_X4 inst_785 ( .A2(net_2304), .ZN(net_2179), .A1(net_2178) );
NOR3_X4 inst_2362 ( .ZN(net_8991), .A2(net_5433), .A1(net_5019), .A3(net_4729) );
AND4_X4 inst_10323 ( .ZN(net_3721), .A2(net_3720), .A3(net_3719), .A4(net_3718), .A1(net_3128) );
NAND3_X2 inst_3299 ( .A3(net_3261), .A1(net_3085), .ZN(net_2550), .A2(net_1912) );
NOR2_X2 inst_2856 ( .A1(net_9621), .ZN(net_2108), .A2(net_1391) );
AOI22_X2 inst_9280 ( .B1(net_9899), .A1(net_5759), .B2(net_5758), .ZN(net_5740), .A2(net_238) );
AND2_X4 inst_10417 ( .A2(net_4408), .ZN(net_4271), .A1(net_2682) );
DFF_X2 inst_7820 ( .QN(net_9177), .D(net_6300), .CK(net_13576) );
INV_X2 inst_7065 ( .A(net_2564), .ZN(net_1260) );
CLKBUF_X2 inst_15717 ( .A(net_15635), .Z(net_15636) );
DFF_X2 inst_7643 ( .D(net_6727), .QN(net_158), .CK(net_13444) );
DFF_X2 inst_7945 ( .QN(net_10336), .D(net_5578), .CK(net_13259) );
DFF_X2 inst_7551 ( .QN(net_9536), .D(net_7717), .CK(net_12747) );
SDFF_X2 inst_527 ( .SI(net_9336), .Q(net_9281), .D(net_9281), .SE(net_7588), .CK(net_14674) );
CLKBUF_X2 inst_12697 ( .A(net_10621), .Z(net_12616) );
NAND2_X2 inst_3567 ( .A2(net_7748), .ZN(net_7680), .A1(net_7679) );
XNOR2_X2 inst_226 ( .ZN(net_4416), .B(net_4172), .A(net_4171) );
OAI22_X2 inst_1180 ( .A1(net_7198), .A2(net_5134), .B2(net_5133), .ZN(net_5079), .B1(net_1286) );
INV_X4 inst_5509 ( .A(net_10124), .ZN(net_976) );
XNOR2_X2 inst_414 ( .B(net_10041), .ZN(net_1414), .A(net_1413) );
CLKBUF_X2 inst_13861 ( .A(net_13779), .Z(net_13780) );
DFF_X2 inst_8223 ( .D(net_4867), .Q(net_228), .CK(net_10833) );
CLKBUF_X2 inst_11232 ( .A(net_11150), .Z(net_11151) );
SDFF_X2 inst_531 ( .SI(net_9341), .Q(net_9286), .D(net_9286), .SE(net_7588), .CK(net_14663) );
CLKBUF_X2 inst_11688 ( .A(net_11606), .Z(net_11607) );
XNOR2_X2 inst_212 ( .ZN(net_4934), .A(net_4393), .B(net_2339) );
NOR2_X2 inst_2732 ( .A2(net_10175), .ZN(net_4220), .A1(net_3872) );
AOI22_X2 inst_9315 ( .B1(net_9720), .A2(net_5755), .B2(net_5754), .ZN(net_5662), .A1(net_257) );
INV_X4 inst_6321 ( .A(net_9533), .ZN(net_7146) );
OAI21_X2 inst_1952 ( .ZN(net_3922), .A(net_3920), .B2(net_3919), .B1(net_3360) );
CLKBUF_X2 inst_15293 ( .A(net_10954), .Z(net_15212) );
AOI22_X2 inst_9323 ( .B1(net_9698), .A2(net_5755), .B2(net_5754), .ZN(net_5653), .A1(net_235) );
AOI21_X2 inst_10013 ( .B2(net_9049), .ZN(net_8598), .A(net_8386), .B1(net_8167) );
DFF_X1 inst_8827 ( .QN(net_9649), .D(net_2900), .CK(net_14122) );
INV_X4 inst_6060 ( .A(net_9213), .ZN(net_2495) );
INV_X4 inst_5431 ( .ZN(net_1492), .A(net_1128) );
INV_X4 inst_5023 ( .ZN(net_2845), .A(net_1969) );
DFF_X2 inst_8330 ( .QN(net_10375), .D(net_3218), .CK(net_12109) );
INV_X4 inst_5617 ( .A(net_5792), .ZN(net_1139) );
NAND2_X2 inst_3698 ( .ZN(net_5941), .A2(net_5939), .A1(net_1038) );
CLKBUF_X2 inst_14638 ( .A(net_10614), .Z(net_14557) );
NAND2_X2 inst_4155 ( .ZN(net_2035), .A1(net_2034), .A2(net_2023) );
INV_X2 inst_6962 ( .ZN(net_1862), .A(net_1861) );
INV_X4 inst_5118 ( .A(net_3399), .ZN(net_1618) );
NOR2_X2 inst_2966 ( .A1(net_10158), .A2(net_3988), .ZN(net_3136) );
CLKBUF_X2 inst_14223 ( .A(net_14141), .Z(net_14142) );
NAND3_X2 inst_3246 ( .ZN(net_4699), .A1(net_4698), .A3(net_4697), .A2(net_2357) );
AOI222_X1 inst_9686 ( .B1(net_9505), .A2(net_8301), .B2(net_8300), .C2(net_8299), .ZN(net_8298), .C1(net_8227), .A1(x2214) );
CLKBUF_X2 inst_15102 ( .A(net_15020), .Z(net_15021) );
AOI21_X2 inst_10208 ( .ZN(net_2531), .A(net_2530), .B2(net_1783), .B1(net_1345) );
INV_X4 inst_4904 ( .ZN(net_4475), .A(net_3072) );
CLKBUF_X2 inst_10699 ( .A(net_10617), .Z(net_10618) );
INV_X4 inst_4887 ( .ZN(net_5320), .A(net_4275) );
CLKBUF_X2 inst_11272 ( .A(net_10712), .Z(net_11191) );
INV_X4 inst_5823 ( .ZN(net_5718), .A(net_2496) );
NOR3_X2 inst_2381 ( .ZN(net_7830), .A1(net_7828), .A3(net_7693), .A2(x3390) );
CLKBUF_X2 inst_11538 ( .A(net_11456), .Z(net_11457) );
INV_X4 inst_5338 ( .ZN(net_2281), .A(net_1254) );
SDFF_X2 inst_570 ( .D(net_9147), .SE(net_933), .CK(net_11020), .SI(x1547), .Q(x1121) );
OAI221_X2 inst_1570 ( .C1(net_10322), .C2(net_9047), .B2(net_7287), .B1(net_7184), .ZN(net_7180), .A(net_6803) );
CLKBUF_X2 inst_11284 ( .A(net_10967), .Z(net_11203) );
CLKBUF_X2 inst_14697 ( .A(net_14615), .Z(net_14616) );
CLKBUF_X2 inst_12055 ( .A(net_11973), .Z(net_11974) );
OAI221_X2 inst_1612 ( .C1(net_10208), .B1(net_7249), .C2(net_5642), .ZN(net_5624), .B2(net_4905), .A(net_3507) );
INV_X4 inst_4645 ( .ZN(net_6014), .A(net_6013) );
XNOR2_X1 inst_454 ( .B(net_9615), .A(net_9614), .ZN(net_1041) );
CLKBUF_X2 inst_13947 ( .A(net_13865), .Z(net_13866) );
CLKBUF_X2 inst_13753 ( .A(net_13608), .Z(net_13672) );
CLKBUF_X2 inst_14299 ( .A(net_12648), .Z(net_14218) );
CLKBUF_X2 inst_12545 ( .A(net_10569), .Z(net_12464) );
DFF_X2 inst_8251 ( .Q(net_10180), .D(net_4835), .CK(net_14529) );
CLKBUF_X2 inst_15649 ( .A(net_15567), .Z(net_15568) );
CLKBUF_X2 inst_15475 ( .A(net_15393), .Z(net_15394) );
DFF_X2 inst_7899 ( .QN(net_10126), .D(net_6023), .CK(net_15520) );
CLKBUF_X2 inst_11419 ( .A(net_11337), .Z(net_11338) );
NAND2_X2 inst_3718 ( .ZN(net_7110), .A2(net_5818), .A1(net_5160) );
CLKBUF_X2 inst_12592 ( .A(net_12510), .Z(net_12511) );
CLKBUF_X2 inst_11130 ( .A(net_10828), .Z(net_11049) );
NAND4_X2 inst_3077 ( .A3(net_5375), .ZN(net_4916), .A2(net_4915), .A4(net_4914), .A1(net_3317) );
CLKBUF_X2 inst_11067 ( .A(net_10749), .Z(net_10986) );
INV_X2 inst_6990 ( .ZN(net_2388), .A(net_1645) );
CLKBUF_X2 inst_13622 ( .A(net_12987), .Z(net_13541) );
CLKBUF_X2 inst_12974 ( .A(net_12892), .Z(net_12893) );
CLKBUF_X2 inst_12599 ( .A(net_11633), .Z(net_12518) );
INV_X4 inst_5224 ( .A(net_4788), .ZN(net_1910) );
DFF_X2 inst_8099 ( .QN(net_9930), .D(net_5045), .CK(net_13613) );
AOI22_X2 inst_9566 ( .B1(net_10003), .A1(net_9738), .A2(net_6442), .ZN(net_3753), .B2(net_2468) );
OAI222_X2 inst_1423 ( .B2(net_7665), .A2(net_7664), .C2(net_7663), .ZN(net_4912), .B1(net_3951), .A1(net_2533), .C1(net_1113) );
CLKBUF_X2 inst_14793 ( .A(net_14711), .Z(net_14712) );
NOR3_X2 inst_2419 ( .A1(net_5101), .ZN(net_5007), .A2(net_4125), .A3(net_3016) );
OAI22_X2 inst_1034 ( .A1(net_9081), .A2(net_8922), .B1(net_8919), .ZN(net_7952), .B2(net_3602) );
CLKBUF_X2 inst_15448 ( .A(net_13451), .Z(net_15367) );
CLKBUF_X2 inst_11612 ( .A(net_10763), .Z(net_11531) );
AOI22_X2 inst_9484 ( .B1(net_9716), .A1(net_9684), .A2(net_5966), .ZN(net_3839), .B2(net_3039) );
AOI221_X2 inst_9855 ( .A(net_6889), .B2(net_6888), .C2(net_6887), .ZN(net_6863), .B1(net_3496), .C1(x4520) );
OAI22_X2 inst_1207 ( .A1(net_7241), .A2(net_5107), .B2(net_5105), .ZN(net_5044), .B1(net_5043) );
CLKBUF_X2 inst_14492 ( .A(net_14410), .Z(net_14411) );
SDFF_X2 inst_613 ( .SE(net_3637), .D(net_3636), .SI(net_313), .Q(net_313), .CK(net_13470) );
AOI221_X2 inst_9945 ( .C1(net_10088), .B1(net_10066), .ZN(net_5321), .B2(net_5320), .C2(net_5319), .A(net_4663) );
NAND2_X2 inst_4275 ( .A1(net_6958), .ZN(net_2305), .A2(net_1350) );
DFF_X1 inst_8694 ( .Q(net_9647), .D(net_6806), .CK(net_12836) );
INV_X4 inst_5041 ( .ZN(net_5491), .A(net_1917) );
INV_X4 inst_6444 ( .ZN(net_7209), .A(x3949) );
OAI222_X2 inst_1428 ( .ZN(net_3156), .C2(net_3155), .B2(net_3155), .A2(net_2311), .A1(net_2309), .B1(net_1580), .C1(net_934) );
CLKBUF_X2 inst_11089 ( .A(net_11007), .Z(net_11008) );
SDFF_X2 inst_483 ( .SE(net_9540), .SI(net_8226), .Q(net_299), .D(net_299), .CK(net_13915) );
INV_X4 inst_5005 ( .ZN(net_5171), .A(net_2610) );
AOI221_X2 inst_9907 ( .B1(net_9891), .B2(net_9101), .A(net_6945), .C2(net_6944), .ZN(net_6787), .C1(net_262) );
AOI22_X2 inst_9456 ( .A2(net_10164), .B2(net_8846), .ZN(net_3936), .A1(net_3736), .B1(net_849) );
NOR2_X2 inst_2739 ( .ZN(net_4241), .A2(net_3690), .A1(net_3298) );
XNOR2_X2 inst_259 ( .B(net_9226), .ZN(net_4002), .A(net_3481) );
CLKBUF_X2 inst_12691 ( .A(net_12054), .Z(net_12610) );
INV_X2 inst_6845 ( .A(net_4468), .ZN(net_3511) );
OAI22_X2 inst_1046 ( .ZN(net_7561), .B2(net_7560), .A1(net_5685), .A2(net_4453), .B1(net_1660) );
INV_X2 inst_6812 ( .A(net_10535), .ZN(net_4790) );
INV_X4 inst_5955 ( .ZN(net_1374), .A(net_555) );
AOI21_X2 inst_10152 ( .ZN(net_4138), .A(net_3660), .B2(net_3281), .B1(net_2625) );
NAND2_X2 inst_4355 ( .A2(net_10117), .ZN(net_2878), .A1(net_756) );
INV_X4 inst_5426 ( .A(net_2016), .ZN(net_1131) );
INV_X4 inst_4707 ( .ZN(net_4740), .A(net_4624) );
INV_X4 inst_6206 ( .A(net_10266), .ZN(net_6958) );
INV_X4 inst_4846 ( .ZN(net_3687), .A(net_3297) );
AOI22_X2 inst_9515 ( .B1(net_9995), .A2(net_6443), .ZN(net_3808), .A1(net_3807), .B2(net_2468) );
DFF_X1 inst_8621 ( .Q(net_9665), .D(net_7255), .CK(net_13279) );
DFF_X2 inst_7592 ( .QN(net_9245), .D(net_7466), .CK(net_11252) );
CLKBUF_X2 inst_13197 ( .A(net_12104), .Z(net_13116) );
AND2_X2 inst_10517 ( .ZN(net_4917), .A1(net_4601), .A2(net_4449) );
OR2_X2 inst_909 ( .ZN(net_4395), .A2(net_4394), .A1(net_1678) );
NOR2_X2 inst_2484 ( .A2(net_8899), .ZN(net_8781), .A1(net_8778) );
AOI221_X2 inst_9927 ( .B2(net_5867), .A(net_5859), .ZN(net_5850), .C1(net_5849), .C2(net_4725), .B1(x5077) );
INV_X4 inst_5758 ( .ZN(net_2279), .A(net_728) );
INV_X4 inst_6494 ( .A(net_10407), .ZN(net_355) );
CLKBUF_X2 inst_10686 ( .A(net_10604), .Z(net_10605) );
NOR2_X2 inst_2919 ( .ZN(net_1441), .A2(net_1440), .A1(net_406) );
OR2_X2 inst_894 ( .A1(net_10398), .ZN(net_5779), .A2(net_5777) );
INV_X4 inst_5039 ( .ZN(net_1929), .A(net_1928) );
NOR3_X2 inst_2425 ( .A1(net_7602), .A3(net_4512), .ZN(net_4315), .A2(net_3917) );
OAI21_X2 inst_1872 ( .ZN(net_5291), .A(net_5290), .B2(net_4366), .B1(x4587) );
CLKBUF_X2 inst_10795 ( .A(net_10696), .Z(net_10714) );
CLKBUF_X2 inst_10827 ( .A(net_10745), .Z(net_10746) );
OAI22_X2 inst_994 ( .B1(net_9267), .A2(net_8962), .B2(net_8659), .ZN(net_8638), .A1(net_7510) );
AOI221_X2 inst_9803 ( .B1(net_9982), .A(net_7090), .B2(net_7089), .C2(net_7088), .ZN(net_6999), .C1(net_6823) );
CLKBUF_X2 inst_12003 ( .A(net_11921), .Z(net_11922) );
NAND2_X2 inst_4028 ( .ZN(net_3267), .A2(net_3027), .A1(net_843) );
DFF_X1 inst_8478 ( .Q(net_9626), .D(net_7952), .CK(net_15030) );
OAI21_X2 inst_1879 ( .B2(net_10133), .ZN(net_5244), .A(net_2105), .B1(net_1586) );
OAI21_X2 inst_1863 ( .ZN(net_5423), .A(net_5259), .B2(net_4984), .B1(net_870) );
OAI211_X2 inst_2135 ( .C2(net_6774), .ZN(net_6713), .A(net_6338), .B(net_6076), .C1(net_525) );
CLKBUF_X2 inst_13556 ( .A(net_13237), .Z(net_13475) );
CLKBUF_X2 inst_14082 ( .A(net_12822), .Z(net_14001) );
NAND4_X2 inst_3119 ( .A1(net_9051), .ZN(net_3626), .A2(net_3625), .A4(net_3624), .A3(net_800) );
INV_X4 inst_5138 ( .ZN(net_3977), .A(net_1592) );
NAND2_X2 inst_3777 ( .ZN(net_5872), .A1(net_4784), .A2(net_4780) );
OR2_X4 inst_764 ( .ZN(net_4734), .A1(net_4323), .A2(net_4322) );
CLKBUF_X2 inst_10961 ( .A(net_10879), .Z(net_10880) );
CLKBUF_X2 inst_14515 ( .A(net_14433), .Z(net_14434) );
CLKBUF_X2 inst_12015 ( .A(net_11933), .Z(net_11934) );
OAI221_X2 inst_1547 ( .B2(net_7295), .C2(net_7293), .ZN(net_7214), .C1(net_7213), .A(net_6815), .B1(net_1589) );
XOR2_X2 inst_29 ( .Z(net_2138), .B(net_2014), .A(net_860) );
AOI221_X2 inst_9900 ( .B1(net_9885), .B2(net_9101), .A(net_6945), .C2(net_6944), .ZN(net_6794), .C1(net_256) );
DFF_X1 inst_8469 ( .QN(net_9590), .D(net_7968), .CK(net_11518) );
INV_X2 inst_6937 ( .ZN(net_1922), .A(net_1921) );
AOI222_X1 inst_9713 ( .C2(net_10452), .B1(net_10451), .ZN(net_7797), .A2(net_7712), .B2(net_7547), .C1(net_7333), .A1(net_7307) );
DFF_X2 inst_7782 ( .Q(net_9815), .D(net_6517), .CK(net_15711) );
CLKBUF_X2 inst_11745 ( .A(net_11663), .Z(net_11664) );
NOR3_X2 inst_2369 ( .A3(net_10383), .A2(net_10382), .ZN(net_8256), .A1(net_1542) );
OAI211_X2 inst_2152 ( .C2(net_6774), .ZN(net_6696), .A(net_6315), .B(net_6055), .C1(net_5051) );
INV_X4 inst_6105 ( .A(net_9751), .ZN(net_4211) );
AND2_X2 inst_10540 ( .A1(net_3917), .ZN(net_3637), .A2(net_3636) );
NAND2_X2 inst_3947 ( .ZN(net_4087), .A2(net_3508), .A1(net_610) );
OAI22_X2 inst_1274 ( .A1(net_9607), .ZN(net_4600), .A2(net_4174), .B2(net_3714), .B1(net_3531) );
CLKBUF_X2 inst_15712 ( .A(net_15630), .Z(net_15631) );
CLKBUF_X2 inst_13270 ( .A(net_13188), .Z(net_13189) );
DFF_X2 inst_7740 ( .QN(net_10158), .D(net_6201), .CK(net_13512) );
NAND2_X2 inst_3838 ( .ZN(net_4680), .A2(net_4308), .A1(net_2232) );
CLKBUF_X2 inst_11152 ( .A(net_11070), .Z(net_11071) );
AND2_X2 inst_10590 ( .ZN(net_2389), .A2(net_2388), .A1(net_2206) );
CLKBUF_X2 inst_12775 ( .A(net_11650), .Z(net_12694) );
INV_X4 inst_5495 ( .ZN(net_5886), .A(net_2607) );
INV_X4 inst_5326 ( .A(net_6813), .ZN(net_1270) );
INV_X4 inst_6207 ( .A(net_10282), .ZN(net_467) );
CLKBUF_X2 inst_11396 ( .A(net_10953), .Z(net_11315) );
CLKBUF_X2 inst_14847 ( .A(net_14765), .Z(net_14766) );
SDFF_X2 inst_538 ( .D(net_9148), .SE(net_933), .CK(net_11029), .SI(x1503), .Q(x1113) );
INV_X2 inst_7237 ( .A(net_9214), .ZN(net_379) );
NOR2_X2 inst_2831 ( .ZN(net_2443), .A2(net_2442), .A1(net_1221) );
CLKBUF_X2 inst_12785 ( .A(net_12149), .Z(net_12704) );
DFF_X2 inst_8344 ( .Q(net_9218), .D(net_2741), .CK(net_11304) );
OAI22_X2 inst_1300 ( .A2(net_10337), .B2(net_8841), .ZN(net_3394), .A1(net_3177), .B1(net_1120) );
INV_X4 inst_5280 ( .ZN(net_1517), .A(net_1327) );
INV_X4 inst_4537 ( .ZN(net_8741), .A(net_8736) );
CLKBUF_X2 inst_12022 ( .A(net_11940), .Z(net_11941) );
XOR2_X2 inst_35 ( .Z(net_1751), .A(net_1750), .B(net_1567) );
INV_X4 inst_5317 ( .ZN(net_2889), .A(net_1280) );
CLKBUF_X2 inst_13698 ( .A(net_13616), .Z(net_13617) );
INV_X4 inst_4765 ( .ZN(net_4473), .A(net_4364) );
CLKBUF_X2 inst_13693 ( .A(net_13611), .Z(net_13612) );
AND2_X2 inst_10599 ( .ZN(net_2832), .A2(net_2164), .A1(net_546) );
CLKBUF_X2 inst_11146 ( .A(net_11037), .Z(net_11065) );
INV_X2 inst_7309 ( .A(net_9086), .ZN(net_9085) );
CLKBUF_X2 inst_15284 ( .A(net_15202), .Z(net_15203) );
OAI211_X2 inst_2279 ( .C1(net_7124), .C2(net_6501), .ZN(net_6221), .B(net_5741), .A(net_3679) );
CLKBUF_X2 inst_12572 ( .A(net_11609), .Z(net_12491) );
NOR2_X2 inst_2600 ( .ZN(net_6664), .A2(net_6663), .A1(net_3202) );
CLKBUF_X2 inst_14158 ( .A(net_12123), .Z(net_14077) );
OAI211_X2 inst_2038 ( .C2(net_8102), .B(net_8098), .ZN(net_8078), .A(net_8004), .C1(net_5189) );
OAI211_X2 inst_2044 ( .C2(net_10381), .B(net_8823), .ZN(net_7886), .A(net_7810), .C1(net_6057) );
DFF_X2 inst_7833 ( .Q(net_9814), .D(net_6518), .CK(net_15685) );
INV_X4 inst_5178 ( .A(net_1949), .ZN(net_1912) );
OAI211_X2 inst_2274 ( .C1(net_7127), .C2(net_6548), .A(net_6546), .ZN(net_6248), .B(net_5714) );
AOI21_X2 inst_10055 ( .B2(net_7175), .ZN(net_7141), .B1(net_5268), .A(net_4316) );
CLKBUF_X2 inst_15820 ( .A(net_15738), .Z(net_15739) );
OR3_X4 inst_695 ( .A2(net_9194), .ZN(net_5449), .A1(net_5101), .A3(net_361) );
CLKBUF_X2 inst_15289 ( .A(net_15207), .Z(net_15208) );
CLKBUF_X2 inst_13630 ( .A(net_13548), .Z(net_13549) );
INV_X4 inst_6249 ( .A(net_9536), .ZN(net_711) );
NAND2_X2 inst_4038 ( .ZN(net_2895), .A1(net_2370), .A2(net_1748) );
CLKBUF_X2 inst_15245 ( .A(net_15163), .Z(net_15164) );
CLKBUF_X2 inst_13711 ( .A(net_13629), .Z(net_13630) );
AND2_X2 inst_10606 ( .ZN(net_2033), .A1(net_2032), .A2(net_2031) );
INV_X4 inst_5492 ( .ZN(net_993), .A(net_992) );
CLKBUF_X2 inst_10663 ( .A(net_10572), .Z(net_10582) );
CLKBUF_X2 inst_14001 ( .A(net_13919), .Z(net_13920) );
CLKBUF_X2 inst_10782 ( .A(net_10700), .Z(net_10701) );
INV_X2 inst_6877 ( .ZN(net_3107), .A(net_2875) );
INV_X4 inst_6610 ( .A(net_10029), .ZN(net_612) );
NOR2_X2 inst_2493 ( .ZN(net_8675), .A2(net_8600), .A1(net_6673) );
CLKBUF_X2 inst_14376 ( .A(net_12951), .Z(net_14295) );
INV_X4 inst_6154 ( .A(net_10429), .ZN(net_671) );
SDFF_X2 inst_511 ( .Q(net_9338), .D(net_9338), .SI(net_9330), .SE(net_7588), .CK(net_14695) );
AOI22_X2 inst_9593 ( .B1(net_10014), .A1(net_9784), .ZN(net_3506), .B2(net_2468), .A2(net_2462) );
DFF_X1 inst_8665 ( .D(net_6775), .Q(net_100), .CK(net_12090) );
CLKBUF_X2 inst_14720 ( .A(net_14638), .Z(net_14639) );
NAND2_X2 inst_3559 ( .ZN(net_7808), .A2(net_7709), .A1(net_685) );
INV_X4 inst_5720 ( .ZN(net_3214), .A(net_762) );
CLKBUF_X2 inst_12277 ( .A(net_12195), .Z(net_12196) );
NOR2_X2 inst_2645 ( .ZN(net_5429), .A1(net_5016), .A2(net_5013) );
OAI22_X2 inst_1164 ( .A1(net_7182), .A2(net_5151), .B2(net_5150), .ZN(net_5109), .B1(net_673) );
AOI22_X2 inst_9449 ( .A1(net_10520), .B1(net_9793), .A2(net_4056), .ZN(net_4045), .B2(net_2556) );
NAND4_X2 inst_3112 ( .ZN(net_4436), .A2(net_4266), .A4(net_4258), .A1(net_4109), .A3(net_2767) );
CLKBUF_X2 inst_14025 ( .A(net_11420), .Z(net_13944) );
INV_X2 inst_7183 ( .A(net_9409), .ZN(net_8222) );
CLKBUF_X2 inst_11772 ( .A(net_10799), .Z(net_11691) );
DFF_X2 inst_8328 ( .QN(net_10061), .D(net_3258), .CK(net_11214) );
CLKBUF_X2 inst_12790 ( .A(net_11453), .Z(net_12709) );
CLKBUF_X2 inst_11410 ( .A(net_11328), .Z(net_11329) );
INV_X2 inst_7276 ( .A(net_8949), .ZN(net_8948) );
CLKBUF_X2 inst_15340 ( .A(net_12143), .Z(net_15259) );
CLKBUF_X2 inst_15501 ( .A(net_15419), .Z(net_15420) );
CLKBUF_X2 inst_14613 ( .A(net_14531), .Z(net_14532) );
INV_X2 inst_7004 ( .A(net_2231), .ZN(net_1619) );
INV_X4 inst_6001 ( .A(net_10227), .ZN(net_1063) );
CLKBUF_X2 inst_12506 ( .A(net_11163), .Z(net_12425) );
CLKBUF_X2 inst_11416 ( .A(net_10663), .Z(net_11335) );
CLKBUF_X2 inst_14596 ( .A(net_14514), .Z(net_14515) );
DFF_X2 inst_8193 ( .Q(net_9848), .D(net_5123), .CK(net_14716) );
OAI22_X2 inst_1242 ( .A1(net_7190), .A2(net_4871), .B2(net_4870), .ZN(net_4868), .B1(net_503) );
CLKBUF_X2 inst_14086 ( .A(net_11393), .Z(net_14005) );
CLKBUF_X2 inst_11646 ( .A(net_11564), .Z(net_11565) );
CLKBUF_X2 inst_11525 ( .A(net_11340), .Z(net_11444) );
CLKBUF_X2 inst_10751 ( .A(net_10567), .Z(net_10670) );
CLKBUF_X2 inst_14915 ( .A(net_14833), .Z(net_14834) );
CLKBUF_X2 inst_14578 ( .A(net_14496), .Z(net_14497) );
CLKBUF_X2 inst_10666 ( .A(net_10583), .Z(net_10585) );
INV_X4 inst_6592 ( .A(net_10111), .ZN(net_5849) );
CLKBUF_X2 inst_14865 ( .A(net_13089), .Z(net_14784) );
INV_X2 inst_7209 ( .A(net_9185), .ZN(net_459) );
CLKBUF_X2 inst_13363 ( .A(net_11360), .Z(net_13282) );
INV_X4 inst_5217 ( .ZN(net_3090), .A(net_1515) );
DFF_X2 inst_8362 ( .QN(net_8846), .D(net_2297), .CK(net_12239) );
DFF_X2 inst_8069 ( .QN(net_10366), .D(net_5308), .CK(net_13622) );
XNOR2_X2 inst_388 ( .ZN(net_2271), .B(net_1482), .A(net_553) );
CLKBUF_X2 inst_15307 ( .A(net_11553), .Z(net_15226) );
INV_X4 inst_4600 ( .A(net_7909), .ZN(net_7647) );
CLKBUF_X2 inst_11574 ( .A(net_11492), .Z(net_11493) );
AOI22_X2 inst_9273 ( .B1(net_9701), .ZN(net_5756), .A1(net_5755), .B2(net_5754), .A2(net_238) );
INV_X2 inst_6923 ( .ZN(net_2067), .A(net_2066) );
NAND2_X2 inst_3872 ( .ZN(net_4357), .A1(net_4077), .A2(net_4076) );
CLKBUF_X2 inst_12374 ( .A(net_12292), .Z(net_12293) );
CLKBUF_X2 inst_15119 ( .A(net_12464), .Z(net_15038) );
SDFF_X2 inst_489 ( .SE(net_9540), .SI(net_8220), .Q(net_305), .D(net_305), .CK(net_13902) );
AOI22_X2 inst_9278 ( .B1(net_10006), .ZN(net_5744), .A1(net_5743), .B2(net_5742), .A2(net_246) );
AOI21_X2 inst_10227 ( .B1(net_2882), .ZN(net_2015), .A(net_2014), .B2(net_1256) );
INV_X4 inst_5502 ( .A(net_10462), .ZN(net_4168) );
INV_X2 inst_7153 ( .A(net_4172), .ZN(net_714) );
NAND2_X2 inst_3622 ( .ZN(net_7104), .A2(net_6874), .A1(net_6590) );
CLKBUF_X2 inst_11625 ( .A(net_11543), .Z(net_11544) );
OAI222_X2 inst_1411 ( .B2(net_7732), .A2(net_7731), .C2(net_7730), .ZN(net_5308), .B1(net_4254), .A1(net_3277), .C1(net_1100) );
XNOR2_X2 inst_149 ( .ZN(net_6914), .B(net_6658), .A(net_6657) );
XOR2_X2 inst_39 ( .A(net_9153), .B(net_9152), .Z(net_2470) );
CLKBUF_X2 inst_11028 ( .A(net_10946), .Z(net_10947) );
CLKBUF_X2 inst_12527 ( .A(net_12445), .Z(net_12446) );
DFF_X1 inst_8854 ( .QN(net_9186), .D(net_2090), .CK(net_13594) );
INV_X2 inst_6924 ( .ZN(net_1974), .A(net_1973) );
NOR2_X2 inst_2627 ( .A2(net_9257), .A1(net_8984), .ZN(net_7461) );
CLKBUF_X1 inst_8987 ( .A(x185142), .Z(x936) );
AOI22_X2 inst_9542 ( .B1(net_10001), .A2(net_6443), .ZN(net_3779), .B2(net_2468), .A1(net_901) );
DFF_X2 inst_7771 ( .Q(net_9722), .D(net_6532), .CK(net_14233) );
CLKBUF_X2 inst_15608 ( .A(net_14254), .Z(net_15527) );
CLKBUF_X2 inst_15203 ( .A(net_11617), .Z(net_15122) );
NOR4_X2 inst_2320 ( .A2(net_9850), .ZN(net_6637), .A4(net_5793), .A1(net_3742), .A3(net_619) );
NAND3_X2 inst_3173 ( .ZN(net_8587), .A1(net_8557), .A3(net_8320), .A2(net_8152) );
XNOR2_X2 inst_125 ( .ZN(net_7544), .A(net_7312), .B(net_2190) );
NOR2_X2 inst_2534 ( .A2(net_9593), .A1(net_9089), .ZN(net_8318) );
INV_X4 inst_4770 ( .ZN(net_7828), .A(net_4135) );
CLKBUF_X2 inst_10775 ( .A(net_10693), .Z(net_10694) );
INV_X4 inst_5377 ( .ZN(net_1201), .A(net_1200) );
CLKBUF_X2 inst_15517 ( .A(net_15435), .Z(net_15436) );
DFF_X2 inst_7696 ( .Q(net_10193), .D(net_6576), .CK(net_15139) );
CLKBUF_X2 inst_15233 ( .A(net_12896), .Z(net_15152) );
NAND2_X2 inst_3737 ( .ZN(net_6191), .A1(net_5405), .A2(net_5402) );
CLKBUF_X2 inst_11919 ( .A(net_11837), .Z(net_11838) );
CLKBUF_X2 inst_14753 ( .A(net_14671), .Z(net_14672) );
OAI221_X2 inst_1636 ( .C1(net_10313), .B1(net_7249), .A(net_5637), .C2(net_5591), .ZN(net_5570), .B2(net_4902) );
XNOR2_X2 inst_430 ( .A(net_9305), .B(net_1406), .ZN(net_1083) );
SDFF_X2 inst_515 ( .Q(net_9330), .D(net_9330), .SI(net_9155), .SE(net_7588), .CK(net_13090) );
DFF_X1 inst_8501 ( .Q(net_9856), .D(net_7745), .CK(net_14418) );
CLKBUF_X2 inst_12242 ( .A(net_12160), .Z(net_12161) );
INV_X2 inst_7278 ( .A(net_8960), .ZN(net_8956) );
OAI221_X2 inst_1501 ( .B2(net_9063), .C2(net_9056), .ZN(net_7360), .B1(net_7221), .A(net_7000), .C1(net_5452) );
CLKBUF_X2 inst_11800 ( .A(net_11718), .Z(net_11719) );
NAND3_X2 inst_3212 ( .A2(net_9539), .A3(net_9515), .ZN(net_6681), .A1(net_797) );
NOR2_X2 inst_2565 ( .ZN(net_7724), .A2(net_7588), .A1(net_3685) );
INV_X2 inst_7061 ( .A(net_1322), .ZN(net_1271) );
NOR2_X2 inst_2945 ( .ZN(net_2424), .A1(net_738), .A2(net_549) );
CLKBUF_X2 inst_14982 ( .A(net_14900), .Z(net_14901) );
OAI221_X2 inst_1584 ( .C1(net_10311), .C2(net_9047), .B2(net_7287), .B1(net_7124), .ZN(net_7121), .A(net_6934) );
SDFF_X2 inst_642 ( .Q(net_9456), .D(net_9456), .SE(net_3293), .CK(net_11883), .SI(x2165) );
CLKBUF_X2 inst_14183 ( .A(net_14101), .Z(net_14102) );
CLKBUF_X2 inst_13035 ( .A(net_12953), .Z(net_12954) );
NOR2_X2 inst_2993 ( .A1(net_10461), .ZN(net_2406), .A2(net_888) );
CLKBUF_X2 inst_14736 ( .A(net_14654), .Z(net_14655) );
AOI22_X2 inst_9361 ( .B1(net_9894), .A1(net_6813), .A2(net_5759), .B2(net_5758), .ZN(net_5561) );
CLKBUF_X2 inst_13168 ( .A(net_13086), .Z(net_13087) );
CLKBUF_X2 inst_11023 ( .A(net_10691), .Z(net_10942) );
DFF_X2 inst_7933 ( .QN(net_10331), .D(net_5461), .CK(net_14364) );
OAI22_X2 inst_1018 ( .ZN(net_8038), .A2(net_7927), .B2(net_7926), .A1(net_7157), .B1(net_360) );
CLKBUF_X2 inst_10726 ( .A(net_10644), .Z(net_10645) );
CLKBUF_X2 inst_15499 ( .A(net_12322), .Z(net_15418) );
CLKBUF_X2 inst_10655 ( .A(net_10573), .Z(net_10574) );
DFF_X2 inst_8129 ( .Q(net_9849), .D(net_5130), .CK(net_14738) );
CLKBUF_X2 inst_14160 ( .A(net_14078), .Z(net_14079) );
NOR2_X2 inst_2933 ( .A2(net_4172), .ZN(net_1485), .A1(net_1108) );
OR3_X4 inst_700 ( .A3(net_10409), .ZN(net_7732), .A1(net_4444), .A2(net_4441) );
CLKBUF_X2 inst_13507 ( .A(net_12761), .Z(net_13426) );
CLKBUF_X2 inst_12295 ( .A(net_11740), .Z(net_12214) );
DFF_X1 inst_8706 ( .Q(net_9143), .D(net_6781), .CK(net_11041) );
INV_X4 inst_6467 ( .A(net_9242), .ZN(net_1507) );
CLKBUF_X2 inst_14641 ( .A(net_14559), .Z(net_14560) );
CLKBUF_X2 inst_13323 ( .A(net_13241), .Z(net_13242) );
DFF_X2 inst_8107 ( .Q(net_9826), .D(net_5131), .CK(net_13394) );
AOI22_X2 inst_9152 ( .A1(net_9749), .A2(net_6420), .ZN(net_6332), .B2(net_5263), .B1(net_2564) );
DFF_X1 inst_8555 ( .Q(net_9988), .D(net_7358), .CK(net_12168) );
CLKBUF_X2 inst_14457 ( .A(net_11371), .Z(net_14376) );
OAI22_X2 inst_979 ( .A2(net_9580), .A1(net_8687), .ZN(net_8678), .B2(net_8677), .B1(net_8200) );
NOR2_X2 inst_2713 ( .A1(net_9613), .ZN(net_4151), .A2(net_3973) );
OAI22_X2 inst_1008 ( .ZN(net_8257), .A2(net_8247), .B2(net_8246), .A1(net_5509), .B1(net_1328) );
DFF_X2 inst_7877 ( .Q(net_10045), .D(net_6149), .CK(net_11955) );
INV_X4 inst_4568 ( .ZN(net_8873), .A(net_8385) );
SDFF_X2 inst_559 ( .D(net_9137), .SE(net_933), .CK(net_10981), .SI(x2165), .Q(x1197) );
DFF_X1 inst_8872 ( .Q(net_97), .CK(net_11857), .D(x3314) );
INV_X4 inst_5989 ( .A(net_9970), .ZN(net_538) );
AOI221_X2 inst_9785 ( .B1(net_9965), .A(net_7090), .B2(net_7089), .C1(net_7088), .ZN(net_7082), .C2(net_237) );
AOI22_X2 inst_9476 ( .B1(net_9952), .A1(net_9691), .B2(net_6443), .A2(net_5966), .ZN(net_3847) );
DFF_X2 inst_7706 ( .Q(net_9708), .D(net_6180), .CK(net_14816) );
INV_X2 inst_6725 ( .ZN(net_7777), .A(net_7743) );
OAI211_X2 inst_2296 ( .C2(net_4661), .ZN(net_4383), .C1(net_4382), .B(net_3913), .A(net_3810) );
CLKBUF_X2 inst_11596 ( .A(net_11514), .Z(net_11515) );
AOI22_X2 inst_9250 ( .A2(net_8042), .B2(net_6120), .ZN(net_6061), .A1(net_6060), .B1(net_619) );
CLKBUF_X2 inst_14940 ( .A(net_14858), .Z(net_14859) );
CLKBUF_X2 inst_13092 ( .A(net_13010), .Z(net_13011) );
CLKBUF_X2 inst_12477 ( .A(net_12395), .Z(net_12396) );
CLKBUF_X2 inst_12012 ( .A(net_10805), .Z(net_11931) );
INV_X4 inst_4964 ( .ZN(net_3027), .A(net_2515) );
AOI22_X2 inst_9587 ( .A1(net_10069), .B1(net_10017), .A2(net_5320), .ZN(net_3573), .B2(net_2468) );
NAND2_X2 inst_3405 ( .ZN(net_8555), .A2(net_8554), .A1(net_8511) );
CLKBUF_X2 inst_14133 ( .A(net_13654), .Z(net_14052) );
CLKBUF_X1 inst_8979 ( .A(x185142), .Z(x890) );
NAND2_X2 inst_3888 ( .A2(net_10490), .ZN(net_4745), .A1(net_4006) );
CLKBUF_X2 inst_14912 ( .A(net_11009), .Z(net_14831) );
CLKBUF_X2 inst_14919 ( .A(net_14837), .Z(net_14838) );
CLKBUF_X2 inst_14802 ( .A(net_13008), .Z(net_14721) );
CLKBUF_X2 inst_12831 ( .A(net_12749), .Z(net_12750) );
NAND2_X2 inst_4258 ( .A2(net_10125), .A1(net_10124), .ZN(net_2068) );
DFF_X2 inst_7889 ( .QN(net_10113), .D(net_6026), .CK(net_13265) );
AOI221_X2 inst_9797 ( .B1(net_9977), .A(net_7090), .B2(net_7089), .C2(net_7088), .ZN(net_7007), .C1(net_249) );
AOI22_X2 inst_9607 ( .A1(net_10082), .B1(net_10008), .A2(net_5319), .ZN(net_3446), .B2(net_2468) );
AOI221_X2 inst_9764 ( .ZN(net_7600), .C2(net_7586), .A(net_7452), .C1(net_2887), .B1(net_2887), .B2(net_2444) );
AOI22_X2 inst_9018 ( .ZN(net_8003), .A1(net_8002), .B2(net_8001), .A2(net_7951), .B1(net_1704) );
NAND2_X2 inst_4040 ( .A1(net_3591), .ZN(net_3299), .A2(net_2887) );
CLKBUF_X2 inst_12221 ( .A(net_12139), .Z(net_12140) );
HA_X1 inst_7366 ( .A(net_9174), .B(net_9173), .S(net_1065), .CO(net_1064) );
CLKBUF_X2 inst_15275 ( .A(net_13066), .Z(net_15194) );
NAND2_X2 inst_4334 ( .ZN(net_2964), .A1(net_1101), .A2(x6531) );
OAI22_X2 inst_1059 ( .ZN(net_7059), .A2(net_7036), .B2(net_7035), .A1(net_3331), .B1(net_2174) );
DFF_X2 inst_8017 ( .QN(net_10326), .D(net_5485), .CK(net_12130) );
OAI22_X2 inst_1075 ( .B2(net_10343), .A1(net_10342), .ZN(net_6836), .A2(net_6587), .B1(net_1830) );
CLKBUF_X2 inst_13987 ( .A(net_13905), .Z(net_13906) );
CLKBUF_X2 inst_14227 ( .A(net_14145), .Z(net_14146) );
AOI21_X2 inst_10215 ( .ZN(net_2309), .B2(net_2308), .A(net_1947), .B1(net_1196) );
CLKBUF_X2 inst_12701 ( .A(net_12619), .Z(net_12620) );
AOI22_X2 inst_9230 ( .A1(net_9871), .B1(net_9772), .B2(net_6129), .A2(net_6109), .ZN(net_6081) );
NAND2_X2 inst_4328 ( .A2(net_2012), .ZN(net_1782), .A1(net_1127) );
CLKBUF_X2 inst_15240 ( .A(net_10577), .Z(net_15159) );
CLKBUF_X2 inst_11504 ( .A(net_11272), .Z(net_11423) );
OAI211_X2 inst_2257 ( .C1(net_7249), .C2(net_6480), .ZN(net_6429), .B(net_5435), .A(net_3507) );
CLKBUF_X2 inst_15698 ( .A(net_15616), .Z(net_15617) );
CLKBUF_X2 inst_11781 ( .A(net_11699), .Z(net_11700) );
NAND2_X2 inst_4173 ( .A2(net_4788), .ZN(net_3696), .A1(net_751) );
INV_X4 inst_6039 ( .A(net_10003), .ZN(net_514) );
CLKBUF_X2 inst_15278 ( .A(net_15196), .Z(net_15197) );
CLKBUF_X2 inst_12454 ( .A(net_12372), .Z(net_12373) );
INV_X4 inst_6425 ( .A(net_9532), .ZN(net_382) );
OAI22_X2 inst_1104 ( .A1(net_7157), .ZN(net_6200), .A2(net_5735), .B2(net_5734), .B1(net_343) );
NOR4_X2 inst_2355 ( .A2(net_9224), .A4(net_9220), .A3(net_9219), .ZN(net_1452), .A1(net_317) );
CLKBUF_X2 inst_15553 ( .A(net_14314), .Z(net_15472) );
CLKBUF_X2 inst_14306 ( .A(net_14224), .Z(net_14225) );
CLKBUF_X2 inst_13641 ( .A(net_13559), .Z(net_13560) );
CLKBUF_X2 inst_15210 ( .A(net_15128), .Z(net_15129) );
CLKBUF_X2 inst_10886 ( .A(net_10804), .Z(net_10805) );
INV_X4 inst_6536 ( .ZN(net_4309), .A(net_127) );
INV_X4 inst_5753 ( .A(net_962), .ZN(net_952) );
INV_X2 inst_7058 ( .A(net_4554), .ZN(net_1284) );
CLKBUF_X2 inst_15794 ( .A(net_15712), .Z(net_15713) );
CLKBUF_X2 inst_12535 ( .A(net_11239), .Z(net_12454) );
AOI221_X2 inst_9742 ( .ZN(net_8726), .A(net_8724), .B1(net_8686), .B2(net_8676), .C2(net_8631), .C1(net_8624) );
INV_X4 inst_6434 ( .A(net_9948), .ZN(net_3576) );
INV_X4 inst_6110 ( .ZN(net_6828), .A(net_232) );
XNOR2_X2 inst_329 ( .B(net_9304), .ZN(net_3641), .A(net_2993) );
SDFF_X2 inst_494 ( .SE(net_9540), .SI(net_8215), .Q(net_311), .D(net_311), .CK(net_11648) );
INV_X2 inst_7287 ( .ZN(net_8980), .A(net_8975) );
SDFF_X2 inst_574 ( .D(net_9127), .SE(net_933), .CK(net_10933), .SI(x2767), .Q(x1290) );
CLKBUF_X2 inst_12446 ( .A(net_11758), .Z(net_12365) );
INV_X4 inst_5552 ( .A(net_8756), .ZN(net_8687) );
INV_X4 inst_5942 ( .ZN(net_826), .A(net_568) );
CLKBUF_X2 inst_13845 ( .A(net_13763), .Z(net_13764) );
NOR4_X2 inst_2347 ( .A3(net_10023), .A4(net_4380), .ZN(net_2748), .A1(net_2747), .A2(net_1841) );
CLKBUF_X2 inst_14349 ( .A(net_14267), .Z(net_14268) );
CLKBUF_X2 inst_13085 ( .A(net_13003), .Z(net_13004) );
DFF_X2 inst_8087 ( .Q(net_10047), .D(net_5095), .CK(net_14748) );
NAND2_X2 inst_4102 ( .ZN(net_8998), .A1(net_3531), .A2(net_1707) );
OAI22_X2 inst_1229 ( .B1(net_7224), .A2(net_4890), .B2(net_4889), .ZN(net_4888), .A1(net_486) );
AND2_X2 inst_10512 ( .ZN(net_5316), .A1(net_4986), .A2(net_4709) );
CLKBUF_X2 inst_14167 ( .A(net_14085), .Z(net_14086) );
CLKBUF_X2 inst_14725 ( .A(net_11228), .Z(net_14644) );
DFF_X2 inst_7545 ( .QN(net_9313), .D(net_7742), .CK(net_15312) );
CLKBUF_X2 inst_13780 ( .A(net_13638), .Z(net_13699) );
CLKBUF_X2 inst_13604 ( .A(net_13522), .Z(net_13523) );
INV_X4 inst_5219 ( .ZN(net_4675), .A(net_1510) );
NOR2_X2 inst_2894 ( .ZN(net_1718), .A2(net_1717), .A1(net_830) );
CLKBUF_X2 inst_15042 ( .A(net_14960), .Z(net_14961) );
NOR4_X2 inst_2358 ( .A4(net_9620), .A3(net_9617), .A2(net_9614), .ZN(net_1296), .A1(net_397) );
CLKBUF_X2 inst_13139 ( .A(net_13057), .Z(net_13058) );
INV_X2 inst_7045 ( .ZN(net_2037), .A(net_1185) );
INV_X4 inst_5949 ( .ZN(net_1371), .A(net_895) );
OAI211_X2 inst_2125 ( .C2(net_6778), .ZN(net_6723), .A(net_6350), .B(net_6085), .C1(net_524) );
INV_X4 inst_6085 ( .A(net_9296), .ZN(net_680) );
CLKBUF_X2 inst_15827 ( .A(net_15745), .Z(net_15746) );
AOI21_X2 inst_10192 ( .ZN(net_3276), .A(net_2837), .B1(net_2624), .B2(net_2177) );
CLKBUF_X2 inst_11572 ( .A(net_11440), .Z(net_11491) );
AND2_X2 inst_10549 ( .A1(net_3668), .A2(net_3486), .ZN(net_3483) );
NOR2_X2 inst_2959 ( .A1(net_10439), .ZN(net_2332), .A2(net_694) );
SDFF_X2 inst_599 ( .QN(net_9267), .SE(net_4297), .SI(net_150), .D(net_116), .CK(net_12542) );
CLKBUF_X2 inst_15130 ( .A(net_15048), .Z(net_15049) );
CLKBUF_X2 inst_13906 ( .A(net_10782), .Z(net_13825) );
OAI221_X2 inst_1683 ( .B1(net_7226), .ZN(net_5481), .C1(net_5480), .C2(net_4477), .B2(net_4455), .A(net_3731) );
CLKBUF_X2 inst_10714 ( .A(net_10632), .Z(net_10633) );
NAND2_X2 inst_3865 ( .A1(net_10533), .ZN(net_4084), .A2(net_3873) );
CLKBUF_X2 inst_13382 ( .A(net_12533), .Z(net_13301) );
SDFF_X2 inst_541 ( .Q(net_9303), .D(net_9303), .SI(net_9154), .SE(net_7553), .CK(net_14047) );
NAND2_X2 inst_4047 ( .A2(net_8830), .A1(net_2824), .ZN(net_2823) );
AND2_X4 inst_10459 ( .A2(net_10356), .ZN(net_2752), .A1(net_1347) );
CLKBUF_X2 inst_13910 ( .A(net_11366), .Z(net_13829) );
CLKBUF_X2 inst_13109 ( .A(net_13027), .Z(net_13028) );
SDFF_X2 inst_505 ( .SE(net_9540), .SI(net_8195), .Q(net_302), .D(net_302), .CK(net_13895) );
INV_X4 inst_6366 ( .A(net_10396), .ZN(net_402) );
OAI222_X2 inst_1365 ( .A2(net_7660), .C2(net_7659), .B2(net_7658), .ZN(net_6302), .C1(net_2294), .A1(net_2277), .B1(net_1188) );
INV_X2 inst_7247 ( .ZN(net_3249), .A(net_131) );
CLKBUF_X2 inst_15722 ( .A(net_15640), .Z(net_15641) );
AOI221_X2 inst_9896 ( .B1(net_9881), .B2(net_9101), .A(net_6945), .C2(net_6944), .ZN(net_6798), .C1(net_252) );
DFF_X2 inst_7936 ( .QN(net_10217), .D(net_5634), .CK(net_15508) );
XNOR2_X2 inst_198 ( .ZN(net_5182), .B(net_4918), .A(net_4917) );
CLKBUF_X2 inst_13624 ( .A(net_13542), .Z(net_13543) );
NAND2_X2 inst_4125 ( .ZN(net_2327), .A2(net_1613), .A1(net_1608) );
OAI222_X2 inst_1371 ( .B2(net_7660), .A2(net_7659), .C2(net_7658), .ZN(net_6201), .B1(net_5209), .A1(net_4132), .C1(net_1330) );
CLKBUF_X2 inst_15099 ( .A(net_12859), .Z(net_15018) );
CLKBUF_X2 inst_10809 ( .A(net_10727), .Z(net_10728) );
INV_X4 inst_5622 ( .ZN(net_6255), .A(net_1111) );
NAND2_X2 inst_4321 ( .A2(net_10462), .ZN(net_2405), .A1(net_1107) );
OAI221_X2 inst_1644 ( .B1(net_10427), .C1(net_7184), .ZN(net_5544), .B2(net_4477), .C2(net_4455), .A(net_3507) );
CLKBUF_X2 inst_15486 ( .A(net_15404), .Z(net_15405) );
INV_X4 inst_6346 ( .A(net_9750), .ZN(net_409) );
NAND2_X2 inst_3543 ( .ZN(net_8996), .A2(net_7989), .A1(net_2895) );
CLKBUF_X2 inst_12645 ( .A(net_11489), .Z(net_12564) );
INV_X2 inst_6712 ( .A(net_8538), .ZN(net_8089) );
CLKBUF_X2 inst_10737 ( .A(net_10655), .Z(net_10656) );
DFF_X2 inst_7529 ( .QN(net_9322), .D(net_7780), .CK(net_13061) );
CLKBUF_X2 inst_13867 ( .A(net_13785), .Z(net_13786) );
CLKBUF_X2 inst_13333 ( .A(net_13251), .Z(net_13252) );
CLKBUF_X2 inst_11361 ( .A(net_11279), .Z(net_11280) );
AOI22_X2 inst_9351 ( .B1(net_9797), .A2(net_5766), .B2(net_5765), .ZN(net_5601), .A1(net_235) );
DFF_X2 inst_8158 ( .QN(net_9736), .D(net_5065), .CK(net_12772) );
CLKBUF_X2 inst_15080 ( .A(net_14998), .Z(net_14999) );
CLKBUF_X2 inst_12423 ( .A(net_12341), .Z(net_12342) );
CLKBUF_X2 inst_10974 ( .A(net_10892), .Z(net_10893) );
NAND2_X2 inst_3461 ( .A1(net_9466), .A2(net_8475), .ZN(net_8463) );
AOI221_X2 inst_9754 ( .ZN(net_7771), .B2(net_7770), .C1(net_7697), .A(net_7673), .B1(net_3369), .C2(net_3066) );
CLKBUF_X2 inst_15071 ( .A(net_12747), .Z(net_14990) );
INV_X4 inst_4969 ( .A(net_3088), .ZN(net_2460) );
NAND2_X2 inst_3511 ( .A2(net_8237), .ZN(net_8142), .A1(net_8141) );
DFF_X1 inst_8546 ( .Q(net_9981), .D(net_7360), .CK(net_14412) );
DFF_X2 inst_8244 ( .Q(net_10077), .D(net_4858), .CK(net_10726) );
INV_X4 inst_4692 ( .ZN(net_4835), .A(net_4651) );
INV_X2 inst_6726 ( .A(net_7797), .ZN(net_7762) );
INV_X4 inst_4883 ( .A(net_3298), .ZN(net_2975) );
AND2_X2 inst_10487 ( .A1(net_8967), .ZN(net_8388), .A2(net_8387) );
AND3_X4 inst_10363 ( .A3(net_9231), .A2(net_9230), .ZN(net_2112), .A1(net_1455) );
DFF_X1 inst_8580 ( .Q(net_9672), .D(net_7103), .CK(net_13885) );
INV_X4 inst_5693 ( .ZN(net_2945), .A(net_1013) );
AOI221_X2 inst_9992 ( .B1(net_3855), .ZN(net_3195), .B2(net_3194), .C2(net_3131), .A(net_2735), .C1(net_2413) );
DFF_X2 inst_7538 ( .QN(net_9512), .D(net_9288), .CK(net_11753) );
OAI211_X2 inst_2178 ( .C1(net_7213), .C2(net_6548), .ZN(net_6531), .B(net_5659), .A(net_3679) );
XNOR2_X2 inst_263 ( .ZN(net_3975), .A(net_3657), .B(net_203) );
CLKBUF_X2 inst_10889 ( .A(net_10807), .Z(net_10808) );
XNOR2_X2 inst_185 ( .ZN(net_5210), .A(net_4556), .B(net_1797) );
CLKBUF_X2 inst_15831 ( .A(net_15749), .Z(net_15750) );
AOI22_X2 inst_9498 ( .B1(net_10284), .A1(net_10179), .B2(net_4774), .A2(net_4217), .ZN(net_3825) );
DFF_X2 inst_7399 ( .Q(net_9577), .D(net_8536), .CK(net_13773) );
INV_X4 inst_5953 ( .ZN(net_796), .A(net_557) );
XNOR2_X2 inst_166 ( .ZN(net_5945), .A(net_5366), .B(net_1481) );
INV_X2 inst_6742 ( .A(net_9378), .ZN(net_6954) );
NAND2_X2 inst_3815 ( .A1(net_10084), .A2(net_4534), .ZN(net_4523) );
INV_X4 inst_4786 ( .A(net_5685), .ZN(net_5168) );
CLKBUF_X2 inst_13822 ( .A(net_10740), .Z(net_13741) );
CLKBUF_X2 inst_12617 ( .A(net_12535), .Z(net_12536) );
INV_X4 inst_6307 ( .ZN(net_4024), .A(net_126) );
DFF_X2 inst_7371 ( .Q(net_9367), .D(net_8690), .CK(net_14192) );
OAI21_X2 inst_1757 ( .ZN(net_8507), .A(net_8448), .B2(net_8447), .B1(net_8012) );
NAND2_X2 inst_3851 ( .A2(net_4640), .ZN(net_4222), .A1(net_4221) );
CLKBUF_X2 inst_10650 ( .A(net_10568), .Z(net_10569) );
AOI21_X2 inst_10121 ( .B2(net_9937), .ZN(net_4781), .A(net_4473), .B1(net_627) );
INV_X2 inst_6772 ( .ZN(net_6029), .A(net_5852) );
INV_X4 inst_6370 ( .A(net_10017), .ZN(net_400) );
CLKBUF_X2 inst_12358 ( .A(net_12276), .Z(net_12277) );
CLKBUF_X2 inst_15683 ( .A(net_15601), .Z(net_15602) );
CLKBUF_X2 inst_11923 ( .A(net_11841), .Z(net_11842) );
INV_X4 inst_6359 ( .ZN(net_7226), .A(x4359) );
NAND2_X2 inst_4118 ( .ZN(net_2346), .A1(net_2345), .A2(net_1628) );
CLKBUF_X2 inst_12026 ( .A(net_10579), .Z(net_11945) );
CLKBUF_X2 inst_13410 ( .A(net_13328), .Z(net_13329) );
OAI221_X2 inst_1605 ( .C1(net_10202), .B1(net_7192), .C2(net_5642), .ZN(net_5631), .B2(net_4905), .A(net_3731) );
INV_X4 inst_5440 ( .ZN(net_1104), .A(net_1103) );
INV_X4 inst_4849 ( .ZN(net_3507), .A(net_3298) );
CLKBUF_X2 inst_14689 ( .A(net_14607), .Z(net_14608) );
AOI21_X2 inst_10206 ( .ZN(net_2535), .A(net_2534), .B2(net_1781), .B1(net_1572) );
CLKBUF_X2 inst_11635 ( .A(net_11182), .Z(net_11554) );
CLKBUF_X2 inst_13593 ( .A(net_13511), .Z(net_13512) );
CLKBUF_X2 inst_14508 ( .A(net_14426), .Z(net_14427) );
INV_X4 inst_4649 ( .ZN(net_6587), .A(net_5783) );
CLKBUF_X2 inst_12904 ( .A(net_12683), .Z(net_12823) );
AND2_X2 inst_10558 ( .ZN(net_3283), .A1(net_3196), .A2(net_2923) );
DFF_X2 inst_8185 ( .Q(net_9954), .D(net_5002), .CK(net_13185) );
CLKBUF_X2 inst_11223 ( .A(net_11141), .Z(net_11142) );
CLKBUF_X2 inst_12922 ( .A(net_10701), .Z(net_12841) );
INV_X4 inst_5308 ( .ZN(net_5482), .A(net_1292) );
DFF_X2 inst_7413 ( .QN(net_9390), .D(net_8356), .CK(net_14022) );
CLKBUF_X2 inst_15770 ( .A(net_15688), .Z(net_15689) );
CLKBUF_X2 inst_15709 ( .A(net_15627), .Z(net_15628) );
CLKBUF_X2 inst_14634 ( .A(net_14552), .Z(net_14553) );
CLKBUF_X2 inst_14263 ( .A(net_11040), .Z(net_14182) );
MUX2_X1 inst_4475 ( .S(net_6041), .A(net_3704), .B(x6401), .Z(x401) );
DFF_X2 inst_7590 ( .QN(net_9302), .D(net_7500), .CK(net_14100) );
DFF_X1 inst_8698 ( .D(net_6746), .Q(net_107), .CK(net_15096) );
INV_X4 inst_5034 ( .A(net_3761), .ZN(net_3533) );
INV_X4 inst_4853 ( .A(net_3456), .ZN(net_3284) );
INV_X4 inst_6322 ( .A(net_10285), .ZN(net_419) );
DFF_X2 inst_7757 ( .Q(net_9654), .D(net_6552), .CK(net_14095) );
CLKBUF_X2 inst_11077 ( .A(net_10995), .Z(net_10996) );
NAND2_X2 inst_3898 ( .ZN(net_4078), .A2(net_3611), .A1(x6599) );
CLKBUF_X2 inst_14831 ( .A(net_14749), .Z(net_14750) );
INV_X4 inst_5254 ( .ZN(net_1850), .A(net_1435) );
INV_X4 inst_5201 ( .ZN(net_1857), .A(net_1533) );
NOR3_X2 inst_2373 ( .A3(net_10173), .A2(net_10172), .ZN(net_8155), .A1(net_1122) );
AOI22_X2 inst_9370 ( .B1(net_10016), .A2(net_5743), .B2(net_5742), .ZN(net_5552), .A1(net_256) );
CLKBUF_X2 inst_11949 ( .A(net_11867), .Z(net_11868) );
CLKBUF_X2 inst_15321 ( .A(net_15239), .Z(net_15240) );
CLKBUF_X2 inst_11436 ( .A(net_10763), .Z(net_11355) );
NAND2_X2 inst_3503 ( .ZN(net_8369), .A1(net_8179), .A2(net_8178) );
CLKBUF_X2 inst_13974 ( .A(net_13892), .Z(net_13893) );
AOI22_X2 inst_9215 ( .A1(net_9908), .B1(net_9809), .A2(net_8042), .B2(net_8041), .ZN(net_6096) );
DFF_X2 inst_7973 ( .QN(net_10307), .D(net_5579), .CK(net_13240) );
OAI222_X2 inst_1331 ( .B1(net_9068), .C2(net_9054), .ZN(net_7977), .A2(net_7974), .B2(net_7973), .A1(net_3061), .C1(net_1584) );
CLKBUF_X2 inst_12322 ( .A(net_12240), .Z(net_12241) );
DFF_X2 inst_7604 ( .Q(net_9350), .D(net_7337), .CK(net_15293) );
NAND2_X2 inst_4138 ( .ZN(net_2982), .A1(net_2712), .A2(net_2066) );
XOR2_X1 inst_52 ( .B(net_9204), .Z(net_2814), .A(net_2511) );
CLKBUF_X2 inst_15779 ( .A(net_15697), .Z(net_15698) );
DFF_X2 inst_7404 ( .QN(net_9637), .D(net_8323), .CK(net_15384) );
CLKBUF_X2 inst_12600 ( .A(net_12518), .Z(net_12519) );
SDFF_X2 inst_668 ( .SI(net_9500), .Q(net_9500), .SE(net_3073), .CK(net_12393), .D(x1459) );
NAND3_X2 inst_3223 ( .A2(net_9534), .A1(net_5353), .A3(net_5351), .ZN(net_5350) );
NAND4_X2 inst_3049 ( .ZN(net_6157), .A4(net_5339), .A3(net_4052), .A1(net_3801), .A2(net_3570) );
CLKBUF_X2 inst_15804 ( .A(net_11224), .Z(net_15723) );
CLKBUF_X2 inst_11987 ( .A(net_11905), .Z(net_11906) );
NAND2_X2 inst_3560 ( .ZN(net_7710), .A2(net_7709), .A1(net_644) );
NAND2_X2 inst_4159 ( .A1(net_4309), .ZN(net_1980), .A2(net_1396) );
NOR2_X2 inst_2683 ( .A2(net_9588), .A1(net_9069), .ZN(net_8927) );
CLKBUF_X2 inst_13736 ( .A(net_13654), .Z(net_13655) );
CLKBUF_X2 inst_12567 ( .A(net_11501), .Z(net_12486) );
NAND2_X2 inst_4223 ( .A2(net_7002), .A1(net_6158), .ZN(net_1660) );
NAND2_X4 inst_3349 ( .ZN(net_8905), .A2(net_8893), .A1(net_8892) );
CLKBUF_X2 inst_11444 ( .A(net_11031), .Z(net_11363) );
CLKBUF_X2 inst_14277 ( .A(net_14195), .Z(net_14196) );
CLKBUF_X2 inst_14152 ( .A(net_14070), .Z(net_14071) );
AOI21_X2 inst_10057 ( .ZN(net_7100), .B2(net_6664), .A(net_3205), .B1(net_2401) );
NOR2_X2 inst_2545 ( .A2(net_9599), .ZN(net_8135), .A1(net_8057) );
DFF_X2 inst_8220 ( .Q(net_10081), .D(net_4854), .CK(net_10683) );
CLKBUF_X2 inst_12390 ( .A(net_12308), .Z(net_12309) );
CLKBUF_X2 inst_10722 ( .A(net_10640), .Z(net_10641) );
DFF_X2 inst_7999 ( .QN(net_10440), .D(net_5514), .CK(net_13721) );
CLKBUF_X2 inst_13283 ( .A(net_13201), .Z(net_13202) );
CLKBUF_X2 inst_13077 ( .A(net_12995), .Z(net_12996) );
NOR2_X2 inst_2768 ( .A1(net_9613), .ZN(net_3269), .A2(net_2520) );
INV_X2 inst_6677 ( .ZN(net_8351), .A(net_8288) );
CLKBUF_X2 inst_14657 ( .A(net_14575), .Z(net_14576) );
AOI221_X2 inst_9878 ( .B1(net_9785), .B2(net_9098), .A(net_6940), .C2(net_6939), .ZN(net_6822), .C1(net_6821) );
OAI21_X2 inst_1835 ( .ZN(net_6290), .B1(net_6289), .A(net_6011), .B2(net_5823) );
OAI21_X2 inst_1910 ( .ZN(net_4664), .B2(net_4661), .A(net_4381), .B1(net_2192) );
CLKBUF_X2 inst_13777 ( .A(net_13695), .Z(net_13696) );
CLKBUF_X2 inst_15614 ( .A(net_15532), .Z(net_15533) );
CLKBUF_X2 inst_14461 ( .A(net_12186), .Z(net_14380) );
CLKBUF_X2 inst_13420 ( .A(net_13338), .Z(net_13339) );
INV_X4 inst_4639 ( .ZN(net_7276), .A(net_6234) );
CLKBUF_X2 inst_12399 ( .A(net_12317), .Z(net_12318) );
AOI22_X2 inst_9670 ( .A2(net_10086), .B2(net_10085), .A1(net_10068), .B1(net_10067), .ZN(net_927) );
DFF_X2 inst_7797 ( .Q(net_9893), .D(net_6496), .CK(net_15429) );
CLKBUF_X2 inst_15410 ( .A(net_14521), .Z(net_15329) );
CLKBUF_X2 inst_15176 ( .A(net_13234), .Z(net_15095) );
SDFF_X2 inst_621 ( .Q(net_9451), .D(net_9451), .SE(net_3293), .CK(net_11369), .SI(x2477) );
AOI211_X2 inst_10272 ( .A(net_7704), .ZN(net_7570), .C2(net_7453), .C1(net_4305), .B(x3390) );
DFF_X2 inst_7764 ( .Q(net_9695), .D(net_6541), .CK(net_15434) );
AOI22_X2 inst_9265 ( .ZN(net_6646), .A2(net_5222), .B1(net_3853), .B2(net_2899), .A1(net_2685) );
INV_X4 inst_5814 ( .A(net_4566), .ZN(net_679) );
NAND4_X2 inst_3115 ( .A3(net_6669), .ZN(net_4242), .A2(net_4241), .A4(net_3626), .A1(net_448) );
NOR2_X2 inst_2560 ( .ZN(net_7752), .A2(net_7653), .A1(net_3355) );
CLKBUF_X2 inst_10867 ( .A(net_10785), .Z(net_10786) );
NAND3_X2 inst_3219 ( .ZN(net_9103), .A2(net_5356), .A1(net_4903), .A3(net_4797) );
INV_X4 inst_5673 ( .A(net_10304), .ZN(net_1495) );
AOI21_X2 inst_10025 ( .B1(net_9365), .A(net_7916), .B2(net_7915), .ZN(net_7854) );
CLKBUF_X2 inst_15224 ( .A(net_15142), .Z(net_15143) );
CLKBUF_X2 inst_12236 ( .A(net_10610), .Z(net_12155) );
AOI22_X2 inst_9651 ( .B2(net_10456), .A2(net_10455), .ZN(net_3151), .B1(net_701), .A1(net_671) );
CLKBUF_X2 inst_14435 ( .A(net_12410), .Z(net_14354) );
OAI222_X2 inst_1387 ( .B1(net_7732), .A2(net_7731), .C2(net_7730), .ZN(net_5958), .B2(net_5204), .A1(net_4131), .C1(net_1149) );
CLKBUF_X2 inst_15138 ( .A(net_11695), .Z(net_15057) );
CLKBUF_X2 inst_14872 ( .A(net_12754), .Z(net_14791) );
OAI21_X2 inst_1991 ( .ZN(net_2599), .B1(net_2598), .A(net_1465), .B2(net_1058) );
CLKBUF_X2 inst_13687 ( .A(net_13605), .Z(net_13606) );
NOR3_X2 inst_2365 ( .A3(net_9587), .A1(net_8848), .ZN(net_8786), .A2(net_8776) );
CLKBUF_X2 inst_13054 ( .A(net_12594), .Z(net_12973) );
NAND4_X2 inst_3066 ( .ZN(net_5690), .A4(net_4736), .A1(net_3782), .A3(net_3771), .A2(net_3754) );
CLKBUF_X2 inst_12094 ( .A(net_12012), .Z(net_12013) );
OAI211_X2 inst_2250 ( .C1(net_7297), .C2(net_6480), .ZN(net_6446), .B(net_5753), .A(net_3679) );
DFF_X2 inst_7861 ( .Q(net_9801), .D(net_6437), .CK(net_12777) );
CLKBUF_X2 inst_14129 ( .A(net_13311), .Z(net_14048) );
CLKBUF_X2 inst_15441 ( .A(net_15359), .Z(net_15360) );
CLKBUF_X2 inst_15190 ( .A(net_15108), .Z(net_15109) );
CLKBUF_X2 inst_11630 ( .A(net_11061), .Z(net_11549) );
INV_X4 inst_6629 ( .A(net_8983), .ZN(net_8982) );
DFF_X2 inst_7419 ( .QN(net_9419), .D(net_8343), .CK(net_11693) );
OAI211_X2 inst_2187 ( .C1(net_7182), .C2(net_6542), .ZN(net_6522), .B(net_5617), .A(net_3679) );
CLKBUF_X2 inst_13221 ( .A(net_13139), .Z(net_13140) );
CLKBUF_X2 inst_11215 ( .A(net_11133), .Z(net_11134) );
INV_X2 inst_6771 ( .ZN(net_6030), .A(net_5855) );
INV_X4 inst_5747 ( .ZN(net_913), .A(net_741) );
CLKBUF_X2 inst_14323 ( .A(net_13182), .Z(net_14242) );
DFF_X2 inst_8173 ( .QN(net_9827), .D(net_5038), .CK(net_14346) );
DFF_X2 inst_7448 ( .QN(net_9292), .D(net_8245), .CK(net_14997) );
INV_X4 inst_6640 ( .ZN(net_9079), .A(net_9078) );
INV_X4 inst_4703 ( .A(net_6677), .ZN(net_5342) );
NOR2_X2 inst_2672 ( .ZN(net_5368), .A2(net_4791), .A1(net_2753) );
XOR2_X2 inst_25 ( .Z(net_2268), .B(net_978), .A(net_672) );
AOI22_X2 inst_9043 ( .A1(net_9155), .A2(net_7155), .B2(net_7154), .ZN(net_7012), .B1(net_1986) );
INV_X4 inst_5239 ( .ZN(net_1885), .A(net_1470) );
NAND2_X2 inst_3527 ( .ZN(net_8238), .A1(net_8091), .A2(net_8090) );
INV_X4 inst_5032 ( .ZN(net_2243), .A(net_2129) );
CLKBUF_X2 inst_13924 ( .A(net_13842), .Z(net_13843) );
INV_X4 inst_5166 ( .ZN(net_1742), .A(net_1566) );
CLKBUF_X2 inst_13637 ( .A(net_13555), .Z(net_13556) );
AOI222_X1 inst_9691 ( .B1(net_9511), .A2(net_8301), .B2(net_8300), .C2(net_8299), .ZN(net_8290), .C1(net_8221), .A1(x1865) );
AOI22_X2 inst_9558 ( .B1(net_10402), .A2(net_6413), .B2(net_4062), .ZN(net_3762), .A1(net_3761) );
NOR2_X2 inst_2500 ( .ZN(net_8601), .A2(net_8535), .A1(net_1166) );
CLKBUF_X2 inst_12119 ( .A(net_11808), .Z(net_12038) );
AOI222_X1 inst_9734 ( .C2(net_10510), .B2(net_10509), .A2(net_10508), .C1(net_10502), .B1(net_10501), .A1(net_10500), .ZN(net_1446) );
INV_X4 inst_6045 ( .A(net_10290), .ZN(net_511) );
NAND2_X2 inst_4395 ( .A2(net_10405), .A1(net_10391), .ZN(net_733) );
NAND2_X2 inst_3434 ( .A1(net_9482), .ZN(net_9017), .A2(net_8490) );
AOI22_X2 inst_9042 ( .A1(net_9154), .A2(net_7155), .B2(net_7154), .ZN(net_7013), .B1(net_1984) );
INV_X4 inst_6408 ( .A(net_9973), .ZN(net_387) );
NAND2_X2 inst_4296 ( .A2(net_2010), .ZN(net_1783), .A1(net_1387) );
NAND2_X2 inst_3764 ( .ZN(net_7658), .A2(net_4979), .A1(net_596) );
DFF_X1 inst_8764 ( .Q(net_10135), .D(net_5010), .CK(net_10782) );
CLKBUF_X2 inst_11912 ( .A(net_11830), .Z(net_11831) );
CLKBUF_X2 inst_13101 ( .A(net_13019), .Z(net_13020) );
HA_X1 inst_7330 ( .S(net_7652), .CO(net_7651), .B(net_7462), .A(net_5792) );
DFF_X2 inst_7581 ( .Q(net_10190), .D(net_7536), .CK(net_12290) );
NOR4_X2 inst_2340 ( .A3(net_9924), .A4(net_6047), .ZN(net_3128), .A1(net_3127), .A2(net_2637) );
NAND3_X2 inst_3204 ( .ZN(net_6936), .A1(net_6417), .A2(net_3806), .A3(net_3805) );
CLKBUF_X2 inst_15492 ( .A(net_12912), .Z(net_15411) );
CLKBUF_X2 inst_14219 ( .A(net_14137), .Z(net_14138) );
NAND2_X2 inst_3421 ( .A2(net_8877), .A1(net_8876), .ZN(net_8513) );
MUX2_X1 inst_4444 ( .S(net_6041), .A(net_302), .B(x4694), .Z(x101) );
CLKBUF_X2 inst_12019 ( .A(net_11937), .Z(net_11938) );
NOR2_X2 inst_2679 ( .ZN(net_4985), .A2(net_4680), .A1(net_1063) );
XOR2_X2 inst_16 ( .Z(net_2790), .A(net_2017), .B(net_1073) );
INV_X2 inst_6935 ( .ZN(net_1927), .A(net_1926) );
CLKBUF_X2 inst_15362 ( .A(net_15280), .Z(net_15281) );
CLKBUF_X2 inst_14173 ( .A(net_14091), .Z(net_14092) );
NAND2_X2 inst_3949 ( .A2(net_9609), .A1(net_9608), .ZN(net_3714) );
CLKBUF_X2 inst_15731 ( .A(net_15519), .Z(net_15650) );
NOR2_X2 inst_2808 ( .A2(net_8866), .ZN(net_5364), .A1(net_2752) );
XNOR2_X2 inst_156 ( .ZN(net_6197), .A(net_5710), .B(net_2183) );
INV_X4 inst_4617 ( .ZN(net_8102), .A(net_7474) );
OAI21_X2 inst_1777 ( .B2(net_7805), .ZN(net_7801), .B1(net_5331), .A(net_833) );
CLKBUF_X2 inst_14971 ( .A(net_14889), .Z(net_14890) );
INV_X4 inst_6239 ( .A(net_9385), .ZN(net_1774) );
OAI22_X2 inst_1068 ( .B2(net_10168), .ZN(net_6909), .A2(net_6634), .A1(net_6633), .B1(net_6305) );
OR2_X2 inst_886 ( .A2(net_7038), .ZN(net_6209), .A1(net_6208) );
CLKBUF_X2 inst_12799 ( .A(net_12717), .Z(net_12718) );
CLKBUF_X2 inst_11799 ( .A(net_10943), .Z(net_11718) );
NAND2_X2 inst_3442 ( .A1(net_9448), .A2(net_8479), .ZN(net_8478) );
CLKBUF_X2 inst_12509 ( .A(net_12427), .Z(net_12428) );
NOR2_X2 inst_2693 ( .ZN(net_4538), .A2(net_4537), .A1(net_4224) );
CLKBUF_X2 inst_14920 ( .A(net_14838), .Z(net_14839) );
CLKBUF_X2 inst_15409 ( .A(net_15327), .Z(net_15328) );
INV_X4 inst_5350 ( .ZN(net_1521), .A(net_1235) );
CLKBUF_X2 inst_15251 ( .A(net_12470), .Z(net_15170) );
AOI211_X2 inst_10307 ( .ZN(net_3164), .A(net_3163), .C2(net_2683), .C1(net_2376), .B(net_619) );
CLKBUF_X2 inst_14838 ( .A(net_13170), .Z(net_14757) );
INV_X4 inst_5380 ( .A(net_2183), .ZN(net_1198) );
CLKBUF_X2 inst_10936 ( .A(net_10854), .Z(net_10855) );
CLKBUF_X2 inst_13319 ( .A(net_13237), .Z(net_13238) );
INV_X4 inst_6473 ( .A(net_9374), .ZN(net_7905) );
MUX2_X1 inst_4468 ( .S(net_6041), .A(net_5972), .B(x6241), .Z(x341) );
CLKBUF_X2 inst_11740 ( .A(net_11658), .Z(net_11659) );
NOR2_X2 inst_3020 ( .A2(net_10513), .A1(net_10512), .ZN(net_659) );
OAI221_X2 inst_1549 ( .B2(net_9047), .C2(net_7287), .ZN(net_7210), .C1(net_7209), .A(net_6788), .B1(net_5518) );
CLKBUF_X2 inst_12894 ( .A(net_12812), .Z(net_12813) );
CLKBUF_X2 inst_11533 ( .A(net_10971), .Z(net_11452) );
AOI22_X2 inst_9239 ( .A1(net_9940), .B1(net_9841), .B2(net_8041), .A2(net_6109), .ZN(net_6072) );
INV_X4 inst_6186 ( .A(net_10463), .ZN(net_4566) );
CLKBUF_X2 inst_14450 ( .A(net_14368), .Z(net_14369) );
CLKBUF_X2 inst_11484 ( .A(net_11402), .Z(net_11403) );
CLKBUF_X2 inst_11270 ( .A(net_11188), .Z(net_11189) );
CLKBUF_X2 inst_12380 ( .A(net_11594), .Z(net_12299) );
CLKBUF_X2 inst_13477 ( .A(net_13395), .Z(net_13396) );
AND2_X2 inst_10576 ( .ZN(net_3309), .A2(net_2832), .A1(net_379) );
DFF_X1 inst_8844 ( .Q(net_9199), .D(net_2445), .CK(net_13596) );
OAI21_X2 inst_1969 ( .B1(net_5454), .ZN(net_3254), .A(net_3013), .B2(net_2810) );
AOI22_X2 inst_9113 ( .A1(net_9666), .A2(net_6404), .ZN(net_6376), .B2(net_5263), .B1(net_104) );
DFF_X2 inst_7837 ( .Q(net_9180), .D(net_6296), .CK(net_13573) );
NOR2_X2 inst_2881 ( .A2(net_10538), .ZN(net_2463), .A1(net_521) );
OR2_X4 inst_821 ( .ZN(net_1859), .A1(net_935), .A2(net_697) );
CLKBUF_X2 inst_11382 ( .A(net_11300), .Z(net_11301) );
DFF_X1 inst_8879 ( .Q(net_92), .CK(net_14110), .D(x3360) );
AOI22_X2 inst_9128 ( .A1(net_9713), .A2(net_6382), .ZN(net_6360), .B2(net_5263), .B1(net_1019) );
CLKBUF_X2 inst_15631 ( .A(net_15549), .Z(net_15550) );
AOI22_X2 inst_9348 ( .B1(net_9823), .A1(net_6811), .A2(net_5766), .B2(net_5765), .ZN(net_5604) );
DFF_X2 inst_8183 ( .Q(net_9951), .D(net_5003), .CK(net_12329) );
INV_X2 inst_6914 ( .A(net_2530), .ZN(net_2177) );
OAI22_X2 inst_980 ( .A2(net_8962), .ZN(net_8661), .B2(net_8659), .B1(net_7043), .A1(net_6317) );
CLKBUF_X2 inst_15004 ( .A(net_14922), .Z(net_14923) );
INV_X4 inst_6540 ( .A(net_9976), .ZN(net_337) );
CLKBUF_X2 inst_15750 ( .A(net_15668), .Z(net_15669) );
CLKBUF_X2 inst_14536 ( .A(net_14454), .Z(net_14455) );
DFF_X1 inst_8486 ( .QN(net_9633), .D(net_7945), .CK(net_11511) );
CLKBUF_X2 inst_13136 ( .A(net_13054), .Z(net_13055) );
OAI21_X2 inst_1785 ( .A(net_9310), .ZN(net_7646), .B2(net_4551), .B1(net_3726) );
AOI21_X2 inst_10104 ( .B1(net_9531), .A(net_4907), .ZN(net_4894), .B2(net_4893) );
CLKBUF_X2 inst_12939 ( .A(net_12857), .Z(net_12858) );
NAND2_X2 inst_4213 ( .ZN(net_4237), .A2(net_2972), .A1(x6599) );
NAND4_X2 inst_3150 ( .ZN(net_2157), .A4(net_1445), .A2(net_964), .A1(net_662), .A3(net_616) );
CLKBUF_X2 inst_15180 ( .A(net_13267), .Z(net_15099) );
AOI22_X2 inst_9341 ( .B1(net_9817), .A1(net_6821), .A2(net_5766), .B2(net_5765), .ZN(net_5611) );
CLKBUF_X2 inst_10761 ( .A(net_10679), .Z(net_10680) );
AOI22_X2 inst_9575 ( .A1(net_6892), .B2(net_6625), .ZN(net_6219), .B1(net_3704), .A2(net_3030) );
CLKBUF_X2 inst_12765 ( .A(net_12683), .Z(net_12684) );
CLKBUF_X2 inst_12118 ( .A(net_11444), .Z(net_12037) );
CLKBUF_X2 inst_10694 ( .A(net_10612), .Z(net_10613) );
DFF_X1 inst_8522 ( .QN(net_9424), .D(net_7411), .CK(net_13780) );
INV_X4 inst_6022 ( .A(net_9641), .ZN(net_1029) );
OAI211_X2 inst_2286 ( .C1(net_7108), .C2(net_6480), .ZN(net_6193), .B(net_5713), .A(net_3679) );
CLKBUF_X2 inst_14741 ( .A(net_14659), .Z(net_14660) );
INV_X4 inst_6216 ( .ZN(net_951), .A(net_179) );
INV_X4 inst_5791 ( .ZN(net_2860), .A(net_693) );
OR2_X2 inst_866 ( .ZN(net_7794), .A1(net_7611), .A2(net_7543) );
DFF_X2 inst_7512 ( .QN(net_9372), .D(net_7942), .CK(net_11916) );
INV_X2 inst_7142 ( .A(net_1702), .ZN(net_816) );
OAI211_X2 inst_2137 ( .C2(net_6778), .ZN(net_6711), .A(net_6403), .B(net_6075), .C1(net_516) );
CLKBUF_X2 inst_11061 ( .A(net_10979), .Z(net_10980) );
AOI22_X2 inst_9406 ( .A1(net_6892), .B2(net_6625), .ZN(net_6293), .B1(net_4910), .A2(net_4302) );
OAI221_X4 inst_1439 ( .B2(net_9630), .B1(net_8971), .ZN(net_8181), .A(net_7955), .C2(net_3526), .C1(net_174) );
INV_X2 inst_7214 ( .ZN(net_725), .A(x6157) );
NAND2_X2 inst_3640 ( .A2(net_7281), .ZN(net_7252), .A1(net_6904) );
INV_X2 inst_7107 ( .A(net_1059), .ZN(net_1019) );
CLKBUF_X2 inst_12367 ( .A(net_12285), .Z(net_12286) );
DFF_X1 inst_8444 ( .Q(net_9435), .D(net_8171), .CK(net_14933) );
INV_X4 inst_5604 ( .A(net_1011), .ZN(net_876) );
XNOR2_X2 inst_248 ( .B(net_9278), .ZN(net_4127), .A(net_3327) );
OAI221_X2 inst_1613 ( .C1(net_10209), .B1(net_7129), .C2(net_5642), .ZN(net_5623), .B2(net_4905), .A(net_3507) );
NAND4_X2 inst_3107 ( .ZN(net_4336), .A1(net_3789), .A3(net_3770), .A2(net_3753), .A4(net_3412) );
INV_X4 inst_6624 ( .A(net_8960), .ZN(net_8959) );
OAI21_X2 inst_1919 ( .B1(net_7785), .ZN(net_4568), .A(net_4140), .B2(net_4139) );
CLKBUF_X2 inst_15508 ( .A(net_11294), .Z(net_15427) );
INV_X4 inst_5659 ( .ZN(net_1218), .A(net_824) );
CLKBUF_X2 inst_15747 ( .A(net_15665), .Z(net_15666) );
INV_X4 inst_5965 ( .ZN(net_4017), .A(net_120) );
CLKBUF_X2 inst_15098 ( .A(net_15016), .Z(net_15017) );
CLKBUF_X2 inst_12222 ( .A(net_11267), .Z(net_12141) );
OAI22_X2 inst_1141 ( .A1(net_7139), .A2(net_5134), .B2(net_5133), .ZN(net_5132), .B1(net_381) );
NAND2_X2 inst_3589 ( .A2(net_8659), .ZN(net_7364), .A1(net_7363) );
NOR2_X2 inst_2488 ( .ZN(net_8734), .A2(net_8728), .A1(net_8168) );
AND2_X2 inst_10528 ( .ZN(net_4165), .A2(net_3964), .A1(net_1303) );
OR2_X2 inst_932 ( .ZN(net_2672), .A1(net_2671), .A2(net_2670) );
CLKBUF_X2 inst_12891 ( .A(net_10570), .Z(net_12810) );
XNOR2_X2 inst_180 ( .ZN(net_5248), .A(net_4693), .B(net_2319) );
CLKBUF_X2 inst_13472 ( .A(net_13390), .Z(net_13391) );
OAI21_X2 inst_1960 ( .A(net_4714), .B2(net_4070), .ZN(net_3592), .B1(net_3591) );
CLKBUF_X2 inst_15675 ( .A(net_15593), .Z(net_15594) );
AOI22_X2 inst_9057 ( .B1(net_9678), .A2(net_6684), .B2(net_6683), .ZN(net_6609), .A1(net_247) );
DFF_X2 inst_8003 ( .QN(net_10115), .D(net_5506), .CK(net_12349) );
CLKBUF_X2 inst_15474 ( .A(net_15392), .Z(net_15393) );
CLKBUF_X2 inst_11995 ( .A(net_11913), .Z(net_11914) );
DFF_X1 inst_8475 ( .QN(net_9600), .D(net_7860), .CK(net_13805) );
DFF_X1 inst_8712 ( .QN(net_10347), .D(net_6942), .CK(net_10647) );
INV_X4 inst_6455 ( .A(net_10013), .ZN(net_374) );
CLKBUF_X2 inst_13273 ( .A(net_13191), .Z(net_13192) );
CLKBUF_X2 inst_12635 ( .A(net_12553), .Z(net_12554) );
CLKBUF_X2 inst_11886 ( .A(net_10983), .Z(net_11805) );
AOI211_X2 inst_10283 ( .ZN(net_5956), .C2(net_5336), .A(net_3615), .B(net_3305), .C1(net_3079) );
CLKBUF_X2 inst_10659 ( .A(net_10577), .Z(net_10578) );
CLKBUF_X2 inst_12654 ( .A(net_12572), .Z(net_12573) );
CLKBUF_X2 inst_10744 ( .A(net_10662), .Z(net_10663) );
INV_X4 inst_4636 ( .ZN(net_7035), .A(net_6436) );
XNOR2_X2 inst_302 ( .B(net_9205), .ZN(net_3274), .A(net_3022) );
CLKBUF_X2 inst_15214 ( .A(net_15132), .Z(net_15133) );
CLKBUF_X2 inst_13527 ( .A(net_13445), .Z(net_13446) );
AND4_X4 inst_10318 ( .ZN(net_8258), .A1(net_8115), .A2(net_8050), .A4(net_7670), .A3(net_7616) );
SDFF_X2 inst_673 ( .SI(net_9479), .Q(net_9479), .SE(net_3073), .CK(net_14134), .D(x2707) );
NAND2_X2 inst_3585 ( .ZN(net_7395), .A2(net_7394), .A1(net_5918) );
NAND3_X2 inst_3287 ( .ZN(net_3109), .A3(net_2361), .A1(net_2050), .A2(net_1778) );
CLKBUF_X2 inst_11628 ( .A(net_10754), .Z(net_11547) );
INV_X4 inst_5892 ( .A(net_7479), .ZN(net_5790) );
XNOR2_X2 inst_211 ( .ZN(net_4935), .A(net_4399), .B(net_2384) );
OAI22_X2 inst_1151 ( .A1(net_7211), .A2(net_5134), .B2(net_5133), .ZN(net_5122), .B1(net_398) );
CLKBUF_X2 inst_14952 ( .A(net_14870), .Z(net_14871) );
CLKBUF_X2 inst_11399 ( .A(net_11317), .Z(net_11318) );
INV_X4 inst_4659 ( .A(net_7721), .ZN(net_6563) );
NAND4_X2 inst_3120 ( .A3(net_6839), .ZN(net_3600), .A2(net_3051), .A4(net_2692), .A1(net_2440) );
INV_X4 inst_5917 ( .ZN(net_4441), .A(net_587) );
INV_X4 inst_5735 ( .ZN(net_2780), .A(net_748) );
SDFF_X2 inst_561 ( .D(net_9136), .SE(net_933), .CK(net_10977), .SI(x2214), .Q(x1206) );
CLKBUF_X2 inst_13417 ( .A(net_13335), .Z(net_13336) );
CLKBUF_X2 inst_11565 ( .A(net_11483), .Z(net_11484) );
CLKBUF_X2 inst_12999 ( .A(net_12917), .Z(net_12918) );
CLKBUF_X2 inst_10903 ( .A(net_10821), .Z(net_10822) );
NOR2_X2 inst_2505 ( .ZN(net_8446), .A2(net_8445), .A1(net_8315) );
INV_X4 inst_6504 ( .A(net_10023), .ZN(net_5106) );
CLKBUF_X2 inst_12253 ( .A(net_12171), .Z(net_12172) );
CLKBUF_X2 inst_15243 ( .A(net_15161), .Z(net_15162) );
OAI221_X2 inst_1641 ( .B1(net_10423), .C1(net_7211), .ZN(net_5547), .B2(net_4477), .C2(net_4455), .A(net_3507) );
CLKBUF_X2 inst_12806 ( .A(net_12724), .Z(net_12725) );
INV_X2 inst_6945 ( .ZN(net_1905), .A(net_1904) );
INV_X2 inst_6765 ( .ZN(net_6168), .A(net_5943) );
NOR2_X2 inst_2736 ( .ZN(net_4198), .A1(net_3706), .A2(net_3705) );
INV_X2 inst_7178 ( .A(net_10472), .ZN(net_530) );
CLKBUF_X2 inst_12524 ( .A(net_12442), .Z(net_12443) );
CLKBUF_X2 inst_14620 ( .A(net_14538), .Z(net_14539) );
CLKBUF_X2 inst_11749 ( .A(net_11667), .Z(net_11668) );
DFF_X2 inst_7636 ( .D(net_6756), .QN(net_127), .CK(net_13449) );
XNOR2_X2 inst_196 ( .ZN(net_5191), .A(net_4544), .B(net_2324) );
OAI221_X2 inst_1567 ( .C1(net_10217), .C2(net_7295), .B2(net_7293), .ZN(net_7185), .B1(net_7184), .A(net_6832) );
CLKBUF_X2 inst_15161 ( .A(net_15079), .Z(net_15080) );
NAND2_X2 inst_3451 ( .A1(net_9487), .A2(net_8476), .ZN(net_8472) );
INV_X8 inst_4489 ( .ZN(net_7090), .A(net_6166) );
NOR3_X2 inst_2417 ( .ZN(net_5366), .A1(net_5365), .A3(net_5364), .A2(net_2237) );
INV_X4 inst_5523 ( .A(net_10140), .ZN(net_1243) );
CLKBUF_X2 inst_13481 ( .A(net_13399), .Z(net_13400) );
CLKBUF_X2 inst_12828 ( .A(net_12746), .Z(net_12747) );
CLKBUF_X2 inst_10637 ( .A(net_10554), .Z(net_10556) );
CLKBUF_X2 inst_14811 ( .A(net_14346), .Z(net_14730) );
DFF_X2 inst_8405 ( .Q(net_9159), .CK(net_15270), .D(x3558) );
INV_X2 inst_7155 ( .A(net_3102), .ZN(net_706) );
OAI222_X2 inst_1403 ( .B2(net_7728), .A2(net_7727), .C2(net_7726), .ZN(net_5327), .B1(net_4388), .A1(net_3671), .C1(net_1918) );
CLKBUF_X2 inst_15100 ( .A(net_15018), .Z(net_15019) );
INV_X4 inst_5606 ( .A(net_10409), .ZN(net_1493) );
CLKBUF_X2 inst_14684 ( .A(net_14602), .Z(net_14603) );
CLKBUF_X2 inst_14371 ( .A(net_13857), .Z(net_14290) );
XNOR2_X2 inst_298 ( .ZN(net_3331), .A(net_3309), .B(net_836) );
OAI211_X2 inst_2180 ( .C1(net_7209), .C2(net_6548), .A(net_6546), .ZN(net_6529), .B(net_5656) );
OAI21_X2 inst_1856 ( .ZN(net_5795), .B1(net_5794), .A(net_5382), .B2(net_1431) );
AOI22_X2 inst_9379 ( .B1(net_9993), .A1(net_6813), .A2(net_5743), .B2(net_5742), .ZN(net_5526) );
INV_X4 inst_5507 ( .ZN(net_1322), .A(net_979) );
XOR2_X2 inst_42 ( .Z(net_1472), .A(net_1417), .B(net_193) );
INV_X4 inst_6594 ( .A(net_10002), .ZN(net_319) );
CLKBUF_X2 inst_13535 ( .A(net_13435), .Z(net_13454) );
AND2_X2 inst_10521 ( .ZN(net_4565), .A1(net_4168), .A2(net_4167) );
NAND2_X2 inst_4084 ( .ZN(net_3356), .A2(net_2182), .A1(net_1471) );
OAI221_X2 inst_1479 ( .ZN(net_7639), .A(net_7549), .B1(net_3514), .C1(net_3512), .C2(net_3301), .B2(net_2723) );
CLKBUF_X2 inst_11390 ( .A(net_11280), .Z(net_11309) );
CLKBUF_X2 inst_11124 ( .A(net_11042), .Z(net_11043) );
INV_X4 inst_6180 ( .ZN(net_1403), .A(net_191) );
NAND2_X2 inst_3529 ( .A2(net_9599), .ZN(net_8119), .A1(net_8057) );
CLKBUF_X2 inst_14548 ( .A(net_14466), .Z(net_14467) );
OAI211_X2 inst_2040 ( .C2(net_8102), .B(net_8098), .ZN(net_8048), .A(net_7943), .C1(net_5801) );
XNOR2_X2 inst_437 ( .B(net_9306), .ZN(net_1043), .A(net_214) );
CLKBUF_X2 inst_10834 ( .A(net_10703), .Z(net_10753) );
CLKBUF_X2 inst_11606 ( .A(net_11159), .Z(net_11525) );
CLKBUF_X2 inst_13307 ( .A(net_13225), .Z(net_13226) );
HA_X1 inst_7327 ( .S(net_7737), .CO(net_7736), .B(net_7566), .A(net_923) );
INV_X4 inst_4742 ( .ZN(net_4844), .A(net_4439) );
DFF_X2 inst_8316 ( .QN(net_10271), .D(net_3950), .CK(net_14437) );
CLKBUF_X2 inst_14489 ( .A(net_13464), .Z(net_14408) );
INV_X4 inst_6527 ( .A(net_9728), .ZN(net_734) );
CLKBUF_X2 inst_14391 ( .A(net_14309), .Z(net_14310) );
CLKBUF_X2 inst_12782 ( .A(net_12700), .Z(net_12701) );
AND2_X4 inst_10451 ( .A1(net_10155), .ZN(net_3117), .A2(net_1756) );
AOI22_X2 inst_9425 ( .A1(net_9755), .B1(net_6834), .ZN(net_4624), .A2(net_4622), .B2(net_4621) );
INV_X4 inst_6099 ( .A(net_9614), .ZN(net_493) );
OAI221_X2 inst_1706 ( .ZN(net_4643), .B1(net_4642), .A(net_4354), .B2(net_2912), .C2(net_2911), .C1(net_831) );
CLKBUF_X2 inst_12687 ( .A(net_12430), .Z(net_12606) );
INV_X2 inst_6733 ( .ZN(net_7542), .A(net_7480) );
INV_X4 inst_4561 ( .ZN(net_8477), .A(net_8415) );
CLKBUF_X2 inst_11315 ( .A(net_11233), .Z(net_11234) );
AOI22_X2 inst_9324 ( .B1(net_9910), .A2(net_5759), .B2(net_5758), .ZN(net_5652), .A1(net_249) );
INV_X2 inst_6778 ( .ZN(net_6020), .A(net_5834) );
AOI22_X2 inst_9611 ( .A1(net_9838), .B1(net_9774), .A2(net_6413), .ZN(net_3442), .B2(net_2462) );
INV_X4 inst_6221 ( .A(net_10334), .ZN(net_640) );
OAI211_X2 inst_2220 ( .C1(net_7209), .C2(net_6501), .ZN(net_6485), .B(net_5560), .A(net_3679) );
NOR2_X2 inst_2743 ( .ZN(net_4139), .A1(net_3685), .A2(x3772) );
OAI211_X2 inst_2083 ( .C2(net_6774), .ZN(net_6765), .A(net_6392), .B(net_6126), .C1(net_469) );
CLKBUF_X2 inst_15144 ( .A(net_13767), .Z(net_15063) );
OAI221_X2 inst_1470 ( .ZN(net_7814), .B2(net_7811), .A(net_5352), .B1(net_4149), .C2(net_3520), .C1(net_3077) );
AOI221_X2 inst_9958 ( .C1(net_10499), .B1(net_10289), .C2(net_6415), .B2(net_4774), .ZN(net_4773), .A(net_4344) );
DFF_X2 inst_8019 ( .QN(net_10227), .D(net_5476), .CK(net_11738) );
OAI211_X2 inst_2247 ( .A(net_8098), .C1(net_7237), .C2(net_6501), .ZN(net_6457), .B(net_5559) );
OAI22_X2 inst_1213 ( .A1(net_7190), .A2(net_5139), .B2(net_5138), .ZN(net_5036), .B1(net_3719) );
CLKBUF_X2 inst_13517 ( .A(net_13435), .Z(net_13436) );
AOI222_X1 inst_9706 ( .B1(net_9511), .A2(net_8295), .B2(net_8294), .C2(net_8293), .ZN(net_8272), .C1(net_8210), .A1(x2826) );
NAND4_X2 inst_3072 ( .ZN(net_5253), .A2(net_4695), .A1(net_4486), .A3(net_3762), .A4(net_3462) );
DFF_X2 inst_7524 ( .QN(net_9317), .D(net_7774), .CK(net_15332) );
CLKBUF_X2 inst_12128 ( .A(net_12046), .Z(net_12047) );
CLKBUF_X2 inst_11852 ( .A(net_10655), .Z(net_11771) );
CLKBUF_X2 inst_14094 ( .A(net_11975), .Z(net_14013) );
NOR3_X2 inst_2452 ( .ZN(net_2763), .A1(net_2318), .A2(net_1591), .A3(x6531) );
CLKBUF_X2 inst_11370 ( .A(net_11288), .Z(net_11289) );
XNOR2_X2 inst_428 ( .ZN(net_2451), .B(net_1450), .A(net_1123) );
CLKBUF_X2 inst_11821 ( .A(net_11739), .Z(net_11740) );
INV_X4 inst_5786 ( .ZN(net_1380), .A(net_931) );
NAND2_X2 inst_3418 ( .ZN(net_8515), .A1(net_8458), .A2(net_8457) );
NAND2_X4 inst_3334 ( .ZN(net_8942), .A1(net_8561), .A2(net_8560) );
XNOR2_X2 inst_407 ( .ZN(net_1692), .B(net_1691), .A(net_629) );
AOI22_X2 inst_9093 ( .A1(net_9709), .A2(net_6420), .ZN(net_6399), .B2(net_5263), .B1(net_149) );
NAND2_X2 inst_3558 ( .A2(net_8919), .ZN(net_7825), .A1(net_7282) );
OAI22_X2 inst_1208 ( .A1(net_7124), .A2(net_5107), .B2(net_5105), .ZN(net_5042), .B1(net_5041) );
XNOR2_X2 inst_97 ( .B(net_8969), .ZN(net_8438), .A(net_5390) );
INV_X4 inst_5843 ( .ZN(net_1379), .A(net_1339) );
CLKBUF_X2 inst_15658 ( .A(net_14645), .Z(net_15577) );
OR2_X4 inst_775 ( .A1(net_9107), .ZN(net_3181), .A2(net_2580) );
DFF_X2 inst_8120 ( .Q(net_9738), .D(net_5148), .CK(net_14298) );
INV_X4 inst_4652 ( .A(net_9254), .ZN(net_7043) );
SDFF_X2 inst_652 ( .SI(net_9473), .Q(net_9473), .SE(net_3073), .CK(net_14653), .D(x3071) );
CLKBUF_X2 inst_15643 ( .A(net_10959), .Z(net_15562) );
DFF_X2 inst_7642 ( .D(net_6728), .QN(net_157), .CK(net_15081) );
CLKBUF_X2 inst_11102 ( .A(net_10573), .Z(net_11021) );
AOI221_X2 inst_9935 ( .B2(net_5867), .A(net_5859), .ZN(net_5834), .C1(net_5833), .C2(net_4725), .B1(x5790) );
CLKBUF_X2 inst_11812 ( .A(net_11730), .Z(net_11731) );
CLKBUF_X2 inst_14281 ( .A(net_14199), .Z(net_14200) );
SDFF_X2 inst_677 ( .SI(net_9481), .Q(net_9481), .SE(net_3073), .CK(net_12384), .D(x2589) );
CLKBUF_X2 inst_12155 ( .A(net_12073), .Z(net_12074) );
XNOR2_X2 inst_130 ( .ZN(net_7451), .B(net_7021), .A(net_6987) );
OAI221_X2 inst_1566 ( .C1(net_10216), .C2(net_7295), .B2(net_7293), .ZN(net_7187), .B1(net_7186), .A(net_6833) );
CLKBUF_X2 inst_12468 ( .A(net_12386), .Z(net_12387) );
CLKBUF_X2 inst_15124 ( .A(net_11282), .Z(net_15043) );
CLKBUF_X2 inst_10829 ( .A(net_10747), .Z(net_10748) );
DFF_X2 inst_7711 ( .Q(net_10020), .D(net_6456), .CK(net_13211) );
CLKBUF_X2 inst_14892 ( .A(net_14810), .Z(net_14811) );
OAI211_X2 inst_2242 ( .C1(net_7190), .C2(net_6480), .ZN(net_6462), .B(net_5648), .A(net_3679) );
AND2_X2 inst_10489 ( .A2(net_9600), .A1(net_8965), .ZN(net_8138) );
OAI22_X2 inst_1054 ( .B1(net_10254), .B2(net_10240), .A1(net_10239), .ZN(net_7460), .A2(net_7459) );
CLKBUF_X2 inst_11420 ( .A(net_10764), .Z(net_11339) );
CLKBUF_X2 inst_12954 ( .A(net_12872), .Z(net_12873) );
OAI22_X2 inst_972 ( .ZN(net_8815), .A1(net_8813), .B2(net_8812), .A2(net_8811), .B1(net_414) );
CLKBUF_X2 inst_15227 ( .A(net_15145), .Z(net_15146) );
OAI221_X2 inst_1671 ( .C1(net_7221), .A(net_6546), .C2(net_5520), .ZN(net_5498), .B2(net_4547), .B1(net_3255) );
CLKBUF_X2 inst_13992 ( .A(net_13853), .Z(net_13911) );
OAI21_X2 inst_1843 ( .ZN(net_6657), .B2(net_5980), .A(net_1743), .B1(net_1388) );
INV_X4 inst_4581 ( .ZN(net_8069), .A(net_8027) );
AOI21_X2 inst_10044 ( .ZN(net_7469), .A(net_7468), .B2(net_7384), .B1(net_1822) );
CLKBUF_X2 inst_13203 ( .A(net_13121), .Z(net_13122) );
CLKBUF_X2 inst_11113 ( .A(net_10907), .Z(net_11032) );
NOR2_X2 inst_2884 ( .ZN(net_4356), .A1(net_2071), .A2(net_1390) );
SDFF_X2 inst_600 ( .QN(net_9191), .D(net_9182), .SI(net_5011), .SE(net_4292), .CK(net_13531) );
CLKBUF_X2 inst_13662 ( .A(net_13580), .Z(net_13581) );
CLKBUF_X2 inst_11951 ( .A(net_11384), .Z(net_11870) );
AOI21_X2 inst_10224 ( .A(net_3988), .ZN(net_2106), .B1(net_2105), .B2(net_1855) );
INV_X4 inst_5319 ( .A(net_1815), .ZN(net_1277) );
INV_X8 inst_4498 ( .ZN(net_6133), .A(net_5298) );
OAI22_X2 inst_1194 ( .A1(net_7136), .A2(net_5151), .B2(net_5150), .ZN(net_5059), .B1(net_1821) );
CLKBUF_X2 inst_14679 ( .A(net_14597), .Z(net_14598) );
CLKBUF_X2 inst_11480 ( .A(net_11398), .Z(net_11399) );
CLKBUF_X2 inst_15392 ( .A(net_15310), .Z(net_15311) );
CLKBUF_X2 inst_12717 ( .A(net_11825), .Z(net_12636) );
CLKBUF_X2 inst_14292 ( .A(net_14210), .Z(net_14211) );
XNOR2_X2 inst_204 ( .ZN(net_4954), .A(net_4418), .B(net_2358) );
XOR2_X2 inst_49 ( .A(net_1413), .Z(net_1077), .B(net_602) );
OAI221_X2 inst_1550 ( .B2(net_7295), .C2(net_7293), .C1(net_7209), .ZN(net_7208), .A(net_6812), .B1(net_5515) );
CLKBUF_X2 inst_14353 ( .A(net_12216), .Z(net_14272) );
CLKBUF_X2 inst_14288 ( .A(net_13447), .Z(net_14207) );
OR2_X2 inst_910 ( .A2(net_5362), .ZN(net_4751), .A1(net_4170) );
CLKBUF_X2 inst_15306 ( .A(net_15224), .Z(net_15225) );
NAND2_X2 inst_4097 ( .ZN(net_2514), .A1(net_2513), .A2(net_2512) );
OR3_X4 inst_693 ( .ZN(net_6548), .A1(net_5171), .A3(net_4779), .A2(net_4625) );
CLKBUF_X2 inst_14816 ( .A(net_14734), .Z(net_14735) );
DFF_X2 inst_7586 ( .QN(net_10511), .D(net_7478), .CK(net_11154) );
AOI21_X2 inst_10134 ( .ZN(net_4252), .B2(net_3623), .B1(net_3132), .A(net_2106) );
CLKBUF_X2 inst_13080 ( .A(net_12998), .Z(net_12999) );
DFF_X1 inst_8772 ( .Q(net_10239), .D(net_4946), .CK(net_10917) );
CLKBUF_X2 inst_12494 ( .A(net_11649), .Z(net_12413) );
DFF_X2 inst_7562 ( .QN(net_10359), .D(net_7626), .CK(net_12228) );
CLKBUF_X2 inst_12344 ( .A(net_12262), .Z(net_12263) );
CLKBUF_X2 inst_11515 ( .A(net_11422), .Z(net_11434) );
AOI21_X2 inst_10119 ( .B2(net_9838), .ZN(net_4785), .A(net_4476), .B1(net_627) );
INV_X4 inst_6217 ( .A(net_10105), .ZN(net_5864) );
DFF_X2 inst_7383 ( .D(net_8658), .QN(net_268), .CK(net_13777) );
DFF_X2 inst_7401 ( .Q(net_9576), .D(net_8438), .CK(net_11507) );
OR2_X2 inst_937 ( .ZN(net_3054), .A2(net_1263), .A1(net_186) );
DFF_X2 inst_7390 ( .D(net_8651), .QN(net_265), .CK(net_13776) );
DFF_X2 inst_8303 ( .QN(net_9380), .D(net_4569), .CK(net_13111) );
CLKBUF_X2 inst_15315 ( .A(net_15233), .Z(net_15234) );
CLKBUF_X2 inst_14987 ( .A(net_13756), .Z(net_14906) );
OR2_X2 inst_908 ( .ZN(net_4692), .A2(net_4406), .A1(net_2754) );
XNOR2_X2 inst_355 ( .ZN(net_2778), .A(net_2777), .B(net_2469) );
CLKBUF_X2 inst_11690 ( .A(net_11608), .Z(net_11609) );
CLKBUF_X2 inst_13731 ( .A(net_13596), .Z(net_13650) );
AOI22_X2 inst_9259 ( .A2(net_6141), .B2(net_6140), .ZN(net_6046), .B1(net_4050), .A1(net_2573) );
AOI22_X2 inst_9227 ( .A1(net_9921), .B1(net_9822), .A2(net_6141), .B2(net_6120), .ZN(net_6084) );
XNOR2_X2 inst_218 ( .ZN(net_4681), .B(net_4446), .A(net_4445) );
INV_X4 inst_6584 ( .A(net_9846), .ZN(net_4659) );
NAND2_X2 inst_3647 ( .ZN(net_7345), .A1(net_6967), .A2(net_6681) );
CLKBUF_X2 inst_14773 ( .A(net_14516), .Z(net_14692) );
NAND2_X2 inst_3498 ( .A1(net_9548), .ZN(net_8242), .A2(net_8241) );
INV_X2 inst_6753 ( .A(net_7248), .ZN(net_6562) );
CLKBUF_X2 inst_11865 ( .A(net_11783), .Z(net_11784) );
CLKBUF_X2 inst_11098 ( .A(net_10647), .Z(net_11017) );
DFF_X2 inst_8226 ( .Q(net_10497), .D(net_4884), .CK(net_13174) );
CLKBUF_X2 inst_10706 ( .A(net_10624), .Z(net_10625) );
INV_X4 inst_6228 ( .ZN(net_7124), .A(x5722) );
NAND2_X2 inst_3693 ( .A2(net_9253), .ZN(net_6651), .A1(net_4687) );
CLKBUF_X2 inst_11309 ( .A(net_11227), .Z(net_11228) );
DFF_X2 inst_7655 ( .D(net_6695), .QN(net_187), .CK(net_12989) );
INV_X2 inst_6806 ( .ZN(net_5083), .A(net_4803) );
CLKBUF_X2 inst_14619 ( .A(net_14537), .Z(net_14538) );
CLKBUF_X2 inst_15655 ( .A(net_10750), .Z(net_15574) );
NAND2_X2 inst_3769 ( .ZN(net_5389), .A1(net_5012), .A2(net_483) );
NAND2_X2 inst_4053 ( .ZN(net_3240), .A2(net_2806), .A1(net_2062) );
OAI21_X2 inst_1747 ( .B1(net_8691), .ZN(net_8673), .B2(net_8645), .A(net_7850) );
INV_X4 inst_5236 ( .ZN(net_3985), .A(net_2301) );
AND2_X2 inst_10477 ( .A2(net_9583), .ZN(net_8769), .A1(net_1977) );
AOI22_X2 inst_9066 ( .B1(net_9686), .A1(net_6821), .A2(net_6684), .B2(net_6683), .ZN(net_6600) );
INV_X4 inst_5109 ( .A(net_2071), .ZN(net_1666) );
CLKBUF_X2 inst_11834 ( .A(net_10683), .Z(net_11753) );
INV_X4 inst_5357 ( .ZN(net_3121), .A(net_1665) );
CLKBUF_X2 inst_12992 ( .A(net_12910), .Z(net_12911) );
CLKBUF_X2 inst_11978 ( .A(net_11896), .Z(net_11897) );
CLKBUF_X2 inst_14204 ( .A(net_13192), .Z(net_14123) );
CLKBUF_X2 inst_13026 ( .A(net_12944), .Z(net_12945) );
CLKBUF_X2 inst_13352 ( .A(net_13270), .Z(net_13271) );
NAND2_X2 inst_3917 ( .A2(net_9055), .ZN(net_7965), .A1(net_470) );
CLKBUF_X2 inst_14104 ( .A(net_11786), .Z(net_14023) );
CLKBUF_X2 inst_13243 ( .A(net_13161), .Z(net_13162) );
AOI22_X2 inst_9467 ( .B1(net_9908), .A1(net_9710), .B2(net_4969), .ZN(net_3860), .A2(net_3039) );
AOI22_X2 inst_9419 ( .A1(net_10183), .A2(net_4656), .B2(net_4655), .ZN(net_4650), .B1(x5003) );
DFF_X2 inst_7601 ( .Q(net_9347), .D(net_7340), .CK(net_15299) );
CLKBUF_X2 inst_12231 ( .A(net_10559), .Z(net_12150) );
NOR2_X2 inst_2682 ( .ZN(net_4782), .A2(net_4639), .A1(net_4368) );
NOR2_X2 inst_2574 ( .ZN(net_7468), .A2(net_7384), .A1(net_4988) );
DFF_X1 inst_8517 ( .QN(net_8817), .D(net_7483), .CK(net_11780) );
CLKBUF_X2 inst_12434 ( .A(net_11318), .Z(net_12353) );
INV_X4 inst_4699 ( .ZN(net_4798), .A(net_4797) );
OAI211_X2 inst_2229 ( .C1(net_7203), .C2(net_6480), .ZN(net_6475), .B(net_5530), .A(net_3679) );
AOI21_X2 inst_10023 ( .ZN(net_8912), .A(net_7916), .B2(net_7915), .B1(net_7856) );
CLKBUF_X2 inst_11456 ( .A(net_11374), .Z(net_11375) );
INV_X4 inst_6252 ( .A(net_9182), .ZN(net_5011) );
INV_X4 inst_4749 ( .ZN(net_4477), .A(net_4369) );
OAI33_X1 inst_964 ( .A1(net_7437), .B1(net_4070), .ZN(net_3599), .B3(net_3598), .A2(net_3598), .A3(net_1959), .B2(net_936) );
CLKBUF_X2 inst_14587 ( .A(net_14505), .Z(net_14506) );
NAND2_X4 inst_3372 ( .ZN(net_3376), .A1(net_3179), .A2(net_2925) );
OAI22_X2 inst_1245 ( .A1(net_7124), .A2(net_4871), .B2(net_4870), .ZN(net_4865), .B1(net_497) );
DFF_X2 inst_7940 ( .QN(net_10231), .D(net_5630), .CK(net_15500) );
AOI21_X2 inst_10165 ( .B1(net_9531), .A(net_7649), .ZN(net_3689), .B2(net_3084) );
NOR4_X2 inst_2313 ( .A3(net_10199), .A1(net_10198), .ZN(net_7414), .A4(net_7066), .A2(net_359) );
CLKBUF_X2 inst_12560 ( .A(net_12478), .Z(net_12479) );
INV_X4 inst_6422 ( .A(net_9930), .ZN(net_676) );
CLKBUF_X2 inst_10649 ( .A(net_10561), .Z(net_10568) );
CLKBUF_X2 inst_14778 ( .A(net_14696), .Z(net_14697) );
CLKBUF_X2 inst_12660 ( .A(net_11384), .Z(net_12579) );
INV_X4 inst_5409 ( .ZN(net_2301), .A(net_1156) );
NAND2_X2 inst_3788 ( .ZN(net_6677), .A2(net_5903), .A1(net_4634) );
CLKBUF_X2 inst_12629 ( .A(net_11994), .Z(net_12548) );
CLKBUF_X2 inst_14030 ( .A(net_13948), .Z(net_13949) );
CLKBUF_X2 inst_12965 ( .A(net_12883), .Z(net_12884) );
INV_X4 inst_6114 ( .A(net_9212), .ZN(net_1750) );
NAND2_X2 inst_3663 ( .A2(net_10485), .ZN(net_6260), .A1(net_1961) );
CLKBUF_X2 inst_15359 ( .A(net_13538), .Z(net_15278) );
CLKBUF_X2 inst_11977 ( .A(net_11895), .Z(net_11896) );
INV_X4 inst_6193 ( .A(net_9835), .ZN(net_839) );
NOR2_X2 inst_3001 ( .A1(net_10430), .ZN(net_1359), .A2(net_879) );
CLKBUF_X2 inst_14111 ( .A(net_14029), .Z(net_14030) );
CLKBUF_X2 inst_13741 ( .A(net_12888), .Z(net_13660) );
NOR2_X2 inst_2818 ( .A2(net_6158), .A1(net_5331), .ZN(net_2603) );
CLKBUF_X2 inst_15526 ( .A(net_15444), .Z(net_15445) );
NOR2_X2 inst_3008 ( .A1(net_9232), .ZN(net_1397), .A2(net_320) );
INV_X4 inst_5515 ( .ZN(net_2943), .A(net_974) );
NAND3_X2 inst_3198 ( .A2(net_9386), .ZN(net_7635), .A1(net_7442), .A3(net_7441) );
INV_X4 inst_5900 ( .ZN(net_845), .A(net_600) );
DFF_X2 inst_8234 ( .Q(net_10493), .D(net_4888), .CK(net_12959) );
DFF_X2 inst_7979 ( .QN(net_10420), .D(net_5549), .CK(net_13322) );
NOR2_X2 inst_2904 ( .A2(net_8687), .A1(net_2849), .ZN(net_1626) );
AOI21_X2 inst_10075 ( .B1(net_7333), .ZN(net_5947), .A(net_5750), .B2(net_1691) );
NOR3_X2 inst_2383 ( .A2(net_8836), .A1(net_8822), .ZN(net_7810), .A3(net_7667) );
OAI221_X2 inst_1701 ( .ZN(net_5387), .C2(net_5375), .A(net_4916), .B2(net_4914), .B1(net_3610), .C1(net_3525) );
CLKBUF_X2 inst_12853 ( .A(net_10686), .Z(net_12772) );
CLKBUF_X2 inst_10640 ( .A(net_10554), .Z(net_10559) );
CLKBUF_X2 inst_13853 ( .A(net_13771), .Z(net_13772) );
AND2_X4 inst_10401 ( .ZN(net_6887), .A2(net_5937), .A1(net_5867) );
CLKBUF_X2 inst_13614 ( .A(net_13299), .Z(net_13533) );
DFF_X1 inst_8738 ( .Q(net_9137), .D(net_5730), .CK(net_10629) );
NAND2_X2 inst_4071 ( .A1(net_2674), .ZN(net_2660), .A2(net_2659) );
CLKBUF_X2 inst_13577 ( .A(net_13495), .Z(net_13496) );
CLKBUF_X2 inst_11363 ( .A(net_11281), .Z(net_11282) );
INV_X4 inst_4987 ( .ZN(net_3088), .A(net_2619) );
DFF_X2 inst_8249 ( .Q(net_10178), .D(net_4837), .CK(net_12860) );
AOI22_X2 inst_9667 ( .B2(net_10507), .A2(net_10506), .B1(net_10500), .A1(net_10499), .ZN(net_958) );
NOR2_X4 inst_2469 ( .ZN(net_8560), .A1(net_8521), .A2(net_8520) );
CLKBUF_X2 inst_12262 ( .A(net_12180), .Z(net_12181) );
AOI22_X2 inst_9287 ( .B1(net_9996), .A1(net_5743), .B2(net_5742), .ZN(net_5713), .A2(net_236) );
DFF_X2 inst_7868 ( .QN(net_10369), .D(net_6000), .CK(net_12208) );
AOI221_X2 inst_9838 ( .A(net_6889), .B2(net_6888), .C2(net_6887), .ZN(net_6880), .B1(net_5847), .C1(x5003) );
AOI22_X2 inst_9627 ( .B1(net_9997), .A2(net_4694), .ZN(net_3416), .B2(net_2468), .A1(net_230) );
AOI22_X2 inst_9163 ( .A1(net_6633), .A2(net_6404), .ZN(net_6310), .B2(net_5263), .B1(net_3107) );
CLKBUF_X2 inst_13405 ( .A(net_13070), .Z(net_13324) );
DFF_X1 inst_8593 ( .Q(net_9684), .D(net_7262), .CK(net_15746) );
CLKBUF_X2 inst_13230 ( .A(net_13101), .Z(net_13149) );
INV_X4 inst_4736 ( .ZN(net_4786), .A(net_4466) );
CLKBUF_X2 inst_14899 ( .A(net_14817), .Z(net_14818) );
INV_X2 inst_7228 ( .A(net_10139), .ZN(net_847) );
CLKBUF_X2 inst_14442 ( .A(net_14360), .Z(net_14361) );
CLKBUF_X2 inst_12503 ( .A(net_12421), .Z(net_12422) );
DFF_X1 inst_8437 ( .Q(net_9578), .D(net_8558), .CK(net_11546) );
CLKBUF_X2 inst_14761 ( .A(net_14429), .Z(net_14680) );
AOI22_X2 inst_9671 ( .A2(net_10077), .B2(net_10076), .A1(net_10068), .B1(net_10067), .ZN(net_817) );
OAI22_X2 inst_1135 ( .A1(net_7201), .A2(net_5151), .B2(net_5150), .ZN(net_5142), .B1(net_763) );
INV_X4 inst_6259 ( .A(net_9640), .ZN(net_685) );
AND4_X4 inst_10330 ( .A2(net_10373), .ZN(net_3340), .A1(net_3100), .A4(net_2259), .A3(net_956) );
INV_X2 inst_6983 ( .A(net_1770), .ZN(net_1670) );
NAND2_X2 inst_3715 ( .A1(net_5903), .ZN(net_5901), .A2(net_5900) );
CLKBUF_X2 inst_10929 ( .A(net_10821), .Z(net_10848) );
DFF_X2 inst_8333 ( .Q(net_9614), .D(net_3146), .CK(net_13547) );
CLKBUF_X2 inst_11871 ( .A(net_11789), .Z(net_11790) );
CLKBUF_X2 inst_14419 ( .A(net_11035), .Z(net_14338) );
NAND4_X2 inst_3127 ( .ZN(net_4047), .A4(net_2288), .A1(net_2282), .A3(net_1419), .A2(net_1375) );
NAND4_X2 inst_3042 ( .ZN(net_7456), .A4(net_6978), .A3(net_4715), .A1(net_4193), .A2(net_2942) );
CLKBUF_X2 inst_10945 ( .A(net_10863), .Z(net_10864) );
DFF_X1 inst_8822 ( .QN(net_10091), .D(net_2933), .CK(net_11205) );
NAND3_X2 inst_3243 ( .ZN(net_4702), .A3(net_4436), .A1(net_4435), .A2(net_2552) );
CLKBUF_X2 inst_14039 ( .A(net_13957), .Z(net_13958) );
DFF_X1 inst_8605 ( .Q(net_9891), .D(net_7238), .CK(net_13292) );
AND2_X2 inst_10564 ( .ZN(net_3502), .A1(net_3026), .A2(net_3025) );
OAI22_X2 inst_981 ( .A2(net_8962), .ZN(net_8660), .B2(net_8659), .A1(net_6288), .B1(net_6233) );
CLKBUF_X2 inst_11940 ( .A(net_11858), .Z(net_11859) );
DFF_X2 inst_7735 ( .Q(net_9998), .D(net_6212), .CK(net_12802) );
DFF_X1 inst_8815 ( .QN(net_10487), .D(net_3346), .CK(net_11130) );
OAI22_X2 inst_1266 ( .B1(net_7224), .A2(net_4842), .B2(net_4841), .ZN(net_4807), .A1(net_385) );
INV_X4 inst_6189 ( .A(net_9236), .ZN(net_2792) );
CLKBUF_X2 inst_12260 ( .A(net_11615), .Z(net_12179) );
CLKBUF_X2 inst_15056 ( .A(net_14974), .Z(net_14975) );
CLKBUF_X2 inst_12064 ( .A(net_11982), .Z(net_11983) );
OAI211_X2 inst_2094 ( .C2(net_6778), .ZN(net_6754), .A(net_6380), .B(net_6114), .C1(net_366) );
INV_X4 inst_5102 ( .ZN(net_2320), .A(net_1688) );
INV_X4 inst_4872 ( .ZN(net_3061), .A(net_3060) );
CLKBUF_X2 inst_15781 ( .A(net_15699), .Z(net_15700) );
INV_X2 inst_7216 ( .ZN(net_447), .A(x6157) );
INV_X4 inst_6287 ( .ZN(net_7203), .A(x4781) );
NAND2_X2 inst_4317 ( .ZN(net_2296), .A1(net_775), .A2(net_719) );
CLKBUF_X2 inst_13310 ( .A(net_13228), .Z(net_13229) );
INV_X4 inst_6279 ( .ZN(net_6808), .A(net_234) );
NAND2_X2 inst_3417 ( .ZN(net_8517), .A1(net_8459), .A2(net_8432) );
CLKBUF_X2 inst_13347 ( .A(net_13003), .Z(net_13266) );
INV_X2 inst_7090 ( .A(net_2007), .ZN(net_1119) );
INV_X2 inst_6794 ( .A(net_9266), .ZN(net_5417) );
CLKBUF_X2 inst_14337 ( .A(net_14255), .Z(net_14256) );
CLKBUF_X2 inst_11379 ( .A(net_10886), .Z(net_11298) );
INV_X4 inst_5406 ( .A(net_1643), .ZN(net_1600) );
CLKBUF_X2 inst_14947 ( .A(net_14865), .Z(net_14866) );
INV_X4 inst_6292 ( .A(net_9964), .ZN(net_434) );
CLKBUF_X2 inst_13959 ( .A(net_13221), .Z(net_13878) );
INV_X4 inst_5324 ( .A(net_2554), .ZN(net_1554) );
NAND2_X2 inst_3491 ( .A2(net_8873), .ZN(net_8383), .A1(net_8330) );
NOR3_X2 inst_2393 ( .ZN(net_7714), .A3(net_7577), .A1(net_7546), .A2(net_3088) );
OAI21_X2 inst_1838 ( .B1(net_8012), .ZN(net_6217), .A(net_5780), .B2(net_5769) );
XNOR2_X2 inst_71 ( .A(net_8928), .ZN(net_8696), .B(net_8390) );
AOI22_X2 inst_9414 ( .A1(net_10176), .ZN(net_4657), .A2(net_4656), .B2(net_4655), .B1(x4449) );
OAI221_X2 inst_1454 ( .ZN(net_7979), .C2(net_7799), .A(net_7796), .B2(net_7761), .B1(net_7711), .C1(net_6210) );
CLKBUF_X2 inst_14787 ( .A(net_14705), .Z(net_14706) );
AOI22_X2 inst_9438 ( .ZN(net_4300), .A1(net_4136), .A2(net_3986), .B2(net_3396), .B1(net_3176) );
AOI21_X2 inst_10114 ( .ZN(net_4559), .B1(net_4558), .B2(net_4557), .A(net_2949) );
NAND2_X2 inst_4079 ( .ZN(net_7521), .A2(net_2615), .A1(net_606) );
NAND3_X2 inst_3231 ( .ZN(net_4944), .A1(net_4943), .A3(net_4942), .A2(net_1796) );
NAND4_X2 inst_3147 ( .ZN(net_2160), .A4(net_1187), .A2(net_972), .A1(net_733), .A3(net_716) );
AOI22_X2 inst_9084 ( .A1(net_9687), .A2(net_6420), .ZN(net_6411), .B2(net_5263), .B1(net_4029) );
OAI21_X2 inst_1945 ( .ZN(net_4209), .B1(net_4070), .A(net_4011), .B2(net_3545) );
INV_X4 inst_5564 ( .A(net_10229), .ZN(net_1551) );
NOR2_X2 inst_2657 ( .A2(net_9161), .ZN(net_7530), .A1(net_4971) );
CLKBUF_X2 inst_12884 ( .A(net_11468), .Z(net_12803) );
CLKBUF_X2 inst_14407 ( .A(net_14325), .Z(net_14326) );
INV_X4 inst_5722 ( .ZN(net_1382), .A(net_1214) );
XNOR2_X2 inst_336 ( .ZN(net_2978), .A(net_2188), .B(net_2146) );
CLKBUF_X2 inst_12129 ( .A(net_12047), .Z(net_12048) );
CLKBUF_X2 inst_14581 ( .A(net_14499), .Z(net_14500) );
DFF_X2 inst_7720 ( .Q(net_9808), .D(net_6543), .CK(net_15609) );
CLKBUF_X2 inst_13239 ( .A(net_13157), .Z(net_13158) );
CLKBUF_X2 inst_13043 ( .A(net_12961), .Z(net_12962) );
CLKBUF_X2 inst_12930 ( .A(net_12254), .Z(net_12849) );
XNOR2_X2 inst_376 ( .ZN(net_2471), .A(net_2470), .B(net_2469) );
INV_X4 inst_6479 ( .ZN(net_365), .A(net_205) );
CLKBUF_X2 inst_10816 ( .A(net_10734), .Z(net_10735) );
INV_X4 inst_5157 ( .ZN(net_1800), .A(net_1578) );
OAI21_X2 inst_1939 ( .ZN(net_4291), .A(net_4120), .B2(net_3969), .B1(net_1834) );
CLKBUF_X2 inst_15356 ( .A(net_15274), .Z(net_15275) );
CLKBUF_X2 inst_14503 ( .A(net_14421), .Z(net_14422) );
NAND3_X2 inst_3268 ( .A1(net_9622), .ZN(net_4155), .A2(net_4154), .A3(net_3043) );
NOR2_X2 inst_2902 ( .A1(net_10473), .ZN(net_2754), .A2(net_1637) );
DFF_X2 inst_7844 ( .Q(net_9996), .D(net_6193), .CK(net_15666) );
CLKBUF_X2 inst_14066 ( .A(net_13984), .Z(net_13985) );
DFF_X1 inst_8726 ( .QN(net_10452), .D(net_6503), .CK(net_11085) );
CLKBUF_X2 inst_11676 ( .A(net_11594), .Z(net_11595) );
CLKBUF_X2 inst_14840 ( .A(net_12406), .Z(net_14759) );
CLKBUF_X2 inst_12167 ( .A(net_12085), .Z(net_12086) );
DFF_X1 inst_8508 ( .QN(net_10373), .D(net_7662), .CK(net_13671) );
INV_X4 inst_5174 ( .ZN(net_3170), .A(net_2279) );
CLKBUF_X2 inst_13450 ( .A(net_13368), .Z(net_13369) );
AOI22_X2 inst_9553 ( .B1(net_9969), .A2(net_6442), .ZN(net_3767), .B2(net_2541), .A1(net_1031) );
DFF_X2 inst_7856 ( .QN(net_10252), .D(net_6331), .CK(net_13922) );
CLKBUF_X2 inst_10991 ( .A(net_10909), .Z(net_10910) );
CLKBUF_X2 inst_11736 ( .A(net_11654), .Z(net_11655) );
INV_X4 inst_6299 ( .A(net_9936), .ZN(net_431) );
DFF_X2 inst_8263 ( .Q(net_10290), .D(net_4817), .CK(net_14511) );
CLKBUF_X2 inst_12627 ( .A(net_12545), .Z(net_12546) );
INV_X4 inst_5870 ( .ZN(net_6847), .A(net_5938) );
CLKBUF_X2 inst_13251 ( .A(net_13169), .Z(net_13170) );
CLKBUF_X2 inst_10852 ( .A(net_10770), .Z(net_10771) );
AOI221_X2 inst_9951 ( .B2(net_7770), .C1(net_7697), .ZN(net_5006), .A(net_4459), .B1(net_3374), .C2(net_2594) );
NAND2_X2 inst_3880 ( .ZN(net_8898), .A2(net_4027), .A1(net_4026) );
NAND4_X2 inst_3100 ( .ZN(net_4343), .A1(net_3777), .A3(net_3765), .A4(net_3584), .A2(net_3406) );
DFF_X2 inst_8359 ( .QN(net_10443), .D(net_2141), .CK(net_11112) );
INV_X4 inst_5998 ( .A(net_9832), .ZN(net_1214) );
NAND2_X2 inst_4052 ( .ZN(net_3238), .A2(net_2807), .A1(net_2661) );
DFF_X1 inst_8552 ( .Q(net_8818), .D(net_7316), .CK(net_12313) );
NAND2_X2 inst_4251 ( .A2(net_10325), .ZN(net_2043), .A1(net_931) );
INV_X8 inst_4487 ( .ZN(net_8235), .A(net_8164) );
OAI221_X2 inst_1596 ( .B1(net_10211), .C1(net_7234), .B2(net_5642), .ZN(net_5641), .C2(net_4905), .A(net_3731) );
NAND2_X2 inst_4364 ( .A2(net_10048), .ZN(net_3748), .A1(net_339) );
CLKBUF_X2 inst_15313 ( .A(net_15231), .Z(net_15232) );
CLKBUF_X2 inst_15788 ( .A(net_15706), .Z(net_15707) );
INV_X4 inst_6400 ( .A(net_10390), .ZN(net_391) );
NAND2_X2 inst_3752 ( .ZN(net_5297), .A2(net_4765), .A1(net_3866) );
INV_X2 inst_7078 ( .ZN(net_3100), .A(net_1195) );
AOI21_X2 inst_10174 ( .ZN(net_3616), .A(net_3615), .B2(net_3120), .B1(net_1979) );
OAI211_X2 inst_2265 ( .C1(net_7139), .C2(net_6542), .ZN(net_6280), .B(net_5706), .A(net_3507) );
XNOR2_X2 inst_284 ( .ZN(net_3643), .A(net_3641), .B(net_2729) );
CLKBUF_X2 inst_13494 ( .A(net_13412), .Z(net_13413) );
OAI221_X2 inst_1555 ( .C2(net_7295), .B2(net_7293), .ZN(net_7202), .B1(net_7201), .A(net_6826), .C1(net_5469) );
CLKBUF_X2 inst_13809 ( .A(net_11098), .Z(net_13728) );
OAI22_X2 inst_1293 ( .B1(net_10040), .A1(net_9941), .A2(net_4274), .B2(net_3588), .ZN(net_3587) );
INV_X2 inst_7132 ( .A(net_1074), .ZN(net_850) );
NAND2_X2 inst_3805 ( .A1(net_10074), .A2(net_4534), .ZN(net_4533) );
NOR2_X2 inst_2579 ( .A1(net_8857), .ZN(net_7080), .A2(net_7079) );
XNOR2_X2 inst_280 ( .ZN(net_3671), .B(net_3670), .A(net_3489) );
CLKBUF_X2 inst_11249 ( .A(net_10915), .Z(net_11168) );
CLKBUF_X2 inst_12668 ( .A(net_12586), .Z(net_12587) );
NAND4_X2 inst_3157 ( .A4(net_9612), .ZN(net_1792), .A1(net_1791), .A2(net_1790), .A3(net_905) );
OAI221_X2 inst_1713 ( .ZN(net_3629), .C1(net_3628), .C2(net_3559), .A(net_3558), .B1(net_3158), .B2(net_2500) );
INV_X2 inst_6970 ( .ZN(net_1730), .A(net_1065) );
INV_X4 inst_5650 ( .A(net_10353), .ZN(net_1102) );
AOI221_X2 inst_9888 ( .B1(net_9765), .B2(net_9097), .A(net_6940), .C2(net_6939), .ZN(net_6807), .C1(net_235) );
INV_X8 inst_4527 ( .A(net_9049), .ZN(net_9048) );
CLKBUF_X2 inst_11657 ( .A(net_11445), .Z(net_11576) );
AOI22_X2 inst_9532 ( .B1(net_9904), .A1(net_9706), .B2(net_4969), .ZN(net_3789), .A2(net_3039) );
NAND4_X2 inst_3137 ( .A4(net_2919), .ZN(net_2910), .A1(net_2909), .A2(net_2908), .A3(net_1032) );
CLKBUF_X2 inst_13648 ( .A(net_13566), .Z(net_13567) );
INV_X4 inst_4676 ( .ZN(net_6190), .A(net_6184) );
CLKBUF_X2 inst_11668 ( .A(net_11586), .Z(net_11587) );
CLKBUF_X2 inst_14071 ( .A(net_13989), .Z(net_13990) );
INV_X4 inst_5437 ( .ZN(net_5949), .A(net_1114) );
DFF_X2 inst_7544 ( .QN(net_9318), .D(net_7739), .CK(net_13039) );
DFF_X2 inst_8110 ( .QN(net_9850), .D(net_5080), .CK(net_14450) );
CLKBUF_X2 inst_11556 ( .A(net_11474), .Z(net_11475) );
CLKBUF_X2 inst_14789 ( .A(net_14707), .Z(net_14708) );
AND4_X2 inst_10344 ( .ZN(net_4612), .A4(net_4611), .A3(net_4332), .A2(net_3335), .A1(net_2808) );
INV_X8 inst_4496 ( .ZN(net_6774), .A(net_5445) );
HA_X1 inst_7357 ( .A(net_9276), .S(net_2458), .CO(net_2457), .B(net_1066) );
INV_X4 inst_6344 ( .ZN(net_7229), .A(x4449) );
OAI33_X1 inst_951 ( .B1(net_7557), .ZN(net_7507), .A1(net_7506), .A3(net_7505), .B2(net_7504), .A2(net_7504), .B3(net_7503) );
CLKBUF_X2 inst_12565 ( .A(net_12483), .Z(net_12484) );
INV_X4 inst_6586 ( .A(net_10042), .ZN(net_720) );
CLKBUF_X2 inst_15332 ( .A(net_15250), .Z(net_15251) );
AOI221_X2 inst_9836 ( .A(net_6889), .B2(net_6888), .C2(net_6887), .ZN(net_6882), .B1(net_5851), .C1(x5143) );
DFF_X2 inst_7727 ( .Q(net_9901), .D(net_6276), .CK(net_15059) );
CLKBUF_X2 inst_15414 ( .A(net_13370), .Z(net_15333) );
CLKBUF_X2 inst_11188 ( .A(net_10671), .Z(net_11107) );
INV_X4 inst_5831 ( .ZN(net_886), .A(net_663) );
NAND2_X2 inst_4393 ( .A2(net_10331), .A1(net_10330), .ZN(net_2704) );
AOI211_X2 inst_10268 ( .A(net_7704), .ZN(net_7703), .C2(net_7601), .C1(net_5269), .B(x3390) );
DFF_X2 inst_8299 ( .QN(net_8828), .D(net_4597), .CK(net_12850) );
CLKBUF_X2 inst_11253 ( .A(net_11122), .Z(net_11172) );
CLKBUF_X2 inst_12743 ( .A(net_12661), .Z(net_12662) );
CLKBUF_X2 inst_14780 ( .A(net_14698), .Z(net_14699) );
OAI222_X2 inst_1359 ( .A1(net_7660), .B2(net_7659), .C2(net_7658), .ZN(net_6930), .A2(net_5979), .B1(net_4430), .C1(net_1271) );
AND4_X2 inst_10345 ( .ZN(net_4263), .A2(net_3643), .A4(net_3642), .A3(net_3389), .A1(net_2994) );
DFF_X2 inst_7499 ( .D(net_8014), .QN(net_202), .CK(net_12512) );
NAND3_X2 inst_3188 ( .ZN(net_7723), .A1(net_7722), .A3(net_7721), .A2(net_7668) );
HA_X1 inst_7358 ( .CO(net_2499), .S(net_1734), .A(net_1733), .B(net_1732) );
CLKBUF_X2 inst_14522 ( .A(net_14440), .Z(net_14441) );
CLKBUF_X2 inst_11545 ( .A(net_10829), .Z(net_11464) );
DFF_X2 inst_7435 ( .QN(net_10090), .D(net_9116), .CK(net_10882) );
HA_X1 inst_7351 ( .S(net_4426), .CO(net_4425), .B(net_4202), .A(net_818) );
NAND4_X2 inst_3129 ( .ZN(net_2933), .A3(net_1991), .A4(net_1989), .A2(net_1987), .A1(net_1985) );
CLKBUF_X2 inst_12590 ( .A(net_12508), .Z(net_12509) );
INV_X4 inst_4674 ( .A(net_7658), .ZN(net_5255) );
CLKBUF_X2 inst_11328 ( .A(net_11246), .Z(net_11247) );
NAND2_X2 inst_3797 ( .ZN(net_4710), .A2(net_4598), .A1(net_950) );
XNOR2_X2 inst_100 ( .B(net_8927), .ZN(net_8409), .A(net_8270) );
INV_X4 inst_5581 ( .ZN(net_5317), .A(net_889) );
NAND2_X2 inst_4352 ( .A2(net_10334), .A1(net_7479), .ZN(net_1009) );
OR2_X2 inst_921 ( .ZN(net_3247), .A1(net_3246), .A2(net_3245) );
XNOR2_X2 inst_279 ( .ZN(net_3674), .A(net_3491), .B(net_1876) );
CLKBUF_X2 inst_14202 ( .A(net_14120), .Z(net_14121) );
CLKBUF_X2 inst_10772 ( .A(net_10690), .Z(net_10691) );
DFF_X2 inst_7618 ( .QN(net_9213), .D(net_6963), .CK(net_11833) );
DFF_X2 inst_7425 ( .QN(net_9396), .D(net_8334), .CK(net_14009) );
NAND2_X2 inst_3970 ( .A1(net_3357), .ZN(net_3334), .A2(net_2691) );
NAND2_X2 inst_3387 ( .ZN(net_8753), .A2(net_8750), .A1(net_1655) );
CLKBUF_X2 inst_11683 ( .A(net_11233), .Z(net_11602) );
CLKBUF_X2 inst_11014 ( .A(net_10932), .Z(net_10933) );
DFF_X2 inst_8271 ( .QN(net_10528), .D(net_4900), .CK(net_10574) );
XNOR2_X2 inst_81 ( .ZN(net_8630), .A(net_8588), .B(net_8261) );
CLKBUF_X2 inst_11499 ( .A(net_11417), .Z(net_11418) );
INV_X4 inst_5806 ( .ZN(net_1073), .A(net_686) );
CLKBUF_X2 inst_13424 ( .A(net_10890), .Z(net_13343) );
AOI221_X2 inst_9761 ( .B2(net_7770), .C1(net_7697), .ZN(net_7693), .A(net_7603), .B1(net_4206), .C2(net_2597) );
INV_X4 inst_6395 ( .A(net_9356), .ZN(net_5392) );
INV_X2 inst_7087 ( .ZN(net_1142), .A(net_1141) );
AOI22_X2 inst_9471 ( .B1(net_9910), .A1(net_9712), .B2(net_4969), .ZN(net_3856), .A2(net_3039) );
DFF_X1 inst_8825 ( .QN(net_9563), .D(net_3248), .CK(net_12081) );
CLKBUF_X2 inst_14411 ( .A(net_11032), .Z(net_14330) );
CLKBUF_X2 inst_12040 ( .A(net_11958), .Z(net_11959) );
OR2_X4 inst_790 ( .ZN(net_2252), .A2(net_908), .A1(net_891) );
AND2_X2 inst_10515 ( .ZN(net_4709), .A1(net_4566), .A2(net_4565) );
OAI22_X2 inst_1009 ( .ZN(net_8248), .A2(net_8247), .B2(net_8246), .A1(net_3568), .B1(net_1795) );
DFF_X2 inst_8024 ( .QN(net_10224), .D(net_5468), .CK(net_14455) );
NOR2_X2 inst_2954 ( .ZN(net_2028), .A2(net_1211), .A1(net_1005) );
AOI222_X1 inst_9711 ( .C2(net_10242), .B1(net_10241), .ZN(net_7878), .A2(net_7794), .B2(net_7611), .C1(net_7481), .A1(net_7460) );
CLKBUF_X2 inst_13217 ( .A(net_13135), .Z(net_13136) );
CLKBUF_X2 inst_12045 ( .A(net_10796), .Z(net_11964) );
CLKBUF_X2 inst_11844 ( .A(net_10661), .Z(net_11763) );
OAI211_X2 inst_2197 ( .C1(net_7198), .C2(net_6542), .ZN(net_6510), .B(net_5608), .A(net_3679) );
DFF_X2 inst_7995 ( .QN(net_10123), .D(net_5521), .CK(net_12364) );
OR2_X4 inst_733 ( .ZN(net_9056), .A2(net_8999), .A1(net_7089) );
INV_X4 inst_5885 ( .ZN(net_2090), .A(net_618) );
CLKBUF_X2 inst_13064 ( .A(net_12982), .Z(net_12983) );
OAI21_X2 inst_1959 ( .ZN(net_3938), .B2(net_3473), .A(net_3110), .B1(net_2051) );
NOR2_X2 inst_2582 ( .ZN(net_7066), .A2(net_6638), .A1(net_3747) );
XNOR2_X2 inst_142 ( .ZN(net_7302), .A(net_6662), .B(net_2323) );
CLKBUF_X2 inst_14294 ( .A(net_10808), .Z(net_14213) );
XNOR2_X2 inst_78 ( .ZN(net_8645), .B(net_8644), .A(net_8611) );
CLKBUF_X2 inst_13182 ( .A(net_12437), .Z(net_13101) );
DFF_X2 inst_8020 ( .QN(net_10435), .D(net_5481), .CK(net_13643) );
DFF_X2 inst_7896 ( .QN(net_10103), .D(net_6017), .CK(net_14799) );
NOR2_X2 inst_2813 ( .ZN(net_2644), .A1(net_2643), .A2(net_2505) );
XNOR2_X2 inst_177 ( .ZN(net_5397), .A(net_4949), .B(net_2642) );
DFF_X2 inst_7892 ( .QN(net_10098), .D(net_6022), .CK(net_15526) );
OR2_X4 inst_783 ( .A1(net_2963), .A2(net_2555), .ZN(net_2461) );
INV_X4 inst_6416 ( .A(net_9847), .ZN(net_4662) );
DFF_X2 inst_7910 ( .QN(net_10262), .D(net_5821), .CK(net_12206) );
DFF_X1 inst_8450 ( .D(net_8085), .Q(net_208), .CK(net_12916) );
INV_X4 inst_5696 ( .A(net_6321), .ZN(net_785) );
OAI21_X2 inst_2014 ( .B1(net_10254), .ZN(net_1703), .A(net_1702), .B2(net_1063) );
CLKBUF_X2 inst_14610 ( .A(net_14528), .Z(net_14529) );
MUX2_X1 inst_4471 ( .S(net_6041), .A(net_5374), .B(x6282), .Z(x366) );
INV_X4 inst_6122 ( .A(net_9316), .ZN(net_7679) );
AOI21_X2 inst_10144 ( .ZN(net_4210), .B2(net_4044), .A(net_3888), .B1(net_3390) );
SDFF_X2 inst_615 ( .QN(net_10446), .SE(net_3268), .D(net_2702), .SI(net_646), .CK(net_11095) );
CLKBUF_X2 inst_12182 ( .A(net_12100), .Z(net_12101) );
CLKBUF_X2 inst_12597 ( .A(net_12052), .Z(net_12516) );
CLKBUF_X2 inst_12821 ( .A(net_12739), .Z(net_12740) );
AOI21_X4 inst_9999 ( .B1(net_8977), .B2(net_8924), .ZN(net_7974), .A(net_3996) );
AOI22_X2 inst_9157 ( .A1(net_9756), .A2(net_6402), .ZN(net_6324), .B2(net_5263), .B1(net_192) );
DFF_X1 inst_8456 ( .Q(net_9528), .D(net_8048), .CK(net_15037) );
NOR2_X2 inst_2822 ( .ZN(net_2557), .A2(net_1762), .A1(net_1757) );
NOR2_X4 inst_2467 ( .A2(net_9113), .A1(net_9112), .ZN(net_9020) );
DFF_X2 inst_7906 ( .QN(net_9351), .D(net_5764), .CK(net_15277) );
INV_X4 inst_6176 ( .A(net_10109), .ZN(net_5854) );
NAND2_X2 inst_3843 ( .ZN(net_4550), .A2(net_4268), .A1(net_1025) );
CLKBUF_X2 inst_11583 ( .A(net_11501), .Z(net_11502) );
AND2_X2 inst_10621 ( .A1(net_9221), .ZN(net_1845), .A2(net_1238) );
AND4_X4 inst_10335 ( .A2(net_10268), .ZN(net_2960), .A4(net_1653), .A1(net_1091), .A3(net_801) );
DFF_X1 inst_8656 ( .Q(net_9761), .D(net_7246), .CK(net_12093) );
OAI211_X2 inst_2031 ( .ZN(net_8105), .C2(net_8102), .B(net_7954), .C1(net_7953), .A(net_3679) );
NAND2_X2 inst_4386 ( .ZN(net_2972), .A2(net_809), .A1(x6531) );
CLKBUF_X2 inst_13632 ( .A(net_13550), .Z(net_13551) );
CLKBUF_X2 inst_15367 ( .A(net_15285), .Z(net_15286) );
INV_X4 inst_5593 ( .ZN(net_2600), .A(net_2246) );
CLKBUF_X2 inst_14797 ( .A(net_14715), .Z(net_14716) );
CLKBUF_X2 inst_11282 ( .A(net_11200), .Z(net_11201) );
AOI211_X2 inst_10255 ( .A(net_8190), .ZN(net_8187), .C2(net_7931), .C1(net_5887), .B(net_3298) );
CLKBUF_X2 inst_11527 ( .A(net_11445), .Z(net_11446) );
DFF_X1 inst_8525 ( .Q(net_9972), .D(net_7347), .CK(net_14864) );
INV_X4 inst_4941 ( .ZN(net_3080), .A(net_2578) );
DFF_X2 inst_7835 ( .Q(net_9894), .D(net_6486), .CK(net_15425) );
INV_X2 inst_7095 ( .A(net_3173), .ZN(net_1087) );
INV_X4 inst_5133 ( .A(net_3121), .ZN(net_1875) );
AOI221_X2 inst_9986 ( .B2(net_7586), .C2(net_7584), .ZN(net_4193), .C1(net_4192), .A(net_3605), .B1(net_1871) );
XNOR2_X2 inst_338 ( .ZN(net_2976), .B(net_2490), .A(net_2336) );
INV_X4 inst_5577 ( .ZN(net_897), .A(net_896) );
NOR3_X2 inst_2412 ( .ZN(net_5382), .A3(net_4674), .A1(net_3211), .A2(net_2431) );
INV_X4 inst_4928 ( .A(net_8867), .ZN(net_2949) );
NAND2_X2 inst_4005 ( .A1(net_9606), .ZN(net_8566), .A2(net_8565) );
AND2_X4 inst_10384 ( .A2(net_9585), .ZN(net_8755), .A1(net_1428) );
INV_X4 inst_5424 ( .A(net_4168), .ZN(net_1132) );
NAND2_X2 inst_4323 ( .A2(net_10368), .ZN(net_2571), .A1(net_1361) );
OAI211_X2 inst_2214 ( .C1(net_7229), .C2(net_6501), .ZN(net_6491), .B(net_5563), .A(net_3679) );
CLKBUF_X2 inst_15212 ( .A(net_15130), .Z(net_15131) );
INV_X4 inst_6468 ( .A(net_9834), .ZN(net_581) );
AOI21_X2 inst_10018 ( .B2(net_8947), .ZN(net_8049), .A(net_7280), .B1(net_6903) );
NOR2_X4 inst_2474 ( .ZN(net_8559), .A1(net_8513), .A2(net_8512) );
CLKBUF_X2 inst_14051 ( .A(net_13969), .Z(net_13970) );
SDFF_X2 inst_579 ( .QN(net_10543), .SE(net_4896), .SI(net_4895), .D(net_3464), .CK(net_11236) );
INV_X4 inst_5247 ( .ZN(net_1454), .A(net_1453) );
NOR2_X2 inst_2495 ( .ZN(net_8579), .A2(net_8570), .A1(net_8319) );
NAND2_X2 inst_4019 ( .ZN(net_7503), .A2(net_2537), .A1(net_564) );
INV_X2 inst_6902 ( .ZN(net_2315), .A(net_2314) );
CLKBUF_X2 inst_11265 ( .A(net_11183), .Z(net_11184) );
DFF_X2 inst_7462 ( .QN(net_9639), .D(net_8121), .CK(net_15376) );
CLKBUF_X2 inst_11697 ( .A(net_11615), .Z(net_11616) );
CLKBUF_X2 inst_11219 ( .A(net_11137), .Z(net_11138) );
NAND3_X2 inst_3236 ( .A1(net_7142), .ZN(net_4721), .A2(net_1643), .A3(net_1507) );
OR3_X4 inst_698 ( .A2(net_10037), .ZN(net_7727), .A3(net_4442), .A1(net_1498) );
CLKBUF_X2 inst_15759 ( .A(net_15677), .Z(net_15678) );
CLKBUF_X2 inst_14378 ( .A(net_14296), .Z(net_14297) );
CLKBUF_X2 inst_11096 ( .A(net_11014), .Z(net_11015) );
AND2_X4 inst_10474 ( .A2(net_9249), .A1(net_9248), .ZN(net_1340) );
NAND2_X2 inst_3964 ( .A2(net_7648), .ZN(net_7525), .A1(net_3385) );
NAND2_X2 inst_3944 ( .A2(net_10232), .ZN(net_3547), .A1(net_3546) );
NAND2_X2 inst_3394 ( .A2(net_9048), .ZN(net_8699), .A1(net_8698) );
NAND2_X2 inst_3408 ( .ZN(net_8532), .A1(net_8531), .A2(net_8530) );
XNOR2_X2 inst_88 ( .A(net_8932), .ZN(net_8610), .B(net_1992) );
INV_X4 inst_5978 ( .A(net_9827), .ZN(net_732) );
INV_X4 inst_6054 ( .A(net_10070), .ZN(net_507) );
AND2_X4 inst_10397 ( .ZN(net_6684), .A2(net_5937), .A1(net_5358) );
NOR2_X2 inst_2863 ( .ZN(net_2719), .A1(net_2098), .A2(net_1180) );
AND3_X4 inst_10356 ( .ZN(net_4693), .A1(net_4692), .A3(net_4691), .A2(net_2651) );
DFF_X2 inst_8401 ( .Q(net_9158), .CK(net_11787), .D(x3565) );
CLKBUF_X2 inst_12882 ( .A(net_12800), .Z(net_12801) );
CLKBUF_X2 inst_11190 ( .A(net_10970), .Z(net_11109) );
XNOR2_X2 inst_360 ( .ZN(net_2729), .A(net_1472), .B(net_1407) );
CLKBUF_X2 inst_15565 ( .A(net_15483), .Z(net_15484) );
CLKBUF_X2 inst_14646 ( .A(net_14564), .Z(net_14565) );
NAND2_X2 inst_3897 ( .ZN(net_4081), .A2(net_3617), .A1(x6599) );
INV_X4 inst_5534 ( .ZN(net_3409), .A(net_947) );
INV_X4 inst_6604 ( .A(net_10011), .ZN(net_316) );
CLKBUF_X2 inst_11458 ( .A(net_11376), .Z(net_11377) );
CLKBUF_X2 inst_10876 ( .A(net_10586), .Z(net_10795) );
CLKBUF_X2 inst_11693 ( .A(net_11611), .Z(net_11612) );
NAND2_X2 inst_3908 ( .A2(net_10175), .ZN(net_4640), .A1(net_4015) );
NAND2_X2 inst_3754 ( .ZN(net_5273), .A1(net_5272), .A2(net_4990) );
INV_X4 inst_6160 ( .A(net_9951), .ZN(net_479) );
CLKBUF_X2 inst_12574 ( .A(net_12438), .Z(net_12493) );
INV_X2 inst_6797 ( .A(net_5950), .ZN(net_5411) );
OAI22_X2 inst_1129 ( .A1(net_7234), .A2(net_5151), .B2(net_5150), .ZN(net_5149), .B1(net_485) );
CLKBUF_X2 inst_15419 ( .A(net_15245), .Z(net_15338) );
AOI21_X2 inst_10229 ( .B1(net_2294), .ZN(net_2011), .A(net_2010), .B2(net_1316) );
OR2_X4 inst_837 ( .A2(net_9291), .A1(net_9290), .ZN(net_1057) );
INV_X4 inst_5716 ( .A(net_1401), .ZN(net_766) );
OR2_X4 inst_744 ( .A1(net_10058), .ZN(net_5895), .A2(net_5894) );
CLKBUF_X2 inst_13116 ( .A(net_13034), .Z(net_13035) );
CLKBUF_X2 inst_13375 ( .A(net_13293), .Z(net_13294) );
NAND2_X2 inst_3827 ( .ZN(net_9088), .A2(net_4178), .A1(net_4020) );
CLKBUF_X2 inst_14425 ( .A(net_12728), .Z(net_14344) );
CLKBUF_X2 inst_12385 ( .A(net_12303), .Z(net_12304) );
INV_X4 inst_6509 ( .A(net_10363), .ZN(net_931) );
INV_X4 inst_5457 ( .A(net_3409), .ZN(net_1577) );
CLKBUF_X2 inst_13492 ( .A(net_13410), .Z(net_13411) );
NAND2_X2 inst_4112 ( .A2(net_2571), .ZN(net_2359), .A1(net_1642) );
INV_X2 inst_7025 ( .A(net_2426), .ZN(net_1513) );
CLKBUF_X2 inst_14997 ( .A(net_12605), .Z(net_14916) );
DFF_X1 inst_8785 ( .QN(net_10483), .D(net_4567), .CK(net_11479) );
DFF_X2 inst_7798 ( .Q(net_9913), .D(net_6494), .CK(net_15701) );
AND2_X2 inst_10497 ( .ZN(net_6986), .A1(net_6658), .A2(net_6657) );
DFF_X2 inst_7664 ( .D(net_6758), .QN(net_125), .CK(net_15716) );
CLKBUF_X2 inst_11002 ( .A(net_10920), .Z(net_10921) );
CLKBUF_X2 inst_15487 ( .A(net_10772), .Z(net_15406) );
XNOR2_X2 inst_65 ( .ZN(net_8723), .A(net_8699), .B(net_8142) );
CLKBUF_X2 inst_12443 ( .A(net_10587), .Z(net_12362) );
SDFF_X2 inst_536 ( .D(net_9146), .SE(net_933), .CK(net_10992), .SI(x1598), .Q(x1129) );
AOI22_X2 inst_9563 ( .B1(net_9808), .A2(net_6443), .ZN(net_3756), .B2(net_2556), .A1(net_1223) );
CLKBUF_X2 inst_12711 ( .A(net_12629), .Z(net_12630) );
NAND2_X2 inst_3592 ( .A2(net_8826), .ZN(net_7327), .A1(net_6191) );
INV_X2 inst_6822 ( .ZN(net_4422), .A(net_4421) );
INV_X4 inst_5121 ( .ZN(net_1612), .A(net_1611) );
NAND2_X2 inst_3732 ( .ZN(net_6298), .A2(net_5447), .A1(net_1398) );
CLKBUF_X2 inst_14931 ( .A(net_14849), .Z(net_14850) );
CLKBUF_X2 inst_11032 ( .A(net_10950), .Z(net_10951) );
INV_X8 inst_4503 ( .ZN(net_6111), .A(net_5296) );
AOI22_X2 inst_9658 ( .A2(net_10245), .ZN(net_3155), .B2(net_1332), .B1(net_1245), .A1(net_1128) );
DFF_X2 inst_8146 ( .Q(net_10039), .D(net_5091), .CK(net_12015) );
INV_X4 inst_4907 ( .ZN(net_3060), .A(net_2201) );
OAI211_X2 inst_2027 ( .ZN(net_8376), .B(net_8375), .C2(net_8155), .C1(net_4764), .A(x1029) );
INV_X4 inst_5882 ( .ZN(net_1366), .A(net_902) );
NOR2_X2 inst_2926 ( .A1(net_10142), .ZN(net_2008), .A2(net_812) );
DFF_X2 inst_7487 ( .D(net_8067), .Q(net_214), .CK(net_15364) );
CLKBUF_X2 inst_15773 ( .A(net_13587), .Z(net_15692) );
XNOR2_X2 inst_416 ( .A(net_9619), .B(net_2928), .ZN(net_1409) );
AOI22_X2 inst_9169 ( .ZN(net_7041), .A2(net_5748), .B2(net_5747), .B1(net_4166), .A1(net_2236) );
OAI22_X2 inst_1158 ( .B1(net_9942), .A1(net_7231), .A2(net_5139), .B2(net_5138), .ZN(net_5115) );
AOI22_X2 inst_9059 ( .B1(net_9680), .A2(net_6684), .B2(net_6683), .ZN(net_6607), .A1(net_249) );
OAI21_X2 inst_1870 ( .ZN(net_5902), .B2(net_5346), .A(net_5342), .B1(net_5341) );
CLKBUF_X2 inst_13445 ( .A(net_13363), .Z(net_13364) );
CLKBUF_X2 inst_10871 ( .A(net_10574), .Z(net_10790) );
INV_X2 inst_7038 ( .ZN(net_1389), .A(net_1388) );
OAI222_X2 inst_1406 ( .B2(net_7732), .A2(net_7731), .C2(net_7730), .ZN(net_5324), .B1(net_4105), .A1(net_3251), .C1(net_1908) );
DFF_X2 inst_8396 ( .Q(net_10409), .D(net_10408), .CK(net_13672) );
INV_X4 inst_5500 ( .ZN(net_6311), .A(net_985) );
INV_X4 inst_5330 ( .A(net_6834), .ZN(net_1264) );
INV_X4 inst_5270 ( .A(net_2513), .ZN(net_1357) );
NAND2_X2 inst_4319 ( .A2(net_10140), .ZN(net_1162), .A1(net_734) );
CLKBUF_X2 inst_10943 ( .A(net_10861), .Z(net_10862) );
AOI22_X2 inst_9520 ( .A1(net_10195), .B1(net_9898), .B2(net_4969), .A2(net_4217), .ZN(net_3802) );
DFF_X1 inst_8436 ( .Q(net_9579), .D(net_8617), .CK(net_11548) );
DFF_X2 inst_8046 ( .QN(net_10311), .D(net_5572), .CK(net_14209) );
NOR3_X2 inst_2445 ( .ZN(net_3500), .A2(net_2956), .A3(net_2791), .A1(net_1591) );
CLKBUF_X2 inst_14704 ( .A(net_14622), .Z(net_14623) );
MUX2_X2 inst_4432 ( .Z(net_8058), .B(net_6379), .A(net_6347), .S(net_4448) );
CLKBUF_X2 inst_11039 ( .A(net_10957), .Z(net_10958) );
CLKBUF_X2 inst_13014 ( .A(net_11352), .Z(net_12933) );
NAND4_X2 inst_3039 ( .ZN(net_8323), .A3(net_8158), .A4(net_7911), .A2(net_6159), .A1(x813) );
INV_X4 inst_5477 ( .ZN(net_1990), .A(net_1383) );
OAI22_X2 inst_973 ( .ZN(net_8814), .A1(net_8813), .B2(net_8812), .A2(net_8810), .B1(net_528) );
CLKBUF_X2 inst_13374 ( .A(net_11340), .Z(net_13293) );
NAND4_X2 inst_3058 ( .ZN(net_5728), .A4(net_4771), .A3(net_4215), .A1(net_3833), .A2(net_3435) );
SDFF_X2 inst_461 ( .D(net_9582), .SE(net_758), .SI(net_593), .Q(net_256), .CK(net_11581) );
INV_X4 inst_6092 ( .A(net_9307), .ZN(net_1406) );
CLKBUF_X2 inst_11258 ( .A(net_10608), .Z(net_11177) );
CLKBUF_X2 inst_11884 ( .A(net_11802), .Z(net_11803) );
DFF_X2 inst_8291 ( .Q(net_10050), .D(net_4750), .CK(net_14501) );
CLKBUF_X2 inst_11771 ( .A(net_10555), .Z(net_11690) );
INV_X4 inst_6387 ( .ZN(net_4190), .A(net_158) );
OAI21_X2 inst_1973 ( .ZN(net_3038), .B1(net_3037), .A(net_2833), .B2(net_2544) );
NAND4_X2 inst_3089 ( .ZN(net_4485), .A4(net_4045), .A1(net_3809), .A2(net_3763), .A3(net_3494) );
NAND4_X2 inst_3051 ( .ZN(net_6155), .A4(net_5394), .A1(net_3840), .A3(net_3839), .A2(net_3581) );
DFF_X2 inst_8326 ( .QN(net_9437), .D(net_3649), .CK(net_12720) );
NOR2_X2 inst_2668 ( .ZN(net_4981), .A2(net_4705), .A1(net_4485) );
CLKBUF_X2 inst_15009 ( .A(net_14927), .Z(net_14928) );
OAI22_X2 inst_1122 ( .A2(net_8116), .ZN(net_5997), .B2(net_3884), .B1(net_680), .A1(net_680) );
CLKBUF_X2 inst_12170 ( .A(net_11318), .Z(net_12089) );
NAND2_X4 inst_3324 ( .A2(net_8875), .A1(net_8874), .ZN(net_8662) );
CLKBUF_X2 inst_14447 ( .A(net_14365), .Z(net_14366) );
CLKBUF_X2 inst_14238 ( .A(net_14156), .Z(net_14157) );
DFF_X2 inst_7987 ( .QN(net_10413), .D(net_5650), .CK(net_14583) );
DFF_X2 inst_7478 ( .D(net_8068), .Q(net_213), .CK(net_15367) );
INV_X4 inst_5742 ( .A(net_2287), .ZN(net_744) );
CLKBUF_X2 inst_14351 ( .A(net_14269), .Z(net_14270) );
INV_X4 inst_5775 ( .ZN(net_925), .A(net_712) );
INV_X4 inst_4808 ( .ZN(net_4227), .A(net_3606) );
INV_X4 inst_4657 ( .A(net_9264), .ZN(net_7378) );
NOR2_X2 inst_2981 ( .A1(net_10221), .ZN(net_2649), .A2(net_615) );
OAI221_X2 inst_1669 ( .B1(net_7216), .A(net_5637), .ZN(net_5500), .C2(net_4477), .B2(net_4455), .C1(net_950) );
DFF_X2 inst_7456 ( .QN(net_9640), .D(net_8189), .CK(net_15381) );
CLKBUF_X2 inst_15677 ( .A(net_13333), .Z(net_15596) );
INV_X4 inst_4998 ( .ZN(net_2854), .A(net_2200) );
CLKBUF_X2 inst_15403 ( .A(net_14879), .Z(net_15322) );
AOI22_X2 inst_9240 ( .A1(net_9925), .B1(net_9826), .B2(net_6133), .A2(net_6109), .ZN(net_6071) );
INV_X4 inst_5390 ( .ZN(net_1186), .A(net_1185) );
NAND2_X2 inst_4406 ( .A1(net_9562), .ZN(net_620), .A2(net_191) );
CLKBUF_X2 inst_12195 ( .A(net_11087), .Z(net_12114) );
INV_X4 inst_6169 ( .A(net_9437), .ZN(net_705) );
INV_X2 inst_6696 ( .ZN(net_8399), .A(net_8369) );
NAND4_X2 inst_3162 ( .A4(net_9312), .A3(net_2524), .ZN(net_1420), .A1(net_468), .A2(net_369) );
NAND2_X2 inst_3956 ( .A1(net_5480), .ZN(net_3648), .A2(net_3479) );
XNOR2_X2 inst_90 ( .A(net_8950), .ZN(net_8576), .B(net_8259) );
CLKBUF_X2 inst_14950 ( .A(net_13256), .Z(net_14869) );
CLKBUF_X2 inst_11166 ( .A(net_11084), .Z(net_11085) );
CLKBUF_X2 inst_10850 ( .A(net_10616), .Z(net_10769) );
INV_X2 inst_6858 ( .A(net_7648), .ZN(net_3553) );
DFF_X1 inst_8860 ( .Q(net_10093), .D(net_3464), .CK(net_10887) );
INV_X4 inst_4650 ( .A(net_9259), .ZN(net_6235) );
INV_X2 inst_7197 ( .A(net_9389), .ZN(net_8231) );
OAI21_X2 inst_1801 ( .B2(net_10452), .A(net_10451), .ZN(net_7334), .B1(net_7333) );
CLKBUF_X2 inst_12777 ( .A(net_12695), .Z(net_12696) );
INV_X4 inst_5093 ( .ZN(net_1739), .A(net_1738) );
DFF_X2 inst_7625 ( .QN(net_10357), .D(net_6921), .CK(net_12218) );
AOI221_X2 inst_9964 ( .C1(net_9703), .B2(net_5173), .ZN(net_4767), .A(net_4338), .C2(net_3039), .B1(net_206) );
NAND2_X2 inst_3833 ( .ZN(net_4607), .A1(net_4331), .A2(net_4320) );
OR3_X2 inst_720 ( .ZN(net_3045), .A1(net_2982), .A2(net_2565), .A3(net_186) );
OAI33_X1 inst_958 ( .ZN(net_4707), .A1(net_4290), .B3(net_3638), .B2(net_3049), .B1(net_3048), .A3(net_1884), .A2(net_1307) );
DFF_X1 inst_8457 ( .Q(net_9527), .D(net_8045), .CK(net_12766) );
NOR3_X1 inst_2460 ( .A1(net_7437), .A2(net_3908), .ZN(net_3522), .A3(net_3348) );
OAI22_X2 inst_1217 ( .A1(net_7129), .A2(net_5151), .B2(net_5150), .ZN(net_5031), .B1(net_2568) );
CLKBUF_X2 inst_12412 ( .A(net_12330), .Z(net_12331) );
AND2_X4 inst_10468 ( .A2(net_10434), .A1(net_10433), .ZN(net_2686) );
CLKBUF_X2 inst_13465 ( .A(net_13383), .Z(net_13384) );
XNOR2_X2 inst_368 ( .ZN(net_2519), .B(net_2495), .A(net_2164) );
CLKBUF_X2 inst_10832 ( .A(net_10690), .Z(net_10751) );
OAI221_X2 inst_1697 ( .B1(net_7224), .A(net_5575), .ZN(net_5458), .C1(net_5457), .C2(net_4477), .B2(net_4455) );
CLKBUF_X2 inst_14909 ( .A(net_14827), .Z(net_14828) );
CLKBUF_X2 inst_14574 ( .A(net_14492), .Z(net_14493) );
CLKBUF_X2 inst_10788 ( .A(net_10706), .Z(net_10707) );
AOI211_X2 inst_10285 ( .ZN(net_5386), .C2(net_4707), .A(net_3368), .C1(net_3300), .B(net_3166) );
INV_X2 inst_6995 ( .ZN(net_1635), .A(net_1634) );
INV_X2 inst_6938 ( .ZN(net_1920), .A(net_1919) );
INV_X2 inst_7126 ( .A(net_10435), .ZN(net_924) );
CLKBUF_X2 inst_15545 ( .A(net_11074), .Z(net_15464) );
AOI21_X2 inst_10187 ( .ZN(net_3418), .A(net_3417), .B1(net_3104), .B2(net_3103) );
INV_X4 inst_5907 ( .ZN(net_844), .A(net_594) );
NOR2_X1 inst_3027 ( .ZN(net_3070), .A1(net_3069), .A2(net_3068) );
NAND2_X2 inst_3689 ( .A2(net_9251), .A1(net_9069), .ZN(net_6937) );
DFF_X1 inst_8614 ( .Q(net_9878), .D(net_7179), .CK(net_14626) );
NAND2_X2 inst_3556 ( .A1(net_8963), .A2(net_8919), .ZN(net_7827) );
CLKBUF_X2 inst_14059 ( .A(net_13977), .Z(net_13978) );
CLKBUF_X2 inst_14016 ( .A(net_13934), .Z(net_13935) );
AOI21_X2 inst_10235 ( .A(net_9110), .B1(net_7953), .ZN(net_1705), .B2(net_1704) );
DFF_X2 inst_7480 ( .D(net_8066), .Q(net_215), .CK(net_15366) );
XNOR2_X2 inst_68 ( .ZN(net_8712), .A(net_8706), .B(net_8400) );
DFF_X1 inst_8811 ( .QN(net_10382), .D(net_3539), .CK(net_10699) );
DFF_X2 inst_8029 ( .QN(net_10226), .D(net_5456), .CK(net_11737) );
OAI21_X2 inst_1966 ( .A(net_9541), .ZN(net_3649), .B2(net_2714), .B1(net_1157) );
NAND2_X2 inst_3914 ( .ZN(net_3886), .A1(net_3885), .A2(net_3059) );
OAI22_X2 inst_1253 ( .B1(net_7213), .A2(net_4826), .B2(net_4825), .ZN(net_4821), .A1(net_422) );
CLKBUF_X2 inst_10913 ( .A(net_10734), .Z(net_10832) );
CLKBUF_X2 inst_11943 ( .A(net_11861), .Z(net_11862) );
CLKBUF_X2 inst_10689 ( .A(net_10607), .Z(net_10608) );
INV_X4 inst_4716 ( .ZN(net_8057), .A(net_7282) );
INV_X2 inst_6838 ( .ZN(net_3874), .A(net_3873) );
NOR2_X2 inst_2793 ( .A2(net_9052), .A1(net_8913), .ZN(net_3263) );
CLKBUF_X2 inst_15647 ( .A(net_15565), .Z(net_15566) );
OAI21_X2 inst_1884 ( .ZN(net_5008), .A(net_4710), .B2(net_4598), .B1(net_950) );
OAI21_X2 inst_2018 ( .ZN(net_8858), .B1(net_2675), .B2(net_2674), .A(net_2673) );
NOR3_X2 inst_2435 ( .A3(net_9039), .A2(net_7504), .A1(net_3512), .ZN(net_3478) );
INV_X4 inst_6488 ( .ZN(net_6349), .A(net_162) );
CLKBUF_X2 inst_13172 ( .A(net_12802), .Z(net_13091) );
DFF_X1 inst_8540 ( .Q(net_9962), .D(net_7368), .CK(net_14634) );
CLKBUF_X2 inst_14078 ( .A(net_13996), .Z(net_13997) );
OAI221_X2 inst_1690 ( .C1(net_7201), .B2(net_5642), .ZN(net_5470), .B1(net_5469), .C2(net_4905), .A(net_3527) );
AOI21_X2 inst_10101 ( .B2(net_10341), .ZN(net_5185), .B1(net_3668), .A(net_3487) );
INV_X4 inst_6413 ( .A(net_10010), .ZN(net_386) );
OAI221_X2 inst_1678 ( .B1(net_7213), .C1(net_5881), .ZN(net_5489), .C2(net_4477), .B2(net_4455), .A(net_3527) );
AOI221_X2 inst_9815 ( .B1(net_9776), .B2(net_9098), .ZN(net_6955), .A(net_6940), .C1(net_6939), .C2(net_246) );
INV_X4 inst_5312 ( .ZN(net_1286), .A(net_619) );
AOI22_X2 inst_9540 ( .B1(net_9809), .A1(net_9678), .A2(net_5966), .ZN(net_3781), .B2(net_2556) );
CLKBUF_X2 inst_11602 ( .A(net_10813), .Z(net_11521) );
CLKBUF_X2 inst_10839 ( .A(net_10757), .Z(net_10758) );
CLKBUF_X2 inst_15424 ( .A(net_15342), .Z(net_15343) );
CLKBUF_X2 inst_13015 ( .A(net_12933), .Z(net_12934) );
OAI22_X2 inst_1287 ( .A2(net_4095), .ZN(net_3918), .A1(net_3917), .B1(net_3916), .B2(net_2245) );
OAI211_X2 inst_2233 ( .C1(net_7211), .C2(net_6548), .ZN(net_6471), .B(net_5438), .A(net_3679) );
NAND2_X2 inst_4231 ( .A2(net_10162), .ZN(net_2538), .A1(net_1543) );
INV_X2 inst_7266 ( .A(net_8917), .ZN(net_8916) );
CLKBUF_X2 inst_14859 ( .A(net_11578), .Z(net_14778) );
CLKBUF_X2 inst_13939 ( .A(net_13857), .Z(net_13858) );
INV_X4 inst_5826 ( .A(net_7331), .ZN(net_5794) );
NAND2_X2 inst_4266 ( .A2(net_10335), .A1(net_10334), .ZN(net_2058) );
OAI22_X2 inst_1169 ( .A1(net_7226), .A2(net_5107), .B2(net_5105), .ZN(net_5095), .B1(net_5094) );
CLKBUF_X2 inst_13870 ( .A(net_10848), .Z(net_13789) );
NAND2_X2 inst_3483 ( .A2(net_8424), .ZN(net_8423), .A1(net_8241) );
INV_X4 inst_5704 ( .ZN(net_885), .A(net_777) );
AOI22_X2 inst_9440 ( .A2(net_10060), .B1(net_9925), .B2(net_6443), .A1(net_5320), .ZN(net_4278) );
DFF_X1 inst_8634 ( .Q(net_9883), .D(net_7220), .CK(net_14389) );
XNOR2_X2 inst_396 ( .ZN(net_1996), .A(net_1995), .B(net_666) );
NAND2_X2 inst_3382 ( .ZN(net_8787), .A2(net_8782), .A1(net_7847) );
CLKBUF_X2 inst_15548 ( .A(net_15466), .Z(net_15467) );
CLKBUF_X2 inst_12251 ( .A(net_12169), .Z(net_12170) );
NAND2_X4 inst_3377 ( .ZN(net_2219), .A2(net_1050), .A1(net_942) );
NOR2_X2 inst_2877 ( .A2(net_9584), .ZN(net_8779), .A1(net_1396) );
CLKBUF_X2 inst_12908 ( .A(net_11603), .Z(net_12827) );
INV_X4 inst_5128 ( .ZN(net_1832), .A(net_1599) );
CLKBUF_X2 inst_15150 ( .A(net_15068), .Z(net_15069) );
CLKBUF_X2 inst_14665 ( .A(net_13946), .Z(net_14584) );
INV_X4 inst_6514 ( .A(net_10492), .ZN(net_349) );
CLKBUF_X2 inst_11221 ( .A(net_10921), .Z(net_11140) );
DFF_X2 inst_7502 ( .Q(net_9544), .D(net_7988), .CK(net_14002) );
CLKBUF_X2 inst_14330 ( .A(net_14150), .Z(net_14249) );
CLKBUF_X2 inst_11709 ( .A(net_11627), .Z(net_11628) );
AND3_X2 inst_10371 ( .ZN(net_4963), .A2(net_4962), .A3(net_4692), .A1(net_4691) );
CLKBUF_X2 inst_11894 ( .A(net_11276), .Z(net_11813) );
CLKBUF_X2 inst_12062 ( .A(net_11980), .Z(net_11981) );
CLKBUF_X2 inst_14992 ( .A(net_10829), .Z(net_14911) );
AOI22_X2 inst_9095 ( .A1(net_9676), .A2(net_6420), .ZN(net_6397), .B2(net_5263), .B1(net_114) );
NOR2_X2 inst_2845 ( .A2(net_2886), .ZN(net_2260), .A1(net_1489) );
OAI222_X2 inst_1418 ( .B2(net_7665), .A2(net_7664), .C2(net_7663), .ZN(net_4926), .B1(net_2775), .A1(net_2278), .C1(net_1266) );
CLKBUF_X2 inst_14124 ( .A(net_14042), .Z(net_14043) );
CLKBUF_X2 inst_14499 ( .A(net_14417), .Z(net_14418) );
AOI21_X2 inst_10171 ( .ZN(net_4108), .B2(net_3467), .A(net_2557), .B1(net_1761) );
DFF_X2 inst_7760 ( .Q(net_9710), .D(net_6549), .CK(net_13271) );
OAI21_X2 inst_1740 ( .B1(net_8928), .ZN(net_8697), .B2(net_8428), .A(net_8340) );
NOR2_X2 inst_2977 ( .ZN(net_1791), .A1(net_1029), .A2(net_1028) );
INV_X4 inst_5663 ( .A(net_3261), .ZN(net_820) );
OAI22_X2 inst_1092 ( .A2(net_9064), .B2(net_6639), .ZN(net_6555), .B1(net_2125), .A1(net_1277) );
CLKBUF_X2 inst_11181 ( .A(net_10640), .Z(net_11100) );
AOI221_X2 inst_9843 ( .A(net_6889), .B2(net_6888), .C2(net_6887), .ZN(net_6875), .B1(net_5837), .C1(x5901) );
DFF_X2 inst_7492 ( .Q(net_10194), .D(net_8009), .CK(net_15169) );
CLKBUF_X2 inst_11176 ( .A(net_11094), .Z(net_11095) );
DFF_X2 inst_7822 ( .Q(net_9653), .D(net_6270), .CK(net_11823) );
INV_X4 inst_4836 ( .A(net_7649), .ZN(net_3342) );
OAI21_X2 inst_2001 ( .ZN(net_2217), .B1(net_2216), .A(net_1709), .B2(net_1424) );
CLKBUF_X2 inst_11784 ( .A(net_10821), .Z(net_11703) );
CLKBUF_X2 inst_15729 ( .A(net_15647), .Z(net_15648) );
AOI21_X2 inst_10011 ( .ZN(net_8637), .A(net_8635), .B2(net_8593), .B1(net_7754) );
AND4_X4 inst_10321 ( .ZN(net_4487), .A4(net_4058), .A1(net_3760), .A2(net_3738), .A3(net_3410) );
OAI221_X2 inst_1657 ( .C1(net_7209), .B2(net_5642), .ZN(net_5516), .B1(net_5515), .C2(net_4905), .A(net_3731) );
CLKBUF_X2 inst_14231 ( .A(net_14149), .Z(net_14150) );
CLKBUF_X2 inst_14385 ( .A(net_11200), .Z(net_14304) );
CLKBUF_X2 inst_12982 ( .A(net_12900), .Z(net_12901) );
CLKBUF_X2 inst_15570 ( .A(net_15488), .Z(net_15489) );
AOI21_X2 inst_10085 ( .ZN(net_5788), .A(net_5361), .B2(net_5280), .B1(net_2518) );
OAI211_X2 inst_2077 ( .C2(net_6778), .ZN(net_6771), .A(net_6398), .B(net_6132), .C1(net_350) );
CLKBUF_X2 inst_14473 ( .A(net_14391), .Z(net_14392) );
CLKBUF_X2 inst_12729 ( .A(net_12647), .Z(net_12648) );
CLKBUF_X2 inst_11356 ( .A(net_11274), .Z(net_11275) );
DFF_X2 inst_8078 ( .QN(net_10468), .D(net_5309), .CK(net_11449) );
DFF_X2 inst_7780 ( .Q(net_9794), .D(net_6520), .CK(net_14613) );
INV_X4 inst_4592 ( .ZN(net_7894), .A(net_7893) );
CLKBUF_X2 inst_15696 ( .A(net_11651), .Z(net_15615) );
XNOR2_X1 inst_451 ( .ZN(net_7042), .A(net_7041), .B(net_2350) );
INV_X4 inst_5478 ( .ZN(net_2617), .A(net_1004) );
OAI211_X2 inst_2166 ( .C1(net_7231), .C2(net_6548), .ZN(net_6544), .B(net_5671), .A(net_3679) );
CLKBUF_X2 inst_13704 ( .A(net_12474), .Z(net_13623) );
CLKBUF_X2 inst_14486 ( .A(net_14404), .Z(net_14405) );
CLKBUF_X2 inst_13930 ( .A(net_11205), .Z(net_13849) );
CLKBUF_X2 inst_15377 ( .A(net_15295), .Z(net_15296) );
INV_X2 inst_6656 ( .A(net_9436), .ZN(net_8492) );
AOI221_X2 inst_9910 ( .B1(net_9775), .B2(net_9098), .A(net_6940), .C1(net_6939), .ZN(net_6687), .C2(net_245) );
CLKBUF_X2 inst_12179 ( .A(net_11754), .Z(net_12098) );
OR2_X4 inst_797 ( .A1(net_10472), .ZN(net_2422), .A2(net_1096) );
OAI221_X2 inst_1495 ( .B1(net_10413), .C2(net_9063), .B2(net_9056), .ZN(net_7368), .C1(net_7190), .A(net_6989) );
INV_X4 inst_5546 ( .ZN(net_937), .A(net_936) );
INV_X4 inst_5051 ( .A(net_4050), .ZN(net_1889) );
DFF_X2 inst_7471 ( .Q(net_9525), .D(net_8044), .CK(net_14967) );
INV_X2 inst_7221 ( .ZN(net_432), .A(net_180) );
AOI22_X2 inst_9310 ( .B1(net_9715), .A2(net_5755), .B2(net_5754), .ZN(net_5667), .A1(net_252) );
NOR2_X1 inst_3032 ( .A1(net_2972), .ZN(net_2541), .A2(net_2540) );
INV_X4 inst_5295 ( .A(net_1345), .ZN(net_1308) );
NAND2_X2 inst_3657 ( .A1(net_9258), .ZN(net_6650), .A2(net_6234) );
DFF_X1 inst_8882 ( .Q(net_90), .CK(net_13587), .D(x3534) );
INV_X2 inst_7319 ( .A(net_9108), .ZN(net_9107) );
INV_X2 inst_6896 ( .ZN(net_2586), .A(net_2585) );
CLKBUF_X2 inst_14529 ( .A(net_14447), .Z(net_14448) );
CLKBUF_X2 inst_12069 ( .A(net_11987), .Z(net_11988) );
OAI21_X2 inst_1998 ( .ZN(net_2467), .A(net_2466), .B1(net_2465), .B2(net_930) );
INV_X2 inst_6856 ( .ZN(net_3368), .A(net_3367) );
CLKBUF_X2 inst_14699 ( .A(net_14617), .Z(net_14618) );
CLKBUF_X2 inst_13195 ( .A(net_13113), .Z(net_13114) );
INV_X2 inst_6787 ( .A(net_9257), .ZN(net_5803) );
NAND3_X2 inst_3302 ( .ZN(net_2194), .A2(net_2193), .A3(net_2192), .A1(net_1020) );
CLKBUF_X2 inst_11157 ( .A(net_11075), .Z(net_11076) );
NOR2_X2 inst_2870 ( .A1(net_2051), .ZN(net_2025), .A2(net_1602) );
NAND2_X2 inst_3583 ( .A2(net_10347), .ZN(net_7403), .A1(net_1351) );
CLKBUF_X2 inst_13242 ( .A(net_12911), .Z(net_13161) );
DFF_X1 inst_8446 ( .Q(net_9116), .D(net_8161), .CK(net_14126) );
CLKBUF_X2 inst_14902 ( .A(net_14820), .Z(net_14821) );
INV_X4 inst_4933 ( .A(net_4719), .ZN(net_3069) );
OAI22_X2 inst_1115 ( .B2(net_8117), .ZN(net_5428), .A1(net_4995), .B1(net_1665), .A2(net_1664) );
INV_X4 inst_6234 ( .A(net_10048), .ZN(net_599) );
OR2_X2 inst_874 ( .A1(net_10188), .ZN(net_6975), .A2(net_6974) );
NOR2_X2 inst_2976 ( .ZN(net_1368), .A2(net_1031), .A1(net_851) );
OAI22_X2 inst_1021 ( .A2(net_8036), .B2(net_8018), .ZN(net_8017), .A1(net_2123), .B1(net_2122) );
OAI221_X2 inst_1681 ( .C1(net_7201), .B2(net_5591), .ZN(net_5485), .B1(net_5484), .C2(net_4902), .A(net_3507) );
AOI21_X2 inst_10222 ( .ZN(net_2802), .B1(net_2773), .B2(net_2047), .A(net_1160) );
AOI22_X2 inst_9140 ( .A1(net_9737), .A2(net_6404), .ZN(net_6346), .B2(net_5263), .B1(net_914) );
NAND2_X2 inst_4204 ( .ZN(net_2540), .A2(net_1779), .A1(x6445) );
CLKBUF_X2 inst_12095 ( .A(net_12013), .Z(net_12014) );
AOI22_X2 inst_9173 ( .A1(net_9870), .B1(net_9771), .B2(net_8041), .ZN(net_6145), .A2(net_6141) );
OAI221_X2 inst_1652 ( .C1(net_10419), .B1(net_7129), .ZN(net_5534), .C2(net_4477), .B2(net_4455), .A(net_3507) );
AOI22_X2 inst_9391 ( .B1(net_9903), .A1(net_5759), .B2(net_5758), .ZN(net_5422), .A2(net_242) );
INV_X4 inst_4827 ( .ZN(net_3679), .A(net_3298) );
CLKBUF_X2 inst_15576 ( .A(net_15494), .Z(net_15495) );
SDFF_X2 inst_572 ( .D(net_9134), .SE(net_933), .CK(net_10951), .SI(x2333), .Q(x1223) );
OAI221_X2 inst_1622 ( .C1(net_10319), .B1(net_7297), .C2(net_5591), .ZN(net_5585), .B2(net_4902), .A(net_3507) );
CLKBUF_X2 inst_13965 ( .A(net_13883), .Z(net_13884) );
CLKBUF_X2 inst_12699 ( .A(net_12617), .Z(net_12618) );
CLKBUF_X2 inst_12392 ( .A(net_12310), .Z(net_12311) );
OAI21_X2 inst_1735 ( .ZN(net_8725), .B2(net_8703), .B1(net_8691), .A(net_7849) );
CLKBUF_X2 inst_15062 ( .A(net_14980), .Z(net_14981) );
INV_X4 inst_5036 ( .ZN(net_2230), .A(net_1263) );
XNOR2_X2 inst_257 ( .ZN(net_4064), .A(net_3854), .B(net_2095) );
OAI211_X2 inst_2050 ( .C2(net_10276), .B(net_8817), .ZN(net_7838), .A(net_7763), .C1(net_6056) );
AOI22_X2 inst_9516 ( .B1(net_10299), .A1(net_9699), .B2(net_4774), .ZN(net_3806), .A2(net_3039) );
CLKBUF_X2 inst_12971 ( .A(net_12030), .Z(net_12890) );
INV_X4 inst_5458 ( .ZN(net_1060), .A(net_1059) );
INV_X4 inst_4555 ( .ZN(net_8549), .A(net_8514) );
SDFF_X2 inst_485 ( .SE(net_9540), .SI(net_8224), .Q(net_282), .D(net_282), .CK(net_12712) );
CLKBUF_X2 inst_10684 ( .A(net_10602), .Z(net_10603) );
DFF_X1 inst_8681 ( .D(net_6738), .Q(net_149), .CK(net_15104) );
CLKBUF_X2 inst_14655 ( .A(net_12643), .Z(net_14574) );
OAI22_X2 inst_1189 ( .A1(net_7127), .A2(net_5151), .B2(net_5150), .ZN(net_5065), .B1(net_1278) );
OAI22_X2 inst_1205 ( .A1(net_7241), .A2(net_5139), .B2(net_5138), .ZN(net_5046), .B1(net_1865) );
CLKBUF_X2 inst_15762 ( .A(net_15680), .Z(net_15681) );
NOR4_X1 inst_2360 ( .ZN(net_7383), .A4(net_6840), .A2(net_3911), .A3(net_3522), .A1(x3390) );
CLKBUF_X2 inst_11052 ( .A(net_10679), .Z(net_10971) );
INV_X4 inst_5085 ( .ZN(net_2501), .A(net_1789) );
CLKBUF_X2 inst_11048 ( .A(net_10827), .Z(net_10967) );
XOR2_X2 inst_33 ( .A(net_9349), .Z(net_1985), .B(net_1984) );
OAI211_X2 inst_2107 ( .C2(net_6774), .ZN(net_6741), .A(net_6368), .B(net_6099), .C1(net_514) );
CLKBUF_X2 inst_12756 ( .A(net_12674), .Z(net_12675) );
XNOR2_X2 inst_232 ( .ZN(net_4314), .A(net_4167), .B(net_1900) );
INV_X4 inst_6253 ( .A(net_9535), .ZN(net_1158) );
DFF_X2 inst_8310 ( .Q(net_9151), .D(net_4288), .CK(net_11308) );
DFF_X2 inst_7575 ( .QN(net_10371), .D(net_7539), .CK(net_12225) );
CLKBUF_X2 inst_15012 ( .A(net_10785), .Z(net_14931) );
DFF_X1 inst_8641 ( .Q(net_9679), .D(net_7269), .CK(net_15552) );
INV_X4 inst_4628 ( .A(net_7519), .ZN(net_7374) );
CLKBUF_X2 inst_14409 ( .A(net_14327), .Z(net_14328) );
NAND2_X2 inst_3794 ( .A2(net_9082), .ZN(net_4728), .A1(net_1384) );
AOI22_X2 inst_9648 ( .A1(net_9568), .B2(net_2849), .ZN(net_2454), .A2(net_1124), .B1(net_192) );
INV_X2 inst_6929 ( .A(net_3202), .ZN(net_1946) );
CLKBUF_X2 inst_14463 ( .A(net_14381), .Z(net_14382) );
NAND2_X2 inst_3716 ( .ZN(net_6013), .A2(net_5824), .A1(net_1589) );
XNOR2_X2 inst_253 ( .ZN(net_4107), .A(net_3472), .B(net_2027) );
AOI22_X2 inst_9608 ( .B1(net_9779), .A2(net_6413), .ZN(net_3445), .B2(net_2462), .A1(net_632) );
DFF_X2 inst_7730 ( .Q(net_9900), .D(net_6432), .CK(net_15056) );
CLKBUF_X2 inst_14080 ( .A(net_13998), .Z(net_13999) );
CLKBUF_X2 inst_13945 ( .A(net_11438), .Z(net_13864) );
NAND2_X2 inst_3652 ( .A2(net_6663), .ZN(net_6662), .A1(net_2655) );
SDFF_X2 inst_589 ( .Q(net_9253), .SE(net_4589), .D(net_136), .SI(net_102), .CK(net_12555) );
INV_X4 inst_5229 ( .A(net_1491), .ZN(net_1490) );
CLKBUF_X2 inst_12428 ( .A(net_12346), .Z(net_12347) );
INV_X4 inst_4868 ( .ZN(net_8899), .A(net_3932) );
CLKBUF_X2 inst_14513 ( .A(net_14431), .Z(net_14432) );
CLKBUF_X2 inst_11969 ( .A(net_11887), .Z(net_11888) );
AOI21_X2 inst_10176 ( .A(net_3748), .ZN(net_3609), .B2(net_2968), .B1(net_1073) );
INV_X4 inst_5043 ( .A(net_6047), .ZN(net_1915) );
NAND2_X2 inst_4273 ( .A2(net_10145), .ZN(net_4553), .A1(net_1213) );
AOI221_X2 inst_9829 ( .B1(net_9869), .B2(net_9101), .A(net_6945), .C1(net_6944), .ZN(net_6915), .C2(net_240) );
CLKBUF_X2 inst_13751 ( .A(net_13669), .Z(net_13670) );
AOI221_X2 inst_9822 ( .B1(net_9766), .B2(net_9098), .A(net_6940), .C1(net_6939), .ZN(net_6929), .C2(net_236) );
INV_X2 inst_6907 ( .A(net_3602), .ZN(net_2590) );
AOI22_X2 inst_9331 ( .B1(net_9793), .A1(net_6834), .A2(net_5766), .B2(net_5765), .ZN(net_5621) );
SDFF_X2 inst_602 ( .SE(net_4040), .SI(net_4039), .CK(net_13472), .Q(x555), .D(x555) );
XOR2_X1 inst_59 ( .B(net_1403), .Z(net_1124), .A(net_192) );
OAI21_X2 inst_1877 ( .ZN(net_5900), .B2(net_5343), .A(net_5342), .B1(net_5341) );
NOR3_X2 inst_2367 ( .ZN(net_8553), .A1(net_8504), .A3(net_8411), .A2(net_8321) );
AOI22_X2 inst_9182 ( .A1(net_9872), .B1(net_9773), .A2(net_8042), .ZN(net_6134), .B2(net_6133) );
XNOR2_X2 inst_135 ( .ZN(net_7402), .A(net_7080), .B(net_2333) );
AND2_X2 inst_10533 ( .ZN(net_4156), .A1(net_3855), .A2(net_3854) );
AOI21_X2 inst_10091 ( .B1(net_10175), .A(net_6679), .ZN(net_5774), .B2(net_5200) );
NAND3_X2 inst_3256 ( .ZN(net_4503), .A3(net_4063), .A2(net_3551), .A1(net_3436) );
CLKBUF_X2 inst_12867 ( .A(net_12785), .Z(net_12786) );
CLKBUF_X2 inst_11711 ( .A(net_11629), .Z(net_11630) );
AOI22_X2 inst_9050 ( .B1(net_9674), .A1(net_6684), .B2(net_6683), .ZN(net_6672), .A2(net_243) );
DFF_X2 inst_7673 ( .D(net_6751), .QN(net_130), .CK(net_14241) );
CLKBUF_X2 inst_15715 ( .A(net_11253), .Z(net_15634) );
OAI21_X2 inst_1865 ( .ZN(net_5914), .A(net_5348), .B1(net_5347), .B2(net_5343) );
CLKBUF_X2 inst_11960 ( .A(net_11878), .Z(net_11879) );
INV_X4 inst_6390 ( .A(net_9732), .ZN(net_555) );
XOR2_X2 inst_37 ( .B(net_9155), .A(net_9154), .Z(net_1725) );
OAI221_X2 inst_1664 ( .C1(net_7201), .C2(net_5520), .ZN(net_5505), .B2(net_4547), .A(net_3731), .B1(net_2794) );
AOI21_X2 inst_10037 ( .A(net_8122), .ZN(net_7755), .B2(net_7637), .B1(net_2970) );
OAI221_X2 inst_1447 ( .ZN(net_8193), .B2(net_8192), .B1(net_8135), .A(net_8134), .C2(net_8119), .C1(net_7994) );
AOI22_X2 inst_9321 ( .B1(net_9725), .A2(net_5755), .B2(net_5754), .ZN(net_5655), .A1(net_262) );
NAND4_X2 inst_3117 ( .A1(net_10057), .A2(net_9958), .ZN(net_4128), .A4(net_3476), .A3(net_2113) );
INV_X4 inst_6072 ( .A(net_8828), .ZN(net_1706) );
NAND2_X2 inst_3770 ( .ZN(net_5278), .A2(net_4511), .A1(net_2799) );
CLKBUF_X2 inst_14881 ( .A(net_12942), .Z(net_14800) );
DFF_X2 inst_8157 ( .QN(net_9938), .D(net_5068), .CK(net_13705) );
AOI22_X2 inst_9601 ( .ZN(net_3959), .B2(net_3234), .B1(net_2880), .A2(net_2485), .A1(net_2484) );
CLKBUF_X2 inst_13863 ( .A(net_13781), .Z(net_13782) );
NOR2_X2 inst_2709 ( .A2(net_4560), .ZN(net_4506), .A1(net_3687) );
XNOR2_X2 inst_224 ( .ZN(net_4541), .A(net_4390), .B(net_205) );
CLKBUF_X2 inst_14756 ( .A(net_11999), .Z(net_14675) );
CLKBUF_X2 inst_14003 ( .A(net_11635), .Z(net_13922) );
AOI22_X2 inst_9661 ( .B2(net_10509), .A2(net_10508), .B1(net_10495), .A1(net_10494), .ZN(net_1052) );
INV_X4 inst_4730 ( .A(net_7732), .ZN(net_4594) );
NAND2_X2 inst_3635 ( .A1(net_10401), .ZN(net_6979), .A2(net_6970) );
INV_X4 inst_5399 ( .ZN(net_1167), .A(net_1166) );
NAND4_X2 inst_3075 ( .ZN(net_5169), .A1(net_5168), .A2(net_5167), .A4(net_5166), .A3(net_685) );
INV_X4 inst_5058 ( .ZN(net_2601), .A(net_1875) );
NOR2_X2 inst_2800 ( .ZN(net_3509), .A2(net_2854), .A1(net_1528) );
AOI22_X2 inst_9487 ( .B1(net_9785), .A1(net_9718), .ZN(net_3836), .A2(net_3039), .B2(net_2462) );
CLKBUF_X2 inst_14297 ( .A(net_14215), .Z(net_14216) );
NOR3_X2 inst_2406 ( .A1(net_7345), .A3(net_7343), .ZN(net_7147), .A2(net_7146) );
OR2_X4 inst_766 ( .ZN(net_4618), .A1(net_4324), .A2(net_4220) );
CLKBUF_X2 inst_14879 ( .A(net_14797), .Z(net_14798) );
DFF_X1 inst_8796 ( .QN(net_10174), .D(net_4008), .CK(net_10864) );
NAND3_X2 inst_3270 ( .A3(net_9037), .ZN(net_4148), .A1(net_4147), .A2(net_957) );
OAI21_X2 inst_1908 ( .B2(net_10384), .ZN(net_4763), .B1(net_4009), .A(x3733) );
NAND3_X2 inst_3273 ( .A3(net_10138), .ZN(net_4142), .A1(net_4141), .A2(net_847) );
OR2_X4 inst_801 ( .ZN(net_2149), .A2(net_1385), .A1(net_1381) );
AND2_X2 inst_10617 ( .ZN(net_2511), .A2(net_1814), .A1(net_722) );
AOI221_X2 inst_9943 ( .ZN(net_5338), .C2(net_5337), .B2(net_5337), .A(net_4643), .B1(net_3096), .C1(net_3082) );
INV_X4 inst_6139 ( .ZN(net_1978), .A(net_123) );
OR2_X2 inst_870 ( .ZN(net_7487), .A2(net_7486), .A1(net_7146) );
CLKBUF_X2 inst_12544 ( .A(net_12462), .Z(net_12463) );
CLKBUF_X2 inst_14282 ( .A(net_11493), .Z(net_14201) );
AOI22_X2 inst_9660 ( .B2(net_10194), .A2(net_10193), .B1(net_10186), .A1(net_10185), .ZN(net_1053) );
XOR2_X2 inst_11 ( .Z(net_3932), .A(net_2930), .B(net_2929) );
CLKBUF_X2 inst_15537 ( .A(net_15455), .Z(net_15456) );
INV_X4 inst_6552 ( .A(net_10501), .ZN(net_332) );
CLKBUF_X2 inst_15344 ( .A(net_15262), .Z(net_15263) );
OAI221_X2 inst_1619 ( .C1(net_10316), .B1(net_7234), .C2(net_5591), .ZN(net_5590), .B2(net_4902), .A(net_3731) );
NAND4_X2 inst_3110 ( .A2(net_9243), .ZN(net_4290), .A4(net_3639), .A3(net_2605), .A1(net_2279) );
XNOR2_X2 inst_441 ( .ZN(net_926), .A(net_218), .B(net_195) );
CLKBUF_X2 inst_13468 ( .A(net_13386), .Z(net_13387) );
DFF_X2 inst_7688 ( .Q(net_10508), .D(net_6578), .CK(net_14557) );
OAI211_X2 inst_2276 ( .C1(net_7136), .C2(net_6548), .ZN(net_6224), .B(net_5756), .A(net_3679) );
DFF_X1 inst_8425 ( .Q(net_9585), .D(net_8733), .CK(net_13819) );
INV_X4 inst_6201 ( .A(net_9978), .ZN(net_469) );
CLKBUF_X2 inst_11414 ( .A(net_11332), .Z(net_11333) );
INV_X4 inst_5228 ( .ZN(net_1804), .A(net_1491) );
OAI211_X2 inst_2301 ( .ZN(net_7648), .B(net_5284), .A(net_5283), .C2(net_3123), .C1(net_183) );
OR2_X4 inst_808 ( .A2(net_9344), .ZN(net_2071), .A1(net_1383) );
DFF_X2 inst_8202 ( .Q(net_9750), .D(net_5147), .CK(net_12873) );
SDFF_X2 inst_557 ( .SI(net_9360), .Q(net_9360), .D(net_9158), .SE(net_7248), .CK(net_15258) );
CLKBUF_X2 inst_13639 ( .A(net_10905), .Z(net_13558) );
NAND2_X2 inst_3859 ( .ZN(net_7663), .A2(net_4169), .A1(net_601) );
AOI222_X1 inst_9683 ( .B1(net_9511), .A2(net_8310), .B2(net_8309), .C2(net_8308), .ZN(net_8304), .C1(net_8194), .A1(x2333) );
CLKBUF_X2 inst_14300 ( .A(net_14218), .Z(net_14219) );
CLKBUF_X2 inst_11154 ( .A(net_11072), .Z(net_11073) );
OAI222_X2 inst_1383 ( .B1(net_7732), .A2(net_7731), .C2(net_7730), .ZN(net_6002), .B2(net_5191), .A1(net_3993), .C1(net_1873) );
NAND3_X2 inst_3279 ( .ZN(net_4196), .A1(net_4047), .A3(net_4046), .A2(net_3556) );
OR2_X4 inst_823 ( .A1(net_10471), .ZN(net_2060), .A2(net_1111) );
OAI221_X2 inst_1461 ( .C1(net_9092), .B2(net_7974), .C2(net_7973), .ZN(net_7962), .A(net_7961), .B1(net_1883) );
DFF_X1 inst_8809 ( .QN(net_10489), .D(net_3609), .CK(net_11158) );
INV_X4 inst_6153 ( .A(net_9997), .ZN(net_481) );
NOR2_X2 inst_2838 ( .A1(net_2731), .ZN(net_2342), .A2(net_1635) );
NAND2_X2 inst_3773 ( .A1(net_8864), .ZN(net_4792), .A2(net_4791) );
NAND2_X2 inst_3423 ( .A2(net_9433), .ZN(net_8510), .A1(net_7363) );
NOR2_X2 inst_2833 ( .ZN(net_2760), .A2(net_2739), .A1(net_2101) );
CLKBUF_X2 inst_15349 ( .A(net_15267), .Z(net_15268) );
INV_X4 inst_4767 ( .ZN(net_5682), .A(net_4173) );
OAI211_X2 inst_2042 ( .C2(net_8102), .ZN(net_8039), .A(net_7978), .B(net_3507), .C1(net_3036) );
AND2_X2 inst_10608 ( .A1(net_4024), .ZN(net_2664), .A2(net_1977) );
DFF_X2 inst_8383 ( .QN(net_9660), .D(net_9659), .CK(net_11165) );
DFF_X2 inst_8248 ( .Q(net_10176), .D(net_4839), .CK(net_12864) );
CLKBUF_X2 inst_13154 ( .A(net_11887), .Z(net_13073) );
INV_X4 inst_5620 ( .A(net_2780), .ZN(net_1145) );
CLKBUF_X2 inst_11409 ( .A(net_11327), .Z(net_11328) );
INV_X2 inst_7104 ( .ZN(net_1026), .A(net_1025) );
CLKBUF_X2 inst_15503 ( .A(net_13575), .Z(net_15422) );
CLKBUF_X2 inst_13361 ( .A(net_12296), .Z(net_13280) );
DFF_X2 inst_7746 ( .QN(net_10461), .D(net_6285), .CK(net_13659) );
INV_X4 inst_5156 ( .ZN(net_2095), .A(net_1579) );
CLKBUF_X2 inst_15383 ( .A(net_15301), .Z(net_15302) );
CLKBUF_X2 inst_10758 ( .A(net_10544), .Z(net_10677) );
INV_X4 inst_6107 ( .A(net_10144), .ZN(net_677) );
AOI221_X2 inst_9976 ( .B1(net_10045), .C1(net_9816), .B2(net_5174), .ZN(net_4384), .A(net_3946), .C2(net_2556) );
DFF_X2 inst_8342 ( .QN(net_9185), .D(net_2787), .CK(net_13543) );
NOR2_X2 inst_2796 ( .A1(net_9108), .ZN(net_3139), .A2(net_2924) );
CLKBUF_X2 inst_14084 ( .A(net_12786), .Z(net_14003) );
AND2_X2 inst_10587 ( .ZN(net_3010), .A2(net_2459), .A1(net_760) );
NOR2_X2 inst_2729 ( .ZN(net_4269), .A2(net_3959), .A1(net_2045) );
OAI222_X2 inst_1413 ( .B2(net_7732), .A2(net_7731), .C2(net_7730), .ZN(net_5306), .B1(net_3957), .A1(net_2529), .C1(net_1941) );
DFF_X2 inst_8364 ( .QN(net_10127), .D(net_2269), .CK(net_10794) );
DFF_X1 inst_8842 ( .Q(net_9610), .D(net_3145), .CK(net_15388) );
CLKBUF_X2 inst_13320 ( .A(net_13238), .Z(net_13239) );
OAI21_X2 inst_1815 ( .B2(net_10345), .ZN(net_6919), .A(net_1433), .B1(net_770) );
NAND2_X2 inst_3993 ( .A2(net_10127), .ZN(net_3174), .A1(net_3173) );
INV_X2 inst_6926 ( .A(net_3177), .ZN(net_1965) );
CLKBUF_X2 inst_13187 ( .A(net_10630), .Z(net_13106) );
INV_X4 inst_5267 ( .A(net_4168), .ZN(net_1468) );
CLKBUF_X2 inst_11140 ( .A(net_11058), .Z(net_11059) );
AND2_X4 inst_10422 ( .A2(net_10385), .ZN(net_4741), .A1(net_4006) );
CLKBUF_X2 inst_13272 ( .A(net_13190), .Z(net_13191) );
INV_X2 inst_7010 ( .ZN(net_1605), .A(net_1604) );
OAI211_X2 inst_2169 ( .C1(net_7203), .C2(net_6548), .ZN(net_6540), .B(net_5669), .A(net_3679) );
CLKBUF_X2 inst_12379 ( .A(net_12297), .Z(net_12298) );
CLKBUF_X2 inst_11903 ( .A(net_11821), .Z(net_11822) );
CLKBUF_X2 inst_15258 ( .A(net_15176), .Z(net_15177) );
OAI22_X2 inst_1326 ( .A2(net_9233), .A1(net_704), .B1(net_416), .B2(x3534), .ZN(x507) );
INV_X2 inst_6708 ( .ZN(net_8131), .A(net_8130) );
CLKBUF_X2 inst_14938 ( .A(net_14856), .Z(net_14857) );
CLKBUF_X2 inst_10840 ( .A(net_10758), .Z(net_10759) );
DFF_X2 inst_8191 ( .QN(net_9835), .D(net_5064), .CK(net_11729) );
CLKBUF_X2 inst_11920 ( .A(net_11838), .Z(net_11839) );
AND4_X4 inst_10319 ( .ZN(net_8190), .A3(net_7937), .A4(net_7646), .A2(net_7615), .A1(net_2126) );
INV_X4 inst_5442 ( .ZN(net_1099), .A(net_1098) );
NAND2_X2 inst_4238 ( .A2(net_10435), .ZN(net_1519), .A1(net_1030) );
AOI22_X2 inst_9496 ( .A1(net_9689), .B2(net_6443), .B1(net_6060), .A2(net_5966), .ZN(net_3827) );
INV_X4 inst_5275 ( .ZN(net_1346), .A(net_1345) );
INV_X4 inst_4758 ( .A(net_7665), .ZN(net_4301) );
AOI221_X2 inst_9857 ( .A(net_6889), .B2(net_6888), .C2(net_6887), .ZN(net_6861), .B1(net_3988), .C1(x4359) );
CLKBUF_X2 inst_15187 ( .A(net_15105), .Z(net_15106) );
NAND2_X2 inst_3875 ( .ZN(net_4034), .A1(net_4033), .A2(net_4021) );
NOR2_X2 inst_2629 ( .ZN(net_5962), .A2(net_5796), .A1(net_279) );
CLKBUF_X1 inst_8989 ( .A(x185142), .Z(x948) );
CLKBUF_X2 inst_14791 ( .A(net_14709), .Z(net_14710) );
CLKBUF_X2 inst_13658 ( .A(net_12284), .Z(net_13577) );
AOI222_X1 inst_9732 ( .B1(net_4188), .C1(net_3897), .C2(net_3121), .ZN(net_3120), .B2(net_2671), .A2(net_2670), .A1(net_1977) );
CLKBUF_X2 inst_14342 ( .A(net_14260), .Z(net_14261) );
CLKBUF_X2 inst_14887 ( .A(net_14661), .Z(net_14806) );
AOI22_X2 inst_9595 ( .A1(net_10541), .B1(net_9993), .ZN(net_3501), .A2(net_3500), .B2(net_2468) );
AOI22_X2 inst_9197 ( .A1(net_9887), .B1(net_9788), .A2(net_8042), .B2(net_8041), .ZN(net_6116) );
INV_X2 inst_7235 ( .A(net_9401), .ZN(net_8232) );
INV_X4 inst_6127 ( .A(net_10493), .ZN(net_486) );
CLKBUF_X2 inst_14867 ( .A(net_14785), .Z(net_14786) );
OAI222_X2 inst_1341 ( .A1(net_7728), .B2(net_7727), .C2(net_7726), .ZN(net_7581), .A2(net_7451), .B1(net_7022), .C1(net_573) );
OAI211_X2 inst_2154 ( .C2(net_6774), .ZN(net_6694), .A(net_6322), .B(net_6061), .C1(net_5073) );
SDFF_X2 inst_587 ( .Q(net_9256), .SE(net_4589), .D(net_139), .SI(net_105), .CK(net_13836) );
SDFF_X2 inst_666 ( .SI(net_9487), .Q(net_9487), .SE(net_3073), .CK(net_11875), .D(x2214) );
CLKBUF_X2 inst_10798 ( .A(net_10716), .Z(net_10717) );
INV_X4 inst_4602 ( .ZN(net_7719), .A(net_7655) );
INV_X4 inst_5937 ( .ZN(net_889), .A(net_571) );
INV_X2 inst_7182 ( .A(net_9416), .ZN(net_8217) );
NOR2_X2 inst_2602 ( .A2(net_6848), .ZN(net_6624), .A1(net_6623) );
OAI21_X2 inst_1829 ( .B1(net_7157), .ZN(net_6453), .B2(net_5657), .A(net_5432) );
XNOR2_X2 inst_109 ( .B(net_9428), .ZN(net_8111), .A(net_6251) );
OAI22_X2 inst_1182 ( .A1(net_7198), .A2(net_5139), .B2(net_5138), .ZN(net_5077), .B1(net_591) );
INV_X2 inst_6875 ( .ZN(net_3378), .A(net_3179) );
INV_X4 inst_6446 ( .ZN(net_3894), .A(net_152) );
NAND2_X2 inst_3983 ( .ZN(net_3241), .A2(net_3240), .A1(net_3118) );
CLKBUF_X2 inst_15066 ( .A(net_14984), .Z(net_14985) );
AOI221_X2 inst_9868 ( .B1(net_9761), .B2(net_9098), .A(net_6940), .C2(net_6939), .ZN(net_6835), .C1(net_6834) );
DFF_X2 inst_7368 ( .D(net_8755), .QN(net_259), .CK(net_11613) );
CLKBUF_X2 inst_12376 ( .A(net_12294), .Z(net_12295) );
CLKBUF_X2 inst_12275 ( .A(net_12193), .Z(net_12194) );
CLKBUF_X2 inst_11019 ( .A(net_10937), .Z(net_10938) );
INV_X4 inst_5984 ( .A(net_10508), .ZN(net_540) );
OAI221_X2 inst_1444 ( .B1(net_8565), .ZN(net_8556), .B2(net_8493), .C2(net_8441), .A(net_3905), .C1(net_2454) );
INV_X4 inst_5252 ( .ZN(net_1586), .A(net_1444) );
CLKBUF_X2 inst_11993 ( .A(net_11077), .Z(net_11912) );
CLKBUF_X2 inst_11217 ( .A(net_11015), .Z(net_11136) );
DFF_X2 inst_7594 ( .Q(net_10506), .D(net_7446), .CK(net_12288) );
INV_X4 inst_5490 ( .A(net_10369), .ZN(net_3706) );
OAI22_X2 inst_1231 ( .B1(net_7216), .A2(net_4890), .B2(net_4889), .ZN(net_4886), .A1(net_532) );
CLKBUF_X2 inst_11939 ( .A(net_11496), .Z(net_11858) );
CLKBUF_X2 inst_12210 ( .A(net_11701), .Z(net_12129) );
CLKBUF_X2 inst_13547 ( .A(net_13465), .Z(net_13466) );
CLKBUF_X2 inst_15557 ( .A(net_15475), .Z(net_15476) );
OR2_X2 inst_904 ( .ZN(net_5158), .A2(net_4638), .A1(net_3649) );
NAND2_X4 inst_3315 ( .ZN(net_8761), .A2(net_8760), .A1(net_8759) );
HA_X1 inst_7347 ( .S(net_4434), .CO(net_4433), .B(net_4198), .A(net_1146) );
CLKBUF_X2 inst_12100 ( .A(net_11816), .Z(net_12019) );
CLKBUF_X2 inst_10628 ( .A(net_10546), .Z(net_10547) );
CLKBUF_X2 inst_13147 ( .A(net_10997), .Z(net_13066) );
OAI211_X2 inst_2159 ( .C2(net_6778), .ZN(net_6689), .A(net_6310), .B(net_6049), .C1(net_5041) );
DFF_X2 inst_7753 ( .Q(net_9181), .D(net_6204), .CK(net_13579) );
INV_X2 inst_7051 ( .A(net_2623), .ZN(net_1330) );
INV_X4 inst_6266 ( .A(net_9173), .ZN(net_1033) );
CLKBUF_X2 inst_15783 ( .A(net_10773), .Z(net_15702) );
NAND2_X2 inst_3923 ( .A2(net_9053), .ZN(net_7955), .A1(net_3884) );
CLKBUF_X2 inst_13094 ( .A(net_13012), .Z(net_13013) );
CLKBUF_X2 inst_11652 ( .A(net_10697), .Z(net_11571) );
INV_X4 inst_4831 ( .ZN(net_4056), .A(net_3188) );
OR2_X4 inst_757 ( .ZN(net_4397), .A2(net_4396), .A1(net_1672) );
CLKBUF_X2 inst_14809 ( .A(net_14727), .Z(net_14728) );
AND2_X4 inst_10431 ( .ZN(net_3489), .A2(net_3010), .A1(net_1156) );
XNOR2_X2 inst_343 ( .ZN(net_2866), .B(net_2865), .A(net_1584) );
OAI221_X2 inst_1627 ( .B1(net_10306), .C1(net_7243), .B2(net_5591), .ZN(net_5580), .C2(net_4902), .A(net_3731) );
INV_X4 inst_4739 ( .ZN(net_5167), .A(net_4454) );
CLKBUF_X2 inst_12670 ( .A(net_12027), .Z(net_12589) );
SDFF_X2 inst_543 ( .Q(net_9305), .D(net_9305), .SI(net_9156), .SE(net_7553), .CK(net_14038) );
OAI22_X2 inst_1106 ( .ZN(net_7641), .A1(net_6192), .A2(net_6191), .B2(net_6190), .B1(net_5249) );
CLKBUF_X2 inst_12131 ( .A(net_12049), .Z(net_12050) );
CLKBUF_X2 inst_14194 ( .A(net_14112), .Z(net_14113) );
CLKBUF_X2 inst_13557 ( .A(net_13475), .Z(net_13476) );
CLKBUF_X2 inst_12994 ( .A(net_12912), .Z(net_12913) );
CLKBUF_X2 inst_13122 ( .A(net_13040), .Z(net_13041) );
INV_X2 inst_6882 ( .A(net_3035), .ZN(net_2844) );
NAND2_X2 inst_3817 ( .A1(net_10086), .A2(net_4534), .ZN(net_4521) );
CLKBUF_X2 inst_15201 ( .A(net_14014), .Z(net_15120) );
DFF_X2 inst_7697 ( .Q(net_9205), .D(net_6556), .CK(net_11326) );
OAI211_X2 inst_2070 ( .C2(net_7167), .ZN(net_7164), .B(net_4722), .A(net_4207), .C1(net_1557) );
CLKBUF_X2 inst_15458 ( .A(net_13197), .Z(net_15377) );
INV_X4 inst_5065 ( .A(net_3807), .ZN(net_1865) );
OAI22_X2 inst_1256 ( .B1(net_7231), .A2(net_4826), .B2(net_4825), .ZN(net_4817), .A1(net_511) );
CLKBUF_X2 inst_15710 ( .A(net_15628), .Z(net_15629) );
INV_X4 inst_5765 ( .A(net_2085), .ZN(net_1177) );
NOR2_X2 inst_2890 ( .ZN(net_2534), .A2(net_1781), .A1(net_748) );
CLKBUF_X2 inst_13858 ( .A(net_10775), .Z(net_13777) );
AOI22_X2 inst_9549 ( .B1(net_9903), .A1(net_9673), .A2(net_5966), .B2(net_4969), .ZN(net_3771) );
CLKBUF_X2 inst_12538 ( .A(net_12456), .Z(net_12457) );
INV_X4 inst_6337 ( .A(net_9842), .ZN(net_632) );
CLKBUF_X2 inst_15752 ( .A(net_15670), .Z(net_15671) );
DFF_X2 inst_7555 ( .QN(net_9354), .D(net_7702), .CK(net_15303) );
OAI21_X2 inst_1903 ( .B1(net_7201), .B2(net_4862), .ZN(net_4849), .A(net_4521) );
CLKBUF_X2 inst_14254 ( .A(net_12928), .Z(net_14173) );
AOI22_X2 inst_9503 ( .A1(net_9889), .B1(net_9790), .ZN(net_3820), .A2(net_2973), .B2(net_2462) );
DFF_X2 inst_8347 ( .QN(net_10374), .D(net_2772), .CK(net_13684) );
CLKBUF_X2 inst_11230 ( .A(net_11148), .Z(net_11149) );
CLKBUF_X2 inst_13716 ( .A(net_11206), .Z(net_13635) );
NAND2_X2 inst_4304 ( .A2(net_10351), .ZN(net_1613), .A1(net_1212) );
NOR2_X2 inst_2554 ( .ZN(net_7860), .A1(net_7859), .A2(net_7827) );
INV_X2 inst_6848 ( .A(net_10374), .ZN(net_3459) );
CLKBUF_X2 inst_13810 ( .A(net_13728), .Z(net_13729) );
NOR2_X2 inst_2745 ( .ZN(net_4145), .A1(net_3685), .A2(x3698) );
AOI22_X2 inst_9423 ( .A1(net_10187), .A2(net_4656), .B2(net_4655), .ZN(net_4646), .B1(x4694) );
CLKBUF_X2 inst_14422 ( .A(net_14340), .Z(net_14341) );
CLKBUF_X2 inst_15295 ( .A(net_15213), .Z(net_15214) );
NOR2_X2 inst_2604 ( .A1(net_9650), .ZN(net_6551), .A2(net_5764) );
CLKBUF_X2 inst_11802 ( .A(net_11720), .Z(net_11721) );
INV_X2 inst_7253 ( .A(net_9215), .ZN(net_342) );
CLKBUF_X2 inst_13125 ( .A(net_13043), .Z(net_13044) );
CLKBUF_X2 inst_11297 ( .A(net_11215), .Z(net_11216) );
CLKBUF_X2 inst_12452 ( .A(net_12370), .Z(net_12371) );
NAND2_X2 inst_4410 ( .A2(net_10119), .A1(net_10118), .ZN(net_3062) );
OAI22_X2 inst_1244 ( .A1(net_7108), .A2(net_4871), .B2(net_4870), .ZN(net_4866), .B1(net_531) );
DFF_X2 inst_8134 ( .Q(net_9947), .D(net_5112), .CK(net_14732) );
CLKBUF_X2 inst_15019 ( .A(net_14937), .Z(net_14938) );
NAND3_X2 inst_3248 ( .A2(net_9243), .ZN(net_5101), .A1(net_4607), .A3(net_4606) );
SDFF_X2 inst_582 ( .QN(net_9193), .D(net_9184), .SI(net_5443), .SE(net_4587), .CK(net_11290) );
INV_X8 inst_4515 ( .A(net_8918), .ZN(net_8915) );
CLKBUF_X2 inst_12329 ( .A(net_12247), .Z(net_12248) );
OAI211_X2 inst_2110 ( .C2(net_6774), .ZN(net_6738), .A(net_6399), .B(net_6097), .C1(net_384) );
OAI21_X2 inst_1850 ( .ZN(net_5882), .B1(net_5881), .A(net_5588), .B2(net_5322) );
NAND2_X2 inst_3477 ( .A1(net_9456), .A2(net_8951), .ZN(net_8435) );
AOI221_X2 inst_9774 ( .B2(net_10170), .ZN(net_7491), .C2(net_7409), .A(net_7074), .C1(net_6909), .B1(net_2227) );
OAI21_X2 inst_1950 ( .A(net_7454), .ZN(net_3927), .B2(net_3291), .B1(net_1858) );
CLKBUF_X2 inst_12057 ( .A(net_11975), .Z(net_11976) );
CLKBUF_X2 inst_13896 ( .A(net_13814), .Z(net_13815) );
DFF_X2 inst_7463 ( .QN(net_9642), .D(net_8157), .CK(net_13138) );
INV_X4 inst_5287 ( .A(net_8687), .ZN(net_1320) );
CLKBUF_X2 inst_15051 ( .A(net_14969), .Z(net_14970) );
AOI22_X2 inst_9402 ( .ZN(net_5976), .A2(net_4701), .B1(net_3712), .B2(net_2698), .A1(net_2364) );
DFF_X2 inst_7690 ( .Q(net_10192), .D(net_6577), .CK(net_12277) );
INV_X2 inst_7292 ( .A(net_9040), .ZN(net_9039) );
CLKBUF_X2 inst_12914 ( .A(net_12832), .Z(net_12833) );
CLKBUF_X2 inst_12673 ( .A(net_11955), .Z(net_12592) );
OAI211_X2 inst_2057 ( .A(net_7783), .C2(net_7782), .ZN(net_7776), .B(net_7682), .C1(net_2478) );
CLKBUF_X2 inst_15217 ( .A(net_15135), .Z(net_15136) );
CLKBUF_X2 inst_14727 ( .A(net_14645), .Z(net_14646) );
CLKBUF_X2 inst_13408 ( .A(net_13326), .Z(net_13327) );
OR2_X4 inst_843 ( .A2(net_10252), .A1(net_10251), .ZN(net_2103) );
OAI21_X2 inst_1779 ( .ZN(net_7786), .B1(net_7785), .A(net_7725), .B2(net_7724) );
CLKBUF_X2 inst_10710 ( .A(net_10628), .Z(net_10629) );
INV_X2 inst_7299 ( .A(net_9062), .ZN(net_9061) );
OAI211_X2 inst_2115 ( .C2(net_6774), .ZN(net_6733), .A(net_6360), .B(net_6147), .C1(net_386) );
INV_X4 inst_5146 ( .ZN(net_2876), .A(net_2198) );
NAND3_X2 inst_3251 ( .ZN(net_4951), .A1(net_4558), .A3(net_4557), .A2(net_2950) );
XNOR2_X2 inst_112 ( .B(net_9427), .ZN(net_8083), .A(net_6427) );
OAI21_X2 inst_1728 ( .ZN(net_8911), .B1(net_8785), .A(net_8783), .B2(net_8781) );
CLKBUF_X2 inst_14974 ( .A(net_11067), .Z(net_14893) );
OR2_X2 inst_916 ( .ZN(net_3468), .A2(net_3467), .A1(net_2265) );
OAI221_X2 inst_1722 ( .B1(net_10460), .ZN(net_2703), .C2(net_2702), .A(net_2070), .C1(net_1544), .B2(net_825) );
CLKBUF_X2 inst_11161 ( .A(net_11079), .Z(net_11080) );
INV_X4 inst_5570 ( .ZN(net_1259), .A(net_910) );
CLKBUF_X2 inst_13799 ( .A(net_11501), .Z(net_13718) );
AOI221_X2 inst_9824 ( .B1(net_9771), .B2(net_9097), .A(net_6940), .C1(net_6939), .ZN(net_6925), .C2(net_241) );
AOI22_X2 inst_9523 ( .B1(net_9769), .A1(net_9670), .A2(net_5966), .ZN(net_3798), .B2(net_2462) );
DFF_X1 inst_8754 ( .D(net_5285), .Q(net_264), .CK(net_15178) );
INV_X2 inst_7300 ( .A(net_9066), .ZN(net_9065) );
INV_X4 inst_6409 ( .A(net_9300), .ZN(net_637) );
NAND2_X2 inst_3665 ( .A2(net_10275), .ZN(net_6258), .A1(net_1960) );
DFF_X2 inst_8376 ( .QN(net_8829), .D(net_1496), .CK(net_12105) );
DFF_X2 inst_7441 ( .QN(net_9300), .D(net_8202), .CK(net_11502) );
NOR2_X2 inst_2724 ( .A2(net_5347), .ZN(net_4621), .A1(net_4170) );
NOR2_X2 inst_2525 ( .ZN(net_8428), .A1(net_8175), .A2(net_8174) );
AOI22_X2 inst_9353 ( .B1(net_10009), .A2(net_5743), .B2(net_5742), .ZN(net_5594), .A1(net_249) );
NOR2_X2 inst_2968 ( .A1(net_10462), .ZN(net_1604), .A2(net_1107) );
CLKBUF_X2 inst_12010 ( .A(net_11703), .Z(net_11929) );
CLKBUF_X2 inst_11334 ( .A(net_10992), .Z(net_11253) );
INV_X2 inst_7067 ( .ZN(net_1257), .A(net_1256) );
CLKBUF_X2 inst_12875 ( .A(net_12793), .Z(net_12794) );
DFF_X2 inst_7916 ( .Q(net_9846), .D(net_5878), .CK(net_11939) );
NOR2_X2 inst_2964 ( .A1(net_10458), .ZN(net_1694), .A2(net_805) );
CLKBUF_X2 inst_11760 ( .A(net_11678), .Z(net_11679) );
NAND2_X2 inst_3721 ( .A2(net_10169), .A1(net_9735), .ZN(net_7070) );
NOR4_X2 inst_2349 ( .A4(net_3712), .ZN(net_2961), .A1(net_2629), .A2(net_2628), .A3(net_2627) );
DFF_X1 inst_8855 ( .Q(net_10526), .D(net_98), .CK(net_10890) );
SDFF_X2 inst_646 ( .Q(net_9452), .D(net_9452), .SE(net_3293), .CK(net_12434), .SI(x2400) );
INV_X4 inst_5751 ( .ZN(net_738), .A(net_737) );
INV_X4 inst_5076 ( .ZN(net_3602), .A(net_2247) );
INV_X2 inst_6667 ( .ZN(net_8361), .A(net_8304) );
NAND2_X2 inst_4032 ( .A2(net_3165), .ZN(net_2969), .A1(net_2086) );
DFF_X2 inst_8062 ( .QN(net_10351), .D(net_5333), .CK(net_13631) );
CLKBUF_X2 inst_14310 ( .A(net_11076), .Z(net_14229) );
AOI21_X2 inst_10213 ( .ZN(net_2431), .B1(net_2430), .B2(net_2181), .A(net_976) );
NAND3_X2 inst_3169 ( .A3(net_9570), .A2(net_9045), .ZN(net_8792), .A1(net_4590) );
AOI22_X2 inst_9387 ( .B1(net_9900), .A1(net_5759), .B2(net_5758), .ZN(net_5436), .A2(net_239) );
XNOR2_X2 inst_382 ( .B(net_9941), .ZN(net_2282), .A(net_2281) );
CLKBUF_X2 inst_13278 ( .A(net_11039), .Z(net_13197) );
AOI221_X2 inst_9841 ( .A(net_6889), .B2(net_6888), .C2(net_6887), .ZN(net_6877), .B1(net_5841), .C1(x5961) );
INV_X4 inst_5344 ( .ZN(net_1568), .A(net_1243) );
NOR4_X2 inst_2329 ( .ZN(net_5221), .A2(net_5220), .A4(net_5219), .A3(net_4540), .A1(net_3354) );
CLKBUF_X2 inst_11119 ( .A(net_11037), .Z(net_11038) );
INV_X4 inst_6101 ( .A(net_10402), .ZN(net_492) );
AND3_X4 inst_10361 ( .ZN(net_4353), .A3(net_4232), .A2(net_4230), .A1(x6599) );
INV_X2 inst_7161 ( .A(net_7031), .ZN(net_628) );
CLKBUF_X2 inst_14248 ( .A(net_14166), .Z(net_14167) );
AOI221_X2 inst_9799 ( .B1(net_9960), .A(net_7090), .B2(net_7089), .C2(net_7088), .ZN(net_7005), .C1(net_6828) );
INV_X4 inst_6067 ( .ZN(net_1995), .A(net_224) );
NOR2_X2 inst_2788 ( .ZN(net_3076), .A1(net_3075), .A2(net_3074) );
AND2_X2 inst_10560 ( .ZN(net_3130), .A1(net_3129), .A2(net_2915) );
INV_X4 inst_6015 ( .A(net_10329), .ZN(net_737) );
CLKBUF_X2 inst_11891 ( .A(net_11809), .Z(net_11810) );
CLKBUF_X2 inst_15040 ( .A(net_14958), .Z(net_14959) );
INV_X4 inst_6565 ( .A(net_10437), .ZN(net_712) );
AND2_X4 inst_10415 ( .ZN(net_4288), .A2(x3638), .A1(x813) );
OAI22_X2 inst_1049 ( .ZN(net_7536), .A1(net_7535), .A2(net_7397), .B2(net_7396), .B1(net_466) );
AOI21_X2 inst_10194 ( .A(net_9107), .ZN(net_3640), .B2(net_2467), .B1(net_1263) );
DFF_X1 inst_8418 ( .Q(net_9570), .D(net_8786), .CK(net_11632) );
XNOR2_X2 inst_168 ( .B(net_6039), .ZN(net_5789), .A(net_5234) );
AOI22_X2 inst_9139 ( .A1(net_9723), .A2(net_6382), .ZN(net_6348), .B1(net_6347), .B2(net_5263) );
INV_X4 inst_5116 ( .ZN(net_2678), .A(net_1629) );
DFF_X2 inst_8085 ( .QN(net_9927), .D(net_5036), .CK(net_12125) );
INV_X4 inst_4575 ( .ZN(net_8338), .A(net_8132) );
INV_X4 inst_6037 ( .A(net_10246), .ZN(net_715) );
CLKBUF_X2 inst_13819 ( .A(net_13737), .Z(net_13738) );
DFF_X1 inst_8688 ( .D(net_6714), .Q(net_140), .CK(net_14250) );
AND2_X2 inst_10547 ( .ZN(net_3965), .A2(net_3485), .A1(net_2378) );
OAI22_X2 inst_991 ( .A2(net_8962), .B2(net_8659), .ZN(net_8641), .B1(net_8403), .A1(net_6586) );
CLKBUF_X2 inst_12258 ( .A(net_12176), .Z(net_12177) );
CLKBUF_X2 inst_10642 ( .A(net_10560), .Z(net_10561) );
INV_X4 inst_5613 ( .ZN(net_6414), .A(net_1367) );
CLKBUF_X2 inst_15113 ( .A(net_15031), .Z(net_15032) );
AOI22_X2 inst_9643 ( .ZN(net_2847), .A1(net_2846), .B2(net_2845), .B1(net_2321), .A2(net_2235) );
AOI22_X2 inst_9249 ( .A2(net_6141), .B2(net_6129), .ZN(net_6062), .B1(net_3433), .A1(net_1228) );
SDFF_X2 inst_580 ( .SE(net_5278), .SI(net_2798), .CK(net_14872), .Q(x480), .D(x480) );
XNOR2_X2 inst_170 ( .ZN(net_5762), .A(net_4919), .B(net_1139) );
CLKBUF_X2 inst_13533 ( .A(net_13451), .Z(net_13452) );
AOI22_X2 inst_9160 ( .A2(net_6420), .ZN(net_6315), .A1(net_6314), .B2(net_5263), .B1(net_2585) );
NAND2_X2 inst_3691 ( .A2(net_9261), .ZN(net_6237), .A1(net_5973) );
CLKBUF_X2 inst_13159 ( .A(net_13077), .Z(net_13078) );
DFF_X2 inst_7823 ( .Q(net_9652), .D(net_6206), .CK(net_11819) );
OAI21_X2 inst_1857 ( .ZN(net_5793), .B1(net_5792), .A(net_5381), .B2(net_1282) );
CLKBUF_X2 inst_12647 ( .A(net_12565), .Z(net_12566) );
CLKBUF_X2 inst_11536 ( .A(net_11033), .Z(net_11455) );
HA_X1 inst_7336 ( .CO(net_7321), .S(net_6959), .A(net_6958), .B(net_5988) );
CLKBUF_X2 inst_11304 ( .A(net_11222), .Z(net_11223) );
SDFF_X2 inst_468 ( .SE(net_8812), .SI(net_8637), .CK(net_11906), .Q(x798), .D(x798) );
OAI22_X2 inst_1099 ( .A1(net_9191), .A2(net_6299), .B2(net_6298), .ZN(net_6272), .B1(net_5011) );
INV_X4 inst_6611 ( .A(net_9934), .ZN(net_901) );
AOI22_X2 inst_9103 ( .A1(net_9683), .A2(net_6420), .ZN(net_6389), .B2(net_5263), .B1(net_1008) );
DFF_X1 inst_8746 ( .Q(net_10240), .D(net_5424), .CK(net_10918) );
MUX2_X2 inst_4428 ( .B(net_9153), .S(net_7553), .Z(net_7500), .A(net_7499) );
NAND2_X2 inst_3616 ( .ZN(net_7116), .A2(net_6877), .A1(net_6594) );
CLKBUF_X2 inst_14762 ( .A(net_14680), .Z(net_14681) );
INV_X4 inst_4889 ( .ZN(net_4239), .A(net_2940) );
CLKBUF_X2 inst_13842 ( .A(net_12672), .Z(net_13761) );
OAI211_X2 inst_2190 ( .C1(net_7203), .C2(net_6542), .ZN(net_6519), .B(net_5615), .A(net_3679) );
XNOR2_X2 inst_429 ( .B(net_10042), .A(net_1417), .ZN(net_1097) );
NOR2_X2 inst_2692 ( .A1(net_9613), .ZN(net_4539), .A2(net_4162) );
CLKBUF_X2 inst_13580 ( .A(net_13498), .Z(net_13499) );
OAI221_X2 inst_1599 ( .C1(net_10214), .B1(net_7297), .C2(net_5642), .ZN(net_5638), .A(net_5637), .B2(net_4905) );
AOI211_X2 inst_10298 ( .ZN(net_3697), .C1(net_3696), .C2(net_3695), .B(net_3294), .A(net_3088) );
DFF_X2 inst_7808 ( .Q(net_10008), .D(net_6479), .CK(net_14311) );
INV_X4 inst_5026 ( .ZN(net_2613), .A(net_1939) );
NAND2_X2 inst_3565 ( .A2(net_7748), .ZN(net_7684), .A1(net_7683) );
HA_X1 inst_7348 ( .S(net_4432), .CO(net_4431), .B(net_4194), .A(net_1190) );
INV_X4 inst_5995 ( .A(net_10193), .ZN(net_534) );
DFF_X2 inst_8055 ( .QN(net_10318), .D(net_5586), .CK(net_15480) );
CLKBUF_X2 inst_14141 ( .A(net_14059), .Z(net_14060) );
DFF_X2 inst_7922 ( .Q(net_9224), .D(net_5817), .CK(net_13002) );
INV_X4 inst_5687 ( .ZN(net_1311), .A(net_967) );
CLKBUF_X2 inst_13824 ( .A(net_13742), .Z(net_13743) );
CLKBUF_X2 inst_13567 ( .A(net_13485), .Z(net_13486) );
INV_X2 inst_6960 ( .A(net_3199), .ZN(net_1869) );
DFF_X1 inst_8629 ( .Q(net_9788), .D(net_7199), .CK(net_13355) );
NAND2_X2 inst_3977 ( .A2(net_5268), .A1(net_3591), .ZN(net_3288) );
NAND2_X2 inst_3467 ( .A1(net_9468), .ZN(net_8877), .A2(net_8475) );
NOR2_X2 inst_2593 ( .ZN(net_7291), .A2(net_6912), .A1(net_2675) );
NAND4_X2 inst_3064 ( .ZN(net_5716), .A4(net_4899), .A1(net_3826), .A2(net_3825), .A3(net_3824) );
CLKBUF_X2 inst_11717 ( .A(net_11635), .Z(net_11636) );
NAND2_X2 inst_3676 ( .A1(net_8117), .ZN(net_6902), .A2(net_6231) );
AOI221_X2 inst_9850 ( .B1(net_9769), .B2(net_9097), .A(net_6940), .C1(net_6939), .ZN(net_6868), .C2(net_239) );
INV_X4 inst_5021 ( .ZN(net_5478), .A(net_1982) );
CLKBUF_X2 inst_13550 ( .A(net_13468), .Z(net_13469) );
XNOR2_X2 inst_318 ( .ZN(net_3217), .B(net_3003), .A(net_2038) );
CLKBUF_X2 inst_15480 ( .A(net_11436), .Z(net_15399) );
DFF_X2 inst_7948 ( .QN(net_10363), .D(net_5700), .CK(net_13646) );
NAND2_X2 inst_4033 ( .ZN(net_2959), .A1(net_2958), .A2(net_2957) );
CLKBUF_X2 inst_14210 ( .A(net_14128), .Z(net_14129) );
DFF_X1 inst_8538 ( .Q(net_9960), .D(net_7350), .CK(net_14637) );
INV_X4 inst_5044 ( .ZN(net_7454), .A(net_1912) );
NOR2_X2 inst_2899 ( .ZN(net_5813), .A1(net_1665), .A2(net_1664) );
NAND2_X2 inst_4065 ( .ZN(net_2722), .A1(net_2721), .A2(net_2720) );
CLKBUF_X2 inst_13790 ( .A(net_13708), .Z(net_13709) );
OAI221_X2 inst_1486 ( .ZN(net_7452), .C2(net_7437), .A(net_7151), .B1(net_4509), .B2(net_4456), .C1(net_3299) );
CLKBUF_X2 inst_13449 ( .A(net_13367), .Z(net_13368) );
OAI211_X2 inst_2281 ( .C1(net_7124), .C2(net_6480), .ZN(net_6215), .B(net_5737), .A(net_3679) );
CLKBUF_X2 inst_15510 ( .A(net_15428), .Z(net_15429) );
OAI22_X2 inst_1175 ( .A1(net_7201), .A2(net_5107), .B2(net_5105), .ZN(net_5086), .B1(net_682) );
CLKBUF_X2 inst_12666 ( .A(net_12584), .Z(net_12585) );
CLKBUF_X2 inst_13929 ( .A(net_13847), .Z(net_13848) );
CLKBUF_X2 inst_14222 ( .A(net_14140), .Z(net_14141) );
INV_X4 inst_5877 ( .ZN(net_1386), .A(net_879) );
INV_X4 inst_5256 ( .A(net_8687), .ZN(net_1428) );
NAND2_X2 inst_4096 ( .ZN(net_2955), .A2(net_2536), .A1(net_2169) );
CLKBUF_X2 inst_12208 ( .A(net_12126), .Z(net_12127) );
CLKBUF_X2 inst_12164 ( .A(net_12082), .Z(net_12083) );
DFF_X2 inst_8305 ( .QN(net_10349), .D(net_4570), .CK(net_11171) );
INV_X8 inst_4509 ( .ZN(net_6404), .A(net_5295) );
XNOR2_X2 inst_395 ( .ZN(net_1998), .B(net_666), .A(net_415) );
CLKBUF_X2 inst_14106 ( .A(net_14024), .Z(net_14025) );
CLKBUF_X2 inst_10927 ( .A(net_10845), .Z(net_10846) );
INV_X2 inst_6808 ( .ZN(net_4996), .A(net_4995) );
OR2_X4 inst_841 ( .A1(net_10158), .A2(net_9734), .ZN(net_2209) );
CLKBUF_X2 inst_15323 ( .A(net_15241), .Z(net_15242) );
NAND2_X2 inst_3963 ( .A2(net_4070), .ZN(net_3896), .A1(net_1246) );
CLKBUF_X2 inst_13682 ( .A(net_13600), .Z(net_13601) );
CLKBUF_X2 inst_12508 ( .A(net_12426), .Z(net_12427) );
HA_X1 inst_7328 ( .S(net_7735), .CO(net_7734), .B(net_7564), .A(net_5790) );
OR4_X2 inst_689 ( .A1(net_5685), .ZN(net_4632), .A4(net_4631), .A3(net_4460), .A2(net_4205) );
CLKBUF_X2 inst_13412 ( .A(net_13330), .Z(net_13331) );
MUX2_X1 inst_4453 ( .S(net_6041), .A(net_293), .B(x5364), .Z(x166) );
NOR2_X2 inst_2689 ( .ZN(net_4544), .A2(net_4543), .A1(net_2393) );
CLKBUF_X2 inst_13538 ( .A(net_13456), .Z(net_13457) );
INV_X4 inst_6361 ( .A(net_9516), .ZN(net_7953) );
INV_X4 inst_4895 ( .A(net_8855), .ZN(net_3135) );
NAND2_X2 inst_3896 ( .ZN(net_3931), .A1(net_3896), .A2(net_3449) );
AOI22_X2 inst_9622 ( .A1(net_10075), .A2(net_5319), .B2(net_5174), .ZN(net_3430), .B1(net_3429) );
OAI221_X2 inst_1558 ( .C2(net_9047), .B2(net_7287), .B1(net_7203), .ZN(net_7197), .A(net_6799), .C1(net_5486) );
NAND2_X2 inst_3679 ( .ZN(net_6589), .A1(net_6205), .A2(net_5802) );
CLKBUF_X2 inst_14212 ( .A(net_14130), .Z(net_14131) );
CLKBUF_X2 inst_12630 ( .A(net_10978), .Z(net_12549) );
NOR2_X2 inst_2906 ( .A1(net_10248), .ZN(net_2330), .A2(net_1393) );
INV_X4 inst_6272 ( .ZN(net_6834), .A(net_231) );
INV_X4 inst_5848 ( .ZN(net_1342), .A(net_649) );
CLKBUF_X2 inst_14622 ( .A(net_13477), .Z(net_14541) );
CLKBUF_X2 inst_14206 ( .A(net_14124), .Z(net_14125) );
CLKBUF_X2 inst_13398 ( .A(net_13316), .Z(net_13317) );
CLKBUF_X2 inst_12836 ( .A(net_12754), .Z(net_12755) );
NAND2_X2 inst_3886 ( .A2(net_10385), .ZN(net_4180), .A1(net_4015) );
CLKBUF_X2 inst_13587 ( .A(net_13505), .Z(net_13506) );
AOI22_X2 inst_9072 ( .B1(net_9664), .A1(net_6813), .A2(net_6684), .B2(net_6683), .ZN(net_6594) );
DFF_X1 inst_8797 ( .QN(net_10384), .D(net_4010), .CK(net_11056) );
DFF_X1 inst_8685 ( .D(net_6718), .QN(net_165), .CK(net_14341) );
OAI221_X2 inst_1615 ( .B1(net_10424), .C1(net_7297), .ZN(net_5596), .B2(net_4477), .C2(net_4455), .A(net_3507) );
CLKBUF_X2 inst_13201 ( .A(net_13119), .Z(net_13120) );
AOI22_X2 inst_9148 ( .A1(net_9741), .A2(net_6382), .ZN(net_6337), .B1(net_5964), .B2(net_5263) );
CLKBUF_X2 inst_11692 ( .A(net_11610), .Z(net_11611) );
CLKBUF_X2 inst_11434 ( .A(net_11352), .Z(net_11353) );
AOI22_X2 inst_9505 ( .B1(net_9862), .A1(net_9696), .ZN(net_3818), .A2(net_3039), .B2(net_2973) );
DFF_X2 inst_7503 ( .Q(net_9540), .D(net_7991), .CK(net_14000) );
CLKBUF_X2 inst_10643 ( .A(net_10561), .Z(net_10562) );
CLKBUF_X2 inst_12406 ( .A(net_12324), .Z(net_12325) );
CLKBUF_X2 inst_11510 ( .A(net_10710), .Z(net_11429) );
CLKBUF_X2 inst_13760 ( .A(net_13678), .Z(net_13679) );
AOI221_X2 inst_9890 ( .B1(net_9876), .B2(net_9101), .A(net_6945), .C2(net_6944), .ZN(net_6804), .C1(net_247) );
DFF_X2 inst_8313 ( .Q(net_10058), .D(net_4091), .CK(net_10852) );
OAI211_X2 inst_2145 ( .C2(net_6778), .ZN(net_6703), .A(net_6328), .B(net_6066), .C1(net_4749) );
OR3_X2 inst_709 ( .A3(net_7519), .ZN(net_7388), .A2(net_6584), .A1(net_2579) );
NOR3_X2 inst_2375 ( .A1(net_8190), .A2(net_8122), .ZN(net_8121), .A3(net_7892) );
CLKBUF_X2 inst_12127 ( .A(net_12045), .Z(net_12046) );
INV_X4 inst_5725 ( .ZN(net_2212), .A(net_759) );
OR2_X2 inst_920 ( .ZN(net_3250), .A1(net_3249), .A2(net_3248) );
NAND2_X2 inst_3454 ( .A1(net_9488), .A2(net_8476), .ZN(net_8470) );
INV_X4 inst_6298 ( .A(net_9203), .ZN(net_722) );
INV_X4 inst_5741 ( .ZN(net_824), .A(net_745) );
CLKBUF_X2 inst_13400 ( .A(net_13318), .Z(net_13319) );
INV_X4 inst_6571 ( .A(net_10101), .ZN(net_5831) );
CLKBUF_X2 inst_12080 ( .A(net_11998), .Z(net_11999) );
AOI221_X2 inst_9956 ( .C1(net_10497), .B1(net_10287), .C2(net_6415), .ZN(net_4776), .B2(net_4774), .A(net_4345) );
CLKBUF_X2 inst_12517 ( .A(net_12435), .Z(net_12436) );
CLKBUF_X2 inst_12331 ( .A(net_12249), .Z(net_12250) );
CLKBUF_X2 inst_12106 ( .A(net_12024), .Z(net_12025) );
DFF_X2 inst_7389 ( .D(net_8656), .QN(net_270), .CK(net_12638) );
INV_X4 inst_4610 ( .ZN(net_7930), .A(net_7560) );
CLKBUF_X2 inst_13350 ( .A(net_13091), .Z(net_13269) );
CLKBUF_X2 inst_11629 ( .A(net_11547), .Z(net_11548) );
INV_X4 inst_6116 ( .ZN(net_4019), .A(net_122) );
NAND2_X2 inst_4403 ( .A2(net_10296), .A1(net_10283), .ZN(net_634) );
CLKBUF_X2 inst_13797 ( .A(net_13715), .Z(net_13716) );
CLKBUF_X2 inst_14203 ( .A(net_14121), .Z(net_14122) );
NOR2_X2 inst_2889 ( .ZN(net_2528), .A2(net_1782), .A1(net_1448) );
CLKBUF_X2 inst_14589 ( .A(net_14507), .Z(net_14508) );
CLKBUF_X2 inst_11432 ( .A(net_11350), .Z(net_11351) );
CLKBUF_X2 inst_11380 ( .A(net_11298), .Z(net_11299) );
AOI21_X2 inst_10109 ( .ZN(net_4627), .B1(net_4626), .A(net_4315), .B2(net_3921) );
AOI221_X2 inst_9885 ( .B1(net_9791), .B2(net_9097), .A(net_6940), .C2(net_6939), .ZN(net_6812), .C1(net_6811) );
CLKBUF_X2 inst_15265 ( .A(net_15183), .Z(net_15184) );
CLKBUF_X2 inst_13743 ( .A(net_13661), .Z(net_13662) );
DFF_X2 inst_8034 ( .Q(net_9228), .D(net_5451), .CK(net_14090) );
OAI211_X2 inst_2189 ( .C1(net_7243), .C2(net_6542), .ZN(net_6520), .B(net_5568), .A(net_3679) );
INV_X4 inst_5448 ( .ZN(net_3204), .A(net_1543) );
NAND2_X2 inst_4198 ( .ZN(net_1803), .A1(net_1802), .A2(net_1337) );
XNOR2_X2 inst_315 ( .ZN(net_3220), .B(net_2802), .A(net_2650) );
NOR2_X2 inst_2935 ( .A2(net_6958), .ZN(net_2304), .A1(net_1350) );
CLKBUF_X2 inst_13176 ( .A(net_13094), .Z(net_13095) );
CLKBUF_X2 inst_14989 ( .A(net_12357), .Z(net_14908) );
DFF_X2 inst_7653 ( .D(net_6706), .QN(net_184), .CK(net_15238) );
XNOR2_X2 inst_216 ( .ZN(net_4683), .A(net_4270), .B(net_2354) );
NAND2_X4 inst_3369 ( .ZN(net_9069), .A1(net_4023), .A2(net_3900) );
AOI22_X2 inst_8992 ( .A2(net_9578), .ZN(net_8693), .A1(net_8685), .B2(net_8675), .B1(net_807) );
CLKBUF_X2 inst_13612 ( .A(net_13530), .Z(net_13531) );
CLKBUF_X2 inst_15126 ( .A(net_15044), .Z(net_15045) );
CLKBUF_X2 inst_10924 ( .A(net_10630), .Z(net_10843) );
CLKBUF_X2 inst_14858 ( .A(net_14776), .Z(net_14777) );
CLKBUF_X2 inst_14444 ( .A(net_14362), .Z(net_14363) );
CLKBUF_X2 inst_13099 ( .A(net_13017), .Z(net_13018) );
CLKBUF_X2 inst_12987 ( .A(net_11924), .Z(net_12906) );
AOI22_X2 inst_9202 ( .A1(net_9891), .B1(net_9792), .B2(net_8041), .ZN(net_6110), .A2(net_6109) );
OAI211_X2 inst_2060 ( .ZN(net_7758), .C2(net_7757), .B(net_7609), .A(net_3679), .C1(net_1312) );
AOI21_X2 inst_10179 ( .B2(net_3891), .ZN(net_3596), .A(net_3595), .B1(net_3594) );
DFF_X1 inst_8771 ( .Q(net_10536), .D(net_4790), .CK(net_10959) );
NOR2_X2 inst_2680 ( .ZN(net_4984), .A2(net_4679), .A1(net_692) );
XNOR2_X2 inst_415 ( .B(net_9745), .A(net_1417), .ZN(net_1412) );
AND2_X2 inst_10592 ( .ZN(net_2382), .A1(net_2381), .A2(net_2380) );
INV_X16 inst_7321 ( .ZN(net_8385), .A(net_8106) );
AOI22_X2 inst_9225 ( .A1(net_9919), .B1(net_9820), .A2(net_8042), .B2(net_6140), .ZN(net_6086) );
CLKBUF_X2 inst_12005 ( .A(net_11896), .Z(net_11924) );
DFF_X2 inst_7866 ( .QN(net_10101), .D(net_6019), .CK(net_15535) );
OAI21_X2 inst_1795 ( .ZN(net_7447), .B1(net_7157), .A(net_6983), .B2(net_6975) );
DFF_X2 inst_7652 ( .D(net_6707), .QN(net_183), .CK(net_15718) );
INV_X2 inst_7291 ( .A(net_9039), .ZN(net_9037) );
OR2_X4 inst_828 ( .A1(net_10366), .ZN(net_2064), .A2(net_1093) );
INV_X4 inst_4697 ( .ZN(net_4830), .A(net_4646) );
CLKBUF_X2 inst_15772 ( .A(net_15690), .Z(net_15691) );
AOI22_X2 inst_9074 ( .B1(net_9693), .A2(net_6684), .B2(net_6683), .ZN(net_6592), .A1(net_262) );
INV_X4 inst_6278 ( .A(net_9925), .ZN(net_2636) );
CLKBUF_X2 inst_13522 ( .A(net_13440), .Z(net_13441) );
INV_X2 inst_7218 ( .A(net_9591), .ZN(net_440) );
CLKBUF_X2 inst_15494 ( .A(net_12561), .Z(net_15413) );
NAND2_X2 inst_4164 ( .A1(net_4177), .ZN(net_2921), .A2(net_807) );
CLKBUF_X2 inst_10869 ( .A(net_10666), .Z(net_10788) );
CLKBUF_X2 inst_14185 ( .A(net_14103), .Z(net_14104) );
AND2_X4 inst_10408 ( .ZN(net_5360), .A2(net_4844), .A1(net_593) );
OAI221_X2 inst_1561 ( .C1(net_10231), .C2(net_7295), .B2(net_7293), .B1(net_7237), .ZN(net_7194), .A(net_6810) );
CLKBUF_X2 inst_13919 ( .A(net_13837), .Z(net_13838) );
OAI211_X2 inst_2104 ( .C2(net_6778), .ZN(net_6744), .A(net_6372), .B(net_6102), .C1(net_509) );
CLKBUF_X2 inst_12190 ( .A(net_12108), .Z(net_12109) );
DFF_X2 inst_8052 ( .QN(net_9561), .D(net_5416), .CK(net_14897) );
CLKBUF_X2 inst_12437 ( .A(net_12355), .Z(net_12356) );
CLKBUF_X2 inst_10854 ( .A(net_10772), .Z(net_10773) );
AOI22_X2 inst_9530 ( .B1(net_9890), .A1(net_9854), .A2(net_6413), .ZN(net_3791), .B2(net_2973) );
NOR2_X2 inst_2573 ( .ZN(net_7470), .A2(net_7385), .A1(net_4986) );
DFF_X1 inst_8762 ( .Q(net_9132), .D(net_5297), .CK(net_10606) );
DFF_X2 inst_7733 ( .Q(net_9898), .D(net_6221), .CK(net_11981) );
DFF_X2 inst_7382 ( .D(net_8660), .QN(net_267), .CK(net_13778) );
INV_X4 inst_6182 ( .ZN(net_7198), .A(x4209) );
DFF_X1 inst_8749 ( .Q(net_10380), .D(net_5397), .CK(net_14375) );
INV_X4 inst_6233 ( .A(net_9727), .ZN(net_1828) );
INV_X4 inst_6240 ( .A(net_9375), .ZN(net_700) );
CLKBUF_X2 inst_14760 ( .A(net_14678), .Z(net_14679) );
CLKBUF_X2 inst_11426 ( .A(net_11344), .Z(net_11345) );
AOI22_X2 inst_9629 ( .A1(net_10080), .B1(net_9999), .A2(net_5319), .ZN(net_3414), .B2(net_2468) );
AOI21_X2 inst_10127 ( .ZN(net_4305), .A(net_4001), .B2(net_2718), .B1(net_2241) );
CLKBUF_X2 inst_14564 ( .A(net_14482), .Z(net_14483) );
CLKBUF_X2 inst_10794 ( .A(net_10712), .Z(net_10713) );
AOI22_X2 inst_9137 ( .A1(net_9721), .A2(net_6418), .ZN(net_6351), .B2(net_5263), .B1(net_4183) );
OAI211_X2 inst_2096 ( .C2(net_6774), .ZN(net_6752), .A(net_6378), .B(net_6113), .C1(net_421) );
AOI21_X2 inst_10169 ( .B2(net_10302), .ZN(net_8449), .A(net_4371), .B1(net_3681) );
SDFF_X2 inst_552 ( .D(net_9154), .SE(net_7248), .SI(net_2285), .Q(net_196), .CK(net_15345) );
CLKBUF_X2 inst_10951 ( .A(net_10869), .Z(net_10870) );
NAND4_X2 inst_3050 ( .ZN(net_6156), .A4(net_5321), .A1(net_3838), .A3(net_3837), .A2(net_3579) );
INV_X4 inst_4793 ( .ZN(net_6575), .A(net_5575) );
CLKBUF_X2 inst_11349 ( .A(net_10690), .Z(net_11268) );
INV_X4 inst_4997 ( .ZN(net_4717), .A(net_2613) );
CLKBUF_X2 inst_13916 ( .A(net_13834), .Z(net_13835) );
DFF_X1 inst_8491 ( .Q(net_9634), .D(net_7900), .CK(net_11508) );
CLKBUF_X2 inst_12483 ( .A(net_12401), .Z(net_12402) );
NAND2_X2 inst_3913 ( .A1(net_4719), .A2(net_3896), .ZN(net_3889) );
OAI221_X2 inst_1564 ( .C1(net_10307), .C2(net_9047), .B2(net_7287), .B1(net_7192), .ZN(net_7189), .A(net_6789) );
INV_X4 inst_5807 ( .ZN(net_945), .A(net_901) );
INV_X2 inst_6985 ( .A(net_2060), .ZN(net_1668) );
CLKBUF_X2 inst_12625 ( .A(net_11091), .Z(net_12544) );
CLKBUF_X2 inst_10995 ( .A(net_10913), .Z(net_10914) );
DFF_X2 inst_7484 ( .Q(net_9275), .D(net_8076), .CK(net_13131) );
OAI21_X2 inst_1941 ( .B1(net_5493), .ZN(net_4285), .A(net_4000), .B2(net_3965) );
INV_X4 inst_6477 ( .A(net_9572), .ZN(net_1581) );
INV_X4 inst_6247 ( .A(net_10160), .ZN(net_851) );
DFF_X2 inst_8064 ( .QN(net_10352), .D(net_5328), .CK(net_13626) );
XOR2_X2 inst_9 ( .Z(net_3948), .B(net_3235), .A(net_2881) );
CLKBUF_X2 inst_15260 ( .A(net_12551), .Z(net_15179) );
AOI22_X2 inst_9492 ( .B1(net_10387), .A1(net_9885), .B2(net_4062), .ZN(net_3831), .A2(net_2973) );
XNOR2_X2 inst_356 ( .ZN(net_2776), .B(net_2502), .A(net_1840) );
AOI22_X2 inst_9311 ( .B1(net_9716), .A2(net_5755), .B2(net_5754), .ZN(net_5666), .A1(net_253) );
NAND2_X4 inst_3358 ( .ZN(net_8415), .A2(net_8385), .A1(net_8379) );
INV_X2 inst_6719 ( .A(net_7878), .ZN(net_7834) );
INV_X4 inst_5587 ( .ZN(net_6314), .A(net_1966) );
CLKBUF_X2 inst_10735 ( .A(net_10653), .Z(net_10654) );
INV_X2 inst_6884 ( .ZN(net_3183), .A(net_2842) );
OAI221_X2 inst_1594 ( .B1(net_10200), .C1(net_7245), .ZN(net_5646), .B2(net_5642), .C2(net_4905), .A(net_3731) );
AOI22_X2 inst_9267 ( .A1(net_6892), .B2(net_6625), .ZN(net_6208), .B1(net_5798), .A2(net_5199) );
OR2_X2 inst_902 ( .A1(net_9527), .ZN(net_5258), .A2(net_4968) );
CLKBUF_X2 inst_15810 ( .A(net_10809), .Z(net_15729) );
AOI22_X2 inst_9105 ( .A1(net_9685), .A2(net_6420), .ZN(net_6387), .B2(net_5263), .B1(net_832) );
CLKBUF_X2 inst_12224 ( .A(net_12142), .Z(net_12143) );
NAND2_X2 inst_3489 ( .ZN(net_8341), .A2(net_8340), .A1(net_8250) );
OR2_X4 inst_778 ( .ZN(net_3942), .A1(net_2956), .A2(net_2955) );
NAND2_X2 inst_4286 ( .A2(net_10355), .ZN(net_2394), .A1(net_1339) );
AOI21_X2 inst_10118 ( .B2(net_10036), .ZN(net_4780), .A(net_4474), .B1(net_627) );
OAI21_X2 inst_1935 ( .B2(net_5344), .A(net_4630), .ZN(net_4467), .B1(net_4360) );
INV_X4 inst_6032 ( .A(net_9239), .ZN(net_728) );
AOI22_X2 inst_9332 ( .B1(net_10018), .A2(net_5743), .B2(net_5742), .ZN(net_5620), .A1(net_258) );
CLKBUF_X2 inst_14949 ( .A(net_14867), .Z(net_14868) );
CLKBUF_X2 inst_14842 ( .A(net_14760), .Z(net_14761) );
DFF_X2 inst_7912 ( .Q(net_9220), .D(net_5922), .CK(net_13015) );
DFF_X1 inst_8678 ( .D(net_6722), .Q(net_145), .CK(net_13880) );
DFF_X2 inst_8235 ( .Q(net_10494), .D(net_4887), .CK(net_15215) );
CLKBUF_X2 inst_11486 ( .A(net_11404), .Z(net_11405) );
CLKBUF_X2 inst_13884 ( .A(net_13802), .Z(net_13803) );
DFF_X1 inst_8845 ( .Q(net_10539), .D(net_2264), .CK(net_12382) );
DFF_X2 inst_7810 ( .Q(net_10011), .D(net_6475), .CK(net_14757) );
OAI211_X2 inst_2140 ( .C2(net_6778), .ZN(net_6708), .A(net_6336), .B(net_6071), .C1(net_5096) );
DFF_X2 inst_8353 ( .QN(net_8844), .D(net_2883), .CK(net_12175) );
CLKBUF_X2 inst_14501 ( .A(net_14419), .Z(net_14420) );
AOI22_X2 inst_9641 ( .B1(net_9802), .A2(net_5174), .ZN(net_3337), .B2(net_2556), .A1(net_1935) );
CLKBUF_X2 inst_12855 ( .A(net_12511), .Z(net_12774) );
CLKBUF_X2 inst_13895 ( .A(net_13813), .Z(net_13814) );
OR2_X4 inst_781 ( .ZN(net_3588), .A1(net_2956), .A2(net_2540) );
CLKBUF_X2 inst_11386 ( .A(net_10736), .Z(net_11305) );
CLKBUF_X2 inst_12033 ( .A(net_11799), .Z(net_11952) );
CLKBUF_X2 inst_12368 ( .A(net_11213), .Z(net_12287) );
NAND2_X2 inst_4042 ( .A2(net_3630), .ZN(net_2843), .A1(net_2744) );
CLKBUF_X2 inst_13409 ( .A(net_11550), .Z(net_13328) );
DFF_X2 inst_7629 ( .D(net_6767), .QN(net_117), .CK(net_14324) );
AOI22_X2 inst_9450 ( .ZN(net_4375), .B2(net_4044), .B1(net_4041), .A2(net_3544), .A1(net_3090) );
NAND2_X2 inst_3696 ( .A2(net_10379), .ZN(net_7286), .A1(net_1365) );
AOI22_X2 inst_9499 ( .B1(net_9986), .A2(net_6442), .A1(net_6321), .ZN(net_3824), .B2(net_2541) );
CLKBUF_X2 inst_15648 ( .A(net_15266), .Z(net_15567) );
CLKBUF_X2 inst_13120 ( .A(net_12189), .Z(net_13039) );
AOI221_X2 inst_9971 ( .C1(net_9962), .ZN(net_4695), .B2(net_4694), .A(net_4276), .C2(net_2541), .B1(net_227) );
INV_X2 inst_7053 ( .ZN(net_1319), .A(net_1318) );
OAI221_X2 inst_1559 ( .C2(net_9047), .B2(net_7287), .B1(net_7201), .ZN(net_7196), .A(net_6798), .C1(net_5484) );
OAI21_X2 inst_1928 ( .ZN(net_4443), .A(net_4155), .B2(net_4154), .B1(net_3984) );
OAI21_X2 inst_1967 ( .B2(net_9531), .A(net_4294), .ZN(net_3264), .B1(net_2854) );
DFF_X1 inst_8830 ( .Q(net_9607), .D(net_3701), .CK(net_12907) );
CLKBUF_X2 inst_13733 ( .A(net_13651), .Z(net_13652) );
INV_X2 inst_6752 ( .A(net_9502), .ZN(net_6985) );
INV_X8 inst_4485 ( .ZN(net_8476), .A(net_8416) );
OR2_X2 inst_927 ( .A2(net_2971), .ZN(net_2965), .A1(net_2964) );
CLKBUF_X2 inst_12944 ( .A(net_12862), .Z(net_12863) );
DFF_X2 inst_7659 ( .D(net_6701), .QN(net_191), .CK(net_13212) );
CLKBUF_X2 inst_13304 ( .A(net_13222), .Z(net_13223) );
DFF_X2 inst_7420 ( .QN(net_9420), .D(net_8344), .CK(net_11691) );
CLKBUF_X2 inst_13258 ( .A(net_13176), .Z(net_13177) );
CLKBUF_X2 inst_10967 ( .A(net_10885), .Z(net_10886) );
XNOR2_X2 inst_73 ( .A(net_9083), .ZN(net_8682), .B(net_8595) );
OAI221_X2 inst_1488 ( .B1(net_10424), .C2(net_9063), .B2(net_9056), .ZN(net_7382), .C1(net_7297), .A(net_7092) );
OAI221_X2 inst_1719 ( .ZN(net_2923), .A(net_2367), .C1(net_2212), .B2(net_2210), .B1(net_1503), .C2(net_906) );
OAI21_X2 inst_1947 ( .B1(net_5480), .ZN(net_3987), .A(net_3648), .B2(net_3479) );
DFF_X2 inst_8030 ( .QN(net_10436), .D(net_5458), .CK(net_13634) );
INV_X2 inst_7318 ( .A(net_9107), .ZN(net_9104) );
INV_X4 inst_6285 ( .A(net_10095), .ZN(net_5866) );
INV_X4 inst_4690 ( .ZN(net_4837), .A(net_4653) );
AOI22_X2 inst_9236 ( .A1(net_9901), .B1(net_9802), .B2(net_6129), .A2(net_6111), .ZN(net_6075) );
OR2_X2 inst_890 ( .A1(net_10272), .ZN(net_6631), .A2(net_5969) );
CLKBUF_X2 inst_12510 ( .A(net_10570), .Z(net_12429) );
CLKBUF_X2 inst_12352 ( .A(net_12270), .Z(net_12271) );
OAI21_X2 inst_1851 ( .ZN(net_5880), .B2(net_5879), .A(net_5287), .B1(net_341) );
INV_X4 inst_5911 ( .A(net_6060), .ZN(net_591) );
INV_X4 inst_4585 ( .ZN(net_8065), .A(net_8023) );
CLKBUF_X2 inst_12896 ( .A(net_12814), .Z(net_12815) );
DFF_X2 inst_8105 ( .QN(net_10048), .D(net_5076), .CK(net_12502) );
INV_X8 inst_4514 ( .ZN(net_8854), .A(net_8853) );
CLKBUF_X2 inst_15143 ( .A(net_15061), .Z(net_15062) );
INV_X2 inst_6903 ( .A(net_7546), .ZN(net_2263) );
AOI22_X2 inst_9539 ( .B1(net_10002), .A1(net_9935), .A2(net_6443), .ZN(net_3782), .B2(net_2468) );
AOI22_X2 inst_9126 ( .A1(net_9711), .A2(net_6382), .ZN(net_6363), .B2(net_5263), .B1(net_3899) );
OAI22_X2 inst_1168 ( .A1(net_7243), .A2(net_5107), .B2(net_5105), .ZN(net_5097), .B1(net_5096) );
CLKBUF_X2 inst_15304 ( .A(net_15222), .Z(net_15223) );
CLKBUF_X2 inst_12963 ( .A(net_12881), .Z(net_12882) );
CLKBUF_X2 inst_11294 ( .A(net_11212), .Z(net_11213) );
DFF_X2 inst_7573 ( .QN(net_9383), .D(net_7590), .CK(net_13115) );
SDFF_X2 inst_659 ( .SI(net_9493), .Q(net_9493), .SE(net_3073), .CK(net_12412), .D(x1865) );
DFF_X2 inst_7681 ( .QN(net_9201), .D(net_8854), .CK(net_11338) );
INV_X2 inst_6890 ( .ZN(net_2691), .A(net_2690) );
CLKBUF_X2 inst_12868 ( .A(net_12786), .Z(net_12787) );
CLKBUF_X2 inst_11747 ( .A(net_10565), .Z(net_11666) );
CLKBUF_X2 inst_15395 ( .A(net_15313), .Z(net_15314) );
CLKBUF_X2 inst_15092 ( .A(net_15010), .Z(net_15011) );
CLKBUF_X2 inst_12883 ( .A(net_11378), .Z(net_12802) );
NAND2_X2 inst_4363 ( .A2(net_10429), .ZN(net_2002), .A1(net_779) );
OAI22_X2 inst_1161 ( .A1(net_7229), .A2(net_5139), .B2(net_5138), .ZN(net_5112), .B1(net_348) );
NAND2_X4 inst_3362 ( .A2(net_9512), .A1(net_9052), .ZN(net_7989) );
INV_X4 inst_5273 ( .ZN(net_2285), .A(net_2283) );
DFF_X2 inst_8094 ( .QN(net_9745), .D(net_5144), .CK(net_12505) );
INV_X4 inst_5505 ( .A(net_2860), .ZN(net_2298) );
AOI211_X2 inst_10289 ( .ZN(net_4674), .C2(net_4252), .A(net_3210), .C1(net_3195), .B(net_2418) );
NAND3_X2 inst_3199 ( .A3(net_9503), .ZN(net_7425), .A1(net_7424), .A2(net_7423) );
INV_X4 inst_6178 ( .ZN(net_617), .A(net_170) );
NAND2_X2 inst_3612 ( .ZN(net_7254), .A2(net_6865), .A1(net_6593) );
CLKBUF_X2 inst_15667 ( .A(net_12157), .Z(net_15586) );
OAI221_X2 inst_1581 ( .C1(net_10312), .C2(net_9047), .B2(net_7287), .B1(net_7136), .ZN(net_7126), .A(net_6933) );
CLKBUF_X2 inst_14096 ( .A(net_14014), .Z(net_14015) );
CLKBUF_X2 inst_10703 ( .A(net_10621), .Z(net_10622) );
NOR3_X2 inst_2388 ( .A1(net_7884), .A3(net_7805), .ZN(net_7802), .A2(net_1963) );
NOR4_X2 inst_2312 ( .ZN(net_7453), .A4(net_7017), .A3(net_4458), .A2(net_4096), .A1(net_3918) );
INV_X4 inst_5633 ( .ZN(net_3171), .A(net_858) );
INV_X4 inst_5336 ( .ZN(net_8747), .A(net_758) );
NAND2_X2 inst_4309 ( .A2(net_9949), .A1(net_6060), .ZN(net_4009) );
CLKBUF_X2 inst_11642 ( .A(net_11560), .Z(net_11561) );
NAND2_X2 inst_3500 ( .ZN(net_8372), .A1(net_8184), .A2(net_8183) );
NOR2_X2 inst_2634 ( .A2(net_5927), .ZN(net_5921), .A1(net_1539) );
AND2_X2 inst_10526 ( .ZN(net_4167), .A2(net_3979), .A1(net_963) );
INV_X4 inst_6381 ( .A(net_10403), .ZN(net_396) );
NAND2_X2 inst_3711 ( .A1(net_5918), .ZN(net_5911), .A2(net_5910) );
INV_X2 inst_7103 ( .A(net_10462), .ZN(net_1030) );
CLKBUF_X2 inst_13419 ( .A(net_11782), .Z(net_13338) );
OAI211_X2 inst_2241 ( .C1(net_7209), .C2(net_6480), .ZN(net_6463), .B(net_5525), .A(net_3679) );
DFF_X2 inst_8165 ( .QN(net_10031), .D(net_5052), .CK(net_13698) );
DFF_X2 inst_7568 ( .QN(net_9241), .D(net_7614), .CK(net_11262) );
OAI211_X2 inst_2182 ( .C1(net_7190), .C2(net_6548), .ZN(net_6527), .B(net_5654), .A(net_3679) );
DFF_X2 inst_8334 ( .Q(net_10490), .D(net_3556), .CK(net_12475) );
SDFF_X2 inst_650 ( .SI(net_9483), .Q(net_9483), .SE(net_3073), .CK(net_11362), .D(x2477) );
XNOR2_X2 inst_289 ( .B(net_4675), .ZN(net_3523), .A(net_3021) );
NOR2_X2 inst_2667 ( .A1(net_8565), .ZN(net_4983), .A2(net_4982) );
DFF_X1 inst_8674 ( .D(net_6747), .Q(net_106), .CK(net_11618) );
NAND2_X2 inst_4194 ( .ZN(net_1840), .A1(net_1839), .A2(net_1200) );
OAI22_X2 inst_987 ( .A2(net_8962), .B2(net_8659), .ZN(net_8653), .B1(net_6238), .A1(net_6183) );
CLKBUF_X2 inst_12467 ( .A(net_11032), .Z(net_12386) );
DFF_X1 inst_8701 ( .D(net_6749), .Q(net_103), .CK(net_13221) );
AOI22_X2 inst_9376 ( .B1(net_10013), .A2(net_5743), .B2(net_5742), .ZN(net_5529), .A1(net_253) );
DFF_X1 inst_8643 ( .Q(net_9881), .D(net_7196), .CK(net_12156) );
SDFF_X2 inst_679 ( .SI(net_9495), .Q(net_9495), .SE(net_3073), .CK(net_11869), .D(x1743) );
INV_X4 inst_5627 ( .A(net_10368), .ZN(net_2621) );
NOR2_X2 inst_3006 ( .ZN(net_4360), .A2(net_627), .A1(net_367) );
CLKBUF_X2 inst_12532 ( .A(net_12450), .Z(net_12451) );
AOI222_X1 inst_9703 ( .B1(net_9508), .A2(net_8295), .B2(net_8294), .C2(net_8293), .ZN(net_8275), .C1(net_8213), .A1(x3022) );
DFF_X2 inst_7689 ( .Q(net_10507), .D(net_6579), .CK(net_14556) );
NAND2_X4 inst_3364 ( .ZN(net_8986), .A2(net_8889), .A1(net_8888) );
OAI222_X2 inst_1351 ( .B1(net_9262), .ZN(net_7284), .A1(net_7283), .C1(net_7282), .C2(net_7281), .B2(net_7281), .A2(net_7057) );
AND2_X4 inst_10443 ( .ZN(net_2544), .A1(net_1843), .A2(net_1842) );
XOR2_X2 inst_44 ( .A(net_2849), .Z(net_1404), .B(net_1403) );
MUX2_X2 inst_4433 ( .Z(net_8960), .B(net_6423), .A(net_6344), .S(net_4448) );
CLKBUF_X2 inst_15350 ( .A(net_15268), .Z(net_15269) );
XNOR2_X2 inst_371 ( .ZN(net_2480), .A(net_2479), .B(net_1726) );
CLKBUF_X2 inst_13994 ( .A(net_10889), .Z(net_13913) );
CLKBUF_X2 inst_12805 ( .A(net_12723), .Z(net_12724) );
XNOR2_X2 inst_435 ( .A(net_9615), .ZN(net_1045), .B(net_313) );
INV_X4 inst_6498 ( .A(net_10533), .ZN(net_354) );
INV_X4 inst_4962 ( .A(net_6165), .ZN(net_2537) );
CLKBUF_X2 inst_11563 ( .A(net_11481), .Z(net_11482) );
CLKBUF_X2 inst_10768 ( .A(net_10686), .Z(net_10687) );
CLKBUF_X2 inst_10791 ( .A(net_10639), .Z(net_10710) );
AOI211_X2 inst_10305 ( .B(net_5813), .C1(net_4029), .C2(net_4024), .ZN(net_3306), .A(net_2665) );
INV_X4 inst_4619 ( .ZN(net_7134), .A(net_7014) );
CLKBUF_X2 inst_13474 ( .A(net_13392), .Z(net_13393) );
NAND2_X2 inst_3787 ( .ZN(net_4637), .A1(net_4358), .A2(net_3924) );
DFF_X2 inst_7470 ( .QN(net_9573), .D(net_8190), .CK(net_15372) );
INV_X4 inst_4982 ( .ZN(net_7697), .A(net_3916) );
SDFF_X2 inst_628 ( .Q(net_9438), .D(net_9438), .SE(net_3293), .CK(net_14658), .SI(x3249) );
NAND2_X2 inst_3684 ( .ZN(net_6665), .A2(net_5992), .A1(net_2548) );
CLKBUF_X2 inst_13633 ( .A(net_11956), .Z(net_13552) );
OAI21_X2 inst_1923 ( .B1(net_7785), .ZN(net_4542), .A(net_4242), .B2(net_4241) );
NOR2_X2 inst_2748 ( .ZN(net_4141), .A1(net_3685), .A2(x3828) );
NOR2_X2 inst_3013 ( .A1(net_9516), .A2(net_1704), .ZN(net_800) );
AOI22_X2 inst_9201 ( .A1(net_9890), .B1(net_9791), .B2(net_6120), .ZN(net_6112), .A2(net_6111) );
INV_X4 inst_4744 ( .A(net_10188), .ZN(net_5915) );
NAND2_X2 inst_3642 ( .ZN(net_9000), .A2(net_7275), .A1(net_6616) );
CLKBUF_X2 inst_11873 ( .A(net_11115), .Z(net_11792) );
INV_X4 inst_5087 ( .A(net_1900), .ZN(net_1777) );
AOI22_X2 inst_9130 ( .A1(net_9714), .A2(net_6404), .ZN(net_6358), .B2(net_5263), .B1(net_3885) );
DFF_X2 inst_7563 ( .QN(net_9246), .D(net_7612), .CK(net_11266) );
CLKBUF_X2 inst_14656 ( .A(net_12263), .Z(net_14575) );
NAND4_X2 inst_3092 ( .ZN(net_4482), .A1(net_4481), .A2(net_4480), .A3(net_4479), .A4(net_4196) );
CLKBUF_X2 inst_14162 ( .A(net_14080), .Z(net_14081) );
INV_X4 inst_6587 ( .A(net_10289), .ZN(net_324) );
CLKBUF_X2 inst_11127 ( .A(net_11045), .Z(net_11046) );
CLKBUF_X2 inst_13931 ( .A(net_13849), .Z(net_13850) );
NOR2_X2 inst_2734 ( .ZN(net_4194), .A1(net_3710), .A2(net_3709) );
INV_X4 inst_4920 ( .ZN(net_2730), .A(net_2456) );
NAND2_X2 inst_3395 ( .A1(net_9083), .A2(net_9042), .ZN(net_8670) );
CLKBUF_X2 inst_14956 ( .A(net_14874), .Z(net_14875) );
OAI22_X2 inst_1130 ( .A1(net_7139), .A2(net_5151), .B2(net_5150), .ZN(net_5148), .B1(net_471) );
CLKBUF_X2 inst_11608 ( .A(net_11526), .Z(net_11527) );
AOI22_X2 inst_9300 ( .B1(net_9908), .A2(net_5759), .B2(net_5758), .ZN(net_5678), .A1(net_247) );
INV_X4 inst_6518 ( .A(net_10099), .ZN(net_5835) );
OR2_X2 inst_855 ( .A2(net_8095), .ZN(net_8094), .A1(net_559) );
OAI211_X2 inst_2039 ( .C2(net_8102), .B(net_8098), .ZN(net_8077), .A(net_7995), .C1(net_4428) );
CLKBUF_X2 inst_15241 ( .A(net_15159), .Z(net_15160) );
CLKBUF_X2 inst_12706 ( .A(net_12624), .Z(net_12625) );
INV_X4 inst_6304 ( .A(net_10018), .ZN(net_427) );
NAND3_X2 inst_3233 ( .A1(net_5167), .A3(net_5166), .ZN(net_4759), .A2(net_613) );
DFF_X2 inst_7851 ( .Q(net_9802), .D(net_6279), .CK(net_15602) );
CLKBUF_X2 inst_15748 ( .A(net_14886), .Z(net_15667) );
AOI22_X2 inst_8996 ( .B2(net_9432), .ZN(net_8572), .A2(net_8542), .A1(net_8510), .B1(net_8412) );
CLKBUF_X2 inst_11823 ( .A(net_10942), .Z(net_11742) );
CLKBUF_X2 inst_15226 ( .A(net_11103), .Z(net_15145) );
INV_X4 inst_5866 ( .A(net_1856), .ZN(net_852) );
INV_X4 inst_5466 ( .A(net_2865), .ZN(net_1175) );
DFF_X2 inst_7588 ( .QN(net_9236), .D(net_7529), .CK(net_11255) );
INV_X4 inst_5425 ( .ZN(net_2612), .A(net_648) );
AOI21_X2 inst_10160 ( .ZN(net_4008), .A(net_4007), .B2(net_3339), .B1(net_1387) );
AOI22_X2 inst_9304 ( .B1(net_9710), .A2(net_5755), .B2(net_5754), .ZN(net_5674), .A1(net_247) );
NAND2_X2 inst_4295 ( .A2(net_10224), .ZN(net_4412), .A1(net_2628) );
SDFF_X2 inst_518 ( .Q(net_9333), .D(net_9333), .SI(net_9158), .SE(net_7588), .CK(net_13078) );
OAI222_X2 inst_1363 ( .B1(net_7660), .A2(net_7659), .C2(net_7658), .ZN(net_6326), .B2(net_5399), .A1(net_4064), .C1(net_1899) );
INV_X4 inst_4851 ( .ZN(net_3872), .A(net_3287) );
INV_X4 inst_5894 ( .ZN(net_875), .A(net_608) );
DFF_X2 inst_8242 ( .Q(net_10072), .D(net_4864), .CK(net_10729) );
NAND2_X2 inst_3863 ( .ZN(net_4112), .A2(net_3938), .A1(net_2019) );
NOR4_X2 inst_2345 ( .A2(net_9179), .ZN(net_2787), .A1(net_2786), .A3(net_2785), .A4(net_2092) );
DFF_X2 inst_8059 ( .D(net_5279), .CK(net_14892), .Q(x494) );
CLKBUF_X2 inst_12157 ( .A(net_12075), .Z(net_12076) );
INV_X4 inst_6538 ( .ZN(net_6408), .A(net_182) );
NAND2_X2 inst_3602 ( .ZN(net_7264), .A1(net_6883), .A2(net_6559) );
AOI22_X2 inst_9614 ( .A1(net_10086), .B1(net_10012), .A2(net_5319), .ZN(net_3439), .B2(net_2468) );
CLKBUF_X2 inst_12388 ( .A(net_11161), .Z(net_12307) );
CLKBUF_X2 inst_14291 ( .A(net_12632), .Z(net_14210) );
DFF_X2 inst_7582 ( .Q(net_10295), .D(net_7534), .CK(net_14563) );
INV_X4 inst_5260 ( .ZN(net_1398), .A(net_1397) );
CLKBUF_X2 inst_12637 ( .A(net_10926), .Z(net_12556) );
CLKBUF_X2 inst_11815 ( .A(net_11733), .Z(net_11734) );
CLKBUF_X2 inst_11372 ( .A(net_11191), .Z(net_11291) );
CLKBUF_X2 inst_12336 ( .A(net_10973), .Z(net_12255) );
INV_X4 inst_5190 ( .A(net_1562), .ZN(net_1547) );
OAI222_X2 inst_1354 ( .B1(net_7665), .A2(net_7664), .C2(net_7663), .ZN(net_7160), .B2(net_6647), .A1(net_4416), .C1(net_714) );
CLKBUF_X2 inst_11806 ( .A(net_11682), .Z(net_11725) );
OAI33_X1 inst_970 ( .B2(net_9172), .ZN(net_3166), .A1(net_3165), .B3(net_2761), .B1(net_2239), .A2(net_1959), .A3(net_1878) );
CLKBUF_X2 inst_15736 ( .A(net_15654), .Z(net_15655) );
CLKBUF_X2 inst_11992 ( .A(net_11910), .Z(net_11911) );
INV_X2 inst_6731 ( .ZN(net_7549), .A(net_7508) );
OAI22_X2 inst_1278 ( .B2(net_7671), .A1(net_7602), .ZN(net_4458), .B1(net_4095), .A2(net_3877) );
NAND2_X2 inst_3763 ( .ZN(net_5259), .A2(net_4984), .A1(net_870) );
AOI21_X2 inst_10136 ( .ZN(net_4250), .B2(net_3620), .B1(net_3130), .A(net_2717) );
OR2_X4 inst_749 ( .ZN(net_5296), .A2(net_5178), .A1(net_4479) );
CLKBUF_X2 inst_15159 ( .A(net_15077), .Z(net_15078) );
CLKBUF_X2 inst_11975 ( .A(net_11742), .Z(net_11894) );
INV_X2 inst_6688 ( .ZN(net_8336), .A(net_8274) );
OAI22_X2 inst_1030 ( .ZN(net_7907), .A2(net_7906), .B1(net_7905), .B2(net_7904), .A1(net_6581) );
OAI211_X2 inst_2127 ( .C2(net_6778), .ZN(net_6721), .A(net_6348), .B(net_6084), .C1(net_333) );
CLKBUF_X2 inst_13689 ( .A(net_13607), .Z(net_13608) );
CLKBUF_X2 inst_13626 ( .A(net_13544), .Z(net_13545) );
AND2_X2 inst_10611 ( .A1(net_4029), .A2(net_3121), .ZN(net_2663) );
NOR2_X2 inst_2649 ( .A2(net_9598), .ZN(net_8192), .A1(net_7846) );
CLKBUF_X2 inst_11441 ( .A(net_11359), .Z(net_11360) );
OAI222_X2 inst_1373 ( .B2(net_7660), .A2(net_7659), .C2(net_7658), .ZN(net_6035), .B1(net_2776), .A1(net_2274), .C1(net_1087) );
OAI211_X2 inst_2268 ( .C1(net_7127), .C2(net_6501), .ZN(net_6277), .B(net_5699), .A(net_3679) );
NOR3_X2 inst_2458 ( .A2(net_3899), .A3(net_3894), .A1(net_1708), .ZN(net_1423) );
NAND2_X2 inst_3828 ( .A1(net_8860), .ZN(net_4447), .A2(net_4440) );
INV_X2 inst_7285 ( .A(net_8979), .ZN(net_8978) );
CLKBUF_X2 inst_14303 ( .A(net_11359), .Z(net_14222) );
DFF_X1 inst_8474 ( .QN(net_10361), .D(net_7842), .CK(net_12235) );
INV_X4 inst_5841 ( .ZN(net_3598), .A(net_653) );
AOI221_X2 inst_9923 ( .B2(net_5867), .ZN(net_5860), .A(net_5859), .C1(net_5858), .C2(net_4725), .B1(x5364) );
INV_X2 inst_6898 ( .ZN(net_3255), .A(net_2582) );
NAND4_X2 inst_3155 ( .ZN(net_1897), .A2(net_977), .A3(net_138), .A4(net_137), .A1(net_134) );
INV_X4 inst_5481 ( .A(net_10145), .ZN(net_1153) );
NAND4_X2 inst_3134 ( .ZN(net_2916), .A4(net_2913), .A3(net_2902), .A2(net_2901), .A1(net_1661) );
OAI22_X2 inst_1006 ( .A1(net_8327), .B2(net_8325), .ZN(net_8324), .A2(net_8235), .B1(net_6626) );
OAI21_X2 inst_1985 ( .ZN(net_2795), .B1(net_2794), .A(net_2118), .B2(net_1859) );
INV_X2 inst_7311 ( .A(net_9090), .ZN(net_9089) );
CLKBUF_X2 inst_14878 ( .A(net_14796), .Z(net_14797) );
CLKBUF_X2 inst_13519 ( .A(net_13437), .Z(net_13438) );
CLKBUF_X2 inst_11787 ( .A(net_11705), .Z(net_11706) );
INV_X2 inst_6710 ( .ZN(net_8114), .A(net_8113) );
NAND2_X2 inst_4043 ( .ZN(net_4275), .A1(net_4080), .A2(net_3630) );
AND2_X4 inst_10473 ( .A2(net_10468), .A1(net_10467), .ZN(net_2017) );
AOI221_X2 inst_9817 ( .B1(net_9875), .B2(net_9101), .ZN(net_6946), .A(net_6945), .C1(net_6944), .C2(net_246) );
INV_X4 inst_5134 ( .A(net_1958), .ZN(net_1878) );
DFF_X1 inst_8407 ( .D(net_8814), .CK(net_11935), .Q(x747) );
INV_X2 inst_7180 ( .A(net_10454), .ZN(net_866) );
CLKBUF_X2 inst_11999 ( .A(net_11917), .Z(net_11918) );
INV_X4 inst_5755 ( .ZN(net_1013), .A(net_732) );
CLKBUF_X2 inst_11933 ( .A(net_10794), .Z(net_11852) );
DFF_X1 inst_8691 ( .D(net_6779), .QN(net_181), .CK(net_12001) );
INV_X4 inst_4753 ( .ZN(net_4905), .A(net_4231) );
CLKBUF_X2 inst_10960 ( .A(net_10878), .Z(net_10879) );
DFF_X2 inst_8122 ( .QN(net_9744), .D(net_5110), .CK(net_12893) );
CLKBUF_X2 inst_11885 ( .A(net_11803), .Z(net_11804) );
AOI21_X2 inst_10082 ( .B1(net_9527), .ZN(net_5403), .A(net_5232), .B2(net_4968) );
CLKBUF_X2 inst_11957 ( .A(net_10728), .Z(net_11876) );
INV_X4 inst_4947 ( .ZN(net_2568), .A(net_2567) );
CLKBUF_X2 inst_15077 ( .A(net_14995), .Z(net_14996) );
CLKBUF_X2 inst_13435 ( .A(net_13353), .Z(net_13354) );
CLKBUF_X2 inst_15728 ( .A(net_15646), .Z(net_15647) );
CLKBUF_X2 inst_11671 ( .A(net_11589), .Z(net_11590) );
CLKBUF_X2 inst_12349 ( .A(net_12267), .Z(net_12268) );
INV_X4 inst_5783 ( .ZN(net_1037), .A(net_702) );
CLKBUF_X2 inst_12490 ( .A(net_12408), .Z(net_12409) );
CLKBUF_X2 inst_15701 ( .A(net_15619), .Z(net_15620) );
CLKBUF_X2 inst_12755 ( .A(net_12673), .Z(net_12674) );
INV_X4 inst_6457 ( .A(net_10126), .ZN(net_5839) );
INV_X4 inst_4588 ( .ZN(net_8062), .A(net_8020) );
CLKBUF_X2 inst_13746 ( .A(net_12640), .Z(net_13665) );
AOI22_X2 inst_9099 ( .A1(net_9680), .A2(net_6420), .ZN(net_6393), .B2(net_5263), .B1(net_4033) );
AOI221_X2 inst_9898 ( .B1(net_9883), .B2(net_9101), .A(net_6945), .C2(net_6944), .C1(net_6823), .ZN(net_6796) );
NAND2_X2 inst_4184 ( .ZN(net_2408), .A1(net_2183), .A2(net_1396) );
NAND2_X2 inst_4049 ( .ZN(net_3014), .A2(net_2811), .A1(net_1597) );
INV_X4 inst_5067 ( .A(net_3085), .ZN(net_1858) );
NOR2_X2 inst_2702 ( .ZN(net_4802), .A2(net_4375), .A1(net_2841) );
CLKBUF_X2 inst_15063 ( .A(net_12376), .Z(net_14982) );
CLKBUF_X2 inst_12820 ( .A(net_12016), .Z(net_12739) );
INV_X4 inst_6531 ( .A(net_9975), .ZN(net_340) );
NOR2_X2 inst_2910 ( .A1(net_3528), .A2(net_2465), .ZN(net_2066) );
CLKBUF_X2 inst_11517 ( .A(net_11435), .Z(net_11436) );
INV_X4 inst_4670 ( .A(net_9270), .ZN(net_6582) );
CLKBUF_X2 inst_15178 ( .A(net_14322), .Z(net_15097) );
INV_X4 inst_5701 ( .ZN(net_780), .A(net_779) );
NAND3_X2 inst_3238 ( .A1(net_7142), .A3(net_4719), .ZN(net_4718), .A2(net_4717) );
XNOR2_X2 inst_145 ( .ZN(net_7032), .B(net_7031), .A(net_6174) );
CLKBUF_X2 inst_13703 ( .A(net_12339), .Z(net_13622) );
NOR2_X2 inst_2854 ( .ZN(net_3453), .A1(net_2169), .A2(net_2168) );
NOR2_X1 inst_3030 ( .ZN(net_2611), .A1(net_2608), .A2(net_1314) );
DFF_X2 inst_7717 ( .Q(net_9905), .D(net_6362), .CK(net_12573) );
INV_X4 inst_4594 ( .ZN(net_7899), .A(net_7827) );
OAI211_X2 inst_2230 ( .A(net_8098), .C1(net_7201), .C2(net_6480), .ZN(net_6474), .B(net_5600) );
AOI222_X1 inst_9689 ( .B1(net_9508), .A2(net_8301), .B2(net_8300), .C2(net_8299), .ZN(net_8292), .C1(net_8222), .A1(x2027) );
INV_X4 inst_5355 ( .ZN(net_5480), .A(net_1637) );
INV_X4 inst_5630 ( .A(net_2862), .ZN(net_2016) );
CLKBUF_X2 inst_15223 ( .A(net_15141), .Z(net_15142) );
CLKBUF_X2 inst_13028 ( .A(net_12946), .Z(net_12947) );
INV_X4 inst_6214 ( .A(net_9317), .ZN(net_7677) );
AOI21_X2 inst_10199 ( .ZN(net_2884), .B1(net_1800), .A(net_1630), .B2(net_1517) );
AND2_X2 inst_10511 ( .ZN(net_4919), .A1(net_4918), .A2(net_4917) );
CLKBUF_X2 inst_12240 ( .A(net_12158), .Z(net_12159) );
INV_X4 inst_5345 ( .ZN(net_1242), .A(net_955) );
OAI222_X1 inst_1437 ( .ZN(net_7788), .A1(net_7665), .B2(net_7664), .C2(net_7663), .A2(net_7652), .B1(net_5762), .C1(net_1140) );
CLKBUF_X2 inst_13820 ( .A(net_10848), .Z(net_13739) );
AND2_X2 inst_10481 ( .A2(net_9577), .ZN(net_8602), .A1(net_1384) );
CLKBUF_X2 inst_14964 ( .A(net_14882), .Z(net_14883) );
AOI22_X2 inst_9292 ( .B1(net_9802), .A1(net_5766), .B2(net_5765), .ZN(net_5705), .A2(net_240) );
AOI22_X2 inst_9119 ( .A1(net_9704), .A2(net_6404), .ZN(net_6370), .B2(net_5263), .B1(net_144) );
CLKBUF_X2 inst_14174 ( .A(net_14092), .Z(net_14093) );
AND2_X2 inst_10557 ( .A1(net_9655), .ZN(net_3650), .A2(net_3307) );
CLKBUF_X2 inst_13661 ( .A(net_13349), .Z(net_13580) );
MUX2_X1 inst_4477 ( .S(net_6041), .A(net_3933), .B(net_1591), .Z(x420) );
NOR2_X2 inst_2533 ( .A2(net_9596), .A1(net_9073), .ZN(net_8317) );
NOR3_X2 inst_2391 ( .A2(net_8837), .A1(net_8816), .ZN(net_7763), .A3(net_7624) );
DFF_X2 inst_7606 ( .QN(net_10253), .D(net_7160), .CK(net_11670) );
CLKBUF_X2 inst_14837 ( .A(net_13305), .Z(net_14756) );
OAI211_X2 inst_2239 ( .C1(net_7216), .C2(net_6480), .ZN(net_6465), .B(net_5527), .A(net_3679) );
CLKBUF_X2 inst_15601 ( .A(net_15519), .Z(net_15520) );
XOR2_X2 inst_27 ( .Z(net_2172), .B(net_1740), .A(net_1294) );
AOI21_X2 inst_10027 ( .B1(net_9367), .A(net_7916), .B2(net_7915), .ZN(net_7852) );
CLKBUF_X2 inst_10741 ( .A(net_10659), .Z(net_10660) );
DFF_X1 inst_8790 ( .Q(net_10448), .D(net_4372), .CK(net_11071) );
INV_X4 inst_6335 ( .A(net_9979), .ZN(net_412) );
OAI221_X2 inst_1639 ( .B1(net_10420), .C1(net_7127), .A(net_5637), .ZN(net_5549), .B2(net_4477), .C2(net_4455) );
CLKBUF_X2 inst_14849 ( .A(net_14767), .Z(net_14768) );
MUX2_X1 inst_4446 ( .S(net_6041), .A(net_300), .B(x4851), .Z(x111) );
CLKBUF_X2 inst_13645 ( .A(net_13563), .Z(net_13564) );
CLKBUF_X2 inst_11468 ( .A(net_10746), .Z(net_11387) );
CLKBUF_X2 inst_10717 ( .A(net_10635), .Z(net_10636) );
CLKBUF_X2 inst_11761 ( .A(net_11380), .Z(net_11680) );
AOI21_X2 inst_10063 ( .ZN(net_7028), .A(net_7027), .B1(net_5187), .B2(net_4930) );
CLKBUF_X2 inst_15443 ( .A(net_15361), .Z(net_15362) );
CLKBUF_X2 inst_14743 ( .A(net_14661), .Z(net_14662) );
INV_X4 inst_5155 ( .ZN(net_1892), .A(net_1396) );
AND3_X2 inst_10365 ( .A1(net_8098), .ZN(net_8075), .A3(net_8074), .A2(net_2458) );
CLKBUF_X2 inst_11071 ( .A(net_10989), .Z(net_10990) );
CLKBUF_X2 inst_15807 ( .A(net_15725), .Z(net_15726) );
CLKBUF_X2 inst_15397 ( .A(net_13237), .Z(net_15316) );
AOI221_X2 inst_9756 ( .ZN(net_7750), .A(net_7749), .B2(net_7748), .C2(net_7747), .C1(net_7683), .B1(net_1450) );
DFF_X2 inst_7403 ( .Q(net_9575), .D(net_8409), .CK(net_11609) );
INV_X4 inst_6420 ( .ZN(net_4029), .A(net_125) );
INV_X4 inst_5230 ( .A(net_1578), .ZN(net_1488) );
AOI22_X2 inst_9045 ( .ZN(net_7170), .A1(net_6892), .B2(net_6625), .B1(net_6040), .A2(net_5948) );
SDFF_X2 inst_639 ( .Q(net_9439), .D(net_9439), .SE(net_3293), .CK(net_14154), .SI(x3194) );
XNOR2_X2 inst_155 ( .ZN(net_6266), .A(net_5990), .B(net_2514) );
CLKBUF_X2 inst_14687 ( .A(net_13794), .Z(net_14606) );
INV_X4 inst_4858 ( .ZN(net_4097), .A(net_3181) );
AOI21_X2 inst_10170 ( .ZN(net_4111), .B2(net_3469), .A(net_2937), .B1(net_2732) );
NAND2_X2 inst_3939 ( .A1(net_9916), .A2(net_4969), .ZN(net_3551) );
INV_X4 inst_6043 ( .A(net_10021), .ZN(net_512) );
INV_X4 inst_5309 ( .A(net_2882), .ZN(net_1291) );
XOR2_X1 inst_55 ( .A(net_9347), .Z(net_1991), .B(net_1990) );
OAI211_X2 inst_2167 ( .C1(net_7294), .ZN(net_6543), .C2(net_6542), .B(net_5767), .A(net_3679) );
OAI211_X2 inst_2280 ( .C1(net_7136), .C2(net_6501), .ZN(net_6218), .B(net_5740), .A(net_3679) );
INV_X2 inst_7008 ( .ZN(net_1608), .A(net_1552) );
CLKBUF_X2 inst_12193 ( .A(net_12111), .Z(net_12112) );
DFF_X2 inst_7412 ( .QN(net_9404), .D(net_8361), .CK(net_13951) );
INV_X4 inst_6328 ( .A(net_9304), .ZN(net_415) );
AOI221_X2 inst_9872 ( .B1(net_9780), .B2(net_9098), .A(net_6940), .C2(net_6939), .ZN(net_6830), .C1(net_250) );
INV_X2 inst_7097 ( .A(net_4918), .ZN(net_1082) );
CLKBUF_X2 inst_12561 ( .A(net_12479), .Z(net_12480) );
NAND2_X2 inst_4248 ( .ZN(net_1434), .A1(net_1433), .A2(net_1432) );
OAI221_X2 inst_1651 ( .C1(net_10418), .B1(net_7249), .ZN(net_5535), .C2(net_4477), .B2(net_4455), .A(net_3507) );
CLKBUF_X2 inst_12176 ( .A(net_11980), .Z(net_12095) );
AOI221_X2 inst_9758 ( .A(net_7749), .B2(net_7748), .C2(net_7747), .ZN(net_7744), .C1(net_7679), .B1(net_430) );
DFF_X2 inst_8281 ( .Q(net_10393), .D(net_4811), .CK(net_13160) );
NAND2_X2 inst_4127 ( .ZN(net_5284), .A2(net_2321), .A1(net_2320) );
CLKBUF_X2 inst_15695 ( .A(net_12760), .Z(net_15614) );
CLKBUF_X2 inst_11634 ( .A(net_11552), .Z(net_11553) );
CLKBUF_X2 inst_11159 ( .A(net_11077), .Z(net_11078) );
INV_X4 inst_6451 ( .A(net_9989), .ZN(net_375) );
OAI22_X2 inst_1137 ( .A1(net_7245), .ZN(net_5140), .A2(net_5139), .B2(net_5138), .B1(net_327) );
CLKBUF_X2 inst_15254 ( .A(net_15172), .Z(net_15173) );
XNOR2_X2 inst_323 ( .B(net_3704), .ZN(net_3030), .A(net_2830) );
OAI222_X2 inst_1389 ( .B1(net_7728), .A2(net_7727), .C2(net_7726), .ZN(net_5822), .B2(net_4938), .A1(net_3418), .C1(net_654) );
AOI22_X2 inst_9032 ( .B2(net_10486), .ZN(net_7625), .A2(net_7494), .A1(net_7408), .B1(net_863) );
CLKBUF_X2 inst_14043 ( .A(net_13961), .Z(net_13962) );
NAND4_X2 inst_3065 ( .ZN(net_5715), .A4(net_4898), .A1(net_3820), .A2(net_3784), .A3(net_3768) );
OR3_X2 inst_715 ( .A3(net_9039), .A1(net_7589), .ZN(net_3991), .A2(net_1010) );
OAI221_X2 inst_1494 ( .B1(net_10441), .C2(net_9063), .B2(net_9056), .ZN(net_7369), .C1(net_7237), .A(net_6990) );
CLKBUF_X2 inst_14936 ( .A(net_14854), .Z(net_14855) );
INV_X4 inst_5206 ( .A(net_1537), .ZN(net_1527) );
HA_X1 inst_7333 ( .S(net_7465), .CO(net_7464), .B(net_7310), .A(net_995) );
INV_X4 inst_6354 ( .A(net_9230), .ZN(net_406) );
INV_X4 inst_5213 ( .A(net_6839), .ZN(net_1522) );
CLKBUF_X2 inst_14113 ( .A(net_14031), .Z(net_14032) );
NAND2_X2 inst_3525 ( .A1(net_9556), .ZN(net_8132), .A2(net_8095) );
CLKBUF_X2 inst_12734 ( .A(net_12228), .Z(net_12653) );
AND2_X2 inst_10479 ( .ZN(net_8715), .A1(net_8714), .A2(net_8713) );
NAND2_X2 inst_3449 ( .A1(net_9462), .ZN(net_8904), .A2(net_8475) );
OAI221_X2 inst_1682 ( .C1(net_7229), .B2(net_5591), .ZN(net_5483), .B1(net_5482), .C2(net_4902), .A(net_3731) );
INV_X4 inst_5077 ( .ZN(net_2163), .A(net_1827) );
OAI222_X2 inst_1340 ( .A1(net_7660), .B2(net_7659), .C2(net_7658), .ZN(net_7607), .A2(net_7465), .B1(net_5183), .C1(net_1224) );
OAI221_X2 inst_1481 ( .B2(net_7671), .ZN(net_7603), .C2(net_7602), .A(net_7513), .C1(net_4512), .B1(net_3543) );
CLKBUF_X2 inst_14275 ( .A(net_14193), .Z(net_14194) );
CLKBUF_X2 inst_13778 ( .A(net_12010), .Z(net_13697) );
CLKBUF_X2 inst_10630 ( .A(net_10548), .Z(net_10549) );
CLKBUF_X2 inst_14785 ( .A(net_10889), .Z(net_14704) );
CLKBUF_X2 inst_13194 ( .A(net_13112), .Z(net_13113) );
AOI21_X2 inst_10191 ( .ZN(net_3277), .A(net_2836), .B1(net_2622), .B2(net_2176) );
DFF_X2 inst_7794 ( .Q(net_9908), .D(net_6500), .CK(net_13269) );
CLKBUF_X2 inst_13349 ( .A(net_13267), .Z(net_13268) );
CLKBUF_X2 inst_15136 ( .A(net_10611), .Z(net_15055) );
XOR2_X2 inst_31 ( .Z(net_2123), .B(net_2122), .A(net_1426) );
NAND2_X2 inst_3505 ( .ZN(net_8340), .A1(net_8175), .A2(net_8174) );
AOI22_X2 inst_9355 ( .B1(net_9909), .A2(net_5759), .B2(net_5758), .ZN(net_5567), .A1(net_248) );
DFF_X1 inst_8788 ( .QN(net_9190), .D(net_4293), .CK(net_13609) );
AOI21_X2 inst_10128 ( .ZN(net_4295), .B1(net_4294), .A(net_4089), .B2(net_3295) );
DFF_X2 inst_7707 ( .Q(net_10002), .D(net_6292), .CK(net_13872) );
CLKBUF_X2 inst_15751 ( .A(net_15669), .Z(net_15670) );
AOI21_X2 inst_10204 ( .B1(net_7583), .ZN(net_2635), .A(net_2634), .B2(net_2612) );
NAND3_X2 inst_3217 ( .ZN(net_5688), .A1(net_5177), .A3(net_3416), .A2(net_3403) );
AOI22_X2 inst_9556 ( .B1(net_10505), .A1(net_9663), .B2(net_6415), .A2(net_5966), .ZN(net_3764) );
CLKBUF_X2 inst_10937 ( .A(net_10855), .Z(net_10856) );
INV_X4 inst_6440 ( .A(net_9943), .ZN(net_1418) );
CLKBUF_X2 inst_14506 ( .A(net_14424), .Z(net_14425) );
CLKBUF_X2 inst_12730 ( .A(net_12648), .Z(net_12649) );
AOI221_X2 inst_9787 ( .B1(net_9964), .A(net_7090), .B2(net_7089), .C1(net_7088), .ZN(net_7076), .C2(net_236) );
NAND2_X2 inst_4376 ( .ZN(net_2072), .A2(net_1031), .A1(net_851) );
NAND2_X2 inst_3537 ( .ZN(net_8997), .A1(net_8047), .A2(net_2369) );
CLKBUF_X2 inst_12606 ( .A(net_12524), .Z(net_12525) );
INV_X4 inst_4556 ( .A(net_9576), .ZN(net_8535) );
CLKBUF_X2 inst_14449 ( .A(net_11895), .Z(net_14368) );
CLKBUF_X2 inst_11778 ( .A(net_11696), .Z(net_11697) );
INV_X4 inst_6023 ( .A(net_9291), .ZN(net_1733) );
OAI21_X2 inst_1833 ( .B2(net_10135), .ZN(net_6329), .A(net_1437), .B1(net_658) );
DFF_X2 inst_8160 ( .QN(net_10033), .D(net_5062), .CK(net_13300) );
INV_X4 inst_5301 ( .ZN(net_5051), .A(net_3799) );
OAI211_X2 inst_2122 ( .C2(net_6778), .ZN(net_6726), .A(net_6353), .B(net_6088), .C1(net_368) );
NAND4_X2 inst_3044 ( .ZN(net_7476), .A2(net_7286), .A4(net_7285), .A3(net_6644), .A1(net_3127) );
INV_X4 inst_5443 ( .A(net_1221), .ZN(net_1095) );
NAND2_X2 inst_3520 ( .A2(net_9593), .A1(net_9089), .ZN(net_8320) );
CLKBUF_X2 inst_14493 ( .A(net_14411), .Z(net_14412) );
CLKBUF_X2 inst_11601 ( .A(net_11519), .Z(net_11520) );
AOI221_X2 inst_9809 ( .B1(net_9988), .A(net_7090), .B2(net_7089), .C2(net_7088), .ZN(net_6993), .C1(net_260) );
CLKBUF_X2 inst_13041 ( .A(net_11364), .Z(net_12960) );
CLKBUF_X2 inst_11914 ( .A(net_11832), .Z(net_11833) );
NAND2_X2 inst_3573 ( .A1(net_8801), .ZN(net_8635), .A2(net_7592) );
CLKBUF_X2 inst_13453 ( .A(net_13371), .Z(net_13372) );
CLKBUF_X2 inst_12324 ( .A(net_11912), .Z(net_12243) );
CLKBUF_X2 inst_11306 ( .A(net_11224), .Z(net_11225) );
SDFF_X2 inst_623 ( .Q(net_9441), .D(net_9441), .SE(net_3293), .CK(net_14162), .SI(x3071) );
CLKBUF_X2 inst_15612 ( .A(net_13090), .Z(net_15531) );
OAI22_X2 inst_1072 ( .ZN(net_6849), .A2(net_6848), .B1(net_6847), .B2(net_6846), .A1(net_6560) );
DFF_X1 inst_8557 ( .Q(net_8836), .D(net_7399), .CK(net_14400) );
OAI221_X2 inst_1621 ( .B1(net_10318), .C1(net_7211), .B2(net_5591), .ZN(net_5586), .C2(net_4902), .A(net_3507) );
OAI21_X2 inst_1993 ( .B1(net_5484), .ZN(net_2493), .A(net_2116), .B2(net_1864) );
AND3_X2 inst_10373 ( .ZN(net_5358), .A1(net_4667), .A3(net_4640), .A2(net_4365) );
CLKBUF_X2 inst_15744 ( .A(net_15662), .Z(net_15663) );
CLKBUF_X2 inst_14877 ( .A(net_13978), .Z(net_14796) );
CLKBUF_X2 inst_14193 ( .A(net_14111), .Z(net_14112) );
AOI221_X2 inst_9791 ( .B1(net_9967), .A(net_7090), .B2(net_7089), .C1(net_7088), .ZN(net_7034), .C2(net_239) );
NAND3_X2 inst_3226 ( .ZN(net_5228), .A3(net_4943), .A1(net_4942), .A2(net_2896) );
CLKBUF_X2 inst_15439 ( .A(net_15357), .Z(net_15358) );
INV_X2 inst_6671 ( .ZN(net_8357), .A(net_8297) );
CLKBUF_X2 inst_10674 ( .A(net_10592), .Z(net_10593) );
DFF_X1 inst_8435 ( .QN(net_9580), .D(net_8618), .CK(net_11553) );
CLKBUF_X2 inst_15580 ( .A(net_15498), .Z(net_15499) );
AOI22_X2 inst_9609 ( .A1(net_10083), .B1(net_10009), .A2(net_5319), .ZN(net_3444), .B2(net_2468) );
CLKBUF_X2 inst_13224 ( .A(net_13142), .Z(net_13143) );
INV_X4 inst_6470 ( .A(net_10361), .ZN(net_7479) );
NAND2_X2 inst_3617 ( .ZN(net_7318), .A2(net_7085), .A1(net_6894) );
CLKBUF_X2 inst_10893 ( .A(net_10811), .Z(net_10812) );
OAI222_X2 inst_1377 ( .B2(net_7660), .A2(net_7659), .C2(net_7658), .ZN(net_6008), .B1(net_3008), .A1(net_2409), .C1(net_1387) );
CLKBUF_X2 inst_15523 ( .A(net_13409), .Z(net_15442) );
CLKBUF_X2 inst_15513 ( .A(net_15431), .Z(net_15432) );
NAND4_X2 inst_3125 ( .ZN(net_3125), .A3(net_2603), .A2(net_2386), .A1(net_1791), .A4(net_1790) );
CLKBUF_X2 inst_14828 ( .A(net_14746), .Z(net_14747) );
AND2_X2 inst_10571 ( .ZN(net_3469), .A2(net_3004), .A1(net_1634) );
OAI211_X2 inst_2201 ( .C1(net_7209), .C2(net_6542), .ZN(net_6506), .B(net_5604), .A(net_3679) );
CLKBUF_X2 inst_14130 ( .A(net_14048), .Z(net_14049) );
AND2_X2 inst_10581 ( .A1(net_2782), .ZN(net_2662), .A2(net_2661) );
CLKBUF_X2 inst_10750 ( .A(net_10668), .Z(net_10669) );
AND2_X2 inst_10562 ( .A1(net_4177), .ZN(net_3083), .A2(net_2225) );
OR2_X4 inst_760 ( .ZN(net_5107), .A1(net_4475), .A2(net_4366) );
CLKBUF_X2 inst_14144 ( .A(net_10768), .Z(net_14063) );
CLKBUF_X2 inst_12842 ( .A(net_10715), .Z(net_12761) );
CLKBUF_X2 inst_10814 ( .A(net_10732), .Z(net_10733) );
DFF_X1 inst_8867 ( .D(net_10519), .CK(net_12658), .Q(x447) );
INV_X4 inst_5671 ( .ZN(net_6956), .A(net_813) );
OAI221_X2 inst_1696 ( .C1(net_7221), .B2(net_5642), .A(net_5575), .ZN(net_5460), .B1(net_5459), .C2(net_4905) );
CLKBUF_X2 inst_14519 ( .A(net_11761), .Z(net_14438) );
AOI22_X2 inst_9347 ( .B1(net_9795), .A1(net_6813), .A2(net_5766), .B2(net_5765), .ZN(net_5605) );
INV_X4 inst_4911 ( .A(net_3101), .ZN(net_2836) );
INV_X8 inst_4525 ( .ZN(net_8966), .A(net_8058) );
NAND2_X2 inst_4115 ( .ZN(net_2351), .A2(net_1603), .A1(net_1104) );
CLKBUF_X2 inst_13264 ( .A(net_13182), .Z(net_13183) );
AOI221_X2 inst_9831 ( .ZN(net_6890), .A(net_6889), .B2(net_6888), .C2(net_6887), .B1(net_5864), .C1(x5498) );
DFF_X2 inst_8174 ( .QN(net_9828), .D(net_5035), .CK(net_14443) );
NAND2_X2 inst_3727 ( .A1(net_8511), .ZN(net_5735), .A2(net_5734) );
CLKBUF_X2 inst_12237 ( .A(net_12155), .Z(net_12156) );
CLKBUF_X2 inst_10812 ( .A(net_10595), .Z(net_10731) );
DFF_X1 inst_8417 ( .QN(net_9377), .D(net_8787), .CK(net_11929) );
INV_X4 inst_5591 ( .ZN(net_1327), .A(net_883) );
INV_X2 inst_7258 ( .A(net_9314), .ZN(net_7683) );
OAI221_X2 inst_1687 ( .C1(net_7229), .ZN(net_5474), .B1(net_5473), .B2(net_4477), .C2(net_4455), .A(net_3507) );
CLKBUF_X2 inst_14983 ( .A(net_14901), .Z(net_14902) );
OAI21_X2 inst_1970 ( .B1(net_5459), .ZN(net_3253), .A(net_3014), .B2(net_2811) );
NAND2_X2 inst_3989 ( .A1(net_9792), .ZN(net_3185), .A2(net_2462) );
INV_X2 inst_7137 ( .A(net_1437), .ZN(net_830) );
CLKBUF_X2 inst_14973 ( .A(net_14891), .Z(net_14892) );
CLKBUF_X2 inst_12211 ( .A(net_12129), .Z(net_12130) );
AOI21_X4 inst_10000 ( .B2(net_8994), .B1(net_8993), .ZN(net_7608), .A(net_7427) );
CLKBUF_X2 inst_12934 ( .A(net_12852), .Z(net_12853) );
INV_X2 inst_6790 ( .ZN(net_5782), .A(net_5396) );
CLKBUF_X2 inst_14100 ( .A(net_14018), .Z(net_14019) );
AOI211_X2 inst_10256 ( .A(net_8190), .ZN(net_8160), .C2(net_8059), .C1(net_5683), .B(net_3298) );
NAND2_X2 inst_3569 ( .A2(net_7748), .ZN(net_7676), .A1(net_2481) );
INV_X2 inst_7268 ( .A(net_8923), .ZN(net_8922) );
NAND2_X2 inst_3411 ( .ZN(net_8525), .A1(net_8471), .A2(net_8470) );
AND2_X4 inst_10436 ( .ZN(net_3023), .A2(net_2509), .A1(net_1218) );
DFF_X2 inst_7417 ( .QN(net_9417), .D(net_8347), .CK(net_11702) );
CLKBUF_X2 inst_12576 ( .A(net_11383), .Z(net_12495) );
NOR2_X2 inst_2524 ( .ZN(net_8398), .A1(net_8179), .A2(net_8178) );
AOI22_X2 inst_9486 ( .B1(net_9717), .A1(net_9685), .A2(net_5966), .ZN(net_3837), .B2(net_3039) );
OAI221_X2 inst_1446 ( .ZN(net_8440), .C1(net_8439), .B1(net_8439), .C2(net_8399), .A(net_8370), .B2(net_8132) );
XNOR2_X2 inst_390 ( .ZN(net_2190), .B(net_1595), .A(net_687) );
NOR3_X2 inst_2421 ( .ZN(net_4897), .A1(net_4483), .A3(net_4298), .A2(net_1569) );
INV_X4 inst_4842 ( .ZN(net_3556), .A(net_3316) );
CLKBUF_X2 inst_14455 ( .A(net_14373), .Z(net_14374) );
DFF_X2 inst_8181 ( .QN(net_9731), .D(net_5023), .CK(net_12256) );
OAI22_X2 inst_1062 ( .A2(net_7036), .B2(net_7035), .ZN(net_6982), .B1(net_5719), .A1(net_3974) );
CLKBUF_X2 inst_13757 ( .A(net_13675), .Z(net_13676) );
DFF_X2 inst_7996 ( .QN(net_10335), .D(net_5519), .CK(net_14357) );
NOR2_X2 inst_2663 ( .ZN(net_7597), .A2(net_5973), .A1(net_4997) );
NAND3_X2 inst_3289 ( .A3(net_3261), .ZN(net_3086), .A1(net_3085), .A2(net_2581) );
DFF_X2 inst_7477 ( .D(net_8070), .Q(net_211), .CK(net_12904) );
CLKBUF_X2 inst_12814 ( .A(net_12732), .Z(net_12733) );
CLKBUF_X2 inst_15597 ( .A(net_15515), .Z(net_15516) );
DFF_X2 inst_7930 ( .QN(net_10206), .D(net_5626), .CK(net_11601) );
CLKBUF_X2 inst_14361 ( .A(net_10643), .Z(net_14280) );
CLKBUF_X2 inst_12650 ( .A(net_12009), .Z(net_12569) );
CLKBUF_X2 inst_12116 ( .A(net_12034), .Z(net_12035) );
AND2_X2 inst_10508 ( .ZN(net_5315), .A1(net_5314), .A2(net_5313) );
CLKBUF_X2 inst_12087 ( .A(net_12005), .Z(net_12006) );
AOI211_X2 inst_10277 ( .A(net_7704), .ZN(net_7466), .C2(net_7178), .C1(net_3992), .B(x3390) );
XNOR2_X2 inst_401 ( .B(net_9652), .ZN(net_1752), .A(net_1564) );
DFF_X2 inst_8086 ( .Q(net_9952), .D(net_5001), .CK(net_12331) );
NAND3_X2 inst_3210 ( .ZN(net_6780), .A1(net_6445), .A3(net_3845), .A2(net_3783) );
CLKBUF_X2 inst_12440 ( .A(net_12358), .Z(net_12359) );
INV_X2 inst_7063 ( .A(net_1819), .ZN(net_1267) );
CLKBUF_X2 inst_12539 ( .A(net_12457), .Z(net_12458) );
INV_X4 inst_5200 ( .ZN(net_1939), .A(net_1537) );
NOR2_X2 inst_2642 ( .ZN(net_5450), .A2(net_5449), .A1(net_1456) );
INV_X4 inst_6145 ( .A(net_9292), .ZN(net_568) );
INV_X4 inst_4653 ( .A(net_9256), .ZN(net_6230) );
INV_X4 inst_6087 ( .ZN(net_498), .A(net_103) );
CLKBUF_X2 inst_12028 ( .A(net_11946), .Z(net_11947) );
CLKBUF_X2 inst_14823 ( .A(net_14741), .Z(net_14742) );
MUX2_X1 inst_4465 ( .S(net_6041), .A(net_281), .B(x6102), .Z(x297) );
CLKBUF_X2 inst_14394 ( .A(net_10724), .Z(net_14313) );
CLKBUF_X2 inst_13107 ( .A(net_13025), .Z(net_13026) );
CLKBUF_X2 inst_12281 ( .A(net_12199), .Z(net_12200) );
INV_X4 inst_4865 ( .ZN(net_4217), .A(net_2953) );
CLKBUF_X2 inst_13479 ( .A(net_13397), .Z(net_13398) );
DFF_X1 inst_8548 ( .Q(net_9984), .D(net_7356), .CK(net_14782) );
INV_X4 inst_5250 ( .ZN(net_2049), .A(net_806) );
XNOR2_X2 inst_123 ( .ZN(net_7551), .A(net_7322), .B(net_7031) );
OR2_X2 inst_930 ( .A2(net_8860), .ZN(net_4947), .A1(net_2755) );
DFF_X2 inst_7634 ( .D(net_6759), .QN(net_124), .CK(net_15727) );
CLKBUF_X2 inst_11908 ( .A(net_11826), .Z(net_11827) );
INV_X2 inst_6801 ( .ZN(net_5234), .A(net_5233) );
OAI211_X2 inst_2160 ( .C2(net_6774), .ZN(net_6688), .A(net_6306), .B(net_6048), .C1(net_5053) );
CLKBUF_X2 inst_15248 ( .A(net_13118), .Z(net_15167) );
DFF_X1 inst_8494 ( .QN(net_10054), .D(net_7819), .CK(net_13747) );
INV_X4 inst_5181 ( .A(net_2192), .ZN(net_1787) );
CLKBUF_X2 inst_10981 ( .A(net_10685), .Z(net_10900) );
OAI211_X2 inst_2298 ( .ZN(net_3560), .A(net_3559), .B(net_3558), .C2(net_2939), .C1(net_1951) );
AND2_X4 inst_10453 ( .A1(net_10159), .A2(net_9735), .ZN(net_1669) );
CLKBUF_X2 inst_14355 ( .A(net_14273), .Z(net_14274) );
INV_X4 inst_6622 ( .A(net_8955), .ZN(net_8954) );
CLKBUF_X2 inst_14546 ( .A(net_14464), .Z(net_14465) );
CLKBUF_X2 inst_11660 ( .A(net_11578), .Z(net_11579) );
XNOR2_X2 inst_167 ( .ZN(net_5807), .A(net_4977), .B(net_208) );
CLKBUF_X2 inst_13138 ( .A(net_13056), .Z(net_13057) );
CLKBUF_X2 inst_11354 ( .A(net_11272), .Z(net_11273) );
CLKBUF_X2 inst_13650 ( .A(net_10559), .Z(net_13569) );
INV_X4 inst_4913 ( .A(net_7095), .ZN(net_6192) );
NAND2_X2 inst_3874 ( .ZN(net_4363), .A2(net_4226), .A1(net_4083) );
DFF_X1 inst_8524 ( .Q(net_9970), .D(net_7353), .CK(net_14868) );
AOI22_X2 inst_9168 ( .A2(net_6418), .ZN(net_6303), .B2(net_5263), .B1(net_2991), .A1(net_2560) );
OAI22_X2 inst_1251 ( .B1(net_7198), .A2(net_4826), .B2(net_4825), .ZN(net_4823), .A1(net_407) );
CLKBUF_X2 inst_12245 ( .A(net_12163), .Z(net_12164) );
INV_X4 inst_4874 ( .ZN(net_6203), .A(net_6165) );
NOR2_X4 inst_2475 ( .A1(net_8931), .ZN(net_8380), .A2(net_8164) );
HA_X1 inst_7360 ( .B(net_9248), .S(net_1460), .CO(net_1459), .A(net_653) );
INV_X2 inst_6824 ( .ZN(net_4197), .A(net_4196) );
CLKBUF_X2 inst_13033 ( .A(net_12951), .Z(net_12952) );
AOI22_X2 inst_9195 ( .A1(net_9885), .B1(net_9786), .A2(net_6141), .B2(net_6120), .ZN(net_6118) );
CLKBUF_X2 inst_13131 ( .A(net_12694), .Z(net_13050) );
CLKBUF_X2 inst_12488 ( .A(net_12406), .Z(net_12407) );
XNOR2_X2 inst_331 ( .ZN(net_2996), .B(net_2995), .A(net_2155) );
AOI211_X2 inst_10300 ( .ZN(net_3619), .C2(net_3046), .B(net_2796), .A(net_2566), .C1(net_2230) );
AOI211_X2 inst_10270 ( .C2(net_7641), .ZN(net_7609), .B(net_7524), .A(net_6784), .C1(net_6623) );
DFF_X2 inst_7433 ( .QN(net_9062), .D(net_8324), .CK(net_11758) );
CLKBUF_X2 inst_10691 ( .A(net_10609), .Z(net_10610) );
AOI221_X2 inst_9937 ( .B2(net_5867), .A(net_5859), .ZN(net_5830), .C1(net_5829), .C2(net_4725), .B1(x5647) );
CLKBUF_X2 inst_13312 ( .A(net_13230), .Z(net_13231) );
CLKBUF_X2 inst_15411 ( .A(net_15329), .Z(net_15330) );
CLKBUF_X2 inst_14317 ( .A(net_14235), .Z(net_14236) );
DFF_X2 inst_7369 ( .QN(net_9370), .D(net_8725), .CK(net_14196) );
OAI211_X2 inst_2172 ( .C1(net_7219), .C2(net_6548), .ZN(net_6537), .B(net_5665), .A(net_3507) );
CLKBUF_X2 inst_11227 ( .A(net_10924), .Z(net_11146) );
NOR4_X2 inst_2353 ( .ZN(net_3455), .A3(net_1728), .A4(net_1727), .A1(net_667), .A2(x6445) );
CLKBUF_X2 inst_11921 ( .A(net_11839), .Z(net_11840) );
DFF_X2 inst_8005 ( .QN(net_10333), .D(net_5503), .CK(net_14472) );
SDFF_X2 inst_667 ( .SI(net_9496), .Q(net_9496), .SE(net_3073), .CK(net_12397), .D(x1660) );
CLKBUF_X2 inst_13483 ( .A(net_13401), .Z(net_13402) );
NOR2_X2 inst_2762 ( .A2(net_3593), .ZN(net_3544), .A1(net_3172) );
CLKBUF_X2 inst_12646 ( .A(net_12564), .Z(net_12565) );
DFF_X1 inst_8870 ( .D(net_10516), .CK(net_12656), .Q(x465) );
NOR2_X2 inst_2896 ( .ZN(net_2386), .A1(net_1280), .A2(net_685) );
OAI22_X2 inst_997 ( .A1(net_8627), .B2(net_8626), .ZN(net_8625), .A2(net_8620), .B1(net_7856) );
OR2_X2 inst_857 ( .ZN(net_8140), .A1(net_8091), .A2(net_8090) );
DFF_X1 inst_8732 ( .QN(net_10451), .D(net_5882), .CK(net_11081) );
INV_X4 inst_4824 ( .A(net_4371), .ZN(net_3678) );
NOR2_X2 inst_2691 ( .A2(net_10166), .A1(net_10165), .ZN(net_5219) );
CLKBUF_X2 inst_14401 ( .A(net_12837), .Z(net_14320) );
INV_X4 inst_6311 ( .A(net_9995), .ZN(net_423) );
OAI221_X2 inst_1511 ( .C1(net_10427), .B2(net_9063), .C2(net_9056), .ZN(net_7349), .B1(net_7184), .A(net_7008) );
INV_X4 inst_6403 ( .A(net_10471), .ZN(net_739) );
DFF_X2 inst_7543 ( .QN(net_9314), .D(net_7740), .CK(net_13042) );
CLKBUF_X2 inst_10777 ( .A(net_10582), .Z(net_10696) );
NAND2_X2 inst_4179 ( .ZN(net_2654), .A2(net_1526), .A1(net_1322) );
CLKBUF_X2 inst_12721 ( .A(net_12639), .Z(net_12640) );
INV_X4 inst_5951 ( .ZN(net_797), .A(net_558) );
DFF_X2 inst_7988 ( .QN(net_10414), .D(net_5541), .CK(net_14752) );
INV_X4 inst_6645 ( .A(net_9107), .ZN(net_9106) );
NAND2_X2 inst_4006 ( .ZN(net_3919), .A2(net_3390), .A1(net_937) );
NAND2_X2 inst_4243 ( .A2(net_10157), .ZN(net_2681), .A1(net_1126) );
NAND3_X2 inst_3203 ( .ZN(net_7406), .A3(net_7405), .A2(net_6632), .A1(net_5985) );
CLKBUF_X2 inst_15368 ( .A(net_15286), .Z(net_15287) );
CLKBUF_X2 inst_14344 ( .A(net_12637), .Z(net_14263) );
CLKBUF_X2 inst_13659 ( .A(net_13577), .Z(net_13578) );
INV_X4 inst_5073 ( .ZN(net_8200), .A(net_1834) );
OAI221_X2 inst_1504 ( .B2(net_9063), .C2(net_9056), .ZN(net_7357), .B1(net_7203), .A(net_7004), .C1(net_978) );
NAND2_X2 inst_3403 ( .ZN(net_8588), .A2(net_8587), .A1(net_8446) );
CLKBUF_X2 inst_13951 ( .A(net_13869), .Z(net_13870) );
INV_X4 inst_5830 ( .ZN(net_1244), .A(net_1031) );
OAI22_X2 inst_1310 ( .ZN(net_3200), .A2(net_2305), .B2(net_2304), .A1(net_2304), .B1(net_1357) );
NAND3_X2 inst_3280 ( .ZN(net_5802), .A2(net_5284), .A3(net_3867), .A1(net_2927) );
AOI221_X2 inst_9802 ( .B1(net_9981), .A(net_7090), .B2(net_7089), .C2(net_7088), .ZN(net_7000), .C1(net_253) );
INV_X8 inst_4491 ( .ZN(net_6940), .A(net_5935) );
AOI22_X2 inst_9006 ( .ZN(net_8032), .A2(net_8030), .B2(net_8029), .B1(net_7499), .A1(net_210) );
DFF_X2 inst_7518 ( .Q(net_9533), .D(net_7882), .CK(net_13988) );
DFF_X2 inst_7397 ( .D(net_8548), .Q(net_221), .CK(net_14618) );
CLKBUF_X2 inst_11594 ( .A(net_11512), .Z(net_11513) );
NOR2_X2 inst_2823 ( .A1(net_2964), .ZN(net_2556), .A2(net_2555) );
INV_X2 inst_7242 ( .A(net_9411), .ZN(net_8223) );
CLKBUF_X2 inst_13981 ( .A(net_13899), .Z(net_13900) );
NAND2_X2 inst_3807 ( .A1(net_10076), .A2(net_4534), .ZN(net_4531) );
CLKBUF_X2 inst_13413 ( .A(net_13331), .Z(net_13332) );
CLKBUF_X2 inst_15171 ( .A(net_15089), .Z(net_15090) );
OAI22_X2 inst_1069 ( .B2(net_10273), .ZN(net_6908), .A2(net_6631), .B1(net_5407), .A1(net_997) );
CLKBUF_X2 inst_12719 ( .A(net_12637), .Z(net_12638) );
CLKBUF_X2 inst_11327 ( .A(net_11245), .Z(net_11246) );
CLKBUF_X2 inst_14464 ( .A(net_14382), .Z(net_14383) );
CLKBUF_X2 inst_14153 ( .A(net_12904), .Z(net_14072) );
XNOR2_X2 inst_136 ( .B(net_9422), .ZN(net_7400), .A(net_6655) );
CLKBUF_X2 inst_13083 ( .A(net_10946), .Z(net_13002) );
CLKBUF_X2 inst_11733 ( .A(net_11651), .Z(net_11652) );
AND4_X4 inst_10326 ( .A4(net_5041), .A3(net_5032), .ZN(net_3351), .A2(net_3350), .A1(net_2748) );
INV_X4 inst_5839 ( .A(net_753), .ZN(net_655) );
NAND2_X2 inst_3541 ( .A2(net_9634), .A1(net_8979), .ZN(net_8095) );
CLKBUF_X2 inst_13837 ( .A(net_13755), .Z(net_13756) );
OAI221_X2 inst_1526 ( .B1(net_10313), .B2(net_9047), .C2(net_7287), .ZN(net_7250), .C1(net_7249), .A(net_6867) );
CLKBUF_X2 inst_11503 ( .A(net_11421), .Z(net_11422) );
CLKBUF_X2 inst_13825 ( .A(net_13743), .Z(net_13744) );
NOR2_X2 inst_2547 ( .A2(net_9635), .A1(net_8978), .ZN(net_8092) );
INV_X4 inst_4637 ( .A(net_7505), .ZN(net_6948) );
CLKBUF_X2 inst_15790 ( .A(net_15708), .Z(net_15709) );
OAI22_X2 inst_1047 ( .ZN(net_7538), .A2(net_7395), .B2(net_7394), .A1(net_7157), .B1(net_465) );
INV_X2 inst_6860 ( .ZN(net_3324), .A(net_3113) );
INV_X4 inst_5167 ( .ZN(net_2739), .A(net_2099) );
NAND2_X2 inst_3850 ( .A2(net_4631), .ZN(net_4223), .A1(net_3553) );
CLKBUF_X2 inst_12582 ( .A(net_10775), .Z(net_12501) );
DFF_X1 inst_8507 ( .QN(net_10163), .D(net_7661), .CK(net_13528) );
CLKBUF_X2 inst_11768 ( .A(net_11686), .Z(net_11687) );
CLKBUF_X2 inst_15519 ( .A(net_10755), .Z(net_15438) );
CLKBUF_X2 inst_14368 ( .A(net_14286), .Z(net_14287) );
CLKBUF_X2 inst_12432 ( .A(net_12350), .Z(net_12351) );
CLKBUF_X2 inst_10972 ( .A(net_10824), .Z(net_10891) );
INV_X2 inst_6744 ( .A(net_7094), .ZN(net_6916) );
NAND2_X2 inst_3700 ( .A1(net_6165), .A2(net_5937), .ZN(net_5936) );
OAI21_X2 inst_1858 ( .ZN(net_5791), .B1(net_5790), .A(net_5380), .B2(net_1069) );
OAI21_X2 inst_1786 ( .B2(net_7659), .ZN(net_7541), .A(net_7429), .B1(net_5241) );
CLKBUF_X2 inst_13668 ( .A(net_13586), .Z(net_13587) );
NAND2_X2 inst_3846 ( .ZN(net_4369), .A1(net_4237), .A2(net_4078) );
CLKBUF_X2 inst_15271 ( .A(net_11403), .Z(net_15190) );
OAI222_X2 inst_1334 ( .ZN(net_7729), .A1(net_7728), .B2(net_7727), .C2(net_7726), .A2(net_7567), .B1(net_5668), .C1(net_1084) );
CLKBUF_X2 inst_15688 ( .A(net_15606), .Z(net_15607) );
SDFF_X2 inst_496 ( .SE(net_9540), .SI(net_8213), .Q(net_285), .D(net_285), .CK(net_12703) );
CLKBUF_X2 inst_10639 ( .A(net_10557), .Z(net_10558) );
INV_X2 inst_7174 ( .A(net_9209), .ZN(net_543) );
CLKBUF_X2 inst_12356 ( .A(net_12274), .Z(net_12275) );
AOI211_X2 inst_10304 ( .C2(net_10082), .C1(net_10064), .B(net_9859), .A(net_9760), .ZN(net_3476) );
INV_X4 inst_5369 ( .A(net_1265), .ZN(net_1207) );
INV_X4 inst_5944 ( .A(net_6960), .ZN(net_565) );
AOI22_X2 inst_9011 ( .B1(net_9306), .A2(net_8030), .B2(net_8029), .ZN(net_8025), .A1(net_214) );
INV_X4 inst_5733 ( .ZN(net_980), .A(net_751) );
INV_X2 inst_6867 ( .ZN(net_3148), .A(net_3147) );
INV_X4 inst_6129 ( .A(net_9737), .ZN(net_485) );
INV_X4 inst_5383 ( .A(net_2132), .ZN(net_1576) );
NAND2_X2 inst_3749 ( .ZN(net_5301), .A2(net_5290), .A1(net_4474) );
CLKBUF_X2 inst_14735 ( .A(net_11489), .Z(net_14654) );
CLKBUF_X2 inst_12130 ( .A(net_11583), .Z(net_12049) );
INV_X2 inst_7273 ( .A(net_8945), .ZN(net_8944) );
NOR2_X2 inst_2620 ( .ZN(net_7642), .A2(net_6205), .A1(net_6188) );
OAI221_X2 inst_1633 ( .C1(net_10310), .B1(net_7108), .C2(net_5591), .A(net_5575), .ZN(net_5573), .B2(net_4902) );
CLKBUF_X2 inst_15567 ( .A(net_13294), .Z(net_15486) );
CLKBUF_X2 inst_12425 ( .A(net_12317), .Z(net_12344) );
CLKBUF_X2 inst_11453 ( .A(net_11371), .Z(net_11372) );
OAI22_X2 inst_1262 ( .B1(net_7184), .A2(net_4842), .B2(net_4841), .ZN(net_4811), .A1(net_388) );
INV_X4 inst_5303 ( .ZN(net_5881), .A(net_1298) );
AOI22_X2 inst_9364 ( .B1(net_9896), .A2(net_5759), .B2(net_5758), .ZN(net_5558), .A1(net_235) );
XNOR2_X2 inst_265 ( .B(net_9620), .ZN(net_3973), .A(net_3653) );
DFF_X2 inst_8048 ( .QN(net_10362), .D(net_5703), .CK(net_13633) );
OAI211_X2 inst_2055 ( .ZN(net_7791), .A(net_7783), .C1(net_7782), .B(net_7687), .C2(net_4956) );
CLKBUF_X2 inst_11702 ( .A(net_11490), .Z(net_11621) );
INV_X2 inst_6799 ( .ZN(net_5373), .A(net_5372) );
NAND2_X2 inst_3856 ( .A2(net_4187), .ZN(net_4179), .A1(net_1847) );
CLKBUF_X2 inst_12453 ( .A(net_11794), .Z(net_12372) );
DFF_X2 inst_7783 ( .Q(net_9816), .D(net_6516), .CK(net_15710) );
INV_X4 inst_5091 ( .ZN(net_2227), .A(net_1747) );
INV_X4 inst_5554 ( .A(net_1708), .ZN(net_1299) );
CLKBUF_X2 inst_14169 ( .A(net_14087), .Z(net_14088) );
CLKBUF_X2 inst_11650 ( .A(net_11568), .Z(net_11569) );
NAND3_X2 inst_3262 ( .A2(net_5335), .ZN(net_4359), .A3(net_3869), .A1(net_2922) );
CLKBUF_X2 inst_12577 ( .A(net_12495), .Z(net_12496) );
CLKBUF_X2 inst_11482 ( .A(net_11400), .Z(net_11401) );
INV_X4 inst_6432 ( .A(net_9290), .ZN(net_663) );
INV_X4 inst_4566 ( .ZN(net_8430), .A(net_8173) );
CLKBUF_X2 inst_10716 ( .A(net_10634), .Z(net_10635) );
CLKBUF_X2 inst_12993 ( .A(net_11504), .Z(net_12912) );
CLKBUF_X2 inst_10653 ( .A(net_10570), .Z(net_10572) );
INV_X4 inst_6301 ( .ZN(net_7224), .A(x4285) );
OAI22_X2 inst_1077 ( .A2(net_9064), .ZN(net_6653), .B2(net_6639), .B1(net_3524), .A1(net_487) );
CLKBUF_X2 inst_15495 ( .A(net_15413), .Z(net_15414) );
DFF_X2 inst_7975 ( .QN(net_10309), .D(net_5576), .CK(net_12138) );
INV_X2 inst_7249 ( .A(net_9232), .ZN(net_361) );
CLKBUF_X2 inst_12956 ( .A(net_11170), .Z(net_12875) );
NAND2_X2 inst_3954 ( .A1(net_10158), .ZN(net_3707), .A2(net_3423) );
AOI22_X2 inst_9367 ( .B1(net_9918), .A2(net_5759), .B2(net_5758), .ZN(net_5555), .A1(net_257) );
INV_X4 inst_6461 ( .A(net_10022), .ZN(net_373) );
NOR2_X2 inst_2757 ( .ZN(net_3873), .A1(net_3604), .A2(net_3386) );
XNOR2_X2 inst_222 ( .ZN(net_4572), .A(net_4414), .B(net_1982) );
OAI21_X2 inst_1932 ( .A(net_4415), .ZN(net_4374), .B1(net_4373), .B2(net_4005) );
CLKBUF_X2 inst_10822 ( .A(net_10740), .Z(net_10741) );
AOI222_X1 inst_9733 ( .B2(net_10297), .C2(net_10295), .A2(net_10294), .B1(net_10290), .C1(net_10288), .A1(net_10287), .ZN(net_1447) );
INV_X4 inst_6372 ( .A(net_9746), .ZN(net_1816) );
DFF_X2 inst_7884 ( .QN(net_10107), .D(net_6033), .CK(net_14910) );
INV_X4 inst_6073 ( .ZN(net_503), .A(net_227) );
NAND2_X2 inst_3704 ( .A1(net_10067), .ZN(net_5925), .A2(net_5896) );
CLKBUF_X2 inst_13903 ( .A(net_11008), .Z(net_13822) );
CLKBUF_X2 inst_13166 ( .A(net_13084), .Z(net_13085) );
CLKBUF_X2 inst_12218 ( .A(net_12136), .Z(net_12137) );
CLKBUF_X2 inst_11828 ( .A(net_11746), .Z(net_11747) );
INV_X2 inst_6728 ( .ZN(net_7738), .A(net_7696) );
OAI22_X2 inst_1052 ( .ZN(net_7532), .A1(net_7531), .B2(net_7530), .A2(net_7389), .B1(net_2998) );
OAI22_X2 inst_1280 ( .A2(net_10061), .ZN(net_4277), .A1(net_4275), .B2(net_4274), .B1(net_1517) );
OAI22_X2 inst_1302 ( .ZN(net_3096), .A1(net_3095), .B2(net_2909), .A2(net_2908), .B1(net_1007) );
CLKBUF_X2 inst_12740 ( .A(net_11553), .Z(net_12659) );
INV_X4 inst_6435 ( .A(net_10114), .ZN(net_749) );
INV_X4 inst_5362 ( .ZN(net_1555), .A(net_1220) );
CLKBUF_X2 inst_13904 ( .A(net_13822), .Z(net_13823) );
AOI22_X2 inst_9578 ( .B1(net_9977), .A2(net_5173), .ZN(net_3586), .B2(net_2541), .A1(net_211) );
INV_X4 inst_6112 ( .ZN(net_1415), .A(net_225) );
AND2_X2 inst_10609 ( .A1(net_4188), .A2(net_3121), .ZN(net_2670) );
OAI221_X2 inst_1648 ( .C1(net_10415), .B1(net_7108), .ZN(net_5540), .C2(net_4477), .B2(net_4455), .A(net_3507) );
CLKBUF_X2 inst_13958 ( .A(net_10682), .Z(net_13877) );
INV_X4 inst_5847 ( .A(net_1755), .ZN(net_812) );
OAI22_X2 inst_1079 ( .A2(net_9064), .B2(net_6639), .ZN(net_6580), .B1(net_4121), .A1(net_1099) );
CLKBUF_X2 inst_13833 ( .A(net_13751), .Z(net_13752) );
INV_X4 inst_6200 ( .A(net_10257), .ZN(net_743) );
NAND2_X2 inst_3925 ( .A2(net_4319), .ZN(net_3882), .A1(net_2111) );
NOR2_X2 inst_2606 ( .ZN(net_6262), .A1(net_5764), .A2(net_3329) );
AOI221_X2 inst_9837 ( .A(net_6889), .B2(net_6888), .C2(net_6887), .ZN(net_6881), .B1(net_5849), .C1(x5077) );
NAND2_X2 inst_4314 ( .ZN(net_2685), .A2(net_919), .A1(net_581) );
NOR2_X2 inst_2523 ( .ZN(net_8252), .A1(net_8182), .A2(net_8181) );
SDFF_X2 inst_506 ( .SE(net_9540), .SI(net_8194), .Q(net_296), .D(net_296), .CK(net_13963) );
CLKBUF_X2 inst_13569 ( .A(net_13487), .Z(net_13488) );
CLKBUF_X2 inst_10662 ( .A(net_10565), .Z(net_10581) );
CLKBUF_X2 inst_14975 ( .A(net_14893), .Z(net_14894) );
CLKBUF_X2 inst_11782 ( .A(net_11700), .Z(net_11701) );
DFF_X1 inst_8572 ( .Q(net_9673), .D(net_7102), .CK(net_14844) );
XNOR2_X2 inst_134 ( .ZN(net_7411), .B(net_7086), .A(net_6895) );
NOR3_X2 inst_2409 ( .A1(net_9087), .ZN(net_6674), .A2(net_6673), .A3(net_6253) );
NAND2_X4 inst_3322 ( .ZN(net_8700), .A1(net_8670), .A2(net_8669) );
CLKBUF_X2 inst_10835 ( .A(net_10753), .Z(net_10754) );
OAI22_X2 inst_1085 ( .A1(net_7157), .ZN(net_6573), .A2(net_5906), .B2(net_5905), .B1(net_489) );
OAI22_X2 inst_1323 ( .B1(net_2780), .B2(net_2643), .A1(net_2302), .ZN(net_1760), .A2(net_1759) );
NAND2_X2 inst_3425 ( .ZN(net_8591), .A1(net_8497), .A2(net_8496) );
CLKBUF_X2 inst_14048 ( .A(net_13966), .Z(net_13967) );
NOR4_X2 inst_2328 ( .ZN(net_5277), .A4(net_5101), .A1(net_5017), .A3(net_2151), .A2(net_894) );
AND2_X4 inst_10464 ( .A2(net_10258), .ZN(net_1682), .A1(net_1342) );
DFF_X1 inst_8791 ( .Q(net_9162), .D(net_4386), .CK(net_10899) );
DFF_X2 inst_8060 ( .QN(net_9167), .D(net_5277), .CK(net_13564) );
NOR2_X2 inst_2655 ( .A1(net_8565), .ZN(net_5257), .A2(net_5256) );
XNOR2_X2 inst_160 ( .ZN(net_5979), .A(net_5978), .B(net_2073) );
OAI221_X2 inst_1720 ( .C1(net_10354), .ZN(net_2915), .A(net_2379), .B1(net_1555), .B2(net_1354), .C2(net_737) );
INV_X4 inst_5779 ( .ZN(net_1381), .A(net_707) );
CLKBUF_X2 inst_14420 ( .A(net_14338), .Z(net_14339) );
CLKBUF_X2 inst_14890 ( .A(net_14808), .Z(net_14809) );
CLKBUF_X2 inst_13541 ( .A(net_13459), .Z(net_13460) );
NOR2_X2 inst_2912 ( .A1(net_4221), .A2(net_2824), .ZN(net_1497) );
AOI22_X2 inst_9243 ( .A1(net_9947), .B1(net_9848), .A2(net_8042), .B2(net_6120), .ZN(net_6068) );
DFF_X2 inst_7450 ( .QN(net_9294), .D(net_8244), .CK(net_14989) );
OR2_X4 inst_762 ( .ZN(net_5151), .A1(net_4475), .A2(net_4363) );
XNOR2_X2 inst_370 ( .ZN(net_2482), .B(net_2481), .A(net_2479) );
AND2_X4 inst_10414 ( .ZN(net_4289), .A2(x3632), .A1(x813) );
DFF_X2 inst_7825 ( .Q(net_9650), .D(net_6551), .CK(net_11817) );
NOR2_X2 inst_3025 ( .A2(net_9275), .A1(net_9274), .ZN(net_592) );
CLKBUF_X2 inst_15472 ( .A(net_13118), .Z(net_15391) );
OAI22_X2 inst_1265 ( .B1(net_7213), .A2(net_4842), .B2(net_4841), .ZN(net_4808), .A1(net_496) );
CLKBUF_X2 inst_14480 ( .A(net_14398), .Z(net_14399) );
CLKBUF_X2 inst_15600 ( .A(net_15518), .Z(net_15519) );
CLKBUF_X2 inst_10669 ( .A(net_10587), .Z(net_10588) );
DFF_X2 inst_7530 ( .QN(net_9323), .D(net_7779), .CK(net_13058) );
AND2_X4 inst_10434 ( .ZN(net_5319), .A1(net_4230), .A2(net_3630) );
DFF_X2 inst_8371 ( .Q(net_9273), .D(net_1469), .CK(net_11425) );
INV_X8 inst_4530 ( .A(net_9100), .ZN(net_9097) );
CLKBUF_X2 inst_11882 ( .A(net_11800), .Z(net_11801) );
DFF_X2 inst_8176 ( .QN(net_10025), .D(net_5034), .CK(net_11441) );
CLKBUF_X2 inst_11288 ( .A(net_11206), .Z(net_11207) );
OAI22_X2 inst_1321 ( .B2(net_9746), .ZN(net_1818), .A1(net_1817), .A2(net_1816), .B1(net_1022) );
CLKBUF_X2 inst_14607 ( .A(net_14525), .Z(net_14526) );
OAI22_X2 inst_1012 ( .A2(net_8247), .B2(net_8246), .ZN(net_8243), .A1(net_2822), .B1(net_1870) );
CLKBUF_X2 inst_12768 ( .A(net_12638), .Z(net_12687) );
INV_X4 inst_5255 ( .ZN(net_1467), .A(net_1431) );
CLKBUF_X2 inst_13843 ( .A(net_13761), .Z(net_13762) );
DFF_X2 inst_8341 ( .Q(net_10175), .D(net_3363), .CK(net_12844) );
OAI21_X2 inst_1956 ( .ZN(net_4253), .A(net_3325), .B2(net_3236), .B1(net_3114) );
DFF_X2 inst_8378 ( .QN(net_8845), .D(net_2295), .CK(net_10789) );
NAND2_X2 inst_3492 ( .A2(net_8385), .ZN(net_8378), .A1(net_8330) );
CLKBUF_X2 inst_10687 ( .A(net_10600), .Z(net_10606) );
CLKBUF_X2 inst_10935 ( .A(net_10853), .Z(net_10854) );
OR2_X4 inst_751 ( .ZN(net_5133), .A2(net_4476), .A1(net_4475) );
CLKBUF_X2 inst_14032 ( .A(net_13950), .Z(net_13951) );
CLKBUF_X2 inst_14724 ( .A(net_14642), .Z(net_14643) );
AOI22_X2 inst_9015 ( .A2(net_8030), .B2(net_8029), .ZN(net_8021), .A1(net_218), .B1(net_195) );
NAND4_X2 inst_3149 ( .ZN(net_2158), .A4(net_1447), .A2(net_953), .A3(net_765), .A1(net_579) );
NAND2_X2 inst_4283 ( .A2(net_10250), .ZN(net_4558), .A1(net_1214) );
NOR2_X4 inst_2471 ( .A2(net_9025), .A1(net_9024), .ZN(net_8881) );
NAND2_X2 inst_4034 ( .ZN(net_4942), .A1(net_2952), .A2(net_2951) );
CLKBUF_X2 inst_13570 ( .A(net_13488), .Z(net_13489) );
XNOR2_X2 inst_377 ( .ZN(net_2453), .A(net_1408), .B(net_1331) );
INV_X2 inst_6993 ( .A(net_3136), .ZN(net_1640) );
AOI21_X2 inst_10157 ( .ZN(net_4089), .B1(net_4088), .B2(net_4087), .A(net_3692) );
INV_X4 inst_4760 ( .ZN(net_4543), .A(net_4112) );
NAND2_X2 inst_3946 ( .A2(net_10539), .ZN(net_4170), .A1(net_2975) );
CLKBUF_X2 inst_15703 ( .A(net_15621), .Z(net_15622) );
NAND3_X2 inst_3244 ( .ZN(net_4701), .A3(net_4581), .A1(net_4580), .A2(net_2699) );
INV_X2 inst_6953 ( .A(net_5161), .ZN(net_1883) );
NAND2_X2 inst_3920 ( .A2(net_9053), .ZN(net_7959), .A1(net_3311) );
INV_X2 inst_6920 ( .A(net_2629), .ZN(net_2097) );
NAND2_X2 inst_3821 ( .ZN(net_4904), .A1(net_4517), .A2(net_3893) );
DFF_X2 inst_7443 ( .QN(net_9298), .D(net_8257), .CK(net_11499) );
INV_X4 inst_5981 ( .A(net_10151), .ZN(net_7331) );
NOR2_X2 inst_3018 ( .A1(net_9639), .A2(net_9279), .ZN(net_7932) );
CLKBUF_X2 inst_13750 ( .A(net_13668), .Z(net_13669) );
NAND4_X2 inst_3078 ( .A3(net_9235), .ZN(net_5361), .A2(net_4349), .A4(net_2740), .A1(net_1673) );
CLKBUF_X2 inst_12779 ( .A(net_11022), .Z(net_12698) );
INV_X4 inst_5792 ( .ZN(net_871), .A(net_691) );
CLKBUF_X2 inst_14554 ( .A(net_12311), .Z(net_14473) );
CLKBUF_X2 inst_12675 ( .A(net_12593), .Z(net_12594) );
CLKBUF_X2 inst_13579 ( .A(net_13497), .Z(net_13498) );
CLKBUF_X2 inst_13330 ( .A(net_12704), .Z(net_13249) );
AOI222_X1 inst_9731 ( .B1(net_4029), .C1(net_4024), .ZN(net_3122), .C2(net_3121), .B2(net_2664), .A2(net_2663), .A1(net_1977) );
INV_X4 inst_4623 ( .ZN(net_7916), .A(net_7700) );
INV_X4 inst_5926 ( .A(net_1950), .ZN(net_974) );
INV_X4 inst_5054 ( .ZN(net_1881), .A(net_1880) );
NAND2_X2 inst_3835 ( .A2(net_4470), .ZN(net_4327), .A1(net_4326) );
INV_X4 inst_4627 ( .ZN(net_7363), .A(net_7040) );
CLKBUF_X2 inst_14429 ( .A(net_14347), .Z(net_14348) );
CLKBUF_X2 inst_13559 ( .A(net_12828), .Z(net_13478) );
CLKBUF_X2 inst_12414 ( .A(net_11999), .Z(net_12333) );
CLKBUF_X2 inst_14191 ( .A(net_14109), .Z(net_14110) );
XNOR2_X2 inst_107 ( .ZN(net_8143), .A(net_8049), .B(net_7049) );
OAI211_X2 inst_2117 ( .C2(net_6778), .ZN(net_6731), .A(net_6358), .B(net_6092), .C1(net_316) );
OAI22_X2 inst_990 ( .A2(net_8962), .B2(net_8659), .ZN(net_8642), .B1(net_7378), .A1(net_7364) );
CLKBUF_X2 inst_12381 ( .A(net_12299), .Z(net_12300) );
AND2_X4 inst_10412 ( .ZN(net_5754), .A1(net_4788), .A2(net_4779) );
INV_X2 inst_7225 ( .A(net_9396), .ZN(net_8210) );
NAND4_X2 inst_3140 ( .ZN(net_2694), .A1(net_2693), .A4(net_2692), .A3(net_1537), .A2(net_1487) );
INV_X4 inst_4710 ( .ZN(net_4737), .A(net_4619) );
CLKBUF_X2 inst_13812 ( .A(net_13730), .Z(net_13731) );
CLKBUF_X2 inst_12035 ( .A(net_11953), .Z(net_11954) );
CLKBUF_X2 inst_14600 ( .A(net_14518), .Z(net_14519) );
NAND2_X2 inst_3628 ( .ZN(net_7093), .A2(net_6670), .A1(net_5413) );
CLKBUF_X2 inst_11941 ( .A(net_10836), .Z(net_11860) );
CLKBUF_X2 inst_15632 ( .A(net_15550), .Z(net_15551) );
CLKBUF_X2 inst_14886 ( .A(net_12879), .Z(net_14805) );
CLKBUF_X2 inst_12308 ( .A(net_12226), .Z(net_12227) );
AOI21_X2 inst_10093 ( .B1(net_9526), .ZN(net_5189), .A(net_4673), .B2(net_4550) );
NOR3_X2 inst_2366 ( .A3(net_9587), .A2(net_9575), .ZN(net_8780), .A1(net_8777) );
CLKBUF_X2 inst_11200 ( .A(net_11118), .Z(net_11119) );
INV_X4 inst_4642 ( .ZN(net_6026), .A(net_5846) );
HA_X1 inst_7340 ( .S(net_6173), .CO(net_6172), .B(net_5240), .A(net_1601) );
INV_X4 inst_5049 ( .ZN(net_2226), .A(net_1894) );
NAND2_X4 inst_3316 ( .A2(net_8896), .A1(net_8895), .ZN(net_8759) );
AOI22_X2 inst_9385 ( .B1(net_9707), .A1(net_5755), .B2(net_5754), .ZN(net_5438), .A2(net_244) );
CLKBUF_X2 inst_11343 ( .A(net_11261), .Z(net_11262) );
CLKBUF_X2 inst_14155 ( .A(net_14073), .Z(net_14074) );
NAND2_X2 inst_4411 ( .ZN(net_1090), .A1(x6496), .A2(x6401) );
CLKBUF_X2 inst_11471 ( .A(net_10778), .Z(net_11390) );
CLKBUF_X2 inst_13998 ( .A(net_13916), .Z(net_13917) );
DFF_X2 inst_7772 ( .Q(net_9723), .D(net_6531), .CK(net_11972) );
NAND2_X2 inst_4014 ( .A1(net_4190), .A2(net_3080), .ZN(net_3079) );
INV_X4 inst_4605 ( .ZN(net_8614), .A(net_7753) );
NAND2_X2 inst_3694 ( .A2(net_9258), .A1(net_8116), .ZN(net_7278) );
CLKBUF_X2 inst_15204 ( .A(net_15122), .Z(net_15123) );
INV_X4 inst_4882 ( .ZN(net_3508), .A(net_3088) );
CLKBUF_X2 inst_11207 ( .A(net_11125), .Z(net_11126) );
AND3_X4 inst_10351 ( .ZN(net_8076), .A3(net_8074), .A1(net_5575), .A2(net_1067) );
NOR2_X2 inst_2698 ( .A2(net_4557), .ZN(net_4393), .A1(net_2344) );
OAI22_X2 inst_1237 ( .B1(net_7203), .A2(net_4890), .B2(net_4889), .ZN(net_4880), .A1(net_332) );
CLKBUF_X2 inst_12873 ( .A(net_12319), .Z(net_12792) );
AOI221_X2 inst_9908 ( .B1(net_9863), .B2(net_9101), .A(net_6945), .C2(net_6944), .C1(net_6808), .ZN(net_6786) );
NOR2_X2 inst_2518 ( .A2(net_8316), .ZN(net_8262), .A1(net_8148) );
NAND2_X2 inst_3460 ( .A1(net_9490), .A2(net_8476), .ZN(net_8464) );
CLKBUF_X2 inst_15196 ( .A(net_15114), .Z(net_15115) );
INV_X4 inst_5152 ( .ZN(net_2629), .A(net_1583) );
INV_X4 inst_5544 ( .ZN(net_1219), .A(net_969) );
INV_X2 inst_7175 ( .A(net_10162), .ZN(net_656) );
OAI211_X2 inst_2075 ( .C2(net_6774), .ZN(net_6773), .A(net_6400), .B(net_6081), .C1(net_538) );
NAND4_X2 inst_3062 ( .ZN(net_5723), .A4(net_4875), .A2(net_3844), .A1(net_3583), .A3(net_3441) );
NAND3_X2 inst_3310 ( .ZN(net_7437), .A3(net_2101), .A1(net_2099), .A2(net_2098) );
OAI21_X2 inst_1911 ( .ZN(net_4663), .B1(net_4662), .B2(net_4661), .A(net_4384) );
INV_X4 inst_6267 ( .A(net_9353), .ZN(net_606) );
INV_X4 inst_5689 ( .A(net_796), .ZN(net_795) );
CLKBUF_X2 inst_14249 ( .A(net_14167), .Z(net_14168) );
CLKBUF_X2 inst_10841 ( .A(net_10592), .Z(net_10760) );
CLKBUF_X2 inst_15528 ( .A(net_15446), .Z(net_15447) );
CLKBUF_X2 inst_13459 ( .A(net_13377), .Z(net_13378) );
SDFF_X2 inst_585 ( .Q(net_9255), .SE(net_4589), .D(net_138), .SI(net_104), .CK(net_13839) );
INV_X4 inst_5100 ( .A(net_4247), .ZN(net_1983) );
DFF_X1 inst_8536 ( .Q(net_9963), .D(net_7351), .CK(net_14788) );
CLKBUF_X2 inst_15239 ( .A(net_15157), .Z(net_15158) );
DFF_X1 inst_8816 ( .QN(net_10129), .D(net_3256), .CK(net_10813) );
CLKBUF_X2 inst_13967 ( .A(net_12690), .Z(net_13886) );
CLKBUF_X2 inst_14745 ( .A(net_13216), .Z(net_14664) );
INV_X4 inst_5435 ( .ZN(net_1491), .A(net_1117) );
INV_X4 inst_5107 ( .ZN(net_4264), .A(net_1674) );
INV_X4 inst_6013 ( .ZN(net_667), .A(x6496) );
INV_X4 inst_5763 ( .ZN(net_933), .A(net_725) );
CLKBUF_X2 inst_11171 ( .A(net_11089), .Z(net_11090) );
XNOR2_X2 inst_383 ( .ZN(net_2280), .B(net_2279), .A(net_1095) );
CLKBUF_X2 inst_15017 ( .A(net_14935), .Z(net_14936) );
CLKBUF_X2 inst_12137 ( .A(net_12055), .Z(net_12056) );
INV_X4 inst_6453 ( .A(net_10025), .ZN(net_584) );
NOR3_X2 inst_2428 ( .ZN(net_4066), .A1(net_3600), .A2(net_2934), .A3(net_1460) );
CLKBUF_X2 inst_11793 ( .A(net_11711), .Z(net_11712) );
CLKBUF_X2 inst_13561 ( .A(net_12145), .Z(net_13480) );
INV_X4 inst_5115 ( .ZN(net_2675), .A(net_1631) );
CLKBUF_X2 inst_14382 ( .A(net_10664), .Z(net_14301) );
DFF_X2 inst_7670 ( .D(net_6734), .QN(net_152), .CK(net_12066) );
INV_X2 inst_7031 ( .A(net_1842), .ZN(net_1465) );
NAND2_X2 inst_4132 ( .ZN(net_2688), .A2(net_2246), .A1(net_1556) );
DFF_X2 inst_7679 ( .Q(net_10068), .D(net_6568), .CK(net_10842) );
AOI221_X2 inst_9765 ( .C1(net_7697), .ZN(net_7599), .A(net_7456), .B2(net_3922), .C2(net_3064), .B1(net_2974) );
DFF_X2 inst_7553 ( .QN(net_9319), .D(net_7692), .CK(net_13038) );
OAI22_X2 inst_1124 ( .A1(net_7211), .ZN(net_5157), .A2(net_5107), .B2(net_5105), .B1(net_328) );
NAND2_X2 inst_4086 ( .ZN(net_2958), .A1(net_2600), .A2(net_1975) );
CLKBUF_X2 inst_11091 ( .A(net_10776), .Z(net_11010) );
CLKBUF_X2 inst_11801 ( .A(net_10806), .Z(net_11720) );
INV_X4 inst_5372 ( .A(net_3855), .ZN(net_1579) );
NOR2_X2 inst_2555 ( .A1(net_7859), .ZN(net_7858), .A2(net_7825) );
NAND2_X4 inst_3375 ( .A2(net_9200), .ZN(net_3390), .A1(net_2751) );
XNOR2_X2 inst_234 ( .B(net_9208), .ZN(net_4303), .A(net_3968) );
CLKBUF_X2 inst_13922 ( .A(net_13840), .Z(net_13841) );
INV_X2 inst_6966 ( .ZN(net_1825), .A(net_1824) );
INV_X4 inst_5293 ( .A(net_5164), .ZN(net_1310) );
CLKBUF_X2 inst_13447 ( .A(net_10922), .Z(net_13366) );
INV_X4 inst_5240 ( .ZN(net_1900), .A(net_1468) );
CLKBUF_X2 inst_12450 ( .A(net_11796), .Z(net_12369) );
INV_X4 inst_5343 ( .ZN(net_1580), .A(net_1245) );
CLKBUF_X2 inst_12398 ( .A(net_12316), .Z(net_12317) );
NAND2_X2 inst_3714 ( .ZN(net_5904), .A1(net_5903), .A2(net_5902) );
CLKBUF_X2 inst_12317 ( .A(net_10760), .Z(net_12236) );
CLKBUF_X2 inst_12269 ( .A(net_12187), .Z(net_12188) );
INV_X4 inst_5285 ( .ZN(net_1323), .A(net_1322) );
CLKBUF_X2 inst_13975 ( .A(net_13893), .Z(net_13894) );
INV_X2 inst_6658 ( .ZN(net_8421), .A(net_8420) );
INV_X4 inst_5611 ( .ZN(net_7928), .A(net_5684) );
OAI22_X2 inst_1304 ( .A1(net_2906), .ZN(net_2903), .A2(net_2902), .B2(net_2901), .B1(net_1059) );
NAND2_X2 inst_3429 ( .A1(net_9471), .ZN(net_8488), .A2(net_8487) );
OAI22_X2 inst_1328 ( .B2(net_9943), .ZN(net_1419), .A2(net_1418), .B1(net_1417), .A1(net_195) );
AOI22_X2 inst_9027 ( .B1(net_9527), .A1(net_8002), .B2(net_8001), .ZN(net_7944), .A2(net_7900) );
DFF_X1 inst_8429 ( .Q(net_9582), .D(net_8694), .CK(net_11559) );
INV_X2 inst_6815 ( .ZN(net_7845), .A(net_5998) );
CLKBUF_X2 inst_15434 ( .A(net_15352), .Z(net_15353) );
NAND3_X2 inst_3292 ( .A3(net_9172), .ZN(net_2888), .A1(net_2887), .A2(net_2886) );
DFF_X1 inst_8575 ( .Q(net_9773), .D(net_7140), .CK(net_14835) );
OAI21_X2 inst_1776 ( .B1(net_7884), .ZN(net_7807), .B2(net_7805), .A(net_4173) );
DFF_X2 inst_7751 ( .Q(net_10189), .D(net_6216), .CK(net_15134) );
INV_X4 inst_5024 ( .ZN(net_1943), .A(net_1942) );
NOR4_X2 inst_2335 ( .A4(net_4631), .ZN(net_4453), .A1(net_4333), .A2(net_4004), .A3(net_3142) );
DFF_X2 inst_7715 ( .Q(net_9804), .D(net_6435), .CK(net_14314) );
CLKBUF_X2 inst_13157 ( .A(net_13075), .Z(net_13076) );
OR2_X2 inst_919 ( .A2(net_9859), .A1(net_9858), .ZN(net_3259) );
AND2_X2 inst_10530 ( .ZN(net_3929), .A2(net_3928), .A1(net_3455) );
CLKBUF_X2 inst_12772 ( .A(net_11491), .Z(net_12691) );
SDFF_X2 inst_598 ( .Q(net_9265), .SE(net_4297), .SI(net_148), .D(net_114), .CK(net_12543) );
OAI21_X2 inst_1916 ( .B1(net_7828), .ZN(net_4571), .A(net_4146), .B2(net_4145) );
AOI222_X1 inst_9705 ( .B1(net_9510), .A2(net_8295), .B2(net_8294), .C2(net_8293), .ZN(net_8273), .C1(net_8199), .A1(x2890) );
OAI221_X2 inst_1624 ( .B1(net_10321), .C1(net_7186), .A(net_5637), .B2(net_5591), .ZN(net_5583), .C2(net_4902) );
CLKBUF_X2 inst_14868 ( .A(net_14786), .Z(net_14787) );
CLKBUF_X2 inst_14057 ( .A(net_11437), .Z(net_13976) );
AND2_X2 inst_10595 ( .ZN(net_2365), .A2(net_2364), .A1(net_2203) );
CLKBUF_X2 inst_12403 ( .A(net_12321), .Z(net_12322) );
OAI21_X2 inst_1797 ( .ZN(net_7445), .B1(net_7157), .A(net_6980), .B2(net_6973) );
CLKBUF_X2 inst_10728 ( .A(net_10646), .Z(net_10647) );
NAND3_X4 inst_3167 ( .ZN(net_8578), .A1(net_8559), .A2(net_8550), .A3(net_8549) );
CLKBUF_X2 inst_13501 ( .A(net_13419), .Z(net_13420) );
NAND2_X2 inst_4408 ( .A2(net_10402), .A1(net_10395), .ZN(net_616) );
NOR2_X2 inst_2708 ( .ZN(net_4534), .A2(net_4238), .A1(net_1910) );
CLKBUF_X2 inst_14029 ( .A(net_11579), .Z(net_13948) );
INV_X4 inst_6197 ( .A(net_9319), .ZN(net_563) );
CLKBUF_X2 inst_14694 ( .A(net_14612), .Z(net_14613) );
AOI221_X2 inst_9866 ( .B1(net_9871), .B2(net_9101), .A(net_6945), .C1(net_6944), .ZN(net_6844), .C2(net_242) );
NAND2_X2 inst_3530 ( .A2(net_9626), .A1(net_8975), .ZN(net_8056) );
INV_X2 inst_7205 ( .A(net_9118), .ZN(net_1038) );
INV_X4 inst_5009 ( .ZN(net_7895), .A(net_2608) );
INV_X4 inst_4785 ( .A(net_10385), .ZN(net_5341) );
CLKBUF_X2 inst_13552 ( .A(net_12273), .Z(net_13471) );
DFF_X2 inst_7785 ( .Q(net_9819), .D(net_6511), .CK(net_15705) );
NOR2_X2 inst_2592 ( .A1(net_9381), .ZN(net_7114), .A2(net_6948) );
XNOR2_X2 inst_325 ( .B(net_9654), .ZN(net_3028), .A(net_2829) );
CLKBUF_X2 inst_14861 ( .A(net_14779), .Z(net_14780) );
INV_X4 inst_6502 ( .A(net_10394), .ZN(net_352) );
CLKBUF_X2 inst_12752 ( .A(net_12670), .Z(net_12671) );
DFF_X1 inst_8858 ( .Q(net_9234), .D(net_1038), .CK(net_13590) );
INV_X4 inst_4769 ( .ZN(net_4448), .A(net_4182) );
HA_X1 inst_7331 ( .S(net_7567), .CO(net_7566), .B(net_7470), .A(net_889) );
OAI22_X2 inst_1197 ( .A1(net_7136), .A2(net_5139), .B2(net_5138), .ZN(net_5056), .B1(net_1915) );
NAND4_X2 inst_3116 ( .A2(net_10056), .A1(net_9957), .ZN(net_4129), .A4(net_3477), .A3(net_2114) );
CLKBUF_X2 inst_15624 ( .A(net_15542), .Z(net_15543) );
NAND2_X2 inst_4378 ( .ZN(net_2956), .A1(net_1392), .A2(net_809) );
CLKBUF_X2 inst_14682 ( .A(net_11456), .Z(net_14601) );
AND2_X2 inst_10544 ( .ZN(net_3979), .A1(net_3490), .A2(net_3489) );
AOI222_X1 inst_9682 ( .B1(net_9510), .A2(net_8310), .B2(net_8309), .C2(net_8308), .ZN(net_8305), .C1(net_8229), .A1(x2400) );
INV_X2 inst_6958 ( .A(net_3741), .ZN(net_1874) );
CLKBUF_X2 inst_15824 ( .A(net_15742), .Z(net_15743) );
CLKBUF_X2 inst_15589 ( .A(net_15507), .Z(net_15508) );
CLKBUF_X2 inst_15552 ( .A(net_15470), .Z(net_15471) );
OAI33_X1 inst_955 ( .A3(net_9170), .ZN(net_6840), .B2(net_6839), .A2(net_6839), .B1(net_4452), .A1(net_4376), .B3(net_2542) );
XNOR2_X2 inst_114 ( .ZN(net_7890), .A(net_7772), .B(net_6896) );
CLKBUF_X2 inst_11767 ( .A(net_11685), .Z(net_11686) );
INV_X2 inst_7116 ( .A(net_1374), .ZN(net_989) );
OAI211_X2 inst_2278 ( .C1(net_7136), .C2(net_6542), .ZN(net_6222), .B(net_5749), .A(net_3679) );
CLKBUF_X2 inst_15793 ( .A(net_13391), .Z(net_15712) );
CLKBUF_X2 inst_11041 ( .A(net_10799), .Z(net_10960) );
INV_X4 inst_4866 ( .ZN(net_4071), .A(net_3593) );
CLKBUF_X2 inst_11415 ( .A(net_11253), .Z(net_11334) );
DFF_X2 inst_7924 ( .Q(net_9226), .D(net_5816), .CK(net_13001) );
DFF_X2 inst_7800 ( .Q(net_9915), .D(net_6492), .CK(net_13408) );
AOI22_X2 inst_9519 ( .B1(net_9767), .A1(net_9668), .A2(net_5966), .ZN(net_3803), .B2(net_2462) );
NAND2_X2 inst_4150 ( .ZN(net_2052), .A2(net_2051), .A1(net_887) );
CLKBUF_X2 inst_15157 ( .A(net_11275), .Z(net_15076) );
AOI22_X2 inst_9630 ( .A1(net_9841), .B1(net_9778), .A2(net_6413), .ZN(net_3413), .B2(net_2462) );
INV_X4 inst_5851 ( .ZN(net_1096), .A(net_921) );
CLKBUF_X2 inst_12371 ( .A(net_12289), .Z(net_12290) );
SDFF_X2 inst_534 ( .D(net_9122), .SE(net_933), .CK(net_10908), .SI(x3071), .Q(x1357) );
CLKBUF_X2 inst_12422 ( .A(net_12340), .Z(net_12341) );
INV_X2 inst_6665 ( .ZN(net_8363), .A(net_8306) );
DFF_X1 inst_8636 ( .Q(net_9886), .D(net_7225), .CK(net_14386) );
CLKBUF_X2 inst_13816 ( .A(net_13734), .Z(net_13735) );
CLKBUF_X2 inst_12502 ( .A(net_12420), .Z(net_12421) );
AOI22_X2 inst_9033 ( .B2(net_10276), .ZN(net_7624), .A2(net_7492), .A1(net_7406), .B1(net_890) );
CLKBUF_X2 inst_10682 ( .A(net_10552), .Z(net_10601) );
INV_X2 inst_7117 ( .ZN(net_1444), .A(net_983) );
INV_X4 inst_5618 ( .ZN(net_1453), .A(net_867) );
CLKBUF_X2 inst_13663 ( .A(net_13581), .Z(net_13582) );
CLKBUF_X2 inst_11142 ( .A(net_11060), .Z(net_11061) );
NOR2_X2 inst_2842 ( .ZN(net_2326), .A1(net_2325), .A2(net_1532) );
CLKBUF_X2 inst_15318 ( .A(net_14686), .Z(net_15237) );
INV_X4 inst_5711 ( .A(net_1507), .ZN(net_772) );
INV_X4 inst_5193 ( .ZN(net_3670), .A(net_1544) );
OAI211_X2 inst_2084 ( .C2(net_6778), .ZN(net_6764), .A(net_6391), .B(net_6125), .C1(net_428) );
NOR2_X2 inst_2836 ( .A2(net_2679), .ZN(net_2360), .A1(net_1641) );
NAND2_X2 inst_3792 ( .ZN(net_5015), .A2(net_4687), .A1(net_1167) );
NAND2_X2 inst_4336 ( .A2(net_10263), .ZN(net_2357), .A1(net_1088) );
CLKBUF_X2 inst_12310 ( .A(net_12205), .Z(net_12229) );
CLKBUF_X2 inst_11534 ( .A(net_11452), .Z(net_11453) );
DFF_X2 inst_8203 ( .Q(net_10073), .D(net_4863), .CK(net_11099) );
AND2_X4 inst_10424 ( .A2(net_10280), .ZN(net_4490), .A1(net_4006) );
NOR2_X2 inst_2770 ( .A1(net_9613), .ZN(net_3244), .A2(net_1754) );
CLKBUF_X2 inst_11735 ( .A(net_11344), .Z(net_11654) );
AOI22_X2 inst_9184 ( .A1(net_9874), .B1(net_9775), .B2(net_8041), .A2(net_6141), .ZN(net_6131) );
CLKBUF_X2 inst_14542 ( .A(net_14038), .Z(net_14461) );
CLKBUF_X2 inst_15010 ( .A(net_14928), .Z(net_14929) );
INV_X4 inst_4573 ( .ZN(net_8250), .A(net_8112) );
NAND2_X2 inst_3444 ( .A1(net_9450), .ZN(net_9023), .A2(net_8479) );
INV_X2 inst_7284 ( .A(net_8978), .ZN(net_8976) );
CLKBUF_X2 inst_10848 ( .A(net_10766), .Z(net_10767) );
OR2_X4 inst_803 ( .A1(net_10263), .A2(net_9833), .ZN(net_2204) );
CLKBUF_X2 inst_12011 ( .A(net_10750), .Z(net_11930) );
AOI22_X2 inst_9295 ( .B1(net_9901), .A1(net_5759), .B2(net_5758), .ZN(net_5697), .A2(net_240) );
CLKBUF_X2 inst_14926 ( .A(net_13960), .Z(net_14845) );
INV_X4 inst_4732 ( .ZN(net_4590), .A(net_4297) );
NOR4_X2 inst_2348 ( .ZN(net_2683), .A2(net_2211), .A4(net_2093), .A1(net_1938), .A3(net_1293) );
CLKBUF_X2 inst_15167 ( .A(net_13652), .Z(net_15086) );
NAND2_X2 inst_4021 ( .ZN(net_4876), .A2(net_3071), .A1(net_955) );
AOI211_X2 inst_10312 ( .ZN(net_2498), .A(net_2497), .B(net_2496), .C1(net_2495), .C2(net_1639) );
CLKBUF_X2 inst_11936 ( .A(net_11854), .Z(net_11855) );
CLKBUF_X2 inst_11059 ( .A(net_10949), .Z(net_10978) );
SDFF_X2 inst_662 ( .SI(net_9492), .Q(net_9492), .SE(net_3073), .CK(net_12410), .D(x1911) );
CLKBUF_X2 inst_15590 ( .A(net_15107), .Z(net_15509) );
INV_X2 inst_7156 ( .A(net_3464), .ZN(net_704) );
OAI221_X2 inst_1533 ( .B1(net_10336), .B2(net_9047), .C2(net_7287), .ZN(net_7238), .C1(net_7237), .A(net_6787) );
NAND2_X2 inst_3495 ( .ZN(net_8968), .A2(net_8127), .A1(net_604) );
AOI221_X2 inst_9827 ( .B1(net_9870), .B2(net_9101), .A(net_6945), .C1(net_6944), .ZN(net_6918), .C2(net_241) );
DFF_X2 inst_7741 ( .Q(net_9656), .D(net_6181), .CK(net_11828) );
DFF_X2 inst_8290 ( .QN(net_9606), .D(net_4897), .CK(net_11593) );
CLKBUF_X2 inst_11046 ( .A(net_10964), .Z(net_10965) );
CLKBUF_X2 inst_11114 ( .A(net_11032), .Z(net_11033) );
CLKBUF_X2 inst_12491 ( .A(net_12409), .Z(net_12410) );
DFF_X2 inst_7713 ( .QN(net_9183), .D(net_6250), .CK(net_13583) );
INV_X4 inst_5080 ( .ZN(net_2182), .A(net_1811) );
INV_X4 inst_4666 ( .ZN(net_8990), .A(net_5419) );
CLKBUF_X2 inst_14115 ( .A(net_14033), .Z(net_14034) );
OAI221_X2 inst_1465 ( .ZN(net_7919), .C2(net_7909), .B1(net_7884), .B2(net_7760), .A(net_7559), .C1(net_1314) );
CLKBUF_X2 inst_12653 ( .A(net_12571), .Z(net_12572) );
INV_X4 inst_5030 ( .ZN(net_2595), .A(net_1936) );
XOR2_X1 inst_53 ( .Z(net_2289), .A(net_1560), .B(net_807) );
INV_X4 inst_5265 ( .ZN(net_4083), .A(net_2956) );
CLKBUF_X2 inst_13009 ( .A(net_12927), .Z(net_12928) );
INV_X4 inst_6550 ( .ZN(net_1417), .A(net_195) );
CLKBUF_X2 inst_15069 ( .A(net_14987), .Z(net_14988) );
NOR2_X2 inst_2614 ( .A1(net_9079), .ZN(net_7274), .A2(net_6233) );
NAND2_X4 inst_3337 ( .A2(net_9029), .A1(net_9028), .ZN(net_8529) );
AND2_X2 inst_10513 ( .ZN(net_5313), .A1(net_4988), .A2(net_4708) );
NAND2_X2 inst_4215 ( .A2(net_9850), .ZN(net_3741), .A1(net_619) );
NAND2_X2 inst_4090 ( .A1(net_10471), .ZN(net_3103), .A2(net_2534) );
CLKBUF_X2 inst_15259 ( .A(net_15177), .Z(net_15178) );
OAI22_X2 inst_999 ( .ZN(net_8573), .A2(net_8555), .B2(net_8554), .A1(net_3994), .B1(net_500) );
DFF_X2 inst_7805 ( .Q(net_9922), .D(net_6485), .CK(net_14226) );
CLKBUF_X2 inst_12378 ( .A(net_12296), .Z(net_12297) );
DFF_X2 inst_8083 ( .QN(net_9194), .D(net_5371), .CK(net_13562) );
CLKBUF_X2 inst_14512 ( .A(net_13663), .Z(net_14431) );
OAI211_X2 inst_2111 ( .C2(net_6778), .ZN(net_6737), .A(net_6376), .B(net_6107), .C1(net_420) );
OAI21_X2 inst_1846 ( .ZN(net_5987), .B2(net_5974), .A(net_2081), .B1(net_1376) );
DFF_X1 inst_8419 ( .D(net_8775), .Q(net_244), .CK(net_12691) );
CLKBUF_X2 inst_13943 ( .A(net_11301), .Z(net_13862) );
OAI211_X2 inst_2139 ( .C2(net_6778), .ZN(net_6709), .A(net_6409), .B(net_6072), .C1(net_5090) );
NAND2_X2 inst_4278 ( .A1(net_6960), .ZN(net_2401), .A2(net_1349) );
OAI221_X2 inst_1463 ( .C1(net_8117), .B2(net_7974), .C2(net_7973), .ZN(net_7958), .A(net_7957), .B1(net_2588) );
CLKBUF_X2 inst_14242 ( .A(net_10576), .Z(net_14161) );
AOI21_X2 inst_10236 ( .B2(net_10439), .ZN(net_1701), .A(net_1700), .B1(net_518) );
XNOR2_X2 inst_186 ( .ZN(net_5209), .A(net_4548), .B(net_1439) );
AOI22_X2 inst_9665 ( .B2(net_10089), .A2(net_10081), .B1(net_10071), .A1(net_10063), .ZN(net_965) );
NAND2_X2 inst_4271 ( .A1(net_4566), .ZN(net_2352), .A2(net_1352) );
CLKBUF_X2 inst_13463 ( .A(net_13381), .Z(net_13382) );
CLKBUF_X2 inst_10756 ( .A(net_10561), .Z(net_10675) );
OR2_X4 inst_759 ( .ZN(net_5134), .A1(net_4475), .A2(net_4367) );
CLKBUF_X2 inst_11655 ( .A(net_11573), .Z(net_11574) );
AOI221_X2 inst_9820 ( .B1(net_9866), .B2(net_9101), .A(net_6945), .C1(net_6944), .ZN(net_6934), .C2(net_237) );
NAND4_X2 inst_3071 ( .ZN(net_5254), .A2(net_4696), .A1(net_4487), .A3(net_3817), .A4(net_3501) );
AND2_X4 inst_10395 ( .ZN(net_7155), .A1(net_6203), .A2(net_6202) );
CLKBUF_X2 inst_13192 ( .A(net_10869), .Z(net_13111) );
CLKBUF_X2 inst_11963 ( .A(net_11881), .Z(net_11882) );
CLKBUF_X2 inst_13536 ( .A(net_13454), .Z(net_13455) );
DFF_X2 inst_8283 ( .QN(net_10247), .D(net_4925), .CK(net_12178) );
OR2_X2 inst_863 ( .A1(net_10398), .ZN(net_7864), .A2(net_7863) );
DFF_X1 inst_8669 ( .D(net_6764), .Q(net_101), .CK(net_13224) );
INV_X4 inst_6315 ( .A(net_10152), .ZN(net_775) );
OAI222_X2 inst_1385 ( .B1(net_7732), .A2(net_7731), .C2(net_7730), .ZN(net_6000), .B2(net_5203), .A1(net_4199), .C1(net_1837) );
CLKBUF_X2 inst_15288 ( .A(net_12892), .Z(net_15207) );
INV_X4 inst_6513 ( .A(net_10268), .ZN(net_7031) );
INV_X4 inst_5921 ( .ZN(net_1478), .A(net_786) );
INV_X4 inst_5770 ( .ZN(net_721), .A(net_720) );
OAI221_X2 inst_1573 ( .C1(net_10318), .C2(net_9047), .B2(net_7287), .B1(net_7211), .ZN(net_7172), .A(net_6843) );
INV_X4 inst_6596 ( .ZN(net_4022), .A(net_117) );
INV_X4 inst_5521 ( .ZN(net_1252), .A(net_1190) );
DFF_X2 inst_8394 ( .Q(net_9155), .CK(net_11799), .D(x3599) );
OAI222_X2 inst_1390 ( .B1(net_7665), .A2(net_7664), .C2(net_7663), .ZN(net_5821), .B2(net_4933), .A1(net_3426), .C1(net_713) );
AOI22_X2 inst_9274 ( .B1(net_10005), .ZN(net_5753), .A1(net_5743), .B2(net_5742), .A2(net_245) );
NAND2_X2 inst_3586 ( .ZN(net_7393), .A2(net_7392), .A1(net_5903) );
CLKBUF_X2 inst_13652 ( .A(net_13570), .Z(net_13571) );
XNOR2_X2 inst_229 ( .ZN(net_4402), .A(net_3954), .B(net_3223) );
CLKBUF_X2 inst_14625 ( .A(net_14543), .Z(net_14544) );
AOI22_X2 inst_9124 ( .A1(net_9708), .A2(net_6404), .ZN(net_6365), .B2(net_5263), .B1(net_148) );
DFF_X2 inst_7744 ( .Q(net_9184), .D(net_6295), .CK(net_11320) );
AOI221_X2 inst_9974 ( .C2(net_10088), .B2(net_10087), .C1(net_10070), .B1(net_10069), .ZN(net_4576), .A(net_4128) );
INV_X2 inst_7203 ( .A(net_9395), .ZN(net_8199) );
OAI211_X2 inst_2282 ( .C1(net_7136), .C2(net_6480), .ZN(net_6212), .B(net_5736), .A(net_3679) );
CLKBUF_X2 inst_12920 ( .A(net_12838), .Z(net_12839) );
AOI22_X2 inst_9596 ( .B1(net_9776), .A2(net_6413), .ZN(net_3498), .B2(net_2462), .A1(net_1165) );
INV_X4 inst_4992 ( .ZN(net_2223), .A(net_2222) );
INV_X4 inst_4689 ( .ZN(net_4838), .A(net_4654) );
CLKBUF_X2 inst_11719 ( .A(net_11637), .Z(net_11638) );
INV_X4 inst_6151 ( .A(net_10469), .ZN(net_686) );
CLKBUF_X2 inst_14594 ( .A(net_14512), .Z(net_14513) );
AOI22_X2 inst_9187 ( .A1(net_9877), .B1(net_9778), .A2(net_8042), .B2(net_6140), .ZN(net_6127) );
OAI211_X2 inst_2131 ( .C2(net_6778), .ZN(net_6717), .A(net_6341), .B(net_6080), .C1(net_449) );
INV_X4 inst_5718 ( .A(net_3385), .ZN(net_905) );
CLKBUF_X2 inst_12007 ( .A(net_11925), .Z(net_11926) );
AOI221_X2 inst_9949 ( .B1(net_6255), .ZN(net_5177), .B2(net_5174), .C2(net_5173), .A(net_4488), .C1(net_203) );
INV_X2 inst_7297 ( .ZN(net_9054), .A(net_9053) );
DFF_X1 inst_8804 ( .QN(net_9530), .D(net_3923), .CK(net_12758) );
XNOR2_X2 inst_169 ( .ZN(net_5763), .A(net_4922), .B(net_1202) );
AOI22_X2 inst_9453 ( .B1(net_10399), .A1(net_9825), .A2(net_6413), .B2(net_4062), .ZN(net_3983) );
INV_X4 inst_6158 ( .A(net_10331), .ZN(net_600) );
XNOR2_X2 inst_421 ( .ZN(net_3223), .B(net_1993), .A(net_1450) );
CLKBUF_X2 inst_12880 ( .A(net_12798), .Z(net_12799) );
CLKBUF_X2 inst_11263 ( .A(net_10655), .Z(net_11182) );
CLKBUF_X2 inst_11748 ( .A(net_10667), .Z(net_11667) );
DFF_X2 inst_8014 ( .QN(net_10229), .D(net_5490), .CK(net_14463) );
SDFF_X2 inst_555 ( .SI(net_9359), .Q(net_9359), .D(net_9157), .SE(net_7248), .CK(net_15337) );
INV_X2 inst_7016 ( .A(net_1756), .ZN(net_1559) );
OR2_X4 inst_816 ( .ZN(net_2148), .A2(net_848), .A1(net_776) );
CLKBUF_X2 inst_11000 ( .A(net_10748), .Z(net_10919) );
CLKBUF_X2 inst_12911 ( .A(net_12829), .Z(net_12830) );
AOI211_X2 inst_10293 ( .C2(net_9197), .A(net_6192), .ZN(net_4537), .B(net_4224), .C1(net_3607) );
CLKBUF_X2 inst_12978 ( .A(net_12896), .Z(net_12897) );
NOR2_X2 inst_2798 ( .A2(net_3111), .ZN(net_2893), .A1(net_2251) );
OAI22_X2 inst_1184 ( .A1(net_7198), .A2(net_5107), .B2(net_5105), .ZN(net_5074), .B1(net_5073) );
CLKBUF_X2 inst_12903 ( .A(net_12821), .Z(net_12822) );
CLKBUF_X2 inst_12692 ( .A(net_12610), .Z(net_12611) );
AOI22_X2 inst_9352 ( .B1(net_10012), .A2(net_5743), .B2(net_5742), .ZN(net_5600), .A1(net_252) );
INV_X4 inst_4685 ( .ZN(net_4992), .A(net_4991) );
CLKBUF_X2 inst_14325 ( .A(net_11369), .Z(net_14244) );
CLKBUF_X2 inst_13694 ( .A(net_13612), .Z(net_13613) );
INV_X4 inst_6157 ( .A(net_9248), .ZN(net_746) );
DFF_X2 inst_7596 ( .Q(net_10296), .D(net_7445), .CK(net_14562) );
CLKBUF_X2 inst_12523 ( .A(net_12441), .Z(net_12442) );
DFF_X2 inst_8197 ( .QN(net_9743), .D(net_5109), .CK(net_12874) );
DFF_X2 inst_7796 ( .Q(net_9911), .D(net_6497), .CK(net_12792) );
CLKBUF_X2 inst_14999 ( .A(net_14854), .Z(net_14918) );
OAI22_X2 inst_1108 ( .A1(net_7219), .ZN(net_6151), .B2(net_5877), .A2(net_5302), .B1(net_4662) );
INV_X4 inst_6580 ( .A(net_10359), .ZN(net_762) );
CLKBUF_X2 inst_11863 ( .A(net_11781), .Z(net_11782) );
AOI22_X2 inst_9480 ( .B1(net_9782), .A1(net_9715), .ZN(net_3843), .A2(net_3039), .B2(net_2462) );
INV_X4 inst_5148 ( .ZN(net_1906), .A(net_1586) );
INV_X4 inst_5140 ( .A(net_4382), .ZN(net_1932) );
CLKBUF_X2 inst_11578 ( .A(net_11496), .Z(net_11497) );
DFF_X1 inst_8756 ( .Q(net_10275), .D(net_5245), .CK(net_11771) );
CLKBUF_X2 inst_12273 ( .A(net_10849), .Z(net_12192) );
INV_X4 inst_4534 ( .ZN(net_8872), .A(net_8778) );
DFF_X2 inst_7521 ( .QN(net_9242), .D(net_7829), .CK(net_13525) );
CLKBUF_X2 inst_12931 ( .A(net_12849), .Z(net_12850) );
NAND2_X2 inst_3991 ( .A2(net_10337), .ZN(net_3178), .A1(net_3177) );
DFF_X2 inst_8286 ( .Q(net_10291), .D(net_4816), .CK(net_12925) );
CLKBUF_X2 inst_13620 ( .A(net_13538), .Z(net_13539) );
AOI22_X2 inst_9546 ( .A1(net_10404), .B1(net_9865), .A2(net_4062), .ZN(net_3775), .B2(net_2973) );
CLKBUF_X2 inst_14812 ( .A(net_14730), .Z(net_14731) );
CLKBUF_X2 inst_11422 ( .A(net_11340), .Z(net_11341) );
CLKBUF_X2 inst_15661 ( .A(net_15579), .Z(net_15580) );
DFF_X1 inst_8604 ( .Q(net_9792), .D(net_7194), .CK(net_13297) );
INV_X4 inst_6203 ( .A(net_9246), .ZN(net_755) );
DFF_X1 inst_8617 ( .Q(net_9680), .D(net_7268), .CK(net_13286) );
NAND2_X4 inst_3343 ( .ZN(net_8523), .A1(net_8468), .A2(net_8467) );
AOI222_X1 inst_9718 ( .A2(net_7142), .ZN(net_5269), .B1(net_5268), .C1(net_3169), .A1(net_3070), .B2(net_2759), .C2(net_2634) );
NAND2_X2 inst_4140 ( .A2(net_9086), .A1(net_3976), .ZN(net_2830) );
CLKBUF_X2 inst_13340 ( .A(net_12033), .Z(net_13259) );
OAI221_X2 inst_1543 ( .B2(net_9047), .C2(net_7287), .ZN(net_7220), .C1(net_7219), .A(net_6796), .B1(net_938) );
CLKBUF_X2 inst_13892 ( .A(net_13810), .Z(net_13811) );
INV_X2 inst_7290 ( .A(net_8985), .ZN(net_8984) );
NAND2_X2 inst_4219 ( .A1(net_8687), .ZN(net_1671), .A2(net_114) );
NOR2_X2 inst_2801 ( .ZN(net_3040), .A2(net_2830), .A1(net_269) );
OAI22_X2 inst_1118 ( .ZN(net_5991), .A2(net_4965), .B2(net_4964), .B1(net_3708), .A1(net_2325) );
AOI22_X2 inst_9153 ( .A1(net_9750), .A2(net_6420), .ZN(net_6330), .B2(net_5263), .B1(net_186) );
NOR4_X2 inst_2303 ( .A1(net_8945), .ZN(net_8708), .A4(net_8695), .A2(net_8136), .A3(net_6160) );
CLKBUF_X2 inst_15341 ( .A(net_15259), .Z(net_15260) );
CLKBUF_X2 inst_13714 ( .A(net_13632), .Z(net_13633) );
INV_X2 inst_6978 ( .A(net_2064), .ZN(net_1678) );
INV_X4 inst_6109 ( .A(net_10033), .ZN(net_1036) );
DFF_X2 inst_8090 ( .QN(net_10531), .D(net_5020), .CK(net_14890) );
CLKBUF_X2 inst_10948 ( .A(net_10866), .Z(net_10867) );
SDFF_X2 inst_473 ( .D(net_9576), .SI(net_2598), .SE(net_758), .Q(net_250), .CK(net_15043) );
CLKBUF_X2 inst_15114 ( .A(net_14038), .Z(net_15033) );
CLKBUF_X2 inst_14765 ( .A(net_11414), .Z(net_14684) );
AOI21_X2 inst_10140 ( .ZN(net_4245), .A(net_3937), .B2(net_3461), .B1(net_1276) );
OAI211_X2 inst_2211 ( .C1(net_7201), .C2(net_6501), .ZN(net_6494), .B(net_5554), .A(net_3527) );
NAND2_X2 inst_3771 ( .A2(net_8511), .A1(net_7095), .ZN(net_5329) );
NAND4_X2 inst_3083 ( .A3(net_10490), .ZN(net_4793), .A4(net_4641), .A2(net_4639), .A1(net_4369) );
AOI22_X2 inst_9170 ( .ZN(net_7052), .A2(net_5746), .B2(net_5745), .B1(net_4168), .A1(net_2405) );
OAI221_X2 inst_1695 ( .B1(net_7224), .C2(net_5591), .A(net_5575), .ZN(net_5461), .B2(net_4902), .C1(net_1512) );
INV_X4 inst_5557 ( .ZN(net_1235), .A(net_925) );
CLKBUF_X2 inst_12609 ( .A(net_10567), .Z(net_12528) );
CLKBUF_X2 inst_15336 ( .A(net_15254), .Z(net_15255) );
AOI221_X2 inst_9917 ( .B1(net_10506), .C1(net_9664), .B2(net_6415), .ZN(net_5968), .C2(net_5966), .A(net_5254) );
CLKBUF_X2 inst_12942 ( .A(net_12249), .Z(net_12861) );
AOI222_X1 inst_9724 ( .C1(net_9869), .B1(net_9770), .A2(net_6413), .ZN(net_4051), .A1(net_4050), .C2(net_2973), .B2(net_2462) );
CLKBUF_X2 inst_15371 ( .A(net_14041), .Z(net_15290) );
CLKBUF_X2 inst_11034 ( .A(net_10952), .Z(net_10953) );
OAI222_X2 inst_1404 ( .B2(net_7732), .A2(net_7731), .C2(net_7730), .ZN(net_5326), .B1(net_4387), .A1(net_3669), .C1(net_1258) );
NOR2_X2 inst_2989 ( .A1(net_10460), .ZN(net_2397), .A2(net_921) );
INV_X4 inst_5880 ( .ZN(net_2862), .A(net_779) );
NAND2_X2 inst_3479 ( .A1(net_9458), .A2(net_8951), .ZN(net_8433) );
OAI222_X2 inst_1339 ( .A1(net_7732), .B2(net_7731), .C2(net_7730), .ZN(net_7626), .A2(net_7469), .B1(net_4989), .C1(net_1823) );
CLKBUF_X2 inst_11235 ( .A(net_11153), .Z(net_11154) );
NAND2_X2 inst_4284 ( .ZN(net_1802), .A2(net_1342), .A1(net_715) );
INV_X4 inst_4971 ( .ZN(net_3630), .A(net_2791) );
INV_X4 inst_4704 ( .A(net_6680), .ZN(net_5363) );
INV_X4 inst_4724 ( .ZN(net_4614), .A(net_4493) );
CLKBUF_X2 inst_13512 ( .A(net_13430), .Z(net_13431) );
MUX2_X1 inst_4467 ( .S(net_6041), .A(net_5953), .B(x6220), .Z(x329) );
NAND2_X2 inst_3575 ( .A1(net_7783), .ZN(net_7690), .A2(net_7556) );
AOI22_X2 inst_9238 ( .A1(net_9939), .B1(net_9840), .B2(net_8041), .A2(net_6111), .ZN(net_6073) );
INV_X8 inst_4493 ( .ZN(net_7089), .A(net_6164) );
NAND2_X2 inst_3654 ( .A2(net_8659), .ZN(net_8327), .A1(net_4413) );
OAI22_X2 inst_977 ( .ZN(net_8799), .A2(net_8796), .B2(net_7648), .B1(net_2809), .A1(net_1314) );
DFF_X1 inst_8484 ( .Q(net_9625), .D(net_7946), .CK(net_15012) );
AOI21_X2 inst_10180 ( .ZN(net_3566), .B1(net_3565), .A(net_3314), .B2(net_2844) );
INV_X2 inst_7251 ( .ZN(net_353), .A(net_183) );
INV_X2 inst_6901 ( .A(net_2720), .ZN(net_2363) );
INV_X4 inst_5669 ( .A(net_10439), .ZN(net_1298) );
INV_X4 inst_4802 ( .ZN(net_4003), .A(net_3648) );
CLKBUF_X2 inst_10941 ( .A(net_10788), .Z(net_10860) );
XNOR2_X2 inst_297 ( .ZN(net_3333), .B(net_3332), .A(net_3312) );
CLKBUF_X2 inst_15402 ( .A(net_15320), .Z(net_15321) );
OAI222_X2 inst_1395 ( .A2(net_7732), .C2(net_7731), .B2(net_7730), .ZN(net_5703), .A1(net_2861), .C1(net_2298), .B1(net_1163) );
NOR2_X4 inst_2477 ( .A2(net_9591), .A1(net_9082), .ZN(net_5383) );
CLKBUF_X2 inst_13933 ( .A(net_13851), .Z(net_13852) );
CLKBUF_X2 inst_13145 ( .A(net_11540), .Z(net_13064) );
CLKBUF_X2 inst_11728 ( .A(net_11646), .Z(net_11647) );
CLKBUF_X2 inst_14660 ( .A(net_14578), .Z(net_14579) );
INV_X4 inst_5460 ( .ZN(net_1263), .A(net_1050) );
CLKBUF_X2 inst_11424 ( .A(net_10947), .Z(net_11343) );
DFF_X2 inst_8322 ( .Q(net_10503), .D(net_3926), .CK(net_12323) );
INV_X4 inst_4838 ( .ZN(net_3527), .A(net_3298) );
OAI211_X2 inst_2188 ( .C1(net_7231), .C2(net_6542), .ZN(net_6521), .B(net_5616), .A(net_3679) );
NAND2_X2 inst_3436 ( .A1(net_9483), .ZN(net_8893), .A2(net_8421) );
OAI21_X2 inst_1875 ( .B2(net_9075), .ZN(net_5267), .A(net_5266), .B1(net_5265) );
NAND2_X4 inst_3351 ( .A2(net_8925), .ZN(net_8505), .A1(net_8387) );
CLKBUF_X2 inst_13057 ( .A(net_12975), .Z(net_12976) );
AND2_X4 inst_10466 ( .ZN(net_2712), .A2(net_914), .A1(net_313) );
AOI21_X2 inst_10005 ( .B2(net_9583), .B1(net_9582), .ZN(net_8746), .A(net_5813) );
NAND3_X2 inst_3190 ( .A1(net_9611), .ZN(net_7909), .A3(net_7605), .A2(net_2460) );
XNOR2_X2 inst_162 ( .ZN(net_5975), .A(net_5974), .B(net_2082) );
DFF_X1 inst_8459 ( .QN(net_10488), .D(net_7980), .CK(net_11139) );
NAND3_X2 inst_3308 ( .ZN(net_1829), .A2(net_1828), .A1(net_1207), .A3(net_985) );
CLKBUF_X2 inst_10873 ( .A(net_10791), .Z(net_10792) );
NAND2_X2 inst_3397 ( .A2(net_9579), .ZN(net_8667), .A1(net_2225) );
CLKBUF_X2 inst_14903 ( .A(net_14821), .Z(net_14822) );
DFF_X2 inst_7373 ( .Q(net_9364), .D(net_8684), .CK(net_11923) );
CLKBUF_X2 inst_13286 ( .A(net_11803), .Z(net_13205) );
INV_X2 inst_7302 ( .A(net_9073), .ZN(net_9070) );
INV_X4 inst_5484 ( .ZN(net_1435), .A(net_999) );
CLKBUF_X2 inst_13387 ( .A(net_13305), .Z(net_13306) );
CLKBUF_X2 inst_11544 ( .A(net_11462), .Z(net_11463) );
NAND2_X1 inst_4421 ( .ZN(net_8456), .A1(net_8455), .A2(net_8454) );
NOR2_X2 inst_2829 ( .A1(net_2964), .A2(net_2540), .ZN(net_2468) );
NAND2_X2 inst_3819 ( .A1(net_10088), .A2(net_4534), .ZN(net_4519) );
CLKBUF_X2 inst_11383 ( .A(net_11112), .Z(net_11302) );
DFF_X1 inst_8448 ( .QN(net_9434), .D(net_8144), .CK(net_12686) );
NAND2_X2 inst_4233 ( .A2(net_10267), .ZN(net_2639), .A1(net_1551) );
NAND2_X2 inst_3668 ( .A2(net_10275), .A1(net_10274), .ZN(net_7067) );
INV_X2 inst_7128 ( .A(net_9196), .ZN(net_1461) );
INV_X4 inst_5905 ( .A(net_2521), .ZN(net_595) );
NAND2_X2 inst_3968 ( .ZN(net_3379), .A2(net_3378), .A1(net_617) );
DFF_X2 inst_8208 ( .Q(net_10533), .D(net_4878), .CK(net_12614) );
CLKBUF_X2 inst_13010 ( .A(net_10664), .Z(net_12929) );
CLKBUF_X2 inst_12086 ( .A(net_12004), .Z(net_12005) );
INV_X4 inst_4633 ( .ZN(net_7054), .A(net_6616) );
DFF_X2 inst_8143 ( .QN(net_9943), .D(net_5114), .CK(net_12490) );
OAI22_X2 inst_1098 ( .A1(net_9193), .A2(net_6299), .B2(net_6298), .ZN(net_6295), .B1(net_5443) );
INV_X2 inst_7077 ( .ZN(net_1203), .A(net_1202) );
NAND2_X2 inst_4149 ( .ZN(net_2057), .A1(net_2056), .A2(net_1373) );
DFF_X2 inst_8113 ( .Q(net_10038), .D(net_5093), .CK(net_11936) );
CLKBUF_X2 inst_14871 ( .A(net_14789), .Z(net_14790) );
AOI21_X2 inst_10051 ( .ZN(net_7309), .A(net_7308), .B2(net_7077), .B1(net_1926) );
NOR3_X2 inst_2443 ( .ZN(net_3245), .A1(net_1897), .A3(net_1736), .A2(net_1049) );
INV_X2 inst_6660 ( .ZN(net_8408), .A(net_8407) );
CLKBUF_X2 inst_10915 ( .A(net_10781), .Z(net_10834) );
DFF_X2 inst_8027 ( .QN(net_10434), .D(net_5474), .CK(net_13637) );
INV_X4 inst_6411 ( .A(net_10438), .ZN(net_1118) );
OR2_X4 inst_723 ( .A2(net_8315), .ZN(net_8267), .A1(net_8266) );
CLKBUF_X2 inst_10990 ( .A(net_10856), .Z(net_10909) );
AOI22_X2 inst_9525 ( .B1(net_9900), .A2(net_6442), .A1(net_6314), .B2(net_4969), .ZN(net_3796) );
DFF_X1 inst_8769 ( .D(net_4972), .CK(net_11061), .Q(x1058) );
SDFF_X2 inst_618 ( .Q(net_9459), .D(net_9459), .SE(net_3293), .CK(net_12458), .SI(x1974) );
NOR3_X2 inst_2444 ( .ZN(net_3248), .A1(net_1909), .A3(net_1735), .A2(net_990) );
CLKBUF_X2 inst_11980 ( .A(net_10937), .Z(net_11899) );
NAND2_X2 inst_3893 ( .ZN(net_4120), .A2(net_3969), .A1(net_680) );
CLKBUF_X2 inst_11616 ( .A(net_11392), .Z(net_11535) );
CLKBUF_X2 inst_11055 ( .A(net_10973), .Z(net_10974) );
NAND4_X2 inst_3057 ( .ZN(net_5729), .A4(net_4772), .A3(net_4216), .A2(net_3849), .A1(net_3466) );
CLKBUF_X2 inst_13274 ( .A(net_11874), .Z(net_13193) );
INV_X4 inst_5777 ( .ZN(net_710), .A(net_709) );
NOR2_X4 inst_2462 ( .A2(net_9011), .A1(net_9010), .ZN(net_8740) );
INV_X2 inst_6706 ( .A(net_8185), .ZN(net_8148) );
SDFF_X2 inst_474 ( .D(net_9575), .SI(net_1175), .SE(net_758), .Q(net_249), .CK(net_11572) );
DFF_X2 inst_7894 ( .QN(net_10100), .D(net_6020), .CK(net_14800) );
OAI211_X2 inst_2067 ( .ZN(net_7440), .C2(net_7439), .C1(net_7435), .A(net_7150), .B(net_2793) );
INV_X4 inst_5561 ( .ZN(net_1664), .A(net_922) );
CLKBUF_X2 inst_14651 ( .A(net_14569), .Z(net_14570) );
SDFF_X2 inst_626 ( .Q(net_9446), .D(net_9446), .SE(net_3293), .CK(net_14161), .SI(x2767) );
CLKBUF_X2 inst_15560 ( .A(net_13668), .Z(net_15479) );
CLKBUF_X2 inst_14497 ( .A(net_11739), .Z(net_14416) );
CLKBUF_X2 inst_13075 ( .A(net_12332), .Z(net_12994) );
DFF_X2 inst_8268 ( .Q(net_10392), .D(net_4809), .CK(net_13171) );
CLKBUF_X2 inst_11539 ( .A(net_11457), .Z(net_11458) );
AOI221_X2 inst_9879 ( .B1(net_9786), .B2(net_9098), .A(net_6940), .C2(net_6939), .ZN(net_6820), .C1(net_256) );
DFF_X2 inst_7476 ( .D(net_8072), .Q(net_210), .CK(net_12905) );
NOR2_X2 inst_2777 ( .ZN(net_4044), .A2(net_3891), .A1(net_3172) );
CLKBUF_X2 inst_12283 ( .A(net_12201), .Z(net_12202) );
INV_X2 inst_6830 ( .ZN(net_4075), .A(net_4074) );
INV_X2 inst_6784 ( .A(net_9252), .ZN(net_5805) );
AOI21_X2 inst_10247 ( .ZN(net_8867), .B1(net_4558), .B2(net_2344), .A(net_2343) );
NOR3_X2 inst_2446 ( .A2(net_5719), .A3(net_5718), .ZN(net_2741), .A1(net_2175) );
CLKBUF_X2 inst_13602 ( .A(net_13520), .Z(net_13521) );
INV_X4 inst_5046 ( .ZN(net_2610), .A(net_1910) );
DFF_X1 inst_8880 ( .D(net_10513), .QN(net_10453), .CK(net_11195) );
DFF_X1 inst_8452 ( .Q(net_9524), .D(net_8077), .CK(net_15041) );
DFF_X2 inst_7840 ( .Q(net_9916), .D(net_6491), .CK(net_13403) );
CLKBUF_X2 inst_14128 ( .A(net_14046), .Z(net_14047) );
CLKBUF_X2 inst_11457 ( .A(net_11375), .Z(net_11376) );
CLKBUF_X2 inst_13070 ( .A(net_12988), .Z(net_12989) );
CLKBUF_X2 inst_12641 ( .A(net_12559), .Z(net_12560) );
CLKBUF_X2 inst_15549 ( .A(net_15467), .Z(net_15468) );
OR2_X4 inst_798 ( .A1(net_10474), .ZN(net_2206), .A2(net_2205) );
CLKBUF_X2 inst_14260 ( .A(net_14178), .Z(net_14179) );
CLKBUF_X2 inst_12648 ( .A(net_10648), .Z(net_12567) );
INV_X4 inst_5210 ( .A(net_5993), .ZN(net_5930) );
INV_X4 inst_6613 ( .ZN(net_8929), .A(net_8643) );
NAND2_X2 inst_4340 ( .ZN(net_2098), .A1(net_892), .A2(net_313) );
CLKBUF_X2 inst_12767 ( .A(net_12685), .Z(net_12686) );
OAI222_X1 inst_1434 ( .ZN(net_7844), .A2(net_7737), .A1(net_7728), .B2(net_7727), .C2(net_7726), .B1(net_6163), .C1(net_1106) );
CLKBUF_X2 inst_12727 ( .A(net_11741), .Z(net_12646) );
INV_X4 inst_5464 ( .A(net_5790), .ZN(net_1399) );
OAI21_X2 inst_1886 ( .B2(net_10236), .A(net_10235), .ZN(net_4930), .B1(net_4929) );
CLKBUF_X2 inst_14089 ( .A(net_14007), .Z(net_14008) );
AOI21_X2 inst_10211 ( .B1(net_2710), .ZN(net_2438), .B2(net_2437), .A(net_924) );
CLKBUF_X2 inst_12889 ( .A(net_12807), .Z(net_12808) );
DFF_X1 inst_8831 ( .QN(net_9608), .D(net_2999), .CK(net_15389) );
DFF_X1 inst_8778 ( .QN(net_10378), .D(net_4683), .CK(net_12149) );
NAND2_X2 inst_4349 ( .A2(net_10225), .ZN(net_1017), .A1(net_1016) );
OAI221_X2 inst_1457 ( .C1(net_9081), .B2(net_7974), .C2(net_7973), .ZN(net_7970), .A(net_7969), .B1(net_2591) );
DFF_X2 inst_8366 ( .QN(net_8843), .D(net_1492), .CK(net_10955) );
DFF_X1 inst_8627 ( .Q(net_9786), .D(net_7223), .CK(net_13361) );
INV_X2 inst_7110 ( .ZN(net_1008), .A(net_1007) );
OAI21_X2 inst_1818 ( .ZN(net_7078), .B2(net_6648), .A(net_2345), .B1(net_1627) );
AND2_X2 inst_10552 ( .ZN(net_3341), .A2(net_3340), .A1(net_3322) );
CLKBUF_X2 inst_10705 ( .A(net_10616), .Z(net_10624) );
CLKBUF_X2 inst_14706 ( .A(net_14624), .Z(net_14625) );
CLKBUF_X2 inst_13244 ( .A(net_13162), .Z(net_13163) );
AOI211_X2 inst_10264 ( .ZN(net_7836), .A(net_7714), .C1(net_7424), .B(net_7342), .C2(net_7329) );
DFF_X2 inst_8209 ( .Q(net_10387), .D(net_4810), .CK(net_15227) );
CLKBUF_X2 inst_11254 ( .A(net_11172), .Z(net_11173) );
NAND2_X2 inst_3662 ( .ZN(net_6912), .A2(net_6261), .A1(net_2659) );
OAI21_X2 inst_1766 ( .B2(net_8246), .ZN(net_8163), .A(net_8109), .B1(net_2570) );
NOR2_X2 inst_2670 ( .ZN(net_5233), .A2(net_4939), .A1(net_274) );
CLKBUF_X2 inst_15726 ( .A(net_15644), .Z(net_15645) );
CLKBUF_X2 inst_13888 ( .A(net_13806), .Z(net_13807) );
CLKBUF_X2 inst_10983 ( .A(net_10901), .Z(net_10902) );
DFF_X2 inst_8380 ( .D(net_10324), .QN(net_8841), .CK(net_11054) );
DFF_X2 inst_8216 ( .Q(net_10499), .D(net_4882), .CK(net_13177) );
NOR2_X2 inst_2974 ( .ZN(net_1388), .A2(net_1036), .A1(net_1035) );
CLKBUF_X2 inst_15398 ( .A(net_15316), .Z(net_15317) );
OAI21_X2 inst_1895 ( .B1(net_7124), .B2(net_4862), .ZN(net_4857), .A(net_4529) );
AOI22_X2 inst_9639 ( .A1(net_10078), .B1(net_9965), .A2(net_5319), .ZN(net_3403), .B2(net_2541) );
DFF_X1 inst_8476 ( .QN(net_9601), .D(net_7862), .CK(net_13800) );
NOR2_X2 inst_2730 ( .A1(net_9238), .ZN(net_4249), .A2(net_3896) );
INV_X4 inst_4548 ( .ZN(net_8620), .A(net_8578) );
OR2_X4 inst_737 ( .A1(net_9099), .ZN(net_7295), .A2(net_4904) );
CLKBUF_X2 inst_11725 ( .A(net_11643), .Z(net_11644) );
OR2_X2 inst_876 ( .A1(net_10398), .ZN(net_6971), .A2(net_6970) );
CLKBUF_X2 inst_11178 ( .A(net_10686), .Z(net_11097) );
NOR2_X2 inst_2979 ( .A1(net_10464), .A2(net_1118), .ZN(net_1018) );
CLKBUF_X1 inst_8990 ( .A(x185142), .Z(x957) );
INV_X4 inst_4727 ( .ZN(net_5998), .A(net_5012) );
SDFF_X2 inst_545 ( .D(net_9140), .SE(net_933), .CK(net_10660), .SI(x1974), .Q(x1179) );
CLKBUF_X2 inst_15819 ( .A(net_14457), .Z(net_15738) );
DFF_X2 inst_8373 ( .D(net_1626), .Q(net_262), .CK(net_12560) );
AOI21_X2 inst_10189 ( .B2(net_7437), .ZN(net_3349), .A(net_3348), .B1(net_3347) );
DFF_X2 inst_8132 ( .QN(net_9844), .D(net_5125), .CK(net_12884) );
NOR3_X2 inst_2433 ( .A3(net_9622), .A1(net_4299), .ZN(net_3525), .A2(net_1356) );
INV_X2 inst_6854 ( .A(net_7439), .ZN(net_3371) );
CLKBUF_X2 inst_11665 ( .A(net_11583), .Z(net_11584) );
CLKBUF_X2 inst_14475 ( .A(net_14393), .Z(net_14394) );
CLKBUF_X2 inst_12188 ( .A(net_12106), .Z(net_12107) );
CLKBUF_X2 inst_11751 ( .A(net_11669), .Z(net_11670) );
INV_X2 inst_6682 ( .ZN(net_8346), .A(net_8280) );
CLKBUF_X2 inst_13595 ( .A(net_13316), .Z(net_13514) );
AOI221_X2 inst_9845 ( .A(net_6889), .B2(net_6888), .C2(net_6887), .ZN(net_6873), .B1(net_5833), .C1(x5790) );
SDFF_X2 inst_562 ( .D(net_9150), .SE(net_933), .CK(net_11053), .SI(x1418), .Q(x1095) );
NOR2_X4 inst_2480 ( .A1(net_9040), .A2(net_8869), .ZN(net_1715) );
DFF_X2 inst_7832 ( .Q(net_10009), .D(net_6478), .CK(net_15234) );
CLKBUF_X2 inst_14714 ( .A(net_14632), .Z(net_14633) );
DFF_X1 inst_8624 ( .Q(net_9782), .D(net_7202), .CK(net_13370) );
INV_X4 inst_5878 ( .A(net_7029), .ZN(net_626) );
CLKBUF_X2 inst_14383 ( .A(net_14214), .Z(net_14302) );
CLKBUF_X2 inst_11445 ( .A(net_11363), .Z(net_11364) );
INV_X4 inst_6385 ( .A(net_10301), .ZN(net_3681) );
CLKBUF_X2 inst_15006 ( .A(net_13163), .Z(net_14925) );
DFF_X2 inst_7615 ( .Q(net_9212), .D(net_6964), .CK(net_11840) );
DFF_X2 inst_8277 ( .Q(net_10496), .D(net_4885), .CK(net_15203) );
INV_X4 inst_4953 ( .A(net_4714), .ZN(net_3917) );
CLKBUF_X2 inst_12404 ( .A(net_12322), .Z(net_12323) );
AOI22_X2 inst_9589 ( .B1(net_9987), .A2(net_5173), .ZN(net_3571), .B2(net_2541), .A1(net_220) );
INV_X2 inst_7164 ( .A(net_7021), .ZN(net_573) );
CLKBUF_X2 inst_13356 ( .A(net_13274), .Z(net_13275) );
NAND2_X2 inst_3659 ( .A2(net_10380), .A1(net_10379), .ZN(net_7285) );
DFF_X2 inst_7465 ( .Q(net_9522), .D(net_8099), .CK(net_14976) );
INV_X4 inst_6573 ( .ZN(net_6347), .A(net_163) );
NAND2_X2 inst_3604 ( .ZN(net_7262), .A2(net_6851), .A1(net_6602) );
CLKBUF_X2 inst_13067 ( .A(net_12985), .Z(net_12986) );
CLKBUF_X2 inst_12347 ( .A(net_11046), .Z(net_12266) );
INV_X4 inst_6487 ( .A(net_9178), .ZN(net_585) );
OAI22_X2 inst_1109 ( .A1(net_7219), .ZN(net_6150), .B2(net_5875), .A2(net_5300), .B1(net_3944) );
CLKBUF_X2 inst_12054 ( .A(net_10689), .Z(net_11973) );
AND2_X2 inst_10559 ( .ZN(net_3132), .A1(net_3131), .A2(net_2835) );
CLKBUF_X2 inst_13879 ( .A(net_13797), .Z(net_13798) );
NAND2_X2 inst_4415 ( .A2(net_10329), .A1(net_10328), .ZN(net_2410) );
NAND2_X2 inst_4209 ( .ZN(net_2983), .A1(net_2565), .A2(net_1763) );
NAND4_X2 inst_3037 ( .ZN(net_8619), .A1(net_8501), .A2(net_8500), .A3(net_8499), .A4(net_8498) );
AOI211_X2 inst_10266 ( .ZN(net_7707), .A(net_7704), .C2(net_7600), .C1(net_4762), .B(x3390) );
INV_X4 inst_6635 ( .ZN(net_9055), .A(net_3376) );
AOI211_X2 inst_10275 ( .ZN(net_7518), .B(net_7169), .C2(net_5004), .A(net_3208), .C1(net_2848) );
CLKBUF_X2 inst_11522 ( .A(net_11440), .Z(net_11441) );
DFF_X1 inst_8561 ( .Q(net_9785), .D(net_7228), .CK(net_13380) );
CLKBUF_X2 inst_14857 ( .A(net_11312), .Z(net_14776) );
DFF_X2 inst_7956 ( .QN(net_10218), .D(net_5633), .CK(net_13254) );
OAI22_X2 inst_1314 ( .ZN(net_2213), .A1(net_2212), .A2(net_2211), .B1(net_2210), .B2(net_1662) );
CLKBUF_X2 inst_12072 ( .A(net_11909), .Z(net_11991) );
INV_X4 inst_5828 ( .ZN(net_5464), .A(net_671) );
NAND2_X2 inst_4260 ( .A1(net_10263), .A2(net_9833), .ZN(net_2827) );
AOI21_X2 inst_10218 ( .ZN(net_2293), .B2(net_2292), .B1(net_1453), .A(net_1443) );
INV_X4 inst_5533 ( .ZN(net_4331), .A(net_1177) );
OAI22_X2 inst_1156 ( .A1(net_7186), .A2(net_5139), .B2(net_5138), .ZN(net_5117), .B1(net_3589) );
DFF_X2 inst_8072 ( .QN(net_9172), .D(net_5281), .CK(net_11310) );
NAND2_X4 inst_3378 ( .A2(net_9060), .A1(net_8954), .ZN(net_1973) );
CLKBUF_X2 inst_11466 ( .A(net_11384), .Z(net_11385) );
INV_X4 inst_5993 ( .A(net_10259), .ZN(net_615) );
CLKBUF_X2 inst_12512 ( .A(net_12430), .Z(net_12431) );
NAND2_X2 inst_3484 ( .ZN(net_8394), .A1(net_8372), .A2(net_8254) );
CLKBUF_X2 inst_13868 ( .A(net_13786), .Z(net_13787) );
CLKBUF_X2 inst_13676 ( .A(net_12382), .Z(net_13595) );
OR2_X2 inst_942 ( .A2(net_10220), .A1(net_10219), .ZN(net_1745) );
CLKBUF_X2 inst_14259 ( .A(net_14177), .Z(net_14178) );
DFF_X2 inst_7755 ( .Q(net_10195), .D(net_6453), .CK(net_15131) );
CLKBUF_X2 inst_12077 ( .A(net_10686), .Z(net_11996) );
DFF_X2 inst_8269 ( .Q(net_10394), .D(net_4813), .CK(net_14509) );
OAI22_X2 inst_1295 ( .B1(net_5094), .A2(net_4274), .B2(net_3588), .ZN(net_3577), .A1(net_3576) );
OAI21_X2 inst_1880 ( .ZN(net_5225), .B1(net_5214), .B2(net_5213), .A(net_1546) );
CLKBUF_X2 inst_13174 ( .A(net_13092), .Z(net_13093) );
DFF_X2 inst_7457 ( .QN(net_9641), .D(net_8188), .CK(net_15380) );
XNOR2_X2 inst_262 ( .ZN(net_3989), .B(net_3988), .A(net_3677) );
INV_X4 inst_6603 ( .A(net_10030), .ZN(net_921) );
NAND2_X2 inst_3630 ( .A2(net_7161), .ZN(net_7016), .A1(net_7015) );
AND4_X4 inst_10333 ( .ZN(net_2900), .A4(net_2109), .A3(net_1261), .A1(net_1072), .A2(net_877) );
HA_X1 inst_7338 ( .S(net_6177), .CO(net_6176), .B(net_5242), .A(net_3400) );
INV_X4 inst_4675 ( .A(net_7660), .ZN(net_5251) );
HA_X1 inst_7353 ( .A(net_9180), .CO(net_4124), .S(net_3518), .B(net_2737) );
INV_X8 inst_4501 ( .ZN(net_6120), .A(net_5298) );
INV_X2 inst_7144 ( .A(net_3194), .ZN(net_1442) );
NAND2_X2 inst_4252 ( .A2(net_9344), .ZN(net_1688), .A1(net_747) );
OAI22_X2 inst_1035 ( .A2(net_9071), .B1(net_8919), .A1(net_8915), .ZN(net_7950), .B2(net_1977) );
DFF_X2 inst_7942 ( .QN(net_10225), .D(net_5477), .CK(net_14474) );
CLKBUF_X2 inst_11758 ( .A(net_11676), .Z(net_11677) );
NAND2_X2 inst_3637 ( .A2(net_7175), .ZN(net_6978), .A1(net_4714) );
CLKBUF_X2 inst_11490 ( .A(net_11408), .Z(net_11409) );
INV_X4 inst_6356 ( .A(net_10364), .ZN(net_589) );
OAI21_X2 inst_1883 ( .ZN(net_5010), .B1(net_5009), .A(net_4711), .B2(net_4599) );
INV_X2 inst_7240 ( .A(net_9408), .ZN(net_8225) );
CLKBUF_X2 inst_12863 ( .A(net_12781), .Z(net_12782) );
AOI22_X2 inst_9580 ( .A1(net_10063), .A2(net_5320), .B2(net_5174), .ZN(net_3583), .B1(net_720) );
DFF_X2 inst_8258 ( .Q(net_10284), .D(net_4823), .CK(net_14524) );
NAND2_X2 inst_3621 ( .ZN(net_7105), .A2(net_6864), .A1(net_6596) );
INV_X4 inst_5451 ( .A(net_1681), .ZN(net_1081) );
INV_X4 inst_6393 ( .A(net_10103), .ZN(net_5827) );
OR2_X2 inst_864 ( .A1(net_8801), .ZN(net_8648), .A2(net_8647) );
XNOR2_X2 inst_418 ( .B(net_9358), .ZN(net_1407), .A(net_1406) );
XNOR2_X2 inst_86 ( .ZN(net_8617), .A(net_8579), .B(net_8264) );
OAI33_X1 inst_949 ( .B1(net_7530), .ZN(net_7524), .A1(net_7522), .B3(net_7521), .A3(net_6624), .A2(net_6245), .B2(net_967) );
NAND3_X2 inst_3283 ( .ZN(net_7671), .A3(net_3593), .A2(net_3448), .A1(net_664) );
NAND2_X2 inst_3961 ( .ZN(net_3611), .A2(net_3456), .A1(net_3454) );
CLKBUF_X2 inst_12580 ( .A(net_12498), .Z(net_12499) );
CLKBUF_X2 inst_15651 ( .A(net_15569), .Z(net_15570) );
CLKBUF_X2 inst_13294 ( .A(net_11765), .Z(net_13213) );
AOI22_X2 inst_9526 ( .B1(net_10000), .A2(net_6443), .ZN(net_3795), .B2(net_2468), .A1(net_1827) );
NAND2_X2 inst_3730 ( .ZN(net_5695), .A2(net_5694), .A1(net_1504) );
AND4_X2 inst_10342 ( .A1(net_5168), .A2(net_5167), .A4(net_5166), .ZN(net_5163), .A3(net_2850) );
NAND2_X2 inst_3598 ( .ZN(net_7268), .A2(net_6879), .A1(net_6607) );
CLKBUF_X2 inst_11851 ( .A(net_11769), .Z(net_11770) );
INV_X4 inst_5871 ( .ZN(net_4997), .A(net_637) );
AOI21_X2 inst_10016 ( .A(net_8190), .ZN(net_8158), .B1(net_7895), .B2(net_7375) );
CLKBUF_X2 inst_12140 ( .A(net_12058), .Z(net_12059) );
OAI21_X2 inst_1826 ( .B1(net_7785), .ZN(net_6567), .A(net_5923), .B2(net_5893) );
OAI211_X2 inst_2109 ( .C2(net_6774), .ZN(net_6739), .A(net_6365), .B(net_6138), .C1(net_536) );
INV_X4 inst_5395 ( .ZN(net_1176), .A(net_1175) );
INV_X4 inst_6192 ( .ZN(net_7127), .A(x5498) );
OAI21_X2 inst_2020 ( .ZN(net_8861), .A(net_2422), .B2(net_2060), .B1(net_1646) );
NAND2_X2 inst_4361 ( .A2(net_10354), .ZN(net_2019), .A1(net_441) );
CLKBUF_X2 inst_13957 ( .A(net_11962), .Z(net_13876) );
OAI22_X2 inst_1177 ( .A1(net_7224), .A2(net_5151), .B2(net_5150), .ZN(net_5082), .B1(net_3536) );
CLKBUF_X2 inst_13721 ( .A(net_13005), .Z(net_13640) );
NOR2_X2 inst_2820 ( .A2(net_3065), .ZN(net_2596), .A1(net_2595) );
NOR2_X2 inst_2548 ( .A2(net_9636), .A1(net_8978), .ZN(net_8090) );
CLKBUF_X2 inst_14417 ( .A(net_14335), .Z(net_14336) );
NOR3_X2 inst_2404 ( .A1(net_7345), .A3(net_7343), .ZN(net_7149), .A2(net_457) );
CLKBUF_X2 inst_14075 ( .A(net_11225), .Z(net_13994) );
CLKBUF_X2 inst_11494 ( .A(net_10676), .Z(net_11413) );
DFF_X2 inst_7994 ( .QN(net_10125), .D(net_5522), .CK(net_12367) );
INV_X4 inst_5127 ( .A(net_3742), .ZN(net_1942) );
CLKBUF_X2 inst_15539 ( .A(net_15457), .Z(net_15458) );
DFF_X2 inst_8022 ( .QN(net_10220), .D(net_5471), .CK(net_14460) );
OAI221_X2 inst_1578 ( .B1(net_10207), .B2(net_7295), .C2(net_7293), .ZN(net_7137), .C1(net_7136), .A(net_6938) );
CLKBUF_X2 inst_12587 ( .A(net_11245), .Z(net_12506) );
AOI22_X2 inst_9051 ( .B1(net_9671), .A1(net_6684), .B2(net_6683), .ZN(net_6671), .A2(net_240) );
DFF_X2 inst_7849 ( .Q(net_10294), .D(net_6214), .CK(net_14540) );
OAI221_X2 inst_1666 ( .C1(net_7216), .B2(net_5591), .ZN(net_5503), .C2(net_4902), .A(net_3731), .B1(net_870) );
DFF_X2 inst_7662 ( .D(net_6690), .QN(net_172), .CK(net_12738) );
OR2_X4 inst_735 ( .ZN(net_9063), .A1(net_7089), .A2(net_4455) );
OAI221_X2 inst_1529 ( .B1(net_10201), .B2(net_7295), .C2(net_7293), .ZN(net_7244), .C1(net_7243), .A(net_6829) );
AOI22_X2 inst_9053 ( .B1(net_9675), .A1(net_6684), .B2(net_6683), .ZN(net_6642), .A2(net_244) );
CLKBUF_X2 inst_12445 ( .A(net_12363), .Z(net_12364) );
INV_X4 inst_4612 ( .ZN(net_7340), .A(net_7158) );
AND2_X4 inst_10426 ( .A1(net_9216), .ZN(net_3656), .A2(net_3655) );
DFF_X2 inst_7890 ( .QN(net_10096), .D(net_6025), .CK(net_13262) );
OAI221_X2 inst_1653 ( .C1(net_7209), .ZN(net_5522), .C2(net_5520), .B2(net_4547), .A(net_3507), .B1(net_1886) );
AOI22_X2 inst_9598 ( .A1(net_10072), .B1(net_10023), .A2(net_5319), .B2(net_5174), .ZN(net_3494) );
CLKBUF_X2 inst_11398 ( .A(net_11316), .Z(net_11317) );
CLKBUF_X2 inst_15676 ( .A(net_15594), .Z(net_15595) );
CLKBUF_X2 inst_13376 ( .A(net_13294), .Z(net_13295) );
DFF_X1 inst_8820 ( .Q(net_10060), .D(net_3259), .CK(net_11106) );
INV_X2 inst_7220 ( .A(net_9410), .ZN(net_8195) );
CLKBUF_X2 inst_11627 ( .A(net_11494), .Z(net_11546) );
NOR2_X2 inst_2984 ( .A1(net_10326), .ZN(net_2646), .A2(net_589) );
XNOR2_X2 inst_175 ( .ZN(net_5399), .A(net_4944), .B(net_2338) );
NAND3_X2 inst_3258 ( .ZN(net_5160), .A1(net_4611), .A3(net_4460), .A2(net_3385) );
CLKBUF_X2 inst_13002 ( .A(net_12920), .Z(net_12921) );
CLKBUF_X2 inst_11989 ( .A(net_11907), .Z(net_11908) );
CLKBUF_X2 inst_12150 ( .A(net_12068), .Z(net_12069) );
AND2_X2 inst_10491 ( .A1(net_9535), .A2(net_9503), .ZN(net_7329) );
INV_X4 inst_5010 ( .ZN(net_2573), .A(net_2163) );
CLKBUF_X2 inst_15764 ( .A(net_15682), .Z(net_15683) );
CLKBUF_X2 inst_10895 ( .A(net_10798), .Z(net_10814) );
OAI21_X2 inst_1737 ( .B2(net_9049), .ZN(net_8988), .B1(net_8711), .A(net_8396) );
DFF_X1 inst_8594 ( .Q(net_9688), .D(net_7259), .CK(net_15741) );
OAI21_X2 inst_1805 ( .ZN(net_7385), .B2(net_7052), .A(net_2352), .B1(net_1622) );
NOR2_X2 inst_2995 ( .A1(net_10352), .ZN(net_1103), .A2(net_902) );
NAND2_X2 inst_3563 ( .A2(net_7748), .ZN(net_7687), .A1(net_326) );
AOI222_X2 inst_9675 ( .ZN(net_3113), .A1(net_3112), .C2(net_3111), .B2(net_3111), .A2(net_2250), .C1(net_1957), .B1(net_611) );
INV_X2 inst_7081 ( .ZN(net_1179), .A(net_1178) );
INV_X4 inst_5513 ( .A(net_10474), .ZN(net_3710) );
DFF_X2 inst_8231 ( .Q(net_10501), .D(net_4880), .CK(net_15223) );
INV_X4 inst_4541 ( .ZN(net_8878), .A(net_8700) );
NOR2_X2 inst_2752 ( .ZN(net_4122), .A2(net_3647), .A1(net_2041) );
AOI21_X2 inst_10095 ( .B2(net_10280), .A(net_6678), .ZN(net_5536), .B1(net_627) );
CLKBUF_X2 inst_14073 ( .A(net_13991), .Z(net_13992) );
OAI22_X2 inst_1149 ( .A1(net_7201), .A2(net_5134), .B2(net_5133), .ZN(net_5124), .B1(net_784) );
AOI21_X2 inst_10146 ( .ZN(net_4203), .A(net_4202), .B1(net_3712), .B2(net_3711) );
CLKBUF_X2 inst_14354 ( .A(net_11518), .Z(net_14273) );
OAI22_X2 inst_1281 ( .A2(net_10062), .ZN(net_4276), .A1(net_4275), .B2(net_4274), .B1(net_4247) );
OAI221_X2 inst_1509 ( .C1(net_10414), .B2(net_9063), .C2(net_9056), .ZN(net_7351), .B1(net_7241), .A(net_6988) );
INV_X4 inst_5640 ( .A(net_852), .ZN(net_846) );
NAND4_X2 inst_3088 ( .ZN(net_4488), .A2(net_4053), .A1(net_3802), .A3(net_3787), .A4(net_3735) );
AND2_X4 inst_10386 ( .ZN(net_8444), .A2(net_8443), .A1(net_5388) );
AOI22_X2 inst_9000 ( .B1(net_9453), .A1(net_9445), .A2(net_8952), .ZN(net_8498), .B2(net_8479) );
CLKBUF_X2 inst_11475 ( .A(net_10787), .Z(net_11394) );
AOI222_X1 inst_9696 ( .B1(net_9507), .A2(net_8286), .B2(net_8285), .C2(net_8284), .ZN(net_8282), .C1(net_8217), .A1(x1598) );
NAND2_X2 inst_3782 ( .A2(net_9088), .A1(net_9078), .ZN(net_5266) );
CLKBUF_X2 inst_15754 ( .A(net_15672), .Z(net_15673) );
INV_X4 inst_4719 ( .A(net_9151), .ZN(net_4971) );
CLKBUF_X2 inst_15026 ( .A(net_14944), .Z(net_14945) );
DFF_X2 inst_7486 ( .D(net_8063), .Q(net_218), .CK(net_12527) );
CLKBUF_X2 inst_15101 ( .A(net_15019), .Z(net_15020) );
CLKBUF_X2 inst_15466 ( .A(net_14041), .Z(net_15385) );
INV_X4 inst_6630 ( .A(net_8986), .ZN(net_8985) );
CLKBUF_X2 inst_15378 ( .A(net_10700), .Z(net_15297) );
INV_X4 inst_6003 ( .A(net_9370), .ZN(net_7848) );
NAND2_X2 inst_4353 ( .A2(net_10222), .ZN(net_2455), .A1(net_1211) );
AOI22_X2 inst_9285 ( .B1(net_9897), .A1(net_5759), .B2(net_5758), .ZN(net_5717), .A2(net_236) );
NAND2_X2 inst_3934 ( .ZN(net_3700), .A1(net_3699), .A2(net_3698) );
AOI222_X1 inst_9716 ( .B2(net_7175), .ZN(net_7165), .C1(net_4723), .B1(net_3591), .A2(net_3076), .A1(net_2887), .C2(net_2616) );
CLKBUF_X2 inst_13302 ( .A(net_13220), .Z(net_13221) );
CLKBUF_X2 inst_12475 ( .A(net_10896), .Z(net_12394) );
DFF_X2 inst_8054 ( .QN(net_9553), .D(net_9259), .CK(net_13750) );
INV_X4 inst_5809 ( .ZN(net_3209), .A(net_683) );
OAI33_X1 inst_948 ( .ZN(net_7563), .B2(net_7562), .B1(net_7560), .A3(net_4631), .A2(net_4318), .A1(net_4176), .B3(net_991) );
OAI22_X2 inst_1140 ( .A1(net_7234), .ZN(net_5135), .A2(net_5134), .B2(net_5133), .B1(net_344) );
CLKBUF_X2 inst_15637 ( .A(net_15555), .Z(net_15556) );
AOI22_X2 inst_9251 ( .B2(net_8041), .A2(net_6141), .ZN(net_6059), .B1(net_1942), .A1(net_1928) );
INV_X4 inst_6140 ( .A(net_9726), .ZN(net_482) );
OAI21_X2 inst_1800 ( .ZN(net_7509), .B1(net_7505), .A(net_7336), .B2(net_7114) );
CLKBUF_X2 inst_14795 ( .A(net_12017), .Z(net_14714) );
INV_X4 inst_4773 ( .ZN(net_4308), .A(net_4119) );
DFF_X1 inst_8463 ( .Q(net_9592), .D(net_7966), .CK(net_11534) );
CLKBUF_X2 inst_11087 ( .A(net_11005), .Z(net_11006) );
INV_X4 inst_6644 ( .A(net_9094), .ZN(net_9093) );
XNOR2_X2 inst_448 ( .A(net_9560), .ZN(net_8849), .B(net_8719) );
INV_X4 inst_5966 ( .A(net_10153), .ZN(net_793) );
CLKBUF_X2 inst_13493 ( .A(net_13411), .Z(net_13412) );
CLKBUF_X2 inst_11407 ( .A(net_11325), .Z(net_11326) );
CLKBUF_X2 inst_11275 ( .A(net_11109), .Z(net_11194) );
INV_X4 inst_5680 ( .A(net_10324), .ZN(net_804) );
AOI211_X2 inst_10253 ( .A(net_8190), .ZN(net_8189), .C2(net_7888), .C1(net_5169), .B(net_3298) );
DFF_X2 inst_8039 ( .Q(net_9560), .D(net_5417), .CK(net_12620) );
INV_X4 inst_6056 ( .ZN(net_6423), .A(net_130) );
INV_X4 inst_4921 ( .ZN(net_2925), .A(net_2220) );
CLKBUF_X2 inst_15579 ( .A(net_15497), .Z(net_15498) );
CLKBUF_X2 inst_14367 ( .A(net_14285), .Z(net_14286) );
CLKBUF_X2 inst_11647 ( .A(net_11565), .Z(net_11566) );
CLKBUF_X2 inst_14671 ( .A(net_10806), .Z(net_14590) );
AOI221_X2 inst_9966 ( .C1(net_9972), .B1(net_9675), .B2(net_5966), .ZN(net_4765), .A(net_4347), .C2(net_2541) );
AOI22_X2 inst_9374 ( .B1(net_10008), .A2(net_5743), .B2(net_5742), .ZN(net_5531), .A1(net_248) );
INV_X4 inst_5444 ( .ZN(net_1589), .A(net_1551) );
INV_X4 inst_6030 ( .A(net_9168), .ZN(net_519) );
NAND2_X2 inst_4380 ( .ZN(net_7884), .A2(net_833), .A1(net_685) );
OAI21_X2 inst_2002 ( .ZN(net_2806), .A(net_2149), .B1(net_2148), .B2(net_1679) );
CLKBUF_X2 inst_10862 ( .A(net_10780), .Z(net_10781) );
AOI21_X2 inst_10053 ( .B2(net_7175), .ZN(net_7151), .A(net_4348), .B1(net_2887) );
CLKBUF_X2 inst_13017 ( .A(net_12935), .Z(net_12936) );
AND2_X4 inst_10471 ( .A2(net_9639), .A1(net_9638), .ZN(net_1023) );
DFF_X1 inst_8430 ( .D(net_8666), .CK(net_11928), .Q(x715) );
DFF_X2 inst_8212 ( .Q(net_10086), .D(net_4849), .CK(net_10752) );
SDFF_X2 inst_608 ( .QN(net_10512), .D(net_4413), .SE(net_3688), .SI(net_659), .CK(net_11140) );
OAI222_X2 inst_1343 ( .B1(net_7732), .A2(net_7731), .C2(net_7730), .ZN(net_7579), .B2(net_7417), .A1(net_6171), .C1(net_1905) );
AOI22_X2 inst_9068 ( .B1(net_9688), .A2(net_6684), .B2(net_6683), .ZN(net_6598), .A1(net_257) );
DFF_X2 inst_8050 ( .QN(net_10313), .D(net_5570), .CK(net_13312) );
OR2_X4 inst_834 ( .ZN(net_1727), .A2(x6351), .A1(x6327) );
CLKBUF_X2 inst_11183 ( .A(net_10946), .Z(net_11102) );
DFF_X1 inst_8729 ( .Q(net_9142), .D(net_6156), .CK(net_11004) );
DFF_X2 inst_7536 ( .QN(net_8824), .D(net_7786), .CK(net_13125) );
NOR2_X2 inst_2920 ( .A2(net_4566), .ZN(net_1622), .A1(net_1352) );
NAND2_X2 inst_4054 ( .ZN(net_3242), .A2(net_2805), .A1(net_2054) );
DFF_X2 inst_7813 ( .Q(net_10016), .D(net_6469), .CK(net_15696) );
INV_X2 inst_6713 ( .A(net_9599), .ZN(net_7994) );
OAI33_X1 inst_966 ( .ZN(net_3216), .B1(net_3215), .A3(net_3215), .B2(net_3214), .A1(net_1721), .B3(net_1344), .A2(net_692) );
CLKBUF_X2 inst_14951 ( .A(net_14869), .Z(net_14870) );
CLKBUF_X2 inst_11833 ( .A(net_11111), .Z(net_11752) );
INV_X2 inst_7189 ( .A(net_9405), .ZN(net_8228) );
OAI22_X2 inst_1246 ( .B1(net_7203), .ZN(net_4845), .A2(net_4842), .B2(net_4841), .A1(net_402) );
NOR2_X2 inst_2961 ( .ZN(net_1798), .A1(net_1387), .A2(net_668) );
NAND3_X2 inst_3185 ( .A3(net_9661), .A2(net_8511), .ZN(net_7926), .A1(net_7832) );
INV_X4 inst_4679 ( .ZN(net_5003), .A(net_4757) );
NOR2_X2 inst_2506 ( .ZN(net_8681), .A1(net_8428), .A2(net_8426) );
CLKBUF_X2 inst_13214 ( .A(net_13132), .Z(net_13133) );
CLKBUF_X2 inst_11699 ( .A(net_11617), .Z(net_11618) );
CLKBUF_X2 inst_11269 ( .A(net_11187), .Z(net_11188) );
INV_X4 inst_5836 ( .ZN(net_5786), .A(net_5392) );
CLKBUF_X2 inst_13163 ( .A(net_13081), .Z(net_13082) );
INV_X4 inst_5976 ( .A(net_10477), .ZN(net_542) );
INV_X4 inst_5647 ( .ZN(net_3173), .A(net_1071) );
AND2_X2 inst_10623 ( .A2(net_9220), .A1(net_9219), .ZN(net_1238) );
INV_X4 inst_5245 ( .ZN(net_2184), .A(net_1464) );
INV_X4 inst_5580 ( .A(net_1020), .ZN(net_890) );
INV_X4 inst_5575 ( .A(net_945), .ZN(net_903) );
INV_X4 inst_4557 ( .ZN(net_8496), .A(net_8431) );
CLKBUF_X2 inst_12180 ( .A(net_12098), .Z(net_12099) );
NAND2_X2 inst_3607 ( .ZN(net_7259), .A2(net_6853), .A1(net_6598) );
DFF_X1 inst_8568 ( .Q(net_9775), .D(net_7298), .CK(net_14852) );
OAI211_X2 inst_2029 ( .C2(net_10055), .ZN(net_8162), .B(net_8079), .A(net_8040), .C1(net_6774) );
CLKBUF_X2 inst_10632 ( .A(net_10550), .Z(net_10551) );
CLKBUF_X2 inst_12812 ( .A(net_12730), .Z(net_12731) );
DFF_X1 inst_8583 ( .Q(net_9769), .D(net_7247), .CK(net_15625) );
AND2_X2 inst_10498 ( .ZN(net_7027), .A1(net_6588), .A2(net_6169) );
DFF_X1 inst_8779 ( .QN(net_10273), .D(net_4684), .CK(net_11767) );
INV_X4 inst_4936 ( .ZN(net_2851), .A(net_2581) );
CLKBUF_X2 inst_13324 ( .A(net_10956), .Z(net_13243) );
CLKBUF_X2 inst_15037 ( .A(net_14955), .Z(net_14956) );
NAND4_X2 inst_3160 ( .ZN(net_1735), .A2(net_874), .A3(net_110), .A4(net_109), .A1(net_105) );
CLKBUF_X2 inst_14022 ( .A(net_13940), .Z(net_13941) );
CLKBUF_X2 inst_14825 ( .A(net_12695), .Z(net_14744) );
NOR2_X2 inst_2861 ( .ZN(net_2069), .A1(net_2068), .A2(net_1436) );
XNOR2_X2 inst_66 ( .ZN(net_8722), .A(net_8697), .B(net_8427) );
INV_X4 inst_4814 ( .ZN(net_4512), .A(net_4319) );
CLKBUF_X2 inst_11139 ( .A(net_11057), .Z(net_11058) );
CLKBUF_X2 inst_11012 ( .A(net_10574), .Z(net_10931) );
AND2_X2 inst_10604 ( .A1(net_3112), .ZN(net_2055), .A2(net_2054) );
DFF_X2 inst_7920 ( .QN(net_10473), .D(net_5799), .CK(net_11386) );
DFF_X1 inst_8807 ( .QN(net_10482), .D(net_3962), .CK(net_11478) );
CLKBUF_X2 inst_12297 ( .A(net_12215), .Z(net_12216) );
XNOR2_X2 inst_273 ( .ZN(net_3952), .A(net_3241), .B(net_2892) );
CLKBUF_X2 inst_13443 ( .A(net_12632), .Z(net_13362) );
CLKBUF_X2 inst_15365 ( .A(net_15283), .Z(net_15284) );
OAI21_X2 inst_1965 ( .ZN(net_3358), .A(net_3357), .B2(net_3356), .B1(net_2689) );
NAND2_X2 inst_3915 ( .A2(net_9055), .ZN(net_7969), .A1(net_1843) );
INV_X4 inst_5419 ( .ZN(net_2292), .A(net_1145) );
XNOR2_X2 inst_366 ( .ZN(net_2522), .B(net_2521), .A(net_2167) );
NOR3_X2 inst_2418 ( .ZN(net_5334), .A3(net_5158), .A2(net_4470), .A1(net_3984) );
INV_X4 inst_6162 ( .A(net_10457), .ZN(net_760) );
DFF_X2 inst_8144 ( .Q(net_9937), .D(net_5111), .CK(net_14281) );
INV_X2 inst_7019 ( .A(net_2757), .ZN(net_2634) );
INV_X4 inst_5743 ( .ZN(net_2272), .A(net_743) );
INV_X4 inst_5422 ( .ZN(net_5061), .A(net_1134) );
CLKBUF_X2 inst_12542 ( .A(net_12460), .Z(net_12461) );
AOI22_X2 inst_9565 ( .B1(net_9970), .A1(net_9737), .A2(net_6442), .ZN(net_3754), .B2(net_2541) );
AOI22_X2 inst_9397 ( .B1(net_9709), .A1(net_5755), .B2(net_5754), .ZN(net_5400), .A2(net_246) );
DFF_X2 inst_7964 ( .QN(net_10209), .D(net_5623), .CK(net_15587) );
CLKBUF_X2 inst_15785 ( .A(net_15703), .Z(net_15704) );
INV_X2 inst_7313 ( .A(net_9094), .ZN(net_9092) );
NAND3_X2 inst_3285 ( .ZN(net_4092), .A3(net_3891), .A2(net_3448), .A1(net_1255) );
INV_X2 inst_6948 ( .A(net_2095), .ZN(net_1899) );
INV_X4 inst_6492 ( .ZN(net_7294), .A(x5143) );
INV_X4 inst_5896 ( .ZN(net_922), .A(net_605) );
INV_X4 inst_4746 ( .A(net_10293), .ZN(net_5908) );
DFF_X2 inst_7950 ( .QN(net_10210), .D(net_5643), .CK(net_11752) );
CLKBUF_X2 inst_14091 ( .A(net_13654), .Z(net_14010) );
CLKBUF_X2 inst_14934 ( .A(net_14212), .Z(net_14853) );
OAI22_X2 inst_1025 ( .A2(net_8036), .B2(net_8018), .ZN(net_8005), .A1(net_4164), .B1(net_346) );
OR3_X2 inst_707 ( .ZN(net_7882), .A1(net_7814), .A3(net_7147), .A2(net_4150) );
INV_X4 inst_4655 ( .A(net_9253), .ZN(net_8326) );
CLKBUF_X2 inst_11931 ( .A(net_11849), .Z(net_11850) );
CLKBUF_X2 inst_11790 ( .A(net_11708), .Z(net_11709) );
DFF_X2 inst_7566 ( .QN(net_9385), .D(net_7639), .CK(net_13029) );
NAND2_X2 inst_3670 ( .A1(net_8964), .ZN(net_7572), .A2(net_6242) );
CLKBUF_X2 inst_11568 ( .A(net_10922), .Z(net_11487) );
MUX2_X1 inst_4460 ( .S(net_6041), .A(net_286), .B(x5790), .Z(x257) );
DFF_X2 inst_8336 ( .QN(net_9562), .D(net_3250), .CK(net_15193) );
DFF_X2 inst_7570 ( .QN(net_10372), .D(net_7579), .CK(net_12227) );
INV_X4 inst_5635 ( .ZN(net_1195), .A(net_1146) );
CLKBUF_X2 inst_12559 ( .A(net_12477), .Z(net_12478) );
DFF_X2 inst_7834 ( .Q(net_9811), .D(net_6522), .CK(net_12043) );
CLKBUF_X2 inst_11681 ( .A(net_11599), .Z(net_11600) );
INV_X2 inst_7002 ( .ZN(net_1623), .A(net_1622) );
NOR2_X2 inst_2804 ( .ZN(net_3234), .A2(net_2801), .A1(net_2645) );
INV_X4 inst_5542 ( .ZN(net_1994), .A(net_941) );
DFF_X1 inst_8654 ( .Q(net_9862), .D(net_7189), .CK(net_15448) );
INV_X4 inst_5131 ( .A(net_2630), .ZN(net_1596) );
AOI21_X2 inst_10080 ( .ZN(net_5683), .B2(net_5682), .A(net_5163), .B1(net_2850) );
CLKBUF_X2 inst_15094 ( .A(net_13645), .Z(net_15013) );
CLKBUF_X2 inst_13710 ( .A(net_13628), .Z(net_13629) );
CLKBUF_X2 inst_13654 ( .A(net_13572), .Z(net_13573) );
INV_X2 inst_7269 ( .A(net_8927), .ZN(net_8926) );
NOR2_X2 inst_2576 ( .ZN(net_7273), .A2(net_6850), .A1(net_3749) );
NOR2_X2 inst_2631 ( .ZN(net_5942), .A2(net_5927), .A1(net_2840) );
OR2_X4 inst_772 ( .A2(net_3344), .A1(net_3161), .ZN(net_3141) );
NAND2_X2 inst_3810 ( .A1(net_10079), .A2(net_4534), .ZN(net_4528) );
DFF_X1 inst_8453 ( .Q(net_9523), .D(net_8097), .CK(net_15039) );
INV_X2 inst_6738 ( .ZN(net_7377), .A(net_7376) );
CLKBUF_X2 inst_13261 ( .A(net_13179), .Z(net_13180) );
NAND2_X2 inst_3682 ( .A2(net_9515), .A1(net_9514), .ZN(net_7505) );
INV_X4 inst_4940 ( .A(net_7895), .ZN(net_2579) );
INV_X8 inst_4523 ( .ZN(net_8951), .A(net_8383) );
INV_X2 inst_7073 ( .ZN(net_3538), .A(net_1228) );
INV_X4 inst_4583 ( .ZN(net_8067), .A(net_8025) );
NOR2_X2 inst_2636 ( .A2(net_9269), .A1(net_6582), .ZN(net_5891) );
CLKBUF_X2 inst_13282 ( .A(net_13200), .Z(net_13201) );
INV_X4 inst_6198 ( .A(net_9520), .ZN(net_576) );
INV_X2 inst_7186 ( .A(net_10466), .ZN(net_518) );
CLKBUF_X2 inst_15141 ( .A(net_10792), .Z(net_15060) );
AND2_X2 inst_10525 ( .ZN(net_4390), .A2(net_3999), .A1(net_204) );
DFF_X2 inst_7579 ( .QN(net_9386), .D(net_7558), .CK(net_13024) );
CLKBUF_X2 inst_14491 ( .A(net_14409), .Z(net_14410) );
CLKBUF_X2 inst_14396 ( .A(net_11797), .Z(net_14315) );
CLKBUF_X2 inst_11561 ( .A(net_10845), .Z(net_11480) );
INV_X4 inst_4870 ( .ZN(net_3503), .A(net_3285) );
CLKBUF_X2 inst_13618 ( .A(net_11683), .Z(net_13537) );
CLKBUF_X2 inst_12961 ( .A(net_11195), .Z(net_12880) );
XNOR2_X2 inst_445 ( .B(net_9303), .ZN(net_856), .A(net_226) );
INV_X4 inst_5454 ( .ZN(net_1070), .A(net_610) );
INV_X4 inst_5192 ( .ZN(net_4281), .A(net_2306) );
INV_X4 inst_6224 ( .A(net_10367), .ZN(net_3102) );
CLKBUF_X2 inst_11566 ( .A(net_11166), .Z(net_11485) );
CLKBUF_X2 inst_11400 ( .A(net_11318), .Z(net_11319) );
INV_X2 inst_6761 ( .ZN(net_6227), .A(net_6226) );
SDFF_X2 inst_606 ( .Q(net_10519), .D(net_10519), .SE(net_4560), .CK(net_11926), .SI(x5901) );
CLKBUF_X2 inst_12350 ( .A(net_12268), .Z(net_12269) );
NOR2_X2 inst_2942 ( .A1(net_10353), .ZN(net_1602), .A2(net_915) );
CLKBUF_X2 inst_15406 ( .A(net_15324), .Z(net_15325) );
AOI221_X2 inst_9929 ( .B2(net_5867), .A(net_5862), .ZN(net_5846), .C1(net_5845), .C2(net_4725), .B1(x4937) );
CLKBUF_X2 inst_13875 ( .A(net_12610), .Z(net_13794) );
AOI21_X2 inst_10138 ( .ZN(net_4248), .B1(net_4247), .A(net_3934), .B2(net_3459) );
INV_X4 inst_5654 ( .ZN(net_1297), .A(net_828) );
INV_X4 inst_5089 ( .ZN(net_1768), .A(net_1767) );
NAND2_X2 inst_3761 ( .ZN(net_5019), .A1(net_5015), .A2(net_4726) );
INV_X4 inst_5864 ( .ZN(net_1250), .A(net_640) );
OR2_X2 inst_853 ( .A1(net_9549), .ZN(net_8397), .A2(net_8145) );
AOI211_X2 inst_10287 ( .C1(net_9896), .ZN(net_4970), .C2(net_4969), .B(net_4383), .A(net_4377) );
DFF_X2 inst_8167 ( .QN(net_9829), .D(net_5048), .CK(net_14446) );
XNOR2_X2 inst_139 ( .ZN(net_7316), .A(net_6927), .B(net_2539) );
CLKBUF_X2 inst_13767 ( .A(net_13685), .Z(net_13686) );
SDFF_X2 inst_657 ( .SI(net_9471), .Q(net_9471), .SE(net_3073), .CK(net_14650), .D(x3194) );
CLKBUF_X2 inst_15813 ( .A(net_15731), .Z(net_15732) );
CLKBUF_X2 inst_10856 ( .A(net_10774), .Z(net_10775) );
INV_X4 inst_4550 ( .A(net_8619), .ZN(net_8596) );
CLKBUF_X2 inst_12803 ( .A(net_12721), .Z(net_12722) );
CLKBUF_X2 inst_12548 ( .A(net_12466), .Z(net_12467) );
OAI22_X2 inst_1316 ( .A2(net_2878), .ZN(net_2135), .B2(net_2134), .A1(net_2129), .B1(net_1346) );
OAI211_X2 inst_2098 ( .C2(net_6778), .ZN(net_6750), .A(net_6342), .B(net_6110), .C1(net_399) );
CLKBUF_X2 inst_12465 ( .A(net_12383), .Z(net_12384) );
DFF_X2 inst_8400 ( .QN(net_9195), .CK(net_11297), .D(x3534) );
NAND2_X2 inst_3551 ( .A1(net_10194), .ZN(net_7873), .A2(net_7867) );
INV_X4 inst_5528 ( .ZN(net_3272), .A(net_2412) );
OAI21_X2 inst_1921 ( .B2(net_10446), .A(net_10445), .ZN(net_4555), .B1(net_4554) );
CLKBUF_X2 inst_13890 ( .A(net_12187), .Z(net_13809) );
CLKBUF_X2 inst_12890 ( .A(net_12808), .Z(net_12809) );
INV_X4 inst_6521 ( .A(net_10064), .ZN(net_343) );
INV_X2 inst_6977 ( .ZN(net_1680), .A(net_1679) );
NAND2_X2 inst_4293 ( .ZN(net_3397), .A2(net_1250), .A1(net_473) );
CLKBUF_X2 inst_13996 ( .A(net_13914), .Z(net_13915) );
XNOR2_X2 inst_191 ( .ZN(net_5204), .A(net_4586), .B(net_2075) );
CLKBUF_X2 inst_14783 ( .A(net_14701), .Z(net_14702) );
CLKBUF_X2 inst_14285 ( .A(net_14203), .Z(net_14204) );
AND3_X4 inst_10357 ( .ZN(net_5766), .A2(net_4788), .A3(net_4630), .A1(net_4467) );
NOR2_X2 inst_2638 ( .A2(net_5927), .ZN(net_5816), .A1(net_4002) );
DFF_X1 inst_8676 ( .D(net_6744), .Q(net_109), .CK(net_15109) );
AOI22_X2 inst_9328 ( .B1(net_10020), .A2(net_5743), .B2(net_5742), .ZN(net_5647), .A1(net_260) );
CLKBUF_X2 inst_13485 ( .A(net_10981), .Z(net_13404) );
INV_X4 inst_4538 ( .ZN(net_9008), .A(net_8728) );
INV_X4 inst_5212 ( .A(net_6839), .ZN(net_2111) );
NAND3_X2 inst_3235 ( .A1(net_7142), .ZN(net_4722), .A2(net_4331), .A3(net_1643) );
CLKBUF_X2 inst_14019 ( .A(net_13937), .Z(net_13938) );
CLKBUF_X2 inst_13988 ( .A(net_13138), .Z(net_13907) );
CLKBUF_X2 inst_14680 ( .A(net_14598), .Z(net_14599) );
DFF_X1 inst_8672 ( .D(net_6737), .Q(net_104), .CK(net_12006) );
CLKBUF_X2 inst_12786 ( .A(net_12704), .Z(net_12705) );
AOI22_X2 inst_9421 ( .A1(net_10185), .A2(net_4656), .B2(net_4655), .ZN(net_4648), .B1(x4851) );
INV_X2 inst_6892 ( .ZN(net_2999), .A(net_2926) );
DFF_X1 inst_8711 ( .QN(net_10242), .D(net_6943), .CK(net_10925) );
NAND2_X2 inst_3879 ( .ZN(net_8889), .A2(net_4027), .A1(net_1978) );
INV_X4 inst_5269 ( .A(net_2655), .ZN(net_1358) );
INV_X4 inst_6544 ( .A(net_9297), .ZN(net_3884) );
CLKBUF_X2 inst_12201 ( .A(net_12119), .Z(net_12120) );
DFF_X2 inst_8125 ( .QN(net_10040), .D(net_5089), .CK(net_12889) );
OAI211_X2 inst_2184 ( .C1(net_7245), .C2(net_6542), .ZN(net_6525), .B(net_5621), .A(net_3527) );
CLKBUF_X2 inst_13296 ( .A(net_13214), .Z(net_13215) );
OR2_X2 inst_892 ( .A1(net_10058), .ZN(net_5893), .A2(net_5892) );
NOR2_X2 inst_2665 ( .A2(net_9091), .ZN(net_5809), .A1(net_641) );
OAI22_X2 inst_1132 ( .A1(net_7186), .A2(net_5151), .B2(net_5150), .ZN(net_5146), .B1(net_477) );
CLKBUF_X2 inst_14415 ( .A(net_14333), .Z(net_14334) );
NAND2_X2 inst_4100 ( .ZN(net_2441), .A1(net_2440), .A2(net_1712) );
OAI33_X1 inst_968 ( .ZN(net_3211), .B1(net_3210), .A3(net_3210), .B2(net_3209), .A1(net_1718), .B3(net_729), .A2(net_614) );
INV_X4 inst_4700 ( .ZN(net_4796), .A(net_4795) );
CLKBUF_X2 inst_13531 ( .A(net_13046), .Z(net_13450) );
MUX2_X1 inst_4441 ( .S(net_6041), .A(net_305), .B(x4449), .Z(x80) );
CLKBUF_X2 inst_15024 ( .A(net_12212), .Z(net_14943) );
INV_X2 inst_6987 ( .ZN(net_2364), .A(net_1656) );
OAI21_X2 inst_1803 ( .B2(net_7175), .ZN(net_7143), .B1(net_7142), .A(net_1643) );
NAND4_X2 inst_3153 ( .A2(net_9208), .A4(net_9202), .A3(net_9201), .ZN(net_1997), .A1(net_1098) );
NOR2_X2 inst_2814 ( .ZN(net_2642), .A1(net_2641), .A2(net_1945) );
INV_X4 inst_6076 ( .ZN(net_602), .A(net_196) );
AOI221_X2 inst_9819 ( .B1(net_9768), .B2(net_9097), .A(net_6940), .C1(net_6939), .ZN(net_6938), .C2(net_238) );
OR2_X2 inst_936 ( .ZN(net_2387), .A2(net_2386), .A1(x589) );
CLKBUF_X2 inst_14957 ( .A(net_14875), .Z(net_14876) );
NAND2_X2 inst_3809 ( .A1(net_10078), .A2(net_4534), .ZN(net_4529) );
CLKBUF_X2 inst_14357 ( .A(net_13521), .Z(net_14276) );
CLKBUF_X2 inst_11990 ( .A(net_11908), .Z(net_11909) );
NAND2_X2 inst_4004 ( .ZN(net_4085), .A2(net_3390), .A1(net_3169) );
CLKBUF_X2 inst_12708 ( .A(net_12626), .Z(net_12627) );
CLKBUF_X2 inst_15352 ( .A(net_14100), .Z(net_15271) );
CLKBUF_X2 inst_11368 ( .A(net_11199), .Z(net_11287) );
CLKBUF_X2 inst_14896 ( .A(net_14814), .Z(net_14815) );
CLKBUF_X2 inst_11838 ( .A(net_11756), .Z(net_11757) );
AOI211_X2 inst_10315 ( .C2(net_10122), .ZN(net_2418), .B(net_1717), .A(net_1438), .C1(net_683) );
INV_X4 inst_6171 ( .A(net_9743), .ZN(net_2000) );
DFF_X1 inst_8887 ( .Q(net_99), .CK(net_15334), .D(x3300) );
CLKBUF_X2 inst_14236 ( .A(net_12575), .Z(net_14155) );
CLKBUF_X2 inst_15300 ( .A(net_15218), .Z(net_15219) );
NAND2_X2 inst_3798 ( .ZN(net_7282), .A1(net_4312), .A2(net_4185) );
INV_X2 inst_6865 ( .A(net_3419), .ZN(net_3229) );
INV_X4 inst_5232 ( .ZN(net_5265), .A(net_1484) );
NAND2_X2 inst_4109 ( .ZN(net_3049), .A1(net_2279), .A2(net_2119) );
NAND2_X2 inst_4192 ( .A1(net_4190), .ZN(net_2917), .A2(net_1850) );
CLKBUF_X2 inst_12948 ( .A(net_12866), .Z(net_12867) );
AOI21_X2 inst_10048 ( .ZN(net_7387), .A(net_7386), .B2(net_6845), .B1(net_6589) );
NOR2_X2 inst_3004 ( .A1(net_8455), .ZN(net_1570), .A2(net_864) );
NAND2_X2 inst_3780 ( .A2(net_7277), .ZN(net_4730), .A1(net_1975) );
CLKBUF_X2 inst_12396 ( .A(net_12314), .Z(net_12315) );
CLKBUF_X2 inst_11305 ( .A(net_10966), .Z(net_11224) );
NOR2_X2 inst_2647 ( .A2(net_7530), .A1(net_5405), .ZN(net_5401) );
INV_X4 inst_4672 ( .ZN(net_5824), .A(net_5260) );
INV_X4 inst_6576 ( .A(net_9208), .ZN(net_1505) );
CLKBUF_X2 inst_14438 ( .A(net_14356), .Z(net_14357) );
CLKBUF_X2 inst_12363 ( .A(net_10916), .Z(net_12282) );
CLKBUF_X2 inst_15464 ( .A(net_15382), .Z(net_15383) );
NOR3_X2 inst_2456 ( .ZN(net_3454), .A1(net_2169), .A3(net_1727), .A2(net_1090) );
CLKBUF_X2 inst_11959 ( .A(net_11877), .Z(net_11878) );
INV_X4 inst_5629 ( .ZN(net_1240), .A(x6599) );
NOR2_X2 inst_2710 ( .A1(net_4876), .ZN(net_4469), .A2(net_3874) );
OAI22_X2 inst_1058 ( .B2(net_10135), .A1(net_10134), .ZN(net_7305), .A2(net_7304), .B1(net_3209) );
NOR2_X2 inst_2887 ( .A2(net_2402), .ZN(net_1784), .A1(net_1353) );
CLKBUF_X2 inst_12162 ( .A(net_11779), .Z(net_12081) );
CLKBUF_X2 inst_12639 ( .A(net_12557), .Z(net_12558) );
CLKBUF_X2 inst_11120 ( .A(net_11038), .Z(net_11039) );
NAND2_X4 inst_3360 ( .A2(net_8997), .A1(net_8996), .ZN(net_8930) );
INV_X2 inst_6821 ( .ZN(net_4424), .A(net_4423) );
INV_X4 inst_4984 ( .ZN(net_3056), .A(net_1959) );
DFF_X1 inst_8805 ( .Q(net_10132), .D(net_3989), .CK(net_10768) );
OAI221_X2 inst_1473 ( .A(net_7783), .C2(net_7782), .ZN(net_7692), .B2(net_7690), .C1(net_3225), .B1(net_2450) );
INV_X4 inst_5334 ( .ZN(net_1487), .A(net_1255) );
CLKBUF_X2 inst_12793 ( .A(net_12711), .Z(net_12712) );
CLKBUF_X2 inst_14098 ( .A(net_14016), .Z(net_14017) );
OAI21_X2 inst_1788 ( .B2(net_7731), .ZN(net_7539), .A(net_7428), .B1(net_5237) );
AOI22_X2 inst_9306 ( .B1(net_9712), .A2(net_5755), .B2(net_5754), .ZN(net_5672), .A1(net_249) );
OAI22_X2 inst_1272 ( .ZN(net_4750), .A1(net_4749), .A2(net_4746), .B2(net_4745), .B1(net_1270) );
NAND2_X2 inst_4182 ( .ZN(net_2512), .A2(net_1566), .A1(net_1141) );
SDFF_X2 inst_632 ( .Q(net_9468), .D(net_9468), .SE(net_3293), .CK(net_12444), .SI(x1459) );
CLKBUF_X2 inst_14566 ( .A(net_12226), .Z(net_14485) );
XOR2_X2 inst_0 ( .Z(net_8404), .B(net_8403), .A(net_8180) );
NOR2_X2 inst_2852 ( .ZN(net_2215), .A1(net_2214), .A2(net_1697) );
CLKBUF_X2 inst_13934 ( .A(net_12710), .Z(net_13853) );
INV_X2 inst_6751 ( .A(net_7275), .ZN(net_6614) );
CLKBUF_X2 inst_11405 ( .A(net_11323), .Z(net_11324) );
CLKBUF_X2 inst_14582 ( .A(net_12622), .Z(net_14501) );
CLKBUF_X2 inst_11199 ( .A(net_11117), .Z(net_11118) );
NAND2_X2 inst_3973 ( .A1(net_9531), .ZN(net_3304), .A2(net_2856) );
CLKBUF_X2 inst_12266 ( .A(net_12184), .Z(net_12185) );
DFF_X2 inst_7584 ( .QN(net_10149), .D(net_7554), .CK(net_12371) );
AOI22_X2 inst_8994 ( .A2(net_8941), .ZN(net_8615), .A1(net_8614), .B2(net_8612), .B1(net_7636) );
XNOR2_X2 inst_433 ( .B(net_9303), .ZN(net_1047), .A(net_211) );
CLKBUF_X2 inst_13520 ( .A(net_13438), .Z(net_13439) );
OAI21_X2 inst_1983 ( .ZN(net_2822), .B1(net_2821), .A(net_2165), .B2(net_1842) );
CLKBUF_X2 inst_13771 ( .A(net_11032), .Z(net_13690) );
CLKBUF_X2 inst_13249 ( .A(net_11489), .Z(net_13168) );
CLKBUF_X2 inst_11817 ( .A(net_11670), .Z(net_11736) );
INV_X4 inst_4939 ( .ZN(net_4966), .A(net_2234) );
CLKBUF_X2 inst_13748 ( .A(net_13503), .Z(net_13667) );
CLKBUF_X2 inst_13772 ( .A(net_13690), .Z(net_13691) );
CLKBUF_X2 inst_11312 ( .A(net_11230), .Z(net_11231) );
INV_X4 inst_6417 ( .ZN(net_1401), .A(net_198) );
CLKBUF_X1 inst_8984 ( .A(x185142), .Z(x921) );
INV_X16 inst_7323 ( .ZN(net_6041), .A(net_5159) );
OAI21_X2 inst_1948 ( .B2(net_10444), .A(net_10443), .ZN(net_3986), .B1(net_3985) );
INV_X2 inst_7158 ( .A(net_4566), .ZN(net_695) );
CLKBUF_X2 inst_11955 ( .A(net_11873), .Z(net_11874) );
DFF_X1 inst_8409 ( .D(net_8806), .CK(net_14205), .Q(x682) );
DFF_X1 inst_8638 ( .Q(net_9888), .D(net_7217), .CK(net_14379) );
AOI22_X2 inst_9269 ( .B1(net_9808), .ZN(net_5767), .A1(net_5766), .B2(net_5765), .A2(net_246) );
CLKBUF_X2 inst_15148 ( .A(net_11824), .Z(net_15067) );
DFF_X2 inst_8266 ( .Q(net_10390), .D(net_4806), .CK(net_15209) );
INV_X4 inst_5781 ( .ZN(net_1691), .A(net_703) );
CLKBUF_X2 inst_14733 ( .A(net_12877), .Z(net_14652) );
CLKBUF_X2 inst_13476 ( .A(net_11049), .Z(net_13395) );
XNOR2_X2 inst_422 ( .A(net_7595), .ZN(net_2154), .B(net_700) );
CLKBUF_X2 inst_15325 ( .A(net_10576), .Z(net_15244) );
INV_X2 inst_7151 ( .A(net_1021), .ZN(net_994) );
OAI211_X2 inst_2243 ( .C1(net_7241), .C2(net_6480), .ZN(net_6461), .B(net_5523), .A(net_3679) );
OAI221_X2 inst_1475 ( .A(net_7783), .B2(net_7782), .C2(net_7690), .ZN(net_7689), .B1(net_2727), .C1(net_1309) );
OAI222_X2 inst_1426 ( .B2(net_8857), .A2(net_8857), .ZN(net_3401), .A1(net_3400), .C2(net_3399), .C1(net_2332), .B1(net_1298) );
AOI22_X2 inst_9021 ( .A1(net_8002), .B2(net_8001), .ZN(net_7998), .A2(net_7948), .B1(net_3565) );
INV_X4 inst_4812 ( .A(net_10175), .ZN(net_5347) );
NAND4_X2 inst_3090 ( .ZN(net_4484), .A4(net_4048), .A1(net_3848), .A2(net_3766), .A3(net_3443) );
OAI221_X2 inst_1637 ( .B1(net_10314), .C1(net_7129), .B2(net_5591), .ZN(net_5569), .C2(net_4902), .A(net_3507) );
CLKBUF_X2 inst_14466 ( .A(net_13147), .Z(net_14385) );
OAI222_X2 inst_1352 ( .B1(net_9260), .ZN(net_7472), .C2(net_7280), .B2(net_7280), .A1(net_7048), .A2(net_6902), .C1(net_6319) );
CLKBUF_X2 inst_12338 ( .A(net_10654), .Z(net_12257) );
CLKBUF_X2 inst_14635 ( .A(net_14553), .Z(net_14554) );
AOI21_X2 inst_10012 ( .B1(net_8968), .ZN(net_8594), .B2(net_8583), .A(net_8496) );
CLKBUF_X2 inst_14624 ( .A(net_14473), .Z(net_14543) );
DFF_X2 inst_8355 ( .Q(net_9227), .D(net_2492), .CK(net_15273) );
OAI211_X2 inst_2261 ( .C1(net_7234), .A(net_6546), .C2(net_6480), .ZN(net_6292), .B(net_5415) );
AOI221_X2 inst_9955 ( .C1(net_9974), .B1(net_9677), .B2(net_5966), .ZN(net_4777), .A(net_4346), .C2(net_2541) );
INV_X4 inst_4879 ( .ZN(net_3485), .A(net_3013) );
CLKBUF_X2 inst_14524 ( .A(net_13515), .Z(net_14443) );
INV_X4 inst_4695 ( .ZN(net_4832), .A(net_4648) );
NAND2_X2 inst_4142 ( .A2(net_2235), .ZN(net_2126), .A1(net_1651) );
NAND2_X2 inst_3390 ( .A2(net_8849), .A1(net_8756), .ZN(net_8750) );
CLKBUF_X2 inst_12125 ( .A(net_10661), .Z(net_12044) );
AOI22_X2 inst_9076 ( .B1(net_9666), .A2(net_6684), .B2(net_6683), .ZN(net_6590), .A1(net_235) );
DFF_X1 inst_8513 ( .QN(net_8823), .D(net_7544), .CK(net_14415) );
CLKBUF_X2 inst_15742 ( .A(net_13613), .Z(net_15661) );
CLKBUF_X2 inst_11260 ( .A(net_11178), .Z(net_11179) );
AOI22_X2 inst_9097 ( .A1(net_9678), .A2(net_6420), .ZN(net_6395), .B2(net_5263), .B1(net_116) );
DFF_X2 inst_8178 ( .QN(net_9933), .D(net_5029), .CK(net_14442) );
DFF_X2 inst_7609 ( .QN(net_9344), .D(net_7134), .CK(net_15289) );
NOR2_X2 inst_2930 ( .ZN(net_2403), .A1(net_843), .A2(net_739) );
CLKBUF_X2 inst_12680 ( .A(net_11563), .Z(net_12599) );
INV_X4 inst_5683 ( .ZN(net_4380), .A(net_1096) );
CLKBUF_X2 inst_12206 ( .A(net_10942), .Z(net_12125) );
INV_X4 inst_4790 ( .ZN(net_3996), .A(net_3526) );
CLKBUF_X2 inst_15267 ( .A(net_14948), .Z(net_15186) );
CLKBUF_X2 inst_14774 ( .A(net_10663), .Z(net_14693) );
AOI221_X2 inst_9851 ( .B1(net_9868), .B2(net_9101), .A(net_6945), .C1(net_6944), .ZN(net_6867), .C2(net_239) );
NAND2_X2 inst_4307 ( .A2(net_10125), .ZN(net_2181), .A1(net_1204) );
NOR2_X2 inst_2859 ( .ZN(net_4499), .A1(net_2071), .A2(net_1687) );
XNOR2_X2 inst_397 ( .ZN(net_2777), .A(net_1994), .B(net_1993) );
SDFF_X2 inst_504 ( .SE(net_9540), .SI(net_8197), .Q(net_309), .D(net_309), .CK(net_11640) );
DFF_X1 inst_8601 ( .Q(net_9691), .D(net_7257), .CK(net_13227) );
NAND3_X2 inst_3192 ( .ZN(net_7576), .A3(net_7575), .A1(net_7573), .A2(net_7423) );
INV_X4 inst_5006 ( .ZN(net_3591), .A(net_1959) );
CLKBUF_X2 inst_14240 ( .A(net_14158), .Z(net_14159) );
AOI22_X2 inst_9026 ( .A1(net_8002), .B2(net_8001), .ZN(net_7954), .B1(net_7953), .A2(net_7920) );
AOI221_X2 inst_9780 ( .C1(net_9348), .B1(net_9157), .A(net_7157), .ZN(net_7156), .B2(net_7155), .C2(net_7154) );
OAI22_X2 inst_1297 ( .B1(net_10048), .A1(net_9949), .A2(net_4274), .B2(net_3588), .ZN(net_3564) );
NAND3_X2 inst_3194 ( .A1(net_7930), .ZN(net_7559), .A2(net_7002), .A3(net_2850) );
CLKBUF_X2 inst_13585 ( .A(net_13503), .Z(net_13504) );
CLKBUF_X2 inst_11129 ( .A(net_11047), .Z(net_11048) );
NAND2_X2 inst_3884 ( .ZN(net_4018), .A1(net_4017), .A2(net_3540) );
CLKBUF_X2 inst_13831 ( .A(net_13749), .Z(net_13750) );
AOI22_X2 inst_9146 ( .A1(net_9700), .A2(net_6402), .ZN(net_6339), .B2(net_5263), .B1(net_140) );
INV_X4 inst_6296 ( .ZN(net_7237), .A(x3889) );
NAND2_X2 inst_4246 ( .A2(net_2767), .A1(net_2209), .ZN(net_1439) );
OAI22_X2 inst_1173 ( .B1(net_10041), .A1(net_7231), .A2(net_5107), .B2(net_5105), .ZN(net_5088) );
NAND2_X2 inst_3904 ( .ZN(net_3901), .A2(net_3059), .A1(net_1972) );
AOI222_X1 inst_9708 ( .B1(net_9505), .A2(net_8310), .B2(net_8309), .C2(net_8308), .ZN(net_8268), .C1(net_8208), .A1(x2707) );
CLKBUF_X2 inst_10634 ( .A(net_10552), .Z(net_10553) );
NOR2_X2 inst_2908 ( .A1(net_10267), .ZN(net_3199), .A2(net_1551) );
INV_X4 inst_6333 ( .A(net_9965), .ZN(net_413) );
INV_X4 inst_5019 ( .ZN(net_2096), .A(net_2095) );
INV_X4 inst_5649 ( .ZN(net_1255), .A(net_835) );
OAI222_X2 inst_1393 ( .B1(net_7728), .A2(net_7727), .C2(net_7726), .ZN(net_5799), .B2(net_5212), .A1(net_4138), .C1(net_1324) );
INV_X4 inst_6276 ( .A(net_10031), .ZN(net_888) );
NAND2_X2 inst_3519 ( .A2(net_9596), .A1(net_9073), .ZN(net_8186) );
NAND2_X2 inst_4075 ( .ZN(net_2640), .A2(net_2639), .A1(net_1869) );
CLKBUF_X2 inst_13402 ( .A(net_13320), .Z(net_13321) );
AOI22_X2 inst_9507 ( .B1(net_9922), .A1(net_9692), .A2(net_5966), .B2(net_4969), .ZN(net_3816) );
CLKBUF_X2 inst_15720 ( .A(net_15638), .Z(net_15639) );
INV_X4 inst_4893 ( .ZN(net_2899), .A(net_2898) );
INV_X4 inst_5875 ( .A(net_7021), .ZN(net_629) );
INV_X4 inst_5153 ( .ZN(net_1895), .A(net_1582) );
INV_X4 inst_5731 ( .ZN(net_996), .A(net_753) );
CLKBUF_X2 inst_11318 ( .A(net_10764), .Z(net_11237) );
CLKBUF_X2 inst_14264 ( .A(net_12408), .Z(net_14183) );
DFF_X1 inst_8514 ( .Q(net_9387), .D(net_7593), .CK(net_13155) );
INV_X2 inst_6717 ( .ZN(net_7939), .A(net_7913) );
DFF_X1 inst_8631 ( .Q(net_9879), .D(net_7232), .CK(net_13461) );
CLKBUF_X2 inst_13118 ( .A(net_13036), .Z(net_13037) );
AOI221_X2 inst_9807 ( .B1(net_9986), .A(net_7090), .B2(net_7089), .C2(net_7088), .ZN(net_6995), .C1(net_258) );
CLKBUF_X2 inst_14446 ( .A(net_12582), .Z(net_14365) );
AOI22_X2 inst_9089 ( .A1(net_9699), .ZN(net_6405), .A2(net_6404), .B2(net_5263), .B1(net_139) );
CLKBUF_X2 inst_13684 ( .A(net_13602), .Z(net_13603) );
INV_X4 inst_6459 ( .A(net_10466), .ZN(net_7333) );
INV_X4 inst_4791 ( .ZN(net_8122), .A(net_4784) );
DFF_X2 inst_8007 ( .QN(net_10328), .D(net_5501), .CK(net_12134) );
AOI22_X2 inst_9302 ( .B1(net_10010), .A2(net_5743), .B2(net_5742), .ZN(net_5676), .A1(net_250) );
INV_X2 inst_7244 ( .ZN(net_367), .A(net_166) );
NOR2_X2 inst_2937 ( .ZN(net_2340), .A1(net_1250), .A2(net_783) );
CLKBUF_X2 inst_12995 ( .A(net_12913), .Z(net_12914) );
INV_X4 inst_6283 ( .A(net_9518), .ZN(net_2139) );
DFF_X2 inst_7380 ( .D(net_8640), .QN(net_275), .CK(net_14924) );
DFF_X2 inst_7864 ( .Q(net_10001), .D(net_6274), .CK(net_12773) );
OR4_X2 inst_687 ( .ZN(net_7628), .A1(net_7507), .A2(net_7157), .A4(net_3515), .A3(net_3478) );
DFF_X2 inst_7387 ( .D(net_8652), .QN(net_274), .CK(net_14917) );
INV_X4 inst_5857 ( .ZN(net_1350), .A(net_1062) );
AOI22_X2 inst_9463 ( .B1(net_10004), .A1(net_9739), .A2(net_6442), .ZN(net_3864), .B2(net_2468) );
OAI21_X2 inst_1774 ( .ZN(net_7822), .B2(net_7816), .B1(net_7815), .A(net_7278) );
NOR4_X2 inst_2319 ( .A2(net_9751), .ZN(net_6638), .A3(net_6321), .A4(net_5795), .A1(net_3746) );
INV_X2 inst_7091 ( .ZN(net_1113), .A(net_1112) );
DFF_X2 inst_8032 ( .Q(net_9230), .D(net_5448), .CK(net_11311) );
CLKBUF_X2 inst_12596 ( .A(net_12514), .Z(net_12515) );
INV_X4 inst_5519 ( .ZN(net_968), .A(net_967) );
OAI22_X2 inst_985 ( .A2(net_8962), .B2(net_8659), .ZN(net_8655), .A1(net_6252), .B1(net_6235) );
DFF_X2 inst_7927 ( .QN(net_10410), .D(net_5550), .CK(net_14606) );
OAI211_X2 inst_2225 ( .C1(net_7184), .C2(net_6480), .ZN(net_6479), .B(net_5531), .A(net_3679) );
CLKBUF_X2 inst_12473 ( .A(net_10975), .Z(net_12392) );
CLKBUF_X2 inst_13805 ( .A(net_13723), .Z(net_13724) );
INV_X2 inst_6943 ( .A(net_4281), .ZN(net_1908) );
NOR2_X2 inst_2513 ( .ZN(net_8531), .A1(net_8398), .A2(net_8338) );
NAND2_X2 inst_4061 ( .A2(net_3347), .ZN(net_2759), .A1(net_2758) );
OAI211_X2 inst_2254 ( .C1(net_7249), .C2(net_6542), .ZN(net_6437), .B(net_5437), .A(net_3679) );
CLKBUF_X2 inst_14690 ( .A(net_14608), .Z(net_14609) );
DFF_X2 inst_7775 ( .Q(net_9697), .D(net_6527), .CK(net_14312) );
INV_X4 inst_6255 ( .A(net_9933), .ZN(net_674) );
AOI21_X2 inst_10111 ( .A(net_8862), .ZN(net_4586), .B2(net_4394), .B1(net_4264) );
CLKBUF_X2 inst_12985 ( .A(net_12903), .Z(net_12904) );
CLKBUF_X2 inst_10627 ( .A(net_10545), .Z(net_10546) );
CLKBUF_X2 inst_14208 ( .A(net_13566), .Z(net_14127) );
CLKBUF_X2 inst_12563 ( .A(net_12481), .Z(net_12482) );
INV_X4 inst_5918 ( .ZN(net_1249), .A(net_737) );
CLKBUF_X2 inst_12969 ( .A(net_12887), .Z(net_12888) );
AOI22_X2 inst_9255 ( .B2(net_8041), .A2(net_6109), .ZN(net_6051), .B1(net_3761), .A1(net_1983) );
OAI21_X2 inst_2007 ( .B1(net_2216), .ZN(net_2115), .A(net_1710), .B2(net_1423) );
CLKBUF_X2 inst_10922 ( .A(net_10840), .Z(net_10841) );
CLKBUF_X2 inst_12519 ( .A(net_12437), .Z(net_12438) );
CLKBUF_X2 inst_15479 ( .A(net_15397), .Z(net_15398) );
NAND2_X2 inst_3644 ( .A2(net_6904), .ZN(net_6897), .A1(net_6237) );
CLKBUF_X2 inst_10965 ( .A(net_10883), .Z(net_10884) );
OR2_X4 inst_805 ( .A1(net_10261), .ZN(net_2078), .A2(net_1367) );
CLKBUF_X2 inst_11755 ( .A(net_11673), .Z(net_11674) );
XNOR2_X2 inst_354 ( .ZN(net_2779), .A(net_2040), .B(net_2002) );
CLKBUF_X2 inst_13794 ( .A(net_11236), .Z(net_13713) );
AOI221_X2 inst_9991 ( .B1(net_3853), .ZN(net_3197), .C2(net_3196), .A(net_2734), .B2(net_2232), .C1(net_2213) );
INV_X4 inst_6005 ( .ZN(net_531), .A(net_229) );
OAI22_X2 inst_1145 ( .A1(net_7184), .A2(net_5134), .B2(net_5133), .ZN(net_5128), .B1(net_403) );
CLKBUF_X2 inst_12859 ( .A(net_12418), .Z(net_12778) );
INV_X4 inst_6235 ( .A(net_9244), .ZN(net_757) );
CLKBUF_X2 inst_12387 ( .A(net_12305), .Z(net_12306) );
CLKBUF_X2 inst_15380 ( .A(net_15298), .Z(net_15299) );
CLKBUF_X2 inst_12664 ( .A(net_12582), .Z(net_12583) );
CLKBUF_X2 inst_13735 ( .A(net_13653), .Z(net_13654) );
INV_X4 inst_5603 ( .ZN(net_2318), .A(net_1101) );
CLKBUF_X2 inst_14257 ( .A(net_14175), .Z(net_14176) );
INV_X4 inst_6569 ( .A(net_10358), .ZN(net_4446) );
XNOR2_X2 inst_373 ( .ZN(net_2475), .A(net_2472), .B(net_1725) );
CLKBUF_X2 inst_14804 ( .A(net_14722), .Z(net_14723) );
DFF_X2 inst_7731 ( .Q(net_9700), .D(net_6236), .CK(net_14238) );
OAI21_X2 inst_1868 ( .ZN(net_5905), .B2(net_5346), .A(net_5345), .B1(net_5344) );
CLKBUF_X2 inst_13672 ( .A(net_10817), .Z(net_13591) );
CLKBUF_X2 inst_11428 ( .A(net_11346), .Z(net_11347) );
AOI22_X2 inst_9537 ( .B1(net_10286), .A1(net_10181), .B2(net_4774), .A2(net_4217), .ZN(net_3784) );
DFF_X1 inst_8414 ( .QN(net_9363), .D(net_8790), .CK(net_11931) );
XOR2_X2 inst_22 ( .B(net_7848), .Z(net_2447), .A(net_2446) );
CLKBUF_X2 inst_13914 ( .A(net_11690), .Z(net_13833) );
OAI221_X2 inst_1717 ( .ZN(net_3620), .A(net_3150), .C2(net_2312), .B1(net_2306), .B2(net_1851), .C1(net_970) );
NAND4_X2 inst_3099 ( .ZN(net_4344), .A1(net_3851), .A3(net_3850), .A4(net_3586), .A2(net_3444) );
CLKBUF_X2 inst_15206 ( .A(net_15124), .Z(net_15125) );
CLKBUF_X2 inst_13289 ( .A(net_12046), .Z(net_13208) );
INV_X2 inst_7034 ( .ZN(net_1426), .A(net_1425) );
NOR2_X2 inst_2901 ( .ZN(net_2119), .A2(net_1643), .A1(net_946) );
OR2_X4 inst_767 ( .ZN(net_4495), .A1(net_4323), .A2(net_4073) );
DFF_X2 inst_7657 ( .D(net_6702), .QN(net_190), .CK(net_14560) );
CLKBUF_X2 inst_14065 ( .A(net_13983), .Z(net_13984) );
INV_X4 inst_6080 ( .A(net_9643), .ZN(net_644) );
NAND2_X4 inst_3356 ( .ZN(net_8418), .A1(net_8382), .A2(net_8381) );
OR3_X2 inst_718 ( .ZN(net_3048), .A2(net_3047), .A1(net_3018), .A3(net_2935) );
AND2_X4 inst_10405 ( .ZN(net_4977), .A2(net_4976), .A1(net_207) );
NAND2_X2 inst_4024 ( .ZN(net_5249), .A2(net_4634), .A1(net_1114) );
DFF_X2 inst_7914 ( .Q(net_9747), .D(net_5880), .CK(net_11947) );
HA_X1 inst_7362 ( .CO(net_2195), .S(net_1457), .A(net_618), .B(net_585) );
CLKBUF_X2 inst_15374 ( .A(net_15292), .Z(net_15293) );
DFF_X2 inst_8100 ( .Q(net_9840), .D(net_5129), .CK(net_14303) );
AOI22_X2 inst_9166 ( .A2(net_6382), .ZN(net_6306), .A1(net_6305), .B2(net_5263), .B1(net_3052) );
INV_X4 inst_5585 ( .ZN(net_4166), .A(net_885) );
DFF_X2 inst_8350 ( .QN(net_10269), .D(net_2774), .CK(net_14430) );
NAND2_X2 inst_4310 ( .ZN(net_1464), .A2(net_1197), .A1(net_974) );
SDFF_X2 inst_526 ( .SI(net_9335), .Q(net_9280), .D(net_9280), .SE(net_7588), .CK(net_13072) );
OAI211_X2 inst_2147 ( .C2(net_6778), .ZN(net_6701), .A(net_6325), .B(net_6064), .C1(net_4755) );
CLKBUF_X2 inst_13171 ( .A(net_13089), .Z(net_13090) );
OAI22_X2 inst_1178 ( .A1(net_7198), .A2(net_5151), .B2(net_5150), .ZN(net_5081), .B1(net_785) );
OAI211_X2 inst_2091 ( .C2(net_6778), .ZN(net_6757), .A(net_6385), .B(net_6117), .C1(net_494) );
NAND4_X2 inst_3104 ( .ZN(net_4339), .A2(net_3797), .A4(net_3796), .A1(net_3750), .A3(net_3414) );
AOI22_X2 inst_9174 ( .A1(net_9914), .B1(net_9815), .A2(net_8042), .B2(net_8041), .ZN(net_6144) );
OAI221_X2 inst_1450 ( .B2(net_9627), .B1(net_8971), .ZN(net_8145), .A(net_7965), .C2(net_3526), .C1(net_171) );
DFF_X1 inst_8423 ( .D(net_8751), .Q(net_245), .CK(net_12688) );
INV_X2 inst_6689 ( .ZN(net_8335), .A(net_8273) );
CLKBUF_X2 inst_12247 ( .A(net_12165), .Z(net_12166) );
CLKBUF_X2 inst_10733 ( .A(net_10651), .Z(net_10652) );
INV_X4 inst_5511 ( .ZN(net_2564), .A(net_1002) );
NAND4_X2 inst_3123 ( .ZN(net_3315), .A1(net_2620), .A3(net_1043), .A4(net_1042), .A2(net_789) );
DFF_X2 inst_8066 ( .QN(net_10458), .D(net_5325), .CK(net_12459) );
CLKBUF_X2 inst_11592 ( .A(net_11510), .Z(net_11511) );
CLKBUF_X2 inst_11149 ( .A(net_10589), .Z(net_11068) );
INV_X4 inst_5863 ( .ZN(net_5493), .A(net_1361) );
CLKBUF_X2 inst_10645 ( .A(net_10563), .Z(net_10564) );
NAND2_X2 inst_3725 ( .A1(net_10189), .ZN(net_5776), .A2(net_5774) );
INV_X4 inst_5400 ( .ZN(net_3742), .A(net_1165) );
SDFF_X2 inst_500 ( .SE(net_9540), .SI(net_8209), .Q(net_289), .D(net_289), .CK(net_11719) );
OAI221_X2 inst_1592 ( .B2(net_10481), .ZN(net_5815), .B1(net_5175), .A(net_4961), .C2(net_4960), .C1(net_4245) );
INV_X4 inst_5348 ( .ZN(net_5356), .A(net_1240) );
OAI21_X2 inst_1770 ( .ZN(net_8009), .A(net_7873), .B2(net_7868), .B1(net_3984) );
CLKBUF_X2 inst_14403 ( .A(net_14321), .Z(net_14322) );
SDFF_X2 inst_550 ( .D(net_9152), .SE(net_7248), .SI(net_194), .Q(net_194), .CK(net_15350) );
NAND2_X2 inst_3413 ( .ZN(net_9113), .A1(net_8469), .A2(net_8435) );
INV_X4 inst_6095 ( .ZN(net_7221), .A(x4587) );
INV_X2 inst_6758 ( .ZN(net_6240), .A(net_6239) );
INV_X8 inst_4483 ( .ZN(net_8487), .A(net_8419) );
CLKBUF_X2 inst_12857 ( .A(net_12775), .Z(net_12776) );
INV_X4 inst_5913 ( .ZN(net_1006), .A(net_696) );
CLKBUF_X2 inst_11972 ( .A(net_11890), .Z(net_11891) );
CLKBUF_X2 inst_13610 ( .A(net_11521), .Z(net_13529) );
DFF_X2 inst_8311 ( .QN(net_9161), .D(net_4287), .CK(net_11808) );
DFF_X1 inst_8702 ( .D(net_6717), .Q(net_137), .CK(net_13217) );
CLKBUF_X2 inst_15617 ( .A(net_11980), .Z(net_15536) );
CLKBUF_X2 inst_15417 ( .A(net_15335), .Z(net_15336) );
CLKBUF_X2 inst_11109 ( .A(net_11027), .Z(net_11028) );
CLKBUF_X2 inst_14132 ( .A(net_14050), .Z(net_14051) );
INV_X4 inst_5471 ( .ZN(net_3067), .A(net_1011) );
OAI222_X2 inst_1419 ( .B2(net_7665), .A2(net_7664), .C2(net_7663), .ZN(net_4925), .B1(net_3221), .A1(net_2172), .C1(net_1267) );
NOR2_X2 inst_2661 ( .A1(net_9073), .ZN(net_5014), .A2(net_4731) );
DFF_X2 inst_8237 ( .Q(net_10498), .D(net_4883), .CK(net_13172) );
INV_X4 inst_6034 ( .ZN(net_2521), .A(net_200) );
CLKBUF_X2 inst_14544 ( .A(net_14462), .Z(net_14463) );
NOR2_X2 inst_2501 ( .A1(net_9066), .ZN(net_8541), .A2(net_8492) );
NAND2_X2 inst_3548 ( .A1(net_9273), .A2(net_9268), .ZN(net_8036) );
CLKBUF_X2 inst_15246 ( .A(net_15164), .Z(net_15165) );
SDFF_X2 inst_594 ( .Q(net_9264), .SE(net_4589), .D(net_147), .SI(net_113), .CK(net_12548) );
CLKBUF_X2 inst_13848 ( .A(net_13766), .Z(net_13767) );
MUX2_X1 inst_4435 ( .S(net_6041), .A(net_311), .B(x3949), .Z(x33) );
CLKBUF_X2 inst_14164 ( .A(net_14082), .Z(net_14083) );
OAI221_X2 inst_1632 ( .B1(net_10422), .C1(net_7139), .A(net_5575), .ZN(net_5574), .B2(net_4477), .C2(net_4455) );
OAI211_X2 inst_2175 ( .C1(net_7224), .C2(net_6548), .ZN(net_6534), .B(net_5662), .A(net_3679) );
NAND2_X2 inst_4241 ( .A1(net_3528), .A2(net_2712), .ZN(net_2083) );
OR2_X2 inst_925 ( .ZN(net_3019), .A2(net_3018), .A1(net_2488) );
CLKBUF_X2 inst_13314 ( .A(net_10585), .Z(net_13233) );
OAI211_X2 inst_2193 ( .C1(net_7219), .C2(net_6542), .ZN(net_6516), .B(net_5612), .A(net_3679) );
NOR3_X2 inst_2378 ( .ZN(net_7981), .A3(net_7831), .A1(net_3315), .A2(net_2932) );
AOI211_X2 inst_10302 ( .B(net_6321), .ZN(net_3537), .A(net_3536), .C2(net_3063), .C1(net_2069) );
INV_X4 inst_6302 ( .A(net_10009), .ZN(net_429) );
CLKBUF_X2 inst_14137 ( .A(net_14055), .Z(net_14056) );
AOI21_X4 inst_9996 ( .ZN(net_8721), .B1(net_8717), .A(net_8192), .B2(net_8118) );
DFF_X1 inst_8734 ( .Q(net_9119), .D(net_5871), .CK(net_10581) );
AOI221_X2 inst_9793 ( .B1(net_9972), .A(net_7090), .B2(net_7089), .C1(net_7088), .ZN(net_7019), .C2(net_244) );
AOI22_X2 inst_8999 ( .B1(net_9469), .A1(net_9461), .A2(net_8951), .ZN(net_8499), .B2(net_8475) );
INV_X4 inst_6147 ( .A(net_10228), .ZN(net_1062) );
CLKBUF_X2 inst_14392 ( .A(net_14310), .Z(net_14311) );
OAI221_X2 inst_1536 ( .B1(net_10324), .B2(net_9047), .C2(net_7287), .ZN(net_7232), .C1(net_7231), .A(net_6801) );
OR2_X2 inst_881 ( .A2(net_7038), .ZN(net_6317), .A1(net_6316) );
CLKBUF_X2 inst_13874 ( .A(net_13792), .Z(net_13793) );
CLKBUF_X2 inst_11300 ( .A(net_11218), .Z(net_11219) );
NAND2_X2 inst_3876 ( .ZN(net_4032), .A2(net_4028), .A1(net_1970) );
NAND2_X2 inst_3848 ( .ZN(net_4656), .A2(net_4236), .A1(net_2891) );
CLKBUF_X2 inst_13164 ( .A(net_11742), .Z(net_13083) );
INV_X2 inst_7001 ( .ZN(net_1625), .A(net_1624) );
CLKBUF_X2 inst_12175 ( .A(net_11086), .Z(net_12094) );
CLKBUF_X2 inst_12079 ( .A(net_11997), .Z(net_11998) );
CLKBUF_X2 inst_15237 ( .A(net_15155), .Z(net_15156) );
NAND2_X2 inst_3706 ( .A1(net_10069), .ZN(net_5923), .A2(net_5892) );
AOI21_X2 inst_10072 ( .ZN(net_6618), .A(net_6617), .B1(net_4931), .B2(net_4676) );
CLKBUF_X2 inst_13979 ( .A(net_13897), .Z(net_13898) );
CLKBUF_X2 inst_11153 ( .A(net_10615), .Z(net_11072) );
AOI22_X2 inst_9219 ( .A1(net_9912), .B1(net_9813), .B2(net_6133), .A2(net_6109), .ZN(net_6092) );
XNOR2_X2 inst_247 ( .ZN(net_4133), .A(net_3964), .B(net_2088) );
CLKBUF_X2 inst_15569 ( .A(net_14700), .Z(net_15488) );
INV_X2 inst_7066 ( .A(net_3668), .ZN(net_1258) );
INV_X4 inst_6089 ( .ZN(net_497), .A(net_230) );
XNOR2_X2 inst_403 ( .A(net_9156), .B(net_9155), .ZN(net_2476) );
CLKBUF_X2 inst_12031 ( .A(net_11949), .Z(net_11950) );
CLKBUF_X2 inst_14560 ( .A(net_14478), .Z(net_14479) );
INV_X2 inst_6740 ( .ZN(net_7163), .A(net_7024) );
AND2_X2 inst_10501 ( .A2(net_10135), .ZN(net_6042), .A1(net_1483) );
NAND2_X2 inst_3446 ( .A1(net_9452), .ZN(net_9014), .A2(net_8477) );
NOR2_X2 inst_2728 ( .A2(net_10165), .ZN(net_5220), .A1(net_3960) );
CLKBUF_X2 inst_10796 ( .A(net_10714), .Z(net_10715) );
DFF_X1 inst_8847 ( .QN(net_9187), .D(net_1457), .CK(net_11348) );
OAI221_X2 inst_1588 ( .B1(net_10310), .B2(net_9047), .C2(net_7287), .C1(net_7108), .ZN(net_7107), .A(net_6928) );
NAND2_X2 inst_3801 ( .ZN(net_4758), .A2(net_4543), .A1(net_2394) );
NAND2_X2 inst_4177 ( .ZN(net_3127), .A1(net_1956), .A2(net_1365) );
AOI22_X2 inst_9350 ( .B1(net_9796), .A1(net_6808), .A2(net_5766), .B2(net_5765), .ZN(net_5602) );
DFF_X2 inst_8002 ( .QN(net_10114), .D(net_5507), .CK(net_12352) );
CLKBUF_X2 inst_14484 ( .A(net_14402), .Z(net_14403) );
CLKBUF_X2 inst_10996 ( .A(net_10914), .Z(net_10915) );
INV_X4 inst_6491 ( .A(net_10389), .ZN(net_357) );
NOR2_X2 inst_2516 ( .A2(net_8317), .ZN(net_8265), .A1(net_8149) );
CLKBUF_X2 inst_13133 ( .A(net_13051), .Z(net_13052) );
AOI22_X2 inst_9193 ( .A1(net_9883), .B1(net_9784), .A2(net_8042), .ZN(net_6121), .B2(net_6120) );
CLKBUF_X2 inst_13901 ( .A(net_12350), .Z(net_13820) );
OAI211_X2 inst_2155 ( .C2(net_6778), .ZN(net_6693), .A(net_6308), .B(net_6052), .C1(net_1577) );
CLKBUF_X2 inst_12927 ( .A(net_11903), .Z(net_12846) );
AOI22_X2 inst_9567 ( .B1(net_10295), .A1(net_10190), .B2(net_4774), .A2(net_4217), .ZN(net_3752) );
INV_X4 inst_6352 ( .A(net_10284), .ZN(net_407) );
OAI221_X2 inst_1506 ( .B2(net_9063), .C2(net_9056), .ZN(net_7355), .B1(net_7198), .A(net_6995), .C1(net_5478) );
CLKBUF_X2 inst_15515 ( .A(net_15433), .Z(net_15434) );
AOI22_X2 inst_9494 ( .B1(net_9819), .A1(net_9688), .A2(net_5966), .ZN(net_3829), .B2(net_2556) );
SDFF_X2 inst_464 ( .SE(net_8812), .SI(net_8650), .CK(net_11911), .Q(x784), .D(x784) );
CLKBUF_X2 inst_13428 ( .A(net_10987), .Z(net_13347) );
INV_X4 inst_5360 ( .A(net_1297), .ZN(net_1222) );
CLKBUF_X2 inst_13392 ( .A(net_13310), .Z(net_13311) );
AND2_X4 inst_10455 ( .A1(net_9242), .ZN(net_2440), .A2(net_1000) );
DFF_X2 inst_7541 ( .QN(net_9356), .D(net_7759), .CK(net_15315) );
INV_X4 inst_6058 ( .A(net_10222), .ZN(net_586) );
XNOR2_X2 inst_341 ( .ZN(net_2868), .B(net_2285), .A(net_219) );
NAND2_X2 inst_3785 ( .A2(net_9591), .A1(net_9082), .ZN(net_4940) );
CLKBUF_X2 inst_15194 ( .A(net_13542), .Z(net_15113) );
CLKBUF_X2 inst_12313 ( .A(net_12231), .Z(net_12232) );
CLKBUF_X2 inst_15800 ( .A(net_14543), .Z(net_15719) );
CLKBUF_X2 inst_14961 ( .A(net_14879), .Z(net_14880) );
CLKBUF_X2 inst_13090 ( .A(net_13008), .Z(net_13009) );
INV_X4 inst_5678 ( .ZN(net_1345), .A(net_808) );
CLKBUF_X2 inst_14006 ( .A(net_13183), .Z(net_13925) );
CLKBUF_X2 inst_11095 ( .A(net_10721), .Z(net_11014) );
NOR4_X2 inst_2359 ( .A4(net_9656), .A3(net_9653), .A2(net_9650), .ZN(net_1261), .A1(net_436) );
NAND2_X2 inst_3702 ( .A2(net_9103), .A1(net_6165), .ZN(net_5934) );
CLKBUF_X2 inst_11229 ( .A(net_11147), .Z(net_11148) );
DFF_X1 inst_8526 ( .Q(net_9973), .D(net_7382), .CK(net_14860) );
CLKBUF_X2 inst_13913 ( .A(net_13831), .Z(net_13832) );
CLKBUF_X2 inst_13031 ( .A(net_12387), .Z(net_12950) );
DFF_X1 inst_8505 ( .Q(net_9288), .D(net_7669), .CK(net_11486) );
DFF_X2 inst_7454 ( .QN(net_9643), .D(net_8191), .CK(net_13146) );
INV_X4 inst_5556 ( .A(net_9172), .ZN(net_3074) );
INV_X2 inst_6826 ( .ZN(net_4181), .A(net_4180) );
OAI222_X2 inst_1361 ( .B1(net_7732), .A2(net_7731), .C2(net_7730), .ZN(net_6921), .B2(net_5945), .A1(net_4313), .C1(net_1833) );
AOI21_X2 inst_10226 ( .ZN(net_2018), .A(net_2017), .B1(net_2016), .B2(net_1318) );
NAND2_X2 inst_3401 ( .A2(net_8932), .A1(net_8614), .ZN(net_8593) );
CLKBUF_X2 inst_13105 ( .A(net_13023), .Z(net_13024) );
CLKBUF_X2 inst_12949 ( .A(net_12867), .Z(net_12868) );
CLKBUF_X2 inst_12688 ( .A(net_12606), .Z(net_12607) );
CLKBUF_X2 inst_12439 ( .A(net_12324), .Z(net_12358) );
CLKBUF_X2 inst_11916 ( .A(net_11834), .Z(net_11835) );
DFF_X2 inst_7525 ( .QN(net_10151), .D(net_7789), .CK(net_12377) );
DFF_X1 inst_8840 ( .Q(net_9760), .D(net_2161), .CK(net_11101) );
INV_X4 inst_4968 ( .ZN(net_2483), .A(net_2130) );
MUX2_X1 inst_4463 ( .S(net_6041), .A(net_283), .B(x5961), .Z(x285) );
OAI211_X2 inst_2208 ( .C1(net_7231), .C2(net_6501), .ZN(net_6497), .B(net_5566), .A(net_3679) );
CLKBUF_X2 inst_14319 ( .A(net_14237), .Z(net_14238) );
INV_X4 inst_5598 ( .ZN(net_3799), .A(net_1961) );
DFF_X1 inst_8789 ( .Q(net_10133), .D(net_4374), .CK(net_10776) );
CLKBUF_X2 inst_10698 ( .A(net_10616), .Z(net_10617) );
AOI21_X2 inst_10122 ( .ZN(net_5155), .A(net_4469), .B1(net_4468), .B2(net_4361) );
NAND2_X2 inst_4162 ( .ZN(net_2912), .A1(net_1978), .A2(net_1975) );
DFF_X2 inst_7873 ( .QN(net_10143), .D(net_6010), .CK(net_13486) );
INV_X4 inst_5171 ( .ZN(net_1917), .A(net_1561) );
CLKBUF_X2 inst_12936 ( .A(net_12854), .Z(net_12855) );
OAI211_X2 inst_2174 ( .C1(net_7226), .C2(net_6548), .ZN(net_6535), .B(net_5663), .A(net_3679) );
INV_X2 inst_6721 ( .ZN(net_7781), .A(net_7751) );
CLKBUF_X2 inst_14363 ( .A(net_12283), .Z(net_14282) );
NAND3_X2 inst_3201 ( .ZN(net_7410), .A3(net_7409), .A2(net_6635), .A1(net_5982) );
CLKBUF_X2 inst_10779 ( .A(net_10697), .Z(net_10698) );
CLKBUF_X2 inst_13089 ( .A(net_11237), .Z(net_13008) );
DFF_X2 inst_7702 ( .Q(net_9906), .D(net_6466), .CK(net_14819) );
XOR2_X2 inst_14 ( .Z(net_2858), .B(net_1580), .A(net_1492) );
AOI22_X2 inst_9366 ( .B1(net_9919), .A2(net_5759), .B2(net_5758), .ZN(net_5556), .A1(net_258) );
DFF_X2 inst_7886 ( .QN(net_10109), .D(net_6030), .CK(net_14804) );
INV_X2 inst_7172 ( .A(net_9588), .ZN(net_545) );
CLKBUF_X2 inst_15774 ( .A(net_15692), .Z(net_15693) );
CLKBUF_X2 inst_15085 ( .A(net_15003), .Z(net_15004) );
CLKBUF_X2 inst_14532 ( .A(net_14410), .Z(net_14451) );
CLKBUF_X2 inst_12068 ( .A(net_11118), .Z(net_11987) );
NOR4_X2 inst_2325 ( .ZN(net_5965), .A1(net_5964), .A2(net_5963), .A4(net_5379), .A3(net_3876) );
CLKBUF_X2 inst_12354 ( .A(net_12272), .Z(net_12273) );
XNOR2_X2 inst_251 ( .ZN(net_4117), .A(net_3958), .B(net_2215) );
CLKBUF_X2 inst_10651 ( .A(net_10569), .Z(net_10570) );
DFF_X2 inst_7983 ( .QN(net_10426), .D(net_5545), .CK(net_14595) );
OAI22_X2 inst_1074 ( .B2(net_10238), .A1(net_10237), .ZN(net_6837), .A2(net_6588), .B1(net_1776) );
DFF_X2 inst_7375 ( .D(net_8678), .QN(net_254), .CK(net_15085) );
AOI21_X2 inst_10149 ( .ZN(net_4195), .A(net_4194), .B1(net_3710), .B2(net_3709) );
OAI221_X2 inst_1552 ( .C2(net_9047), .B2(net_7287), .B1(net_7213), .ZN(net_7206), .A(net_6790), .C1(net_6289) );
OAI221_X2 inst_1524 ( .B1(net_10320), .B2(net_9047), .C1(net_7294), .ZN(net_7288), .C2(net_7287), .A(net_6946) );
CLKBUF_X2 inst_13983 ( .A(net_13901), .Z(net_13902) );
AOI22_X2 inst_9369 ( .B1(net_9917), .A2(net_5759), .B2(net_5758), .ZN(net_5553), .A1(net_256) );
INV_X4 inst_4789 ( .A(net_4332), .ZN(net_3717) );
INV_X4 inst_4977 ( .A(net_3696), .ZN(net_2254) );
CLKBUF_X2 inst_14944 ( .A(net_14862), .Z(net_14863) );
CLKBUF_X2 inst_15481 ( .A(net_15399), .Z(net_15400) );
CLKBUF_X2 inst_11100 ( .A(net_11018), .Z(net_11019) );
AOI221_X2 inst_9892 ( .B1(net_9878), .B2(net_9101), .A(net_6945), .C2(net_6944), .ZN(net_6802), .C1(net_249) );
AOI221_X2 inst_9883 ( .B1(net_9790), .B2(net_9097), .A(net_6940), .C2(net_6939), .ZN(net_6815), .C1(net_260) );
DFF_X2 inst_7781 ( .Q(net_9813), .D(net_6519), .CK(net_13420) );
OAI221_X2 inst_1602 ( .B1(net_10217), .C1(net_7184), .B2(net_5642), .ZN(net_5634), .C2(net_4905), .A(net_3527) );
OAI33_X1 inst_969 ( .ZN(net_3167), .A2(net_3054), .A1(net_2983), .A3(net_2084), .B3(net_1263), .B2(net_1003), .B1(net_928) );
CLKBUF_X2 inst_14569 ( .A(net_14487), .Z(net_14488) );
CLKBUF_X2 inst_15734 ( .A(net_15079), .Z(net_15653) );
DFF_X1 inst_8567 ( .Q(net_9873), .D(net_7172), .CK(net_15566) );
INV_X4 inst_6463 ( .ZN(net_372), .A(net_228) );
CLKBUF_X2 inst_13081 ( .A(net_12999), .Z(net_13000) );
CLKBUF_X2 inst_12487 ( .A(net_10804), .Z(net_12406) );
NOR2_X2 inst_2528 ( .ZN(net_8139), .A2(net_8138), .A1(net_8089) );
AOI221_X2 inst_9749 ( .C1(net_9367), .C2(net_8783), .A(net_7916), .B2(net_7915), .ZN(net_7914), .B1(net_700) );
INV_X4 inst_4917 ( .ZN(net_6415), .A(net_2765) );
CLKBUF_X2 inst_13628 ( .A(net_13546), .Z(net_13547) );
OR2_X2 inst_898 ( .A1(net_10293), .ZN(net_5693), .A2(net_5536) );
INV_X2 inst_7049 ( .A(net_2732), .ZN(net_1335) );
OAI21_X2 inst_1977 ( .ZN(net_2881), .A(net_2880), .B2(net_2527), .B1(net_2224) );
OAI21_X2 inst_1793 ( .B2(net_10347), .A(net_10346), .ZN(net_7480), .B1(net_7479) );
NAND2_X2 inst_4227 ( .A2(net_10473), .ZN(net_2651), .A1(net_1637) );
DFF_X2 inst_8012 ( .QN(net_10334), .D(net_5495), .CK(net_14353) );
INV_X2 inst_6840 ( .ZN(net_3869), .A(net_3603) );
AOI221_X2 inst_9800 ( .B1(net_9979), .A(net_7090), .B2(net_7089), .C2(net_7088), .ZN(net_7004), .C1(net_251) );
AOI22_X2 inst_9223 ( .A1(net_9917), .B1(net_9818), .B2(net_8041), .A2(net_6111), .ZN(net_6088) );
AOI221_X2 inst_9747 ( .C1(net_9364), .C2(net_8783), .ZN(net_7918), .A(net_7916), .B2(net_7915), .B1(net_7632) );
CLKBUF_X2 inst_11804 ( .A(net_11722), .Z(net_11723) );
INV_X4 inst_5299 ( .A(net_6956), .ZN(net_1301) );
CLKBUF_X2 inst_10824 ( .A(net_10742), .Z(net_10743) );
CLKBUF_X2 inst_10805 ( .A(net_10693), .Z(net_10724) );
INV_X4 inst_5697 ( .A(net_2021), .ZN(net_784) );
CLKBUF_X2 inst_12290 ( .A(net_11985), .Z(net_12209) );
OAI211_X2 inst_2291 ( .ZN(net_5184), .C1(net_4671), .B(net_4498), .C2(net_3723), .A(net_3157) );
NOR4_X2 inst_2343 ( .A3(net_5954), .A2(net_3529), .ZN(net_2989), .A1(net_2988), .A4(net_2982) );
DFF_X2 inst_8230 ( .QN(net_10249), .D(net_4924), .CK(net_12189) );
CLKBUF_X2 inst_11500 ( .A(net_10986), .Z(net_11419) );
NOR2_X2 inst_2538 ( .ZN(net_8295), .A2(net_8293), .A1(net_8081) );
INV_X4 inst_5708 ( .A(net_1972), .ZN(net_1059) );
INV_X4 inst_4822 ( .ZN(net_3969), .A(net_3516) );
NAND4_X2 inst_3132 ( .ZN(net_2922), .A1(net_2921), .A2(net_2920), .A4(net_2919), .A3(net_1027) );
CLKBUF_X2 inst_13835 ( .A(net_13753), .Z(net_13754) );
DFF_X2 inst_7395 ( .D(net_8543), .Q(net_223), .CK(net_14621) );
INV_X4 inst_4999 ( .A(net_7584), .ZN(net_3907) );
INV_X4 inst_6071 ( .A(net_9966), .ZN(net_504) );
INV_X4 inst_5819 ( .ZN(net_1108), .A(net_839) );
NAND2_X2 inst_3910 ( .ZN(net_3895), .A1(net_3894), .A2(net_3059) );
CLKBUF_X2 inst_12303 ( .A(net_12221), .Z(net_12222) );
OAI222_X2 inst_1332 ( .B1(net_7823), .A2(net_7811), .ZN(net_7768), .C1(net_3695), .B2(net_3693), .C2(net_3303), .A1(net_3302) );
CLKBUF_X2 inst_12427 ( .A(net_12345), .Z(net_12346) );
OAI21_X2 inst_1841 ( .B1(net_7157), .ZN(net_6213), .B2(net_5779), .A(net_5778) );
CLKBUF_X2 inst_11929 ( .A(net_11401), .Z(net_11848) );
NAND2_X4 inst_3345 ( .A2(net_8880), .A1(net_8879), .ZN(net_8520) );
NAND3_X2 inst_3264 ( .ZN(net_4352), .A3(net_3786), .A2(net_3785), .A1(net_3189) );
CLKBUF_X2 inst_15599 ( .A(net_15517), .Z(net_15518) );
CLKBUF_X2 inst_12584 ( .A(net_11317), .Z(net_12503) );
INV_X4 inst_5169 ( .ZN(net_1876), .A(net_1563) );
INV_X4 inst_4945 ( .ZN(net_2574), .A(net_2573) );
DFF_X1 inst_8782 ( .Q(net_9270), .D(net_4637), .CK(net_15395) );
NOR4_X2 inst_2332 ( .ZN(net_5408), .A2(net_5161), .A4(net_5160), .A3(net_3138), .A1(net_1892) );
CLKBUF_X2 inst_15497 ( .A(net_11972), .Z(net_15416) );
AOI221_X2 inst_9982 ( .C1(net_10177), .B1(net_9750), .B2(net_6442), .C2(net_4217), .ZN(net_4215), .A(net_3577) );
CLKBUF_X2 inst_13415 ( .A(net_13333), .Z(net_13334) );
AOI22_X2 inst_9082 ( .A1(net_9696), .ZN(net_6419), .A2(net_6418), .B2(net_5263), .B1(net_136) );
CLKBUF_X2 inst_13431 ( .A(net_12308), .Z(net_13350) );
CLKBUF_X2 inst_13908 ( .A(net_13826), .Z(net_13827) );
CLKBUF_X2 inst_10970 ( .A(net_10888), .Z(net_10889) );
INV_X4 inst_5946 ( .ZN(net_2450), .A(net_563) );
NOR4_X2 inst_2310 ( .ZN(net_7527), .A4(net_7166), .A1(net_4633), .A2(net_4513), .A3(net_3906) );
AOI222_X1 inst_9720 ( .C1(net_10491), .B1(net_10386), .A1(net_9686), .C2(net_6415), .A2(net_5966), .ZN(net_4063), .B2(net_4062) );
OAI22_X2 inst_1089 ( .B1(net_6847), .ZN(net_6561), .A1(net_6560), .A2(net_6190), .B2(net_6184) );
AOI211_X2 inst_10251 ( .C2(net_9309), .ZN(net_8804), .C1(net_8803), .B(net_8625), .A(net_7903) );
INV_X4 inst_6537 ( .A(net_9169), .ZN(net_648) );
CLKBUF_X2 inst_14327 ( .A(net_14245), .Z(net_14246) );
INV_X4 inst_6430 ( .ZN(net_6040), .A(net_278) );
INV_X4 inst_5017 ( .A(net_6044), .ZN(net_2110) );
INV_X2 inst_6932 ( .A(net_2527), .ZN(net_1941) );
OAI22_X2 inst_1290 ( .B1(net_5090), .A2(net_4274), .ZN(net_3645), .A1(net_3644), .B2(net_3588) );
DFF_X2 inst_7939 ( .QN(net_10441), .D(net_5542), .CK(net_15503) );
CLKBUF_X2 inst_11451 ( .A(net_11272), .Z(net_11370) );
INV_X4 inst_6342 ( .A(net_9828), .ZN(net_649) );
INV_X4 inst_5367 ( .ZN(net_4382), .A(net_2249) );
AOI22_X2 inst_9092 ( .A1(net_9673), .A2(net_6420), .ZN(net_6400), .B2(net_5263), .B1(net_111) );
INV_X4 inst_5845 ( .A(net_3311), .ZN(net_1011) );
INV_X4 inst_5038 ( .ZN(net_1933), .A(net_1932) );
CLKBUF_X2 inst_13399 ( .A(net_11108), .Z(net_13318) );
INV_X4 inst_5142 ( .ZN(net_4283), .A(net_2308) );
INV_X4 inst_5757 ( .ZN(net_730), .A(net_729) );
CLKBUF_X2 inst_12614 ( .A(net_12532), .Z(net_12533) );
INV_X4 inst_4899 ( .A(net_7343), .ZN(net_2856) );
OAI211_X2 inst_2046 ( .C1(net_10344), .ZN(net_7877), .A(net_7876), .B(net_7457), .C2(net_6667) );
CLKBUF_X2 inst_12021 ( .A(net_11930), .Z(net_11940) );
INV_X4 inst_6041 ( .ZN(net_7190), .A(x5901) );
CLKBUF_X2 inst_12604 ( .A(net_12522), .Z(net_12523) );
INV_X4 inst_5079 ( .A(net_6305), .ZN(net_1821) );
NAND2_X2 inst_4129 ( .A2(net_2612), .ZN(net_2248), .A1(net_1939) );
CLKBUF_X2 inst_11632 ( .A(net_11550), .Z(net_11551) );
DFF_X2 inst_7505 ( .Q(net_10404), .D(net_8007), .CK(net_15156) );
INV_X4 inst_6340 ( .A(net_10046), .ZN(net_5084) );
INV_X4 inst_6429 ( .A(net_10465), .ZN(net_571) );
NAND2_X2 inst_3861 ( .ZN(net_4406), .A2(net_4122), .A1(net_2404) );
CLKBUF_X2 inst_15809 ( .A(net_10691), .Z(net_15728) );
NAND2_X2 inst_4399 ( .A2(net_10224), .A1(net_10223), .ZN(net_2211) );
CLKBUF_X2 inst_14176 ( .A(net_14094), .Z(net_14095) );
CLKBUF_X2 inst_11547 ( .A(net_11465), .Z(net_11466) );
AOI221_X2 inst_9847 ( .A(net_6889), .B2(net_6888), .C2(net_6887), .ZN(net_6871), .B1(net_5829), .C1(x5647) );
AOI221_X2 inst_9840 ( .A(net_6889), .B2(net_6888), .C2(net_6887), .ZN(net_6878), .B1(net_5843), .C1(x6028) );
CLKBUF_X2 inst_14835 ( .A(net_14753), .Z(net_14754) );
CLKBUF_X2 inst_14224 ( .A(net_14142), .Z(net_14143) );
CLKBUF_X2 inst_13783 ( .A(net_13701), .Z(net_13702) );
INV_X4 inst_6533 ( .A(net_10470), .ZN(net_748) );
NAND2_X2 inst_4196 ( .A2(net_2673), .ZN(net_1835), .A1(net_1631) );
NAND2_X2 inst_3524 ( .ZN(net_8113), .A2(net_8006), .A1(net_4043) );
CLKBUF_X2 inst_12333 ( .A(net_12203), .Z(net_12252) );
CLKBUF_X2 inst_10672 ( .A(net_10590), .Z(net_10591) );
MUX2_X1 inst_4479 ( .S(net_6041), .B(net_3631), .A(net_792), .Z(x437) );
OAI22_X2 inst_1014 ( .A2(net_8247), .B2(net_8246), .ZN(net_8207), .B1(net_8206), .A1(net_4596) );
NOR2_X2 inst_2531 ( .A2(net_9594), .A1(net_8983), .ZN(net_8315) );
AOI21_X2 inst_10009 ( .B1(net_9579), .B2(net_9578), .ZN(net_8676), .A(net_8675) );
INV_X2 inst_6781 ( .ZN(net_6017), .A(net_5828) );
CLKBUF_X2 inst_14918 ( .A(net_14836), .Z(net_14837) );
CLKBUF_X2 inst_11879 ( .A(net_11797), .Z(net_11798) );
CLKBUF_X2 inst_10882 ( .A(net_10800), .Z(net_10801) );
DFF_X2 inst_7719 ( .Q(net_9807), .D(net_6553), .CK(net_14811) );
CLKBUF_X2 inst_15283 ( .A(net_15201), .Z(net_15202) );
INV_X4 inst_4782 ( .ZN(net_8098), .A(net_7704) );
OAI222_X2 inst_1347 ( .B1(net_7728), .A2(net_7727), .C2(net_7726), .ZN(net_7497), .B2(net_7138), .A1(net_6177), .C1(net_1924) );
CLKBUF_X2 inst_11073 ( .A(net_10991), .Z(net_10992) );
SDFF_X2 inst_509 ( .SI(net_9338), .Q(net_9283), .D(net_9283), .SE(net_7588), .CK(net_14699) );
CLKBUF_X2 inst_12299 ( .A(net_12217), .Z(net_12218) );
NOR2_X2 inst_2687 ( .A2(net_10271), .ZN(net_4549), .A1(net_2249) );
OAI221_X2 inst_1680 ( .B1(net_7203), .C2(net_5591), .ZN(net_5487), .C1(net_5486), .B2(net_4902), .A(net_3731) );
CLKBUF_X2 inst_15221 ( .A(net_14646), .Z(net_15140) );
CLKBUF_X2 inst_11775 ( .A(net_11128), .Z(net_11694) );
CLKBUF_X2 inst_11473 ( .A(net_11391), .Z(net_11392) );
INV_X2 inst_7139 ( .A(net_2419), .ZN(net_822) );
OAI221_X2 inst_1626 ( .B1(net_10323), .C1(net_7182), .A(net_5637), .B2(net_5591), .ZN(net_5581), .C2(net_4902) );
NOR2_X2 inst_2622 ( .ZN(net_6179), .A1(net_5764), .A2(net_1040) );
XNOR2_X2 inst_153 ( .ZN(net_6268), .A(net_5992), .B(net_2549) );
CLKBUF_X2 inst_12834 ( .A(net_12752), .Z(net_12753) );
INV_X4 inst_4856 ( .ZN(net_4299), .A(net_3503) );
AOI221_X2 inst_9751 ( .C1(net_9368), .C2(net_8783), .A(net_7916), .B2(net_7915), .ZN(net_7912), .B1(net_7595) );
CLKBUF_X2 inst_12271 ( .A(net_11795), .Z(net_12190) );
OAI221_X2 inst_1459 ( .C1(net_9075), .B2(net_7974), .C2(net_7973), .ZN(net_7966), .A(net_7965), .B1(net_3001) );
NAND2_X2 inst_4094 ( .ZN(net_2764), .A2(net_2463), .A1(x6157) );
AND2_X2 inst_10483 ( .A2(net_8950), .ZN(net_8583), .A1(net_8397) );
INV_X4 inst_6528 ( .A(net_9376), .ZN(net_7595) );
AOI221_X2 inst_9789 ( .B1(net_9971), .A(net_7090), .B2(net_7089), .C1(net_7088), .ZN(net_7062), .C2(net_243) );
AOI22_X2 inst_9117 ( .A1(net_9671), .A2(net_6420), .ZN(net_6372), .B2(net_5263), .B1(net_109) );
XNOR2_X2 inst_209 ( .ZN(net_4937), .A(net_4395), .B(net_2390) );
NAND2_X2 inst_3894 ( .ZN(net_4000), .A2(net_3965), .A1(net_774) );
INV_X4 inst_6068 ( .A(net_10118), .ZN(net_3496) );
DFF_X2 inst_8037 ( .QN(net_9557), .D(net_9263), .CK(net_12630) );
AOI21_X2 inst_10132 ( .B2(net_10234), .ZN(net_4421), .A(net_1820), .B1(net_1819) );
INV_X4 inst_5385 ( .ZN(net_2873), .A(net_680) );
OAI22_X2 inst_1087 ( .A1(net_6575), .ZN(net_6571), .A2(net_5904), .B2(net_5902), .B1(net_396) );
INV_X4 inst_6365 ( .A(net_9841), .ZN(net_403) );
OAI21_X2 inst_1781 ( .ZN(net_7754), .A(net_7753), .B1(net_7719), .B2(net_7631) );
CLKBUF_X2 inst_13701 ( .A(net_13619), .Z(net_13620) );
NOR2_X2 inst_2769 ( .A1(net_3496), .A2(net_3266), .ZN(net_3265) );
CLKBUF_X2 inst_14453 ( .A(net_14371), .Z(net_14372) );
AOI21_X2 inst_10061 ( .ZN(net_7074), .B1(net_7070), .B2(net_7069), .A(net_6314) );
OAI222_X2 inst_1375 ( .B2(net_7660), .A2(net_7659), .C2(net_7658), .ZN(net_6015), .B1(net_4260), .A1(net_3273), .C1(net_1268) );
CLKBUF_X2 inst_11353 ( .A(net_10701), .Z(net_11272) );
INV_X4 inst_6230 ( .A(net_9537), .ZN(net_462) );
CLKBUF_X2 inst_15797 ( .A(net_15715), .Z(net_15716) );
CLKBUF_X2 inst_12199 ( .A(net_12117), .Z(net_12118) );
CLKBUF_X2 inst_15693 ( .A(net_15611), .Z(net_15612) );
DFF_X2 inst_7966 ( .QN(net_10316), .D(net_5590), .CK(net_15489) );
NAND2_X2 inst_3982 ( .ZN(net_3243), .A2(net_3242), .A1(net_3112) );
INV_X4 inst_4564 ( .ZN(net_8429), .A(net_8251) );
INV_X4 inst_6482 ( .A(net_10472), .ZN(net_3104) );
CLKBUF_X2 inst_15134 ( .A(net_13557), .Z(net_15053) );
CLKBUF_X2 inst_14273 ( .A(net_11274), .Z(net_14192) );
AOI22_X2 inst_9290 ( .B1(net_9803), .A1(net_5766), .B2(net_5765), .ZN(net_5708), .A2(net_241) );
INV_X4 inst_5258 ( .ZN(net_3400), .A(net_1411) );
NAND3_X2 inst_3215 ( .ZN(net_6164), .A2(net_5356), .A1(net_5179), .A3(net_4793) );
CLKBUF_X2 inst_12235 ( .A(net_12153), .Z(net_12154) );
INV_X4 inst_5810 ( .A(net_2284), .ZN(net_682) );
CLKBUF_X2 inst_11209 ( .A(net_11127), .Z(net_11128) );
NOR2_X2 inst_2564 ( .ZN(net_7766), .A2(net_7715), .A1(net_7054) );
DFF_X1 inst_8462 ( .Q(net_9594), .D(net_7964), .CK(net_11539) );
CLKBUF_X2 inst_15173 ( .A(net_15091), .Z(net_15092) );
OAI22_X2 inst_1082 ( .ZN(net_6577), .A1(net_6575), .A2(net_5916), .B2(net_5914), .B1(net_515) );
NAND2_X2 inst_4167 ( .ZN(net_2908), .A1(net_1970), .A2(net_1846) );
CLKBUF_X2 inst_15185 ( .A(net_15103), .Z(net_15104) );
AOI22_X2 inst_9204 ( .A1(net_9864), .B1(net_9765), .B2(net_6120), .A2(net_6111), .ZN(net_6107) );
NOR2_X2 inst_2677 ( .ZN(net_4762), .A2(net_4457), .A1(net_4093) );
NAND2_X2 inst_4374 ( .A1(net_9183), .A2(net_5443), .ZN(net_3016) );
OAI21_X2 inst_1995 ( .ZN(net_3004), .B1(net_2631), .A(net_1802), .B2(net_1338) );
AOI21_X2 inst_10068 ( .B1(net_10175), .ZN(net_6974), .A(net_6679), .B2(net_264) );
XNOR2_X2 inst_105 ( .ZN(net_8170), .A(net_8169), .B(net_6897) );
CLKBUF_X2 inst_15031 ( .A(net_14949), .Z(net_14950) );
AOI22_X2 inst_9145 ( .A1(net_9698), .A2(net_6382), .ZN(net_6340), .B2(net_5263), .B1(net_138) );
NAND2_X2 inst_3518 ( .A2(net_9592), .A1(net_9077), .ZN(net_8150) );
OAI211_X2 inst_2161 ( .C1(net_7297), .ZN(net_6553), .C2(net_6542), .B(net_5772), .A(net_3679) );
DFF_X2 inst_8294 ( .Q(net_9852), .D(net_4614), .CK(net_14580) );
SDFF_X2 inst_625 ( .Q(net_9453), .D(net_9453), .SE(net_3293), .CK(net_12453), .SI(x2333) );
DFF_X2 inst_7405 ( .QN(net_9250), .D(net_8322), .CK(net_14771) );
CLKBUF_X2 inst_12736 ( .A(net_12654), .Z(net_12655) );
NAND2_X4 inst_3367 ( .ZN(net_6319), .A1(net_4025), .A2(net_3898) );
INV_X2 inst_6747 ( .ZN(net_6968), .A(net_6681) );
CLKBUF_X2 inst_14041 ( .A(net_13959), .Z(net_13960) );
SDFF_X2 inst_568 ( .D(net_9135), .SE(net_933), .CK(net_10974), .SI(x2278), .Q(x1215) );
CLKBUF_X2 inst_15445 ( .A(net_14903), .Z(net_15364) );
OAI221_X2 inst_1483 ( .ZN(net_7558), .C2(net_7557), .B1(net_7115), .B2(net_7113), .A(net_3991), .C1(net_3700) );
SDFF_X2 inst_523 ( .Q(net_9340), .D(net_9340), .SI(net_9332), .SE(net_7588), .CK(net_14683) );
DFF_X2 inst_8119 ( .Q(net_9737), .D(net_5149), .CK(net_14299) );
AOI21_X2 inst_10202 ( .ZN(net_2717), .B1(net_2716), .B2(net_2705), .A(net_1361) );
OAI221_X2 inst_1492 ( .B1(net_10426), .C2(net_9063), .B2(net_9056), .ZN(net_7371), .C1(net_7186), .A(net_7009) );
XNOR2_X2 inst_181 ( .ZN(net_5246), .A(net_4690), .B(net_2326) );
CLKBUF_X2 inst_13212 ( .A(net_13130), .Z(net_13131) );
DFF_X2 inst_8329 ( .QN(net_10480), .D(net_3227), .CK(net_11433) );
INV_X4 inst_5215 ( .A(net_2131), .ZN(net_1520) );
NAND2_X2 inst_4234 ( .ZN(net_2684), .A2(net_981), .A1(net_900) );
INV_X2 inst_6722 ( .ZN(net_7780), .A(net_7750) );
CLKBUF_X2 inst_11982 ( .A(net_11900), .Z(net_11901) );
CLKBUF_X2 inst_10885 ( .A(net_10803), .Z(net_10804) );
AOI222_X1 inst_9738 ( .B2(net_10402), .C2(net_10400), .A2(net_10399), .B1(net_10389), .C1(net_10387), .A1(net_10386), .ZN(net_1187) );
OR3_X2 inst_713 ( .ZN(net_4689), .A1(net_4409), .A3(net_4408), .A2(net_3136) );
AOI21_X2 inst_10125 ( .B1(net_4713), .ZN(net_4321), .A(net_4320), .B2(net_4319) );
NOR2_X2 inst_2898 ( .A2(net_6658), .ZN(net_1667), .A1(net_798) );
INV_X2 inst_6918 ( .A(net_2532), .ZN(net_2136) );
AOI211_X2 inst_10280 ( .A(net_9115), .ZN(net_6265), .C2(net_5998), .B(net_4727), .C1(net_1554) );
DFF_X1 inst_8875 ( .D(net_10518), .CK(net_12652), .Q(x454) );
CLKBUF_X2 inst_11508 ( .A(net_11426), .Z(net_11427) );
OAI222_X2 inst_1368 ( .B2(net_7660), .A2(net_7659), .C2(net_7658), .ZN(net_6282), .B1(net_5210), .A1(net_3675), .C1(net_1907) );
CLKBUF_X2 inst_13708 ( .A(net_10580), .Z(net_13627) );
CLKBUF_X2 inst_15665 ( .A(net_15583), .Z(net_15584) );
INV_X2 inst_7282 ( .A(net_8975), .ZN(net_8971) );
CLKBUF_X2 inst_15256 ( .A(net_14480), .Z(net_15175) );
CLKBUF_X2 inst_15199 ( .A(net_15117), .Z(net_15118) );
INV_X2 inst_6775 ( .ZN(net_6023), .A(net_5840) );
OAI211_X2 inst_2088 ( .C2(net_6774), .ZN(net_6760), .A(net_6387), .B(net_6121), .C1(net_510) );
DFF_X2 inst_7768 ( .Q(net_9718), .D(net_6536), .CK(net_13428) );
CLKBUF_X2 inst_14062 ( .A(net_11999), .Z(net_13981) );
NAND3_X2 inst_3208 ( .A3(net_9649), .ZN(net_7519), .A1(net_7060), .A2(net_797) );
DFF_X2 inst_7410 ( .QN(net_9402), .D(net_8363), .CK(net_14023) );
INV_X2 inst_6673 ( .ZN(net_8355), .A(net_8292) );
NAND2_X2 inst_4134 ( .A1(net_3289), .ZN(net_2245), .A2(net_2244) );
NAND2_X2 inst_3507 ( .ZN(net_8239), .A2(net_8129), .A1(net_356) );
OAI222_X2 inst_1379 ( .B2(net_7660), .A2(net_7659), .C2(net_7658), .ZN(net_6006), .B1(net_4259), .A1(net_3276), .C1(net_1226) );
XNOR2_X2 inst_271 ( .ZN(net_3956), .B(net_3955), .A(net_3224) );
CLKBUF_X2 inst_11918 ( .A(net_11836), .Z(net_11837) );
CLKBUF_X2 inst_12326 ( .A(net_12244), .Z(net_12245) );
AOI22_X2 inst_9582 ( .B1(net_9981), .A2(net_5173), .ZN(net_3581), .B2(net_2541), .A1(net_215) );
INV_X2 inst_6705 ( .A(net_8320), .ZN(net_8263) );
OAI22_X2 inst_1230 ( .B1(net_7198), .A2(net_4890), .B2(net_4889), .ZN(net_4887), .A1(net_380) );
CLKBUF_X2 inst_15739 ( .A(net_15657), .Z(net_15658) );
CLKBUF_X2 inst_10844 ( .A(net_10762), .Z(net_10763) );
DFF_X2 inst_7691 ( .Q(net_10297), .D(net_6574), .CK(net_14554) );
INV_X2 inst_7262 ( .A(net_9639), .ZN(net_652) );
NAND2_X2 inst_3535 ( .ZN(net_9002), .A1(net_8954), .A2(net_8047) );
CLKBUF_X2 inst_12217 ( .A(net_12135), .Z(net_12136) );
AOI22_X2 inst_9344 ( .B1(net_9820), .A2(net_5766), .B2(net_5765), .ZN(net_5608), .A1(net_258) );
CLKBUF_X2 inst_15582 ( .A(net_14710), .Z(net_15501) );
AOI22_X2 inst_9221 ( .A1(net_9915), .B1(net_9816), .B2(net_8041), .A2(net_6141), .ZN(net_6090) );
CLKBUF_X2 inst_14685 ( .A(net_14603), .Z(net_14604) );
NAND2_X2 inst_3497 ( .A1(net_9547), .ZN(net_8387), .A2(net_8131) );
INV_X4 inst_6131 ( .ZN(net_4910), .A(net_272) );
OAI22_X2 inst_1064 ( .A2(net_7036), .B2(net_7035), .ZN(net_6965), .A1(net_1536), .B1(net_1534) );
INV_X4 inst_5416 ( .ZN(net_1594), .A(net_1148) );
CLKBUF_X2 inst_14875 ( .A(net_10580), .Z(net_14794) );
CLKBUF_X2 inst_13643 ( .A(net_13561), .Z(net_13562) );
CLKBUF_X2 inst_14229 ( .A(net_14147), .Z(net_14148) );
CLKBUF_X2 inst_11110 ( .A(net_11028), .Z(net_11029) );
INV_X4 inst_5796 ( .ZN(net_1960), .A(net_690) );
NAND2_X2 inst_3599 ( .ZN(net_7267), .A2(net_6859), .A1(net_6606) );
CLKBUF_X2 inst_14335 ( .A(net_14253), .Z(net_14254) );
CLKBUF_X2 inst_14539 ( .A(net_11047), .Z(net_14458) );
CLKBUF_X2 inst_14924 ( .A(net_14842), .Z(net_14843) );
CLKBUF_X2 inst_14654 ( .A(net_14572), .Z(net_14573) );
AOI22_X2 inst_9571 ( .B2(net_6442), .A2(net_5173), .ZN(net_3737), .B1(net_3736), .A1(net_2521) );
CLKBUF_X2 inst_13727 ( .A(net_13645), .Z(net_13646) );
SDFF_X2 inst_583 ( .Q(net_9252), .SE(net_4589), .D(net_135), .SI(net_101), .CK(net_13846) );
CLKBUF_X2 inst_12124 ( .A(net_12042), .Z(net_12043) );
OAI21_X2 inst_1904 ( .B1(net_7221), .B2(net_4862), .ZN(net_4848), .A(net_4520) );
CLKBUF_X2 inst_13970 ( .A(net_13888), .Z(net_13889) );
INV_X4 inst_5208 ( .ZN(net_2631), .A(net_1184) );
NAND2_X2 inst_3581 ( .ZN(net_7548), .A2(net_7118), .A1(net_2430) );
CLKBUF_X2 inst_10732 ( .A(net_10650), .Z(net_10651) );
AOI221_X2 inst_9930 ( .B2(net_5867), .A(net_5862), .ZN(net_5844), .C1(net_5843), .C2(net_4725), .B1(x6028) );
CLKBUF_X2 inst_14146 ( .A(net_14064), .Z(net_14065) );
CLKBUF_X2 inst_10932 ( .A(net_10699), .Z(net_10851) );
NAND2_X2 inst_4325 ( .ZN(net_5272), .A1(net_174), .A2(net_173) );
AND2_X4 inst_10441 ( .A2(net_3062), .ZN(net_2077), .A1(net_2076) );
INV_X4 inst_4833 ( .ZN(net_7514), .A(net_3373) );
OAI211_X2 inst_2065 ( .C2(net_7757), .ZN(net_7708), .B(net_7569), .A(net_7135), .C1(net_6847) );
CLKBUF_X2 inst_10765 ( .A(net_10673), .Z(net_10684) );
OAI211_X2 inst_2251 ( .C1(net_7234), .C2(net_6548), .ZN(net_6440), .B(net_5440), .A(net_3679) );
NAND2_X2 inst_3987 ( .A1(net_9772), .ZN(net_3189), .A2(net_2462) );
INV_X2 inst_6913 ( .A(net_3908), .ZN(net_2191) );
CLKBUF_X2 inst_12825 ( .A(net_11373), .Z(net_12744) );
CLKBUF_X2 inst_13720 ( .A(net_13638), .Z(net_13639) );
INV_X2 inst_6788 ( .A(net_9263), .ZN(net_6242) );
INV_X4 inst_5124 ( .ZN(net_1824), .A(net_1601) );
CLKBUF_X2 inst_14346 ( .A(net_13313), .Z(net_14265) );
DFF_X2 inst_7709 ( .Q(net_9903), .D(net_6309), .CK(net_12578) );
CLKBUF_X2 inst_13226 ( .A(net_13144), .Z(net_13145) );
INV_X4 inst_4863 ( .ZN(net_6442), .A(net_3942) );
CLKBUF_X2 inst_12513 ( .A(net_12431), .Z(net_12432) );
INV_X4 inst_4910 ( .A(net_3015), .ZN(net_2837) );
OAI21_X2 inst_1899 ( .B1(net_7184), .B2(net_4862), .ZN(net_4853), .A(net_4525) );
CLKBUF_X2 inst_14667 ( .A(net_14585), .Z(net_14586) );
INV_X2 inst_7200 ( .A(net_9393), .ZN(net_8213) );
AOI22_X2 inst_9349 ( .B1(net_9824), .A2(net_5766), .B2(net_5765), .ZN(net_5603), .A1(net_262) );
CLKBUF_X2 inst_14985 ( .A(net_14903), .Z(net_14904) );
CLKBUF_X2 inst_12113 ( .A(net_12031), .Z(net_12032) );
NOR2_X2 inst_2569 ( .A2(net_9542), .A1(net_9531), .ZN(net_7488) );
AND2_X2 inst_10573 ( .ZN(net_2968), .A1(net_2967), .A2(net_2966) );
AOI221_X2 inst_9811 ( .B1(net_9989), .A(net_7090), .B2(net_7089), .C2(net_7088), .ZN(net_6991), .C1(net_6811) );
AOI21_X2 inst_10197 ( .ZN(net_2939), .B1(net_2938), .A(net_2499), .B2(net_2201) );
AOI22_X2 inst_9048 ( .B1(net_9667), .A1(net_6684), .B2(net_6683), .ZN(net_6676), .A2(net_236) );
CLKBUF_X2 inst_14504 ( .A(net_10709), .Z(net_14423) );
NOR2_X2 inst_2716 ( .A2(net_10375), .A1(net_5983), .ZN(net_5214) );
DFF_X1 inst_8693 ( .D(net_6770), .Q(net_114), .CK(net_12592) );
INV_X4 inst_6025 ( .A(net_9926), .ZN(net_582) );
NAND3_X2 inst_3228 ( .A3(net_10091), .A2(net_8511), .A1(net_7832), .ZN(net_5734) );
AOI22_X2 inst_9212 ( .A1(net_9904), .B1(net_9805), .B2(net_6129), .A2(net_6109), .ZN(net_6099) );
OAI211_X2 inst_2124 ( .C2(net_6774), .ZN(net_6724), .A(net_6351), .B(net_6086), .C1(net_427) );
CLKBUF_X2 inst_13268 ( .A(net_12889), .Z(net_13187) );
OAI211_X2 inst_2289 ( .ZN(net_5750), .C2(net_4668), .A(net_3493), .C1(net_2436), .B(net_1844) );
OAI222_X1 inst_1435 ( .ZN(net_7842), .A2(net_7735), .A1(net_7732), .B2(net_7731), .C2(net_7730), .B1(net_6162), .C1(net_1400) );
CLKBUF_X2 inst_11582 ( .A(net_11142), .Z(net_11501) );
NAND2_X2 inst_3746 ( .ZN(net_5304), .A2(net_4767), .A1(net_4051) );
CLKBUF_X2 inst_15610 ( .A(net_15528), .Z(net_15529) );
CLKBUF_X2 inst_12288 ( .A(net_10913), .Z(net_12207) );
NOR2_X2 inst_2750 ( .ZN(net_4143), .A1(net_3685), .A2(x3733) );
CLKBUF_X2 inst_10810 ( .A(net_10728), .Z(net_10729) );
NAND2_X2 inst_4121 ( .ZN(net_2336), .A2(net_1611), .A1(net_1550) );
INV_X4 inst_5800 ( .A(net_1344), .ZN(net_870) );
OAI221_X2 inst_1467 ( .ZN(net_7881), .A(net_7878), .C2(net_7162), .B2(net_7027), .B1(net_5933), .C1(net_5276) );
NOR2_X2 inst_2640 ( .A1(net_9354), .ZN(net_6854), .A2(net_5391) );
CLKBUF_X2 inst_14313 ( .A(net_13405), .Z(net_14232) );
AOI211_X2 inst_10258 ( .ZN(net_8059), .A(net_7928), .B(net_7919), .C1(net_7887), .C2(net_6564) );
INV_X4 inst_5772 ( .ZN(net_1071), .A(net_717) );
CLKBUF_X2 inst_12732 ( .A(net_10746), .Z(net_12651) );
DFF_X2 inst_8162 ( .QN(net_9832), .D(net_5058), .CK(net_11734) );
DFF_X2 inst_7908 ( .QN(net_10250), .D(net_5819), .CK(net_11662) );
CLKBUF_X2 inst_10803 ( .A(net_10721), .Z(net_10722) );
MUX2_X1 inst_4448 ( .S(net_6041), .A(net_298), .B(x5003), .Z(x121) );
CLKBUF_X2 inst_14102 ( .A(net_10569), .Z(net_14021) );
CLKBUF_X2 inst_13227 ( .A(net_13145), .Z(net_13146) );
INV_X4 inst_6317 ( .A(net_9829), .ZN(net_1015) );
NOR2_X2 inst_2834 ( .A1(net_3487), .ZN(net_2379), .A2(net_2378) );
CLKBUF_X2 inst_15067 ( .A(net_10993), .Z(net_14986) );
INV_X4 inst_4784 ( .A(net_10490), .ZN(net_5362) );
CLKBUF_X2 inst_15155 ( .A(net_15073), .Z(net_15074) );
DFF_X2 inst_8130 ( .Q(net_9841), .D(net_5128), .CK(net_12018) );
INV_X2 inst_7207 ( .A(net_9658), .ZN(net_464) );
CLKBUF_X2 inst_12256 ( .A(net_12174), .Z(net_12175) );
OAI221_X2 inst_1513 ( .C1(net_10423), .B2(net_9063), .C2(net_9056), .ZN(net_7347), .B1(net_7211), .A(net_7019) );
AOI221_X2 inst_9864 ( .B1(net_9774), .B2(net_9097), .A(net_6940), .C1(net_6939), .ZN(net_6852), .C2(net_244) );
CLKBUF_X2 inst_11756 ( .A(net_10826), .Z(net_11675) );
CLKBUF_X2 inst_14716 ( .A(net_12075), .Z(net_14635) );
CLKBUF_X2 inst_10916 ( .A(net_10701), .Z(net_10835) );
NAND2_X4 inst_3321 ( .A2(net_8901), .A1(net_8900), .ZN(net_8701) );
NAND2_X2 inst_4080 ( .A1(net_9531), .ZN(net_7343), .A2(net_2610) );
CLKBUF_X2 inst_10846 ( .A(net_10648), .Z(net_10765) );
DFF_X2 inst_7667 ( .D(net_6762), .QN(net_121), .CK(net_12804) );
CLKBUF_X2 inst_12750 ( .A(net_12668), .Z(net_12669) );
OAI221_X2 inst_1545 ( .B2(net_9047), .C2(net_7287), .ZN(net_7217), .C1(net_7216), .A(net_6791), .B1(net_870) );
XNOR2_X2 inst_333 ( .ZN(net_2981), .A(net_2385), .B(net_2142) );
NAND2_X4 inst_3338 ( .A2(net_8904), .A1(net_8903), .ZN(net_8528) );
DFF_X2 inst_7684 ( .Q(net_10067), .D(net_6569), .CK(net_10837) );
INV_X4 inst_5988 ( .A(net_9524), .ZN(net_539) );
DFF_X2 inst_8368 ( .QN(net_8840), .D(net_2003), .CK(net_11428) );
INV_X4 inst_5279 ( .ZN(net_1328), .A(net_593) );
XNOR2_X2 inst_406 ( .A(net_9305), .ZN(net_2728), .B(net_193) );
CLKBUF_X2 inst_14696 ( .A(net_12314), .Z(net_14615) );
CLKBUF_X2 inst_11934 ( .A(net_11831), .Z(net_11853) );
INV_X4 inst_5933 ( .ZN(net_2122), .A(net_572) );
INV_X4 inst_4579 ( .ZN(net_8071), .A(net_8031) );
CLKBUF_X2 inst_13818 ( .A(net_13736), .Z(net_13737) );
XNOR2_X2 inst_328 ( .ZN(net_3006), .B(net_2805), .A(net_2055) );
CLKBUF_X2 inst_11394 ( .A(net_10960), .Z(net_11313) );
AOI22_X2 inst_9335 ( .B1(net_9811), .A2(net_5766), .B2(net_5765), .ZN(net_5617), .A1(net_249) );
CLKBUF_X2 inst_10953 ( .A(net_10871), .Z(net_10872) );
CLKBUF_X2 inst_10897 ( .A(net_10815), .Z(net_10816) );
NAND2_X2 inst_4217 ( .A1(net_8687), .ZN(net_1677), .A2(net_116) );
NOR2_X2 inst_2764 ( .ZN(net_4046), .A1(net_3363), .A2(net_3191) );
DFF_X1 inst_8496 ( .Q(net_9758), .D(net_7839), .CK(net_15185) );
OR2_X4 inst_818 ( .A2(net_10159), .A1(net_9735), .ZN(net_2208) );
CLKBUF_X2 inst_12373 ( .A(net_12291), .Z(net_12292) );
INV_X4 inst_6246 ( .A(net_10120), .ZN(net_3988) );
CLKBUF_X2 inst_13755 ( .A(net_13673), .Z(net_13674) );
CLKBUF_X2 inst_11065 ( .A(net_10860), .Z(net_10984) );
INV_X4 inst_6155 ( .A(net_9323), .ZN(net_1123) );
INV_X4 inst_5774 ( .A(net_840), .ZN(net_818) );
AOI22_X2 inst_9664 ( .B2(net_10404), .A2(net_10403), .B1(net_10390), .A1(net_10389), .ZN(net_972) );
DFF_X1 inst_8719 ( .QN(net_10346), .D(net_6290), .CK(net_10643) );
AOI221_X2 inst_9902 ( .B1(net_9887), .B2(net_9101), .A(net_6945), .C2(net_6944), .ZN(net_6792), .C1(net_258) );
CLKBUF_X2 inst_11610 ( .A(net_11528), .Z(net_11529) );
AOI221_X2 inst_9825 ( .B1(net_9773), .B2(net_9097), .A(net_6940), .C1(net_6939), .ZN(net_6924), .C2(net_243) );
DFF_X2 inst_7561 ( .QN(net_10464), .D(net_7627), .CK(net_11406) );
AOI21_X2 inst_10172 ( .ZN(net_3639), .A(net_3638), .B2(net_3019), .B1(net_2489) );
NAND3_X2 inst_3178 ( .ZN(net_8174), .A1(net_8053), .A3(net_7975), .A2(net_3730) );
NAND3_X2 inst_3274 ( .A3(net_10243), .ZN(net_4140), .A1(net_4139), .A2(net_904) );
CLKBUF_X2 inst_13920 ( .A(net_12445), .Z(net_13839) );
NAND2_X2 inst_4203 ( .A1(net_10353), .A2(net_2051), .ZN(net_1780) );
CLKBUF_X2 inst_11776 ( .A(net_11694), .Z(net_11695) );
CLKBUF_X2 inst_12643 ( .A(net_12561), .Z(net_12562) );
AOI221_X2 inst_9972 ( .ZN(net_4672), .C1(net_4671), .A(net_4240), .B1(net_4239), .B2(net_3358), .C2(net_2959) );
NOR2_X2 inst_2840 ( .ZN(net_2333), .A2(net_2332), .A1(net_1618) );
CLKBUF_X2 inst_12521 ( .A(net_12102), .Z(net_12440) );
CLKBUF_X2 inst_10939 ( .A(net_10724), .Z(net_10858) );
AOI22_X2 inst_9178 ( .A1(net_9906), .B1(net_9807), .B2(net_8041), .A2(net_6141), .ZN(net_6138) );
AOI21_X2 inst_10066 ( .ZN(net_6784), .A(net_6188), .B1(net_5955), .B2(net_5952) );
CLKBUF_X2 inst_14214 ( .A(net_14132), .Z(net_14133) );
DFF_X2 inst_8360 ( .QN(net_9232), .D(net_2112), .CK(net_13540) );
NOR2_X2 inst_2781 ( .A1(net_9613), .ZN(net_3144), .A2(net_1041) );
CLKBUF_X2 inst_15622 ( .A(net_13753), .Z(net_15541) );
AOI22_X2 inst_9544 ( .B1(net_9812), .A1(net_9681), .A2(net_5966), .ZN(net_3777), .B2(net_2556) );
INV_X4 inst_6442 ( .A(net_9573), .ZN(net_5283) );
CLKBUF_X2 inst_13190 ( .A(net_13108), .Z(net_13109) );
INV_X2 inst_7146 ( .ZN(net_792), .A(net_791) );
OR2_X2 inst_906 ( .A1(net_9526), .ZN(net_4968), .A2(net_4550) );
NAND2_X2 inst_4276 ( .A2(net_10335), .ZN(net_2186), .A1(net_1351) );
INV_X4 inst_5222 ( .ZN(net_6044), .A(net_1957) );
CLKBUF_X2 inst_13600 ( .A(net_11129), .Z(net_13519) );
INV_X4 inst_5098 ( .ZN(net_1695), .A(net_1694) );
CLKBUF_X2 inst_11043 ( .A(net_10961), .Z(net_10962) );
OAI22_X2 inst_1248 ( .B1(net_7224), .ZN(net_4828), .A2(net_4826), .B2(net_4825), .A1(net_537) );
NOR2_X2 inst_2598 ( .ZN(net_7557), .A2(net_7505), .A1(net_1716) );
CLKBUF_X2 inst_12780 ( .A(net_12698), .Z(net_12699) );
NOR3_X2 inst_2402 ( .A3(net_9379), .A2(net_9378), .ZN(net_7501), .A1(net_345) );
DFF_X1 inst_8877 ( .D(net_10198), .QN(net_10138), .CK(net_10857) );
NOR2_X2 inst_2616 ( .A1(net_9087), .ZN(net_7050), .A2(net_6230) );
CLKBUF_X2 inst_14627 ( .A(net_14545), .Z(net_14546) );
DFF_X2 inst_8095 ( .D(net_4983), .QN(net_166), .CK(net_13192) );
NAND2_X2 inst_3998 ( .ZN(net_7439), .A2(net_3390), .A1(net_3171) );
AOI22_X2 inst_9035 ( .ZN(net_7556), .A2(net_7386), .A1(net_7015), .B2(net_6205), .B1(net_5392) );
NAND2_X2 inst_4300 ( .A2(net_10158), .A1(net_3988), .ZN(net_2355) );
OAI211_X2 inst_2113 ( .C2(net_6778), .ZN(net_6735), .A(net_6363), .B(net_6095), .C1(net_488) );
CLKBUF_X2 inst_12000 ( .A(net_11918), .Z(net_11919) );
DFF_X2 inst_7645 ( .D(net_6724), .QN(net_161), .CK(net_13441) );
INV_X4 inst_5249 ( .ZN(net_1449), .A(net_1448) );
OAI21_X2 inst_1820 ( .ZN(net_6632), .A(net_6631), .B1(net_6414), .B2(net_5969) );
CLKBUF_X2 inst_15674 ( .A(net_15592), .Z(net_15593) );
XNOR2_X2 inst_183 ( .ZN(net_5212), .A(net_4579), .B(net_2080) );
DFF_X2 inst_8253 ( .Q(net_10183), .D(net_4834), .CK(net_12949) );
INV_X2 inst_6998 ( .A(net_2305), .ZN(net_2178) );
DFF_X2 inst_7748 ( .QN(net_10146), .D(net_6282), .CK(net_13504) );
INV_X2 inst_6703 ( .ZN(net_8151), .A(net_8150) );
DFF_X1 inst_8471 ( .Q(net_9529), .D(net_7925), .CK(net_15032) );
CLKBUF_X2 inst_15822 ( .A(net_15740), .Z(net_15741) );
INV_X4 inst_6065 ( .A(net_9293), .ZN(net_1843) );
INV_X4 inst_4729 ( .A(net_7730), .ZN(net_4595) );
OAI211_X2 inst_2271 ( .C1(net_7139), .C2(net_6480), .ZN(net_6271), .B(net_5692), .A(net_3679) );
INV_X4 inst_6209 ( .A(net_10190), .ZN(net_466) );
DFF_X2 inst_7793 ( .Q(net_9892), .D(net_6502), .CK(net_13202) );
AOI211_X2 inst_10314 ( .C2(net_10332), .ZN(net_2421), .B(net_1720), .A(net_1434), .C1(net_762) );
DFF_X2 inst_8081 ( .QN(net_10529), .D(net_5355), .CK(net_14790) );
NAND2_X2 inst_3779 ( .A2(net_8986), .ZN(net_4993), .A1(net_174) );
OAI21_X2 inst_1848 ( .B1(net_7823), .ZN(net_5890), .B2(net_5889), .A(net_5350) );
CLKBUF_X2 inst_12694 ( .A(net_12612), .Z(net_12613) );
MUX2_X1 inst_4451 ( .S(net_6041), .A(net_295), .B(x5225), .Z(x143) );
CLKBUF_X2 inst_11644 ( .A(net_11162), .Z(net_11563) );
OR3_X4 inst_697 ( .ZN(net_7731), .A3(net_4444), .A2(net_4441), .A1(net_1493) );
CLKBUF_X2 inst_11150 ( .A(net_11068), .Z(net_11069) );
CLKBUF_X2 inst_14035 ( .A(net_13953), .Z(net_13954) );
SDFF_X2 inst_487 ( .SE(net_9540), .SI(net_8222), .Q(net_301), .D(net_301), .CK(net_13908) );
INV_X4 inst_5159 ( .ZN(net_1851), .A(net_1576) );
CLKBUF_X2 inst_14540 ( .A(net_14458), .Z(net_14459) );
CLKBUF_X2 inst_11338 ( .A(net_10550), .Z(net_11257) );
AND4_X2 inst_10350 ( .ZN(net_977), .A4(net_150), .A1(net_148), .A2(net_136), .A3(net_135) );
DFF_X2 inst_7527 ( .QN(net_9312), .D(net_7791), .CK(net_15330) );
CLKBUF_X2 inst_13941 ( .A(net_13859), .Z(net_13860) );
INV_X4 inst_5315 ( .ZN(net_1482), .A(net_1282) );
CLKBUF_X2 inst_11512 ( .A(net_11430), .Z(net_11431) );
CLKBUF_X2 inst_13696 ( .A(net_10838), .Z(net_13615) );
OAI211_X2 inst_2133 ( .C2(net_6778), .ZN(net_6715), .A(net_6405), .B(net_6078), .C1(net_517) );
OAI211_X2 inst_2163 ( .C1(net_7186), .ZN(net_6549), .C2(net_6548), .A(net_6546), .B(net_5674) );
CLKBUF_X2 inst_12307 ( .A(net_11954), .Z(net_12226) );
AOI221_X2 inst_9947 ( .C2(net_10339), .B1(net_10338), .ZN(net_5275), .A(net_4592), .B2(net_4420), .C1(net_4281) );
INV_X4 inst_6051 ( .A(net_9320), .ZN(net_590) );
INV_X4 inst_4668 ( .ZN(net_5961), .A(net_5247) );
DFF_X1 inst_8758 ( .QN(net_9602), .D(net_5387), .CK(net_15175) );
CLKBUF_X2 inst_12975 ( .A(net_12382), .Z(net_12894) );
INV_X4 inst_5497 ( .ZN(net_7002), .A(net_991) );
CLKBUF_X2 inst_14853 ( .A(net_11506), .Z(net_14772) );
CLKBUF_X2 inst_13972 ( .A(net_13890), .Z(net_13891) );
OAI21_X2 inst_1861 ( .ZN(net_5509), .A(net_5143), .B2(net_4844), .B1(net_593) );
CLKBUF_X2 inst_15165 ( .A(net_15083), .Z(net_15084) );
NAND2_X2 inst_3570 ( .A1(net_8801), .ZN(net_8627), .A2(net_8614) );
AOI22_X2 inst_9133 ( .A1(net_9717), .A2(net_6420), .ZN(net_6355), .B2(net_5263), .B1(net_1056) );
CLKBUF_X2 inst_14198 ( .A(net_14116), .Z(net_14117) );
DFF_X2 inst_7598 ( .QN(net_10358), .D(net_7432), .CK(net_12223) );
INV_X4 inst_4835 ( .ZN(net_4326), .A(net_3649) );
CLKBUF_X2 inst_15050 ( .A(net_10936), .Z(net_14969) );
OAI21_X2 inst_2004 ( .ZN(net_2804), .A(net_2145), .B1(net_2144), .B2(net_1658) );
DFF_X1 inst_8667 ( .D(net_6771), .Q(net_113), .CK(net_12601) );
NOR2_X2 inst_2857 ( .A2(net_9660), .A1(net_9659), .ZN(net_2107) );
CLKBUF_X2 inst_15116 ( .A(net_15034), .Z(net_15035) );
XNOR2_X2 inst_220 ( .ZN(net_4602), .B(net_4601), .A(net_4449) );
OAI221_X2 inst_1585 ( .B1(net_10314), .B2(net_9047), .C2(net_7287), .C1(net_7129), .ZN(net_7120), .A(net_6915) );
CLKBUF_X2 inst_11412 ( .A(net_11120), .Z(net_11331) );
CLKBUF_X2 inst_10754 ( .A(net_10672), .Z(net_10673) );
XNOR2_X2 inst_245 ( .B(net_9657), .ZN(net_4161), .A(net_3651) );
INV_X2 inst_6991 ( .A(net_2755), .ZN(net_1642) );
CLKBUF_X2 inst_11965 ( .A(net_11292), .Z(net_11884) );
AOI221_X2 inst_9779 ( .C1(net_9347), .B1(net_9156), .ZN(net_7158), .A(net_7157), .B2(net_7155), .C2(net_7154) );
OAI21_X2 inst_1873 ( .ZN(net_5289), .A(net_5288), .B2(net_4364), .B1(x4587) );
CLKBUF_X2 inst_15584 ( .A(net_15502), .Z(net_15503) );
NAND2_X2 inst_4111 ( .ZN(net_2361), .A2(net_1695), .A1(net_1186) );
DFF_X2 inst_8388 ( .Q(net_10408), .D(net_857), .CK(net_13109) );
DFF_X1 inst_8768 ( .Q(net_9269), .D(net_4909), .CK(net_15398) );
DFF_X2 inst_7854 ( .Q(net_9657), .D(net_6246), .CK(net_11815) );
XNOR2_X2 inst_147 ( .ZN(net_7026), .B(net_7025), .A(net_6170) );
INV_X4 inst_6135 ( .ZN(net_6816), .A(net_259) );
XNOR2_X2 inst_313 ( .ZN(net_3222), .B(net_3005), .A(net_2266) );
OAI221_X2 inst_1676 ( .C1(net_7198), .B2(net_5591), .ZN(net_5492), .B1(net_5491), .C2(net_4902), .A(net_3507) );
NAND2_X2 inst_4170 ( .A2(net_9735), .ZN(net_2749), .A1(net_1966) );
CLKBUF_X2 inst_11765 ( .A(net_11683), .Z(net_11684) );
DFF_X1 inst_8480 ( .Q(net_9631), .D(net_7950), .CK(net_15025) );
OAI22_X2 inst_1041 ( .B2(net_8918), .A2(net_8917), .A1(net_8117), .ZN(net_7893), .B1(net_2562) );
INV_X4 inst_5263 ( .ZN(net_4230), .A(net_2972) );
OAI211_X2 inst_2086 ( .C2(net_6778), .ZN(net_6762), .A(net_6389), .B(net_6123), .C1(net_439) );
NAND4_X2 inst_3114 ( .ZN(net_4563), .A2(net_4264), .A4(net_4253), .A1(net_4110), .A3(net_2768) );
NAND2_X2 inst_3577 ( .ZN(net_7610), .A2(net_7403), .A1(net_2432) );
AOI22_X2 inst_9451 ( .A1(net_10524), .B2(net_6442), .A2(net_4056), .ZN(net_4038), .B1(net_4037) );
CLKBUF_X2 inst_15035 ( .A(net_14953), .Z(net_14954) );
CLKBUF_X2 inst_12918 ( .A(net_12514), .Z(net_12837) );
DFF_X1 inst_8743 ( .Q(net_9149), .D(net_5681), .CK(net_11033) );
DFF_X1 inst_8570 ( .Q(net_9776), .D(net_7296), .CK(net_15636) );
DFF_X2 inst_8195 ( .Q(net_10023), .D(net_5108), .CK(net_14713) );
CLKBUF_X2 inst_12789 ( .A(net_12707), .Z(net_12708) );
INV_X4 inst_4754 ( .ZN(net_4455), .A(net_4353) );
SDFF_X2 inst_553 ( .SI(net_9357), .Q(net_9357), .D(net_9155), .SE(net_7248), .CK(net_15263) );
AOI22_X2 inst_9271 ( .B1(net_9907), .ZN(net_5760), .A1(net_5759), .B2(net_5758), .A2(net_246) );
AOI21_X2 inst_10216 ( .ZN(net_2307), .B2(net_2306), .B1(net_2132), .A(net_1948) );
NAND2_X4 inst_3331 ( .ZN(net_8939), .A1(net_8563), .A2(net_8562) );
CLKBUF_X2 inst_11554 ( .A(net_11472), .Z(net_11473) );
XNOR2_X2 inst_242 ( .ZN(net_4164), .A(net_3999), .B(net_204) );
INV_X4 inst_6589 ( .A(net_9216), .ZN(net_5719) );
INV_X4 inst_4680 ( .ZN(net_5002), .A(net_4744) );
CLKBUF_X2 inst_14592 ( .A(net_14510), .Z(net_14511) );
CLKBUF_X2 inst_14759 ( .A(net_11944), .Z(net_14678) );
OAI22_X2 inst_1186 ( .A1(net_7294), .A2(net_5134), .B2(net_5133), .ZN(net_5069), .B1(net_1943) );
OAI21_X2 inst_1753 ( .ZN(net_8631), .A(net_8603), .B2(net_8571), .B1(net_8551) );
OAI21_X2 inst_1727 ( .B2(net_9567), .ZN(net_8794), .A(net_8793), .B1(net_5256) );
AOI22_X2 inst_9513 ( .B1(net_10403), .A1(net_9864), .B2(net_4062), .ZN(net_3810), .A2(net_2973) );
AND2_X2 inst_10542 ( .ZN(net_3854), .A2(net_3502), .A1(net_1444) );
OAI22_X2 inst_1166 ( .A1(net_7234), .A2(net_5107), .B2(net_5105), .ZN(net_5104), .B1(net_5103) );
OAI21_X2 inst_1739 ( .ZN(net_8713), .B2(net_8698), .A(net_8598), .B1(net_8249) );
XNOR2_X2 inst_116 ( .ZN(net_7843), .A(net_7767), .B(net_7051) );
CLKBUF_X2 inst_15183 ( .A(net_15101), .Z(net_15102) );
CLKBUF_X2 inst_13712 ( .A(net_13630), .Z(net_13631) );
INV_X4 inst_6559 ( .A(net_10499), .ZN(net_329) );
INV_X4 inst_5498 ( .A(net_2607), .ZN(net_988) );
AOI21_X2 inst_10142 ( .ZN(net_4243), .A(net_4076), .B2(net_3619), .B1(net_3055) );
CLKBUF_X2 inst_14863 ( .A(net_14781), .Z(net_14782) );
CLKBUF_X2 inst_12430 ( .A(net_12348), .Z(net_12349) );
SDFF_X2 inst_471 ( .D(net_9578), .SI(net_3037), .SE(net_758), .Q(net_252), .CK(net_15049) );
NAND2_X2 inst_4087 ( .A2(net_3602), .ZN(net_3558), .A1(net_2554) );
CLKBUF_X2 inst_10680 ( .A(net_10598), .Z(net_10599) );
INV_X4 inst_5446 ( .A(net_1141), .ZN(net_1091) );
CLKBUF_X2 inst_12104 ( .A(net_12022), .Z(net_12023) );
INV_X4 inst_6557 ( .A(net_10012), .ZN(net_330) );
INV_X4 inst_4956 ( .A(net_4717), .ZN(net_4376) );
CLKBUF_X2 inst_11081 ( .A(net_10999), .Z(net_11000) );
NAND2_X2 inst_3609 ( .ZN(net_7257), .A2(net_6862), .A1(net_6595) );
OR2_X2 inst_896 ( .A1(net_10293), .ZN(net_5771), .A2(net_5770) );
DFF_X1 inst_8619 ( .Q(net_9664), .D(net_7116), .CK(net_13281) );
CLKBUF_X2 inst_12315 ( .A(net_10680), .Z(net_12234) );
INV_X4 inst_6649 ( .A(net_9540), .ZN(net_9114) );
CLKBUF_X2 inst_13338 ( .A(net_13256), .Z(net_13257) );
CLKBUF_X2 inst_14552 ( .A(net_14470), .Z(net_14471) );
AOI22_X2 inst_9276 ( .B1(net_9799), .A1(net_5766), .B2(net_5765), .ZN(net_5751), .A2(net_237) );
DFF_X2 inst_8221 ( .Q(net_10079), .D(net_4856), .CK(net_10746) );
NOR2_X2 inst_2608 ( .A2(net_6253), .ZN(net_6249), .A1(net_5810) );
INV_X4 inst_6008 ( .ZN(net_528), .A(x747) );
CLKBUF_X2 inst_15021 ( .A(net_14939), .Z(net_14940) );
AOI22_X2 inst_9317 ( .B1(net_9722), .A1(net_6816), .A2(net_5755), .B2(net_5754), .ZN(net_5660) );
CLKBUF_X2 inst_11840 ( .A(net_11200), .Z(net_11759) );
DFF_X2 inst_7445 ( .QN(net_9296), .D(net_8201), .CK(net_15005) );
CLKBUF_X2 inst_12659 ( .A(net_10864), .Z(net_12578) );
DFF_X1 inst_8577 ( .Q(net_9872), .D(net_7123), .CK(net_14830) );
CLKBUF_X2 inst_14766 ( .A(net_14684), .Z(net_14685) );
DFF_X2 inst_7438 ( .QN(net_9409), .D(net_8355), .CK(net_13924) );
NOR2_X2 inst_2557 ( .ZN(net_7819), .A2(net_7736), .A1(net_3351) );
NOR2_X2 inst_2521 ( .A1(net_9271), .ZN(net_8377), .A2(net_8203) );
XNOR2_X2 inst_385 ( .ZN(net_2277), .A(net_2276), .B(net_2275) );
CLKBUF_X2 inst_15639 ( .A(net_10700), .Z(net_15558) );
CLKBUF_X2 inst_15718 ( .A(net_14556), .Z(net_15637) );
NAND2_X4 inst_3319 ( .A1(net_8987), .ZN(net_8728), .A2(net_8237) );
CLKBUF_X2 inst_14110 ( .A(net_13080), .Z(net_14029) );
NOR2_X2 inst_2653 ( .ZN(net_5279), .A2(net_5278), .A1(net_472) );
CLKBUF_X2 inst_11062 ( .A(net_10618), .Z(net_10981) );
CLKBUF_X2 inst_14827 ( .A(net_14745), .Z(net_14746) );
INV_X4 inst_4621 ( .ZN(net_7132), .A(net_7012) );
CLKBUF_X2 inst_11519 ( .A(net_11102), .Z(net_11438) );
CLKBUF_X2 inst_11324 ( .A(net_10906), .Z(net_11243) );
NOR2_X2 inst_2550 ( .A1(net_9513), .ZN(net_8046), .A2(net_7986) );
CLKBUF_X2 inst_15799 ( .A(net_15717), .Z(net_15718) );
CLKBUF_X2 inst_14966 ( .A(net_14884), .Z(net_14885) );
CLKBUF_X2 inst_10696 ( .A(net_10598), .Z(net_10615) );
CLKBUF_X2 inst_13150 ( .A(net_13068), .Z(net_13069) );
DFF_X2 inst_7559 ( .QN(net_10255), .D(net_7606), .CK(net_11689) );
NAND2_X2 inst_4281 ( .ZN(net_2673), .A1(net_1344), .A2(net_813) );
SDFF_X2 inst_596 ( .Q(net_9260), .SE(net_4589), .D(net_143), .SI(net_109), .CK(net_13824) );
NOR2_X2 inst_2771 ( .ZN(net_3235), .A2(net_3234), .A1(net_2646) );
DFF_X1 inst_8835 ( .Q(net_9759), .D(net_2423), .CK(net_10810) );
INV_X4 inst_4687 ( .ZN(net_4840), .A(net_4658) );
OAI211_X2 inst_2142 ( .C2(net_6774), .ZN(net_6706), .A(net_6333), .C1(net_6148), .B(net_6069) );
AOI22_X2 inst_9245 ( .A1(net_9951), .B1(net_9852), .A2(net_6141), .B2(net_6140), .ZN(net_6066) );
CLKBUF_X2 inst_12810 ( .A(net_12728), .Z(net_12729) );
OAI221_X2 inst_1705 ( .ZN(net_4644), .B1(net_4642), .A(net_4359), .B2(net_2918), .C2(net_2917), .C1(net_1055) );
CLKBUF_X2 inst_11286 ( .A(net_11204), .Z(net_11205) );
INV_X4 inst_5110 ( .ZN(net_3024), .A(net_1662) );
INV_X4 inst_4664 ( .ZN(net_5589), .A(net_5588) );
CLKBUF_X2 inst_14601 ( .A(net_13800), .Z(net_14520) );
INV_X2 inst_6817 ( .A(net_9161), .ZN(net_4706) );
INV_X4 inst_5003 ( .ZN(net_2581), .A(net_1515) );
MUX2_X1 inst_4458 ( .S(net_6041), .A(net_288), .B(x5647), .Z(x233) );
CLKBUF_X2 inst_12215 ( .A(net_10827), .Z(net_12134) );
AOI22_X2 inst_9407 ( .B1(net_9175), .ZN(net_4803), .A2(net_4802), .B2(net_4801), .A1(net_2087) );
CLKBUF_X2 inst_15454 ( .A(net_13518), .Z(net_15373) );
INV_X4 inst_5798 ( .A(net_1970), .ZN(net_1007) );
NAND3_X2 inst_3253 ( .ZN(net_4943), .A1(net_4553), .A3(net_4552), .A2(net_2952) );
INV_X4 inst_5321 ( .ZN(net_4247), .A(net_1275) );
CLKBUF_X2 inst_14250 ( .A(net_12935), .Z(net_14169) );
CLKBUF_X2 inst_14055 ( .A(net_13973), .Z(net_13974) );
AND2_X2 inst_10518 ( .ZN(net_4708), .A1(net_4446), .A2(net_4445) );
INV_X4 inst_5184 ( .ZN(net_4723), .A(net_1000) );
INV_X4 inst_4596 ( .ZN(net_7900), .A(net_7825) );
AOI22_X2 inst_9013 ( .A2(net_8030), .B2(net_8029), .ZN(net_8023), .B1(net_7495), .A1(net_216) );
DFF_X1 inst_8427 ( .Q(net_9584), .D(net_8718), .CK(net_13812) );
CLKBUF_X2 inst_15767 ( .A(net_14173), .Z(net_15686) );
SDFF_X2 inst_637 ( .Q(net_9465), .D(net_9465), .SE(net_3293), .CK(net_11891), .SI(x1598) );
SDFF_X2 inst_547 ( .D(net_9126), .SE(net_933), .CK(net_10597), .SI(x2826), .Q(x1298) );
AOI22_X2 inst_9107 ( .A1(net_9688), .A2(net_6402), .ZN(net_6385), .B2(net_5263), .B1(net_4024) );
CLKBUF_X2 inst_13572 ( .A(net_13490), .Z(net_13491) );
OAI221_X2 inst_1607 ( .C1(net_10203), .B1(net_7190), .C2(net_5642), .ZN(net_5629), .B2(net_4905), .A(net_3507) );
CLKBUF_X2 inst_13148 ( .A(net_13066), .Z(net_13067) );
CLKBUF_X2 inst_11847 ( .A(net_11765), .Z(net_11766) );
INV_X2 inst_7033 ( .ZN(net_4373), .A(net_1442) );
CLKBUF_X2 inst_15787 ( .A(net_13566), .Z(net_15706) );
DFF_X2 inst_8152 ( .QN(net_9949), .D(net_5078), .CK(net_13710) );
AOI21_X2 inst_10159 ( .ZN(net_4010), .A(net_4009), .B2(net_3341), .B1(net_1127) );
AND3_X2 inst_10367 ( .A2(net_9538), .A1(net_5353), .A3(net_5351), .ZN(net_5349) );
INV_X4 inst_4762 ( .ZN(net_4225), .A(net_4090) );
XNOR2_X2 inst_164 ( .B(net_6040), .ZN(net_5948), .A(net_5373) );
CLKBUF_X2 inst_11623 ( .A(net_11541), .Z(net_11542) );
DFF_X1 inst_8534 ( .Q(net_9964), .D(net_7313), .CK(net_15751) );
AOI22_X2 inst_9002 ( .ZN(net_8386), .B1(net_8238), .A1(net_8238), .B2(net_8237), .A2(net_8110) );
OAI21_X2 inst_1854 ( .ZN(net_5874), .B1(net_5873), .B2(net_5872), .A(net_5291) );
CLKBUF_X2 inst_12676 ( .A(net_12594), .Z(net_12595) );
INV_X4 inst_5922 ( .ZN(net_947), .A(net_584) );
OAI221_X2 inst_1710 ( .C2(net_4274), .ZN(net_3946), .B1(net_3945), .C1(net_3944), .B2(net_3942), .A(net_3506) );
INV_X2 inst_7295 ( .A(net_9046), .ZN(net_9045) );
NOR3_X2 inst_2407 ( .ZN(net_7474), .A2(net_7110), .A3(net_7094), .A1(net_3044) );
CLKBUF_X2 inst_13814 ( .A(net_11801), .Z(net_13733) );
DFF_X1 inst_8467 ( .Q(net_9597), .D(net_7958), .CK(net_11524) );
INV_X4 inst_4884 ( .ZN(net_4378), .A(net_2974) );
DFF_X2 inst_7516 ( .Q(net_9534), .D(net_7923), .CK(net_13993) );
NAND4_X2 inst_3142 ( .ZN(net_2508), .A3(net_1458), .A4(net_1451), .A1(net_1421), .A2(net_1068) );
NOR4_X2 inst_2305 ( .A1(net_8963), .A2(net_8960), .ZN(net_7983), .A3(net_7841), .A4(net_7598) );
OR2_X4 inst_753 ( .ZN(net_5138), .A1(net_4475), .A2(net_4473) );
AOI21_X2 inst_10079 ( .B1(net_9528), .ZN(net_5801), .A(net_5800), .B2(net_5258) );
AOI22_X2 inst_9647 ( .B2(net_2641), .ZN(net_2572), .A1(net_2571), .A2(net_1944), .B1(net_1512) );
OAI211_X2 inst_2150 ( .C2(net_6778), .ZN(net_6698), .A(net_6312), .B(net_6058), .C1(net_5061) );
INV_X4 inst_5486 ( .ZN(net_1411), .A(net_998) );
NAND2_X2 inst_3427 ( .A2(net_9470), .ZN(net_8884), .A1(net_8482) );
CLKBUF_X2 inst_10930 ( .A(net_10848), .Z(net_10849) );
INV_X4 inst_6262 ( .A(net_10121), .ZN(net_1233) );
INV_X4 inst_5768 ( .ZN(net_984), .A(net_722) );
AOI221_X2 inst_9770 ( .C2(net_7586), .B2(net_7584), .ZN(net_7513), .C1(net_7512), .B1(net_7512), .A(net_7164) );
INV_X2 inst_6946 ( .ZN(net_1903), .A(net_1345) );
OAI33_X1 inst_946 ( .B2(net_9638), .A2(net_9638), .A3(net_9612), .B3(net_9279), .ZN(net_7837), .A1(net_7808), .B1(net_7562) );
OAI21_X2 inst_1954 ( .ZN(net_3716), .A(net_3664), .B2(net_3485), .B1(net_938) );
OAI211_X2 inst_2260 ( .C1(net_7234), .C2(net_6501), .ZN(net_6309), .B(net_5422), .A(net_3679) );
DFF_X2 inst_8141 ( .QN(net_9941), .D(net_5154), .CK(net_12879) );
CLKBUF_X2 inst_13276 ( .A(net_13194), .Z(net_13195) );
NAND2_X2 inst_3941 ( .A1(net_9919), .A2(net_4969), .ZN(net_3549) );
CLKBUF_X2 inst_13543 ( .A(net_13350), .Z(net_13462) );
DFF_X2 inst_7815 ( .Q(net_10019), .D(net_6465), .CK(net_11963) );
CLKBUF_X2 inst_12746 ( .A(net_12513), .Z(net_12665) );
AND2_X2 inst_10588 ( .A2(net_4267), .A1(net_2422), .ZN(net_2391) );
INV_X2 inst_7014 ( .ZN(net_1575), .A(net_1574) );
NAND2_X2 inst_3858 ( .A2(net_5168), .ZN(net_4176), .A1(net_4175) );
CLKBUF_X2 inst_13129 ( .A(net_11914), .Z(net_13048) );
CLKBUF_X2 inst_11700 ( .A(net_11299), .Z(net_11619) );
INV_X4 inst_4625 ( .ZN(net_7459), .A(net_6920) );
INV_X2 inst_6951 ( .A(net_3708), .ZN(net_1890) );
NAND2_X2 inst_3922 ( .A2(net_9055), .ZN(net_7961), .A1(net_377) );
OAI211_X2 inst_2053 ( .C1(net_10449), .ZN(net_7798), .A(net_7797), .B(net_7306), .C2(net_6043) );
CLKBUF_X2 inst_13949 ( .A(net_12759), .Z(net_13868) );
AND2_X2 inst_10539 ( .A1(net_9656), .ZN(net_3651), .A2(net_3650) );
AOI21_X2 inst_10038 ( .ZN(net_7696), .A(net_7630), .B2(net_7629), .B1(net_438) );
OAI22_X2 inst_1325 ( .B2(net_2265), .A2(net_1761), .ZN(net_1757), .A1(net_1756), .B1(net_1755) );
DFF_X1 inst_8859 ( .D(net_3464), .CK(net_11196), .Q(x871) );
CLKBUF_X2 inst_13503 ( .A(net_13421), .Z(net_13422) );
CLKBUF_X2 inst_13008 ( .A(net_12926), .Z(net_12927) );
INV_X2 inst_6873 ( .ZN(net_3001), .A(net_3000) );
CLKBUF_X2 inst_14087 ( .A(net_14005), .Z(net_14006) );
HA_X1 inst_7342 ( .S(net_5243), .CO(net_5242), .B(net_4431), .A(net_913) );
DFF_X1 inst_8818 ( .QN(net_10339), .D(net_3254), .CK(net_10695) );
INV_X4 inst_5105 ( .ZN(net_4266), .A(net_1686) );
NAND3_X2 inst_3312 ( .ZN(net_1707), .A1(net_1706), .A3(net_1502), .A2(net_187) );
CLKBUF_X2 inst_15432 ( .A(net_12431), .Z(net_15351) );
AOI22_X2 inst_9207 ( .A1(net_9867), .B1(net_9768), .B2(net_6133), .A2(net_6111), .ZN(net_6104) );
CLKBUF_X2 inst_12725 ( .A(net_12643), .Z(net_12644) );
CLKBUF_X2 inst_12143 ( .A(net_11129), .Z(net_12062) );
OAI22_X2 inst_1235 ( .B1(net_7182), .A2(net_4890), .B2(net_4889), .ZN(net_4882), .A1(net_329) );
NAND2_X2 inst_3561 ( .ZN(net_7741), .A1(net_7700), .A2(net_7699) );
CLKBUF_X2 inst_15015 ( .A(net_10901), .Z(net_14934) );
CLKBUF_X2 inst_14107 ( .A(net_14025), .Z(net_14026) );
INV_X2 inst_7233 ( .ZN(net_3541), .A(x3653) );
CLKBUF_X2 inst_14286 ( .A(net_14204), .Z(net_14205) );
CLKBUF_X2 inst_13143 ( .A(net_11476), .Z(net_13062) );
NAND4_X2 inst_3046 ( .ZN(net_7407), .A2(net_7072), .A4(net_7071), .A3(net_6260), .A1(net_2747) );
DFF_X1 inst_8751 ( .Q(net_9128), .D(net_5304), .CK(net_10944) );
NAND2_X2 inst_3626 ( .ZN(net_7099), .A1(net_6884), .A2(net_6642) );
NAND2_X2 inst_4036 ( .A2(net_9198), .ZN(net_3593), .A1(net_2501) );
INV_X4 inst_4644 ( .ZN(net_6024), .A(net_5842) );
INV_X4 inst_5244 ( .ZN(net_1466), .A(net_1396) );
CLKBUF_X2 inst_14994 ( .A(net_14912), .Z(net_14913) );
INV_X4 inst_4844 ( .A(net_3482), .ZN(net_3314) );
NAND2_X2 inst_3757 ( .A1(net_6039), .ZN(net_5250), .A2(net_5233) );
OR2_X2 inst_917 ( .ZN(net_3677), .A2(net_3266), .A1(net_3062) );
NAND2_X2 inst_3712 ( .ZN(net_5909), .A1(net_5908), .A2(net_5907) );
CLKBUF_X2 inst_14942 ( .A(net_13262), .Z(net_14861) );
CLKBUF_X2 inst_13457 ( .A(net_13375), .Z(net_13376) );
OAI21_X2 inst_1743 ( .B1(net_8691), .ZN(net_8690), .B2(net_8671), .A(net_7852) );
CLKBUF_X2 inst_11713 ( .A(net_11631), .Z(net_11632) );
CLKBUF_X2 inst_13403 ( .A(net_13321), .Z(net_13322) );
OAI221_X2 inst_1600 ( .B1(net_10215), .C1(net_7294), .B2(net_5642), .ZN(net_5636), .C2(net_4905), .A(net_3731) );
INV_X4 inst_5022 ( .ZN(net_2291), .A(net_1981) );
XNOR2_X2 inst_215 ( .ZN(net_4684), .A(net_4272), .B(net_2360) );
NOR2_X2 inst_2850 ( .A2(net_5175), .ZN(net_3350), .A1(net_2255) );
CLKBUF_X2 inst_14884 ( .A(net_14802), .Z(net_14803) );
CLKBUF_X2 inst_14268 ( .A(net_12579), .Z(net_14187) );
INV_X4 inst_5163 ( .ZN(net_2491), .A(net_1571) );
NOR2_X2 inst_2624 ( .A1(net_9270), .A2(net_6581), .ZN(net_6153) );
AOI22_X2 inst_9590 ( .B1(net_10079), .B2(net_5319), .A2(net_5173), .ZN(net_3570), .A1(net_204) );
DFF_X2 inst_7677 ( .QN(net_10475), .D(net_6953), .CK(net_11399) );
OR2_X2 inst_849 ( .ZN(net_8584), .A2(net_8583), .A1(net_8430) );
DFF_X2 inst_7393 ( .D(net_8567), .QN(net_233), .CK(net_14334) );
INV_X4 inst_6258 ( .A(net_9945), .ZN(net_452) );
DFF_X2 inst_7550 ( .QN(net_9243), .D(net_7703), .CK(net_11347) );
XOR2_X2 inst_3 ( .Z(net_6515), .B(net_6514), .A(net_5598) );
CLKBUF_X2 inst_14517 ( .A(net_14435), .Z(net_14436) );
CLKBUF_X2 inst_11293 ( .A(net_11211), .Z(net_11212) );
NAND4_X2 inst_3060 ( .ZN(net_5726), .A4(net_4776), .A3(net_4219), .A2(net_3860), .A1(net_3404) );
INV_X4 inst_5812 ( .A(net_2792), .ZN(net_1074) );
AOI21_X2 inst_10041 ( .B2(net_9503), .ZN(net_7811), .A(net_7619), .B1(net_7618) );
SDFF_X2 inst_566 ( .D(net_9123), .SE(net_933), .CK(net_10904), .SI(x3022), .Q(x1343) );
OAI222_X2 inst_1399 ( .B2(net_7728), .A2(net_7727), .C2(net_7726), .ZN(net_5340), .B1(net_2976), .A1(net_2864), .C1(net_1931) );
CLKBUF_X2 inst_12301 ( .A(net_12219), .Z(net_12220) );
AND2_X2 inst_10613 ( .A2(net_4109), .ZN(net_1771), .A1(net_1770) );
NAND2_X2 inst_4357 ( .A2(net_10436), .ZN(net_2437), .A1(net_963) );
INV_X4 inst_4819 ( .ZN(net_5862), .A(net_3678) );
CLKBUF_X2 inst_15437 ( .A(net_15355), .Z(net_15356) );
NAND2_X2 inst_4327 ( .A2(net_10350), .ZN(net_1571), .A1(net_582) );
CLKBUF_X2 inst_12997 ( .A(net_12915), .Z(net_12916) );
CLKBUF_X2 inst_11375 ( .A(net_11293), .Z(net_11294) );
INV_X4 inst_4774 ( .ZN(net_4470), .A(net_4361) );
DFF_X1 inst_8622 ( .Q(net_9780), .D(net_7205), .CK(net_13462) );
AND2_X4 inst_10419 ( .ZN(net_4396), .A2(net_4255), .A1(net_4114) );
NOR4_X2 inst_2333 ( .ZN(net_4960), .A2(net_4959), .A4(net_4958), .A3(net_4389), .A1(net_3350) );
CLKBUF_X2 inst_14844 ( .A(net_12579), .Z(net_14763) );
CLKBUF_X2 inst_12401 ( .A(net_12319), .Z(net_12320) );
CLKBUF_X2 inst_15291 ( .A(net_12329), .Z(net_15210) );
CLKBUF_X2 inst_14632 ( .A(net_11438), .Z(net_14551) );
INV_X2 inst_7047 ( .A(net_2455), .ZN(net_1341) );
CLKBUF_X2 inst_11345 ( .A(net_10845), .Z(net_11264) );
INV_X4 inst_5928 ( .ZN(net_2275), .A(net_775) );
INV_X4 inst_5056 ( .A(net_3289), .ZN(net_2240) );
NAND2_X2 inst_4016 ( .A1(net_9533), .A2(net_3084), .ZN(net_3077) );
INV_X4 inst_5370 ( .A(net_3736), .ZN(net_1558) );
OAI21_X2 inst_1732 ( .ZN(net_8757), .A(net_8756), .B1(net_8740), .B2(net_8735) );
NOR2_X2 inst_2914 ( .A2(net_2824), .ZN(net_1494), .A1(net_1493) );
DFF_X2 inst_7648 ( .D(net_6710), .QN(net_167), .CK(net_12820) );
NAND3_X2 inst_3294 ( .A1(net_3630), .ZN(net_2745), .A3(net_2744), .A2(net_222) );
INV_X2 inst_7256 ( .A(net_9312), .ZN(net_326) );
NOR2_X2 inst_2741 ( .ZN(net_3688), .A1(net_3687), .A2(net_3686) );
CLKBUF_X2 inst_15262 ( .A(net_15180), .Z(net_15181) );
CLKBUF_X2 inst_11825 ( .A(net_11685), .Z(net_11744) );
CLKBUF_X2 inst_11966 ( .A(net_11884), .Z(net_11885) );
INV_X4 inst_6119 ( .A(net_9733), .ZN(net_1213) );
CLKBUF_X2 inst_14380 ( .A(net_10765), .Z(net_14299) );
OAI221_X2 inst_1522 ( .B1(net_10215), .ZN(net_7296), .B2(net_7295), .C1(net_7294), .C2(net_7293), .A(net_6955) );
CLKBUF_X2 inst_15461 ( .A(net_15379), .Z(net_15380) );
CLKBUF_X2 inst_12135 ( .A(net_11130), .Z(net_12054) );
CLKBUF_X2 inst_11455 ( .A(net_10899), .Z(net_11374) );
INV_X4 inst_6269 ( .ZN(net_7108), .A(x5790) );
CLKBUF_X2 inst_13955 ( .A(net_13873), .Z(net_13874) );
CLKBUF_X2 inst_13247 ( .A(net_11891), .Z(net_13166) );
AOI22_X2 inst_9481 ( .A1(net_10187), .B1(net_9814), .A2(net_4217), .ZN(net_3842), .B2(net_2556) );
INV_X4 inst_5858 ( .ZN(net_1190), .A(net_1035) );
NAND4_X2 inst_3069 ( .ZN(net_5444), .A2(net_4712), .A4(net_4450), .A3(net_3592), .A1(net_3391) );
DFF_X1 inst_8645 ( .Q(net_9889), .D(net_7206), .CK(net_13349) );
NAND2_X2 inst_3631 ( .ZN(net_7003), .A1(net_7002), .A2(net_6565) );
INV_X4 inst_5761 ( .ZN(net_948), .A(net_726) );
INV_X2 inst_6964 ( .A(net_3706), .ZN(net_1837) );
CLKBUF_X2 inst_12809 ( .A(net_12727), .Z(net_12728) );
CLKBUF_X2 inst_12520 ( .A(net_12438), .Z(net_12439) );
OAI22_X2 inst_1101 ( .B2(net_10448), .A1(net_10447), .ZN(net_6211), .A2(net_5961), .B1(net_1777) );
DFF_X1 inst_8596 ( .Q(net_9682), .D(net_7265), .CK(net_15255) );
AOI22_X2 inst_9528 ( .B1(net_9968), .A2(net_6442), .ZN(net_3793), .B2(net_2541), .A1(net_1747) );
INV_X2 inst_6652 ( .ZN(net_8748), .A(net_8744) );
NOR2_X2 inst_2950 ( .A1(net_10351), .ZN(net_1552), .A2(net_1212) );
CLKBUF_X2 inst_11889 ( .A(net_11807), .Z(net_11808) );
DFF_X1 inst_8584 ( .Q(net_9670), .D(net_7233), .CK(net_11626) );
DFF_X2 inst_7902 ( .QN(net_10153), .D(net_6007), .CK(net_13479) );
INV_X4 inst_5691 ( .A(net_7562), .ZN(net_1280) );
CLKBUF_X2 inst_15777 ( .A(net_15695), .Z(net_15696) );
DFF_X2 inst_8392 ( .Q(net_10514), .D(net_10513), .CK(net_11420) );
OR2_X2 inst_861 ( .A1(net_10188), .ZN(net_7868), .A2(net_7867) );
CLKBUF_X2 inst_11549 ( .A(net_10555), .Z(net_11468) );
DFF_X2 inst_7431 ( .QN(net_9411), .D(net_8354), .CK(net_13931) );
CLKBUF_X2 inst_12013 ( .A(net_10781), .Z(net_11932) );
NOR2_X2 inst_2990 ( .A1(net_1728), .ZN(net_1181), .A2(x6496) );
DFF_X2 inst_7495 ( .D(net_7985), .Q(net_203), .CK(net_12515) );
OAI22_X2 inst_1283 ( .A1(net_4456), .ZN(net_4093), .A2(net_4092), .B1(net_3916), .B2(net_3262) );
CLKBUF_X2 inst_15572 ( .A(net_15490), .Z(net_15491) );
NOR3_X2 inst_2451 ( .ZN(net_2416), .A3(net_2375), .A1(net_1703), .A2(net_1474) );
CLKBUF_X2 inst_11225 ( .A(net_10699), .Z(net_11144) );
CLKBUF_X2 inst_10625 ( .A(x3675), .Z(net_10544) );
OAI22_X2 inst_1202 ( .A1(net_7124), .A2(net_5151), .B2(net_5150), .ZN(net_5049), .B1(net_3352) );
NAND2_X2 inst_4290 ( .A2(net_10124), .A1(net_7331), .ZN(net_1302) );
CLKBUF_X2 inst_15106 ( .A(net_15024), .Z(net_15025) );
INV_X2 inst_7020 ( .ZN(net_1532), .A(net_1531) );
OAI211_X2 inst_2227 ( .C1(net_7231), .C2(net_6480), .ZN(net_6477), .B(net_5676), .A(net_3679) );
CLKBUF_X2 inst_12594 ( .A(net_11844), .Z(net_12513) );
SDFF_X2 inst_660 ( .SI(net_9497), .Q(net_9497), .SE(net_3073), .CK(net_12411), .D(x1598) );
NOR2_X2 inst_2490 ( .ZN(net_8709), .A1(net_8708), .A2(net_8539) );
CLKBUF_X2 inst_15104 ( .A(net_11447), .Z(net_15023) );
CLKBUF_X2 inst_11027 ( .A(net_10697), .Z(net_10946) );
AOI21_X2 inst_10238 ( .ZN(net_8850), .A(net_8724), .B1(net_8693), .B2(net_8667) );
CLKBUF_X2 inst_14526 ( .A(net_10909), .Z(net_14445) );
CLKBUF_X2 inst_14701 ( .A(net_14619), .Z(net_14620) );
AOI21_X2 inst_10150 ( .B1(net_9523), .A(net_4268), .ZN(net_4191), .B2(net_3727) );
INV_X4 inst_5195 ( .ZN(net_1861), .A(net_1541) );
OAI221_X2 inst_1576 ( .B2(net_7437), .C2(net_7167), .ZN(net_7166), .A(net_4716), .B1(net_2852), .C1(net_1515) );
CLKBUF_X2 inst_11532 ( .A(net_11450), .Z(net_11451) );
NAND2_X2 inst_3462 ( .A1(net_9499), .ZN(net_8462), .A2(net_8461) );
DFF_X2 inst_8288 ( .Q(net_10283), .D(net_4828), .CK(net_12921) );
NAND2_X2 inst_4254 ( .ZN(net_2963), .A2(net_1392), .A1(net_718) );
INV_X4 inst_5642 ( .ZN(net_1116), .A(net_845) );
NAND2_X2 inst_4330 ( .ZN(net_2676), .A1(net_1118), .A2(net_742) );
DFF_X2 inst_7459 ( .QN(net_9541), .D(net_8166), .CK(net_12753) );
CLKBUF_X2 inst_11898 ( .A(net_11816), .Z(net_11817) );
AOI21_X2 inst_10031 ( .A(net_7916), .B2(net_7915), .ZN(net_7847), .B1(net_623) );
DFF_X2 inst_8390 ( .QN(net_9196), .CK(net_11301), .D(x3507) );
CLKBUF_X2 inst_14220 ( .A(net_12968), .Z(net_14139) );
CLKBUF_X2 inst_11925 ( .A(net_11843), .Z(net_11844) );
INV_X2 inst_6659 ( .ZN(net_8461), .A(net_8418) );
DFF_X2 inst_7828 ( .Q(net_10300), .D(net_6452), .CK(net_14542) );
NAND2_X2 inst_4368 ( .A2(net_10353), .ZN(net_916), .A1(net_915) );
AND4_X4 inst_10331 ( .A2(net_10163), .ZN(net_3338), .A4(net_2256), .A1(net_1323), .A3(net_882) );
CLKBUF_X2 inst_12204 ( .A(net_11666), .Z(net_12123) );
CLKBUF_X2 inst_11137 ( .A(net_10895), .Z(net_11056) );
AOI22_X2 inst_9388 ( .B1(net_9999), .A1(net_5743), .B2(net_5742), .ZN(net_5435), .A2(net_239) );
CLKBUF_X2 inst_14577 ( .A(net_10733), .Z(net_14496) );
OR2_X4 inst_794 ( .A1(net_10473), .ZN(net_2207), .A2(net_1961) );
NOR2_X2 inst_2754 ( .ZN(net_3610), .A2(net_3167), .A1(net_2009) );
HA_X1 inst_7354 ( .A(net_9277), .S(net_3328), .CO(net_3327), .B(net_2457) );
CLKBUF_X2 inst_12049 ( .A(net_10607), .Z(net_11968) );
NOR2_X2 inst_2759 ( .ZN(net_3554), .A1(net_3364), .A2(net_3148) );
CLKBUF_X2 inst_12092 ( .A(net_12010), .Z(net_12011) );
OAI22_X2 inst_1147 ( .A1(net_7231), .A2(net_5134), .B2(net_5133), .ZN(net_5126), .B1(net_670) );
OAI21_X2 inst_1768 ( .ZN(net_8044), .B1(net_7924), .B2(net_7894), .A(net_7475) );
INV_X4 inst_6410 ( .ZN(net_929), .A(net_185) );
CLKBUF_X2 inst_12865 ( .A(net_12055), .Z(net_12784) );
CLKBUF_X2 inst_11165 ( .A(net_11083), .Z(net_11084) );
DFF_X2 inst_8256 ( .Q(net_10281), .D(net_4827), .CK(net_12947) );
NOR2_X2 inst_2917 ( .ZN(net_9086), .A2(net_1462), .A1(net_267) );
NOR3_X2 inst_2423 ( .A1(net_7602), .A2(net_7454), .A3(net_4512), .ZN(net_4317) );
OAI222_X2 inst_1408 ( .B2(net_7732), .A2(net_7731), .C2(net_7730), .ZN(net_5311), .B1(net_3226), .A1(net_2789), .C1(net_1127) );
OAI22_X2 inst_996 ( .B1(net_9366), .A2(net_8953), .ZN(net_8628), .A1(net_8627), .B2(net_8626) );
CLKBUF_X2 inst_10963 ( .A(net_10644), .Z(net_10882) );
INV_X4 inst_5889 ( .ZN(net_1111), .A(net_612) );
CLKBUF_X2 inst_12074 ( .A(net_11992), .Z(net_11993) );
CLKBUF_X2 inst_13563 ( .A(net_13481), .Z(net_13482) );
OAI21_X2 inst_1889 ( .B1(net_7245), .ZN(net_4864), .B2(net_4862), .A(net_4536) );
OAI221_X2 inst_1527 ( .C1(net_10208), .C2(net_7295), .B2(net_7293), .B1(net_7249), .ZN(net_7247), .A(net_6868) );
INV_X4 inst_6142 ( .A(net_10372), .ZN(net_783) );
OAI21_X2 inst_2011 ( .A(net_10439), .ZN(net_1844), .B2(net_1700), .B1(net_822) );
CLKBUF_X2 inst_13495 ( .A(net_11343), .Z(net_13414) );
OAI21_X2 inst_1761 ( .B2(net_8852), .ZN(net_8539), .A(net_8193), .B1(net_8120) );
OR2_X4 inst_740 ( .A1(net_9102), .ZN(net_7287), .A2(net_4902) );
INV_X4 inst_6582 ( .A(net_10328), .ZN(net_1354) );
AOI22_X2 inst_9418 ( .A1(net_10180), .A2(net_4656), .B2(net_4655), .ZN(net_4651), .B1(x4117) );
DFF_X2 inst_7803 ( .Q(net_9919), .D(net_6488), .CK(net_13404) );
INV_X4 inst_5474 ( .A(net_2721), .ZN(net_1307) );
NAND2_X2 inst_4189 ( .A1(net_4019), .ZN(net_2909), .A2(net_807) );
XNOR2_X2 inst_84 ( .ZN(net_8621), .A(net_8620), .B(net_8619) );
INV_X2 inst_6803 ( .ZN(net_5188), .A(net_5187) );
INV_X4 inst_5974 ( .A(net_9176), .ZN(net_752) );
CLKBUF_X2 inst_15756 ( .A(net_15674), .Z(net_15675) );
OAI21_X2 inst_1937 ( .B2(net_5341), .A(net_4629), .ZN(net_4462), .B1(net_4360) );
XNOR2_X2 inst_173 ( .ZN(net_5668), .B(net_5317), .A(net_5316) );
DFF_X2 inst_7660 ( .D(net_6691), .QN(net_171), .CK(net_12743) );
INV_X4 inst_5568 ( .ZN(net_2626), .A(net_912) );
NAND2_X2 inst_4405 ( .A2(net_10195), .A1(net_10181), .ZN(net_624) );
SDFF_X2 inst_611 ( .QN(net_10341), .SE(net_3665), .D(net_1292), .SI(net_1249), .CK(net_10649) );
AND2_X2 inst_10550 ( .A1(net_9225), .ZN(net_3481), .A2(net_3480) );
NOR2_X2 inst_2487 ( .A1(net_9561), .ZN(net_8735), .A2(net_8727) );
CLKBUF_X2 inst_12417 ( .A(net_12231), .Z(net_12336) );
INV_X4 inst_5821 ( .ZN(net_672), .A(net_671) );
INV_X2 inst_7187 ( .A(net_9397), .ZN(net_8209) );
INV_X4 inst_5713 ( .A(net_4446), .ZN(net_770) );
CLKBUF_X2 inst_12462 ( .A(net_11212), .Z(net_12381) );
AND2_X2 inst_10493 ( .ZN(net_6950), .A1(net_6949), .A2(net_6948) );
CLKBUF_X2 inst_12549 ( .A(net_11353), .Z(net_12468) );
DFF_X1 inst_8723 ( .D(net_6426), .CK(net_10986), .Q(x1074) );
CLKBUF_X2 inst_13047 ( .A(net_12965), .Z(net_12966) );
DFF_X2 inst_7802 ( .Q(net_9918), .D(net_6489), .CK(net_13405) );
OAI21_X2 inst_1943 ( .B2(net_10339), .A(net_10338), .ZN(net_4282), .B1(net_4281) );
DFF_X2 inst_7847 ( .Q(net_10010), .D(net_6477), .CK(net_11957) );
SDFF_X2 inst_490 ( .SE(net_9540), .SI(net_8219), .Q(net_306), .D(net_306), .CK(net_13898) );
INV_X4 inst_5573 ( .A(net_10224), .ZN(net_906) );
INV_X2 inst_7305 ( .A(net_9074), .ZN(net_9073) );
CLKBUF_X2 inst_13378 ( .A(net_13296), .Z(net_13297) );
DFF_X2 inst_8375 ( .QN(net_8830), .D(net_1494), .CK(net_13674) );
OAI211_X2 inst_2218 ( .C1(net_7216), .C2(net_6501), .ZN(net_6487), .B(net_5562), .A(net_3679) );
OAI22_X2 inst_1309 ( .ZN(net_3203), .A2(net_2401), .B2(net_2400), .A1(net_2400), .B1(net_1358) );
OAI221_X2 inst_1531 ( .B1(net_10305), .B2(net_9047), .C2(net_7287), .C1(net_7245), .ZN(net_7240), .A(net_6805) );
DFF_X2 inst_7640 ( .D(net_6731), .QN(net_154), .CK(net_13448) );
INV_X2 inst_7083 ( .ZN(net_1171), .A(net_1170) );
CLKBUF_X2 inst_15045 ( .A(net_14963), .Z(net_14964) );
CLKBUF_X2 inst_11706 ( .A(net_11624), .Z(net_11625) );
CLKBUF_X2 inst_15075 ( .A(net_14993), .Z(net_14994) );
CLKBUF_X2 inst_15049 ( .A(net_10629), .Z(net_14968) );
INV_X4 inst_4938 ( .ZN(net_5747), .A(net_2238) );
NOR2_X2 inst_2922 ( .A1(net_10355), .ZN(net_2392), .A2(net_1339) );
NAND2_X2 inst_3803 ( .A1(net_10072), .ZN(net_4536), .A2(net_4534) );
CLKBUF_X2 inst_13234 ( .A(net_10799), .Z(net_13153) );
CLKBUF_X2 inst_11831 ( .A(net_11749), .Z(net_11750) );
CLKBUF_X2 inst_11649 ( .A(net_11567), .Z(net_11568) );
AOI21_X2 inst_10242 ( .ZN(net_8860), .B1(net_2426), .B2(net_2425), .A(net_2424) );
NAND3_X2 inst_3183 ( .ZN(net_8088), .A1(net_8087), .A3(net_8086), .A2(net_7379) );
AND2_X4 inst_10410 ( .ZN(net_5765), .A1(net_4788), .A2(net_4787) );
CLKBUF_X2 inst_15095 ( .A(net_15013), .Z(net_15014) );
CLKBUF_X2 inst_10860 ( .A(net_10778), .Z(net_10779) );
CLKBUF_X2 inst_13301 ( .A(net_13219), .Z(net_13220) );
CLKBUF_X2 inst_11256 ( .A(net_11174), .Z(net_11175) );
NAND2_X2 inst_4312 ( .A2(net_10324), .ZN(net_2299), .A1(net_693) );
CLKBUF_X2 inst_12950 ( .A(net_12868), .Z(net_12869) );
INV_X4 inst_5328 ( .A(net_2255), .ZN(net_1470) );
DFF_X1 inst_8410 ( .Q(net_9308), .D(net_8800), .CK(net_14202) );
CLKBUF_X2 inst_13161 ( .A(net_13079), .Z(net_13080) );
INV_X4 inst_6226 ( .ZN(net_7216), .A(x4117) );
OAI22_X2 inst_1037 ( .B1(net_8919), .A2(net_8915), .ZN(net_7946), .A1(net_7845), .B2(net_2871) );
DFF_X2 inst_7777 ( .Q(net_9809), .D(net_6524), .CK(net_15430) );
DFF_X1 inst_8652 ( .Q(net_9685), .D(net_7261), .CK(net_15734) );
XNOR2_X2 inst_300 ( .B(net_9655), .ZN(net_3329), .A(net_3307) );
NAND2_X2 inst_3596 ( .ZN(net_7270), .A2(net_6881), .A1(net_6609) );
OAI22_X2 inst_1250 ( .B1(net_7226), .A2(net_4826), .B2(net_4825), .ZN(net_4824), .A1(net_467) );
CLKBUF_X2 inst_15407 ( .A(net_15325), .Z(net_15326) );
OAI22_X2 inst_1226 ( .A2(net_5155), .ZN(net_5020), .B1(net_4067), .B2(net_3871), .A1(net_562) );
INV_X2 inst_7071 ( .ZN(net_5009), .A(net_1232) );
AOI21_X2 inst_10240 ( .ZN(net_8852), .B2(net_8317), .A(net_8316), .B1(net_8185) );
INV_X4 inst_5964 ( .A(net_9326), .ZN(net_786) );
CLKBUF_X2 inst_15619 ( .A(net_15537), .Z(net_15538) );
DFF_X1 inst_8802 ( .QN(net_10340), .D(net_3716), .CK(net_10665) );
XNOR2_X2 inst_446 ( .B(net_9307), .ZN(net_802), .A(net_230) );
OAI21_X2 inst_1979 ( .B2(net_5420), .ZN(net_3158), .B1(net_2871), .A(net_2602) );
XNOR2_X2 inst_364 ( .ZN(net_2525), .B(net_2524), .A(net_2470) );
CLKBUF_X2 inst_11586 ( .A(net_11504), .Z(net_11505) );
AOI22_X2 inst_9253 ( .B2(net_6140), .A2(net_6109), .ZN(net_6055), .A1(net_6054), .B1(net_6053) );
INV_X4 inst_4923 ( .ZN(net_2699), .A(net_2698) );
AOI22_X2 inst_9283 ( .B1(net_9699), .A1(net_5755), .B2(net_5754), .ZN(net_5724), .A2(net_236) );
OR2_X4 inst_824 ( .A2(net_10145), .ZN(net_2076), .A1(net_609) );
NOR2_X2 inst_2997 ( .A1(net_10142), .ZN(net_2265), .A2(net_895) );
NAND2_X2 inst_3533 ( .A2(net_9631), .A1(net_8974), .ZN(net_8053) );
DFF_X2 inst_7839 ( .Q(net_9698), .D(net_6526), .CK(net_15676) );
INV_X4 inst_4712 ( .ZN(net_4729), .A(net_4728) );
XNOR2_X2 inst_411 ( .B(net_9312), .ZN(net_1479), .A(net_1478) );
CLKBUF_X2 inst_12897 ( .A(net_12815), .Z(net_12816) );
AOI22_X2 inst_9055 ( .ZN(net_8412), .A1(net_6892), .B2(net_6625), .B1(net_6039), .A2(net_5789) );
CLKBUF_X2 inst_14678 ( .A(net_14596), .Z(net_14597) );
AND2_X4 inst_10393 ( .A2(net_7046), .ZN(net_7044), .A1(net_7043) );
AND3_X2 inst_10380 ( .ZN(net_2102), .A1(net_2101), .A3(net_2098), .A2(net_819) );
INV_X4 inst_6600 ( .A(net_9383), .ZN(net_564) );
CLKBUF_X2 inst_13691 ( .A(net_11905), .Z(net_13610) );
AOI22_X2 inst_9007 ( .ZN(net_8031), .A2(net_8030), .B2(net_8029), .B1(net_2285), .A1(net_219) );
NAND2_X2 inst_3750 ( .ZN(net_5300), .A2(net_5288), .A1(net_4473) );
NAND2_X2 inst_4026 ( .A2(net_4067), .ZN(net_3604), .A1(net_2764) );
CLKBUF_X2 inst_14722 ( .A(net_14640), .Z(net_14641) );
CLKBUF_X2 inst_14649 ( .A(net_14567), .Z(net_14568) );
CLKBUF_X2 inst_11173 ( .A(net_11091), .Z(net_11092) );
CLKBUF_X2 inst_15286 ( .A(net_15204), .Z(net_15205) );
AOI22_X2 inst_9395 ( .B1(net_10004), .A1(net_5743), .B2(net_5742), .ZN(net_5412), .A2(net_244) );
CLKBUF_X2 inst_11333 ( .A(net_11251), .Z(net_11252) );
CLKBUF_X2 inst_10668 ( .A(net_10562), .Z(net_10587) );
NAND2_X2 inst_4056 ( .A2(net_8862), .ZN(net_4562), .A1(net_2768) );
CLKBUF_X2 inst_11010 ( .A(net_10928), .Z(net_10929) );
NAND2_X2 inst_4382 ( .ZN(net_2081), .A2(net_901), .A1(net_823) );
CLKBUF_X2 inst_10908 ( .A(net_10826), .Z(net_10827) );
NAND2_X2 inst_4401 ( .A2(net_10121), .A1(net_10120), .ZN(net_1854) );
CLKBUF_X2 inst_14426 ( .A(net_14344), .Z(net_14345) );
AND2_X4 inst_10388 ( .A2(net_9272), .ZN(net_8030), .A1(net_3286) );
NAND2_X2 inst_3430 ( .A1(net_9472), .A2(net_8487), .ZN(net_8486) );
CLKBUF_X2 inst_13480 ( .A(net_11500), .Z(net_13399) );
DFF_X1 inst_8708 ( .Q(net_9124), .D(net_6936), .CK(net_10586) );
CLKBUF_X2 inst_15400 ( .A(net_15318), .Z(net_15319) );
CLKBUF_X2 inst_13297 ( .A(net_13215), .Z(net_13216) );
CLKBUF_X2 inst_14020 ( .A(net_13938), .Z(net_13939) );
CLKBUF_X2 inst_13368 ( .A(net_10766), .Z(net_13287) );
AOI221_X2 inst_9874 ( .B1(net_9781), .B2(net_9097), .A(net_6940), .C2(net_6939), .ZN(net_6827), .C1(net_251) );
INV_X4 inst_5538 ( .A(net_10159), .ZN(net_3708) );
INV_X4 inst_5462 ( .ZN(net_1183), .A(net_1037) );
NAND2_X2 inst_3439 ( .A1(net_9484), .A2(net_8490), .ZN(net_8480) );
CLKBUF_X2 inst_13968 ( .A(net_13886), .Z(net_13887) );
DFF_X2 inst_8308 ( .QN(net_9572), .D(net_4561), .CK(net_12848) );
INV_X4 inst_5412 ( .ZN(net_1510), .A(net_1153) );
XNOR2_X2 inst_61 ( .ZN(net_8733), .A(net_8721), .B(net_8137) );
XNOR2_X2 inst_203 ( .ZN(net_4955), .A(net_4410), .B(net_2356) );
INV_X4 inst_5834 ( .ZN(net_1961), .A(net_888) );
CLKBUF_X2 inst_10901 ( .A(net_10819), .Z(net_10820) );
CLKBUF_X2 inst_14077 ( .A(net_13995), .Z(net_13996) );
AOI21_X2 inst_10014 ( .ZN(net_8571), .B2(net_8534), .A(net_2216), .B1(net_1857) );
OAI22_X2 inst_1139 ( .A1(net_7245), .ZN(net_5136), .A2(net_5134), .B2(net_5133), .B1(net_2193) );
AND2_X2 inst_10597 ( .ZN(net_2834), .A2(net_2167), .A1(net_315) );
CLKBUF_X2 inst_12459 ( .A(net_12364), .Z(net_12378) );
DFF_X1 inst_8852 ( .Q(net_10523), .D(net_95), .CK(net_10860) );
DFF_X1 inst_8520 ( .QN(net_10196), .D(net_7414), .CK(net_10867) );
INV_X4 inst_6601 ( .A(net_9166), .ZN(net_892) );
INV_X8 inst_4507 ( .ZN(net_6382), .A(net_5295) );
CLKBUF_X2 inst_14558 ( .A(net_13448), .Z(net_14477) );
AOI221_X2 inst_9968 ( .C1(net_9990), .B1(net_9756), .B2(net_6442), .ZN(net_4760), .A(net_4350), .C2(net_2541) );
CLKBUF_X2 inst_15540 ( .A(net_10757), .Z(net_15459) );
OAI221_X2 inst_1571 ( .C1(net_10323), .C2(net_9047), .B2(net_7287), .B1(net_7182), .ZN(net_7179), .A(net_6802) );
DFF_X2 inst_7631 ( .D(net_6763), .QN(net_120), .CK(net_15728) );
CLKBUF_X2 inst_14669 ( .A(net_14587), .Z(net_14588) );
CLKBUF_X2 inst_12009 ( .A(net_11927), .Z(net_11928) );
INV_X4 inst_6607 ( .A(net_10053), .ZN(net_4753) );
SDFF_X2 inst_456 ( .D(net_9570), .SI(net_9569), .Q(net_9568), .SE(net_4299), .CK(net_11585) );
OR2_X4 inst_832 ( .A2(net_10256), .A1(net_10255), .ZN(net_2428) );
DFF_X2 inst_8214 ( .Q(net_10082), .D(net_4853), .CK(net_10687) );
CLKBUF_X2 inst_11246 ( .A(net_11164), .Z(net_11165) );
INV_X4 inst_6511 ( .A(net_9972), .ZN(net_350) );
OAI222_X2 inst_1402 ( .B2(net_7732), .A2(net_7731), .C2(net_7730), .ZN(net_5328), .B1(net_3219), .A1(net_2770), .C1(net_1237) );
DFF_X2 inst_8102 ( .QN(net_9839), .D(net_5069), .CK(net_13308) );
XNOR2_X2 inst_275 ( .ZN(net_3950), .A(net_3233), .B(net_2029) );
CLKBUF_X2 inst_11492 ( .A(net_10705), .Z(net_11411) );
NAND4_X2 inst_3106 ( .ZN(net_4337), .A2(net_3779), .A3(net_3774), .A4(net_3767), .A1(net_3447) );
INV_X2 inst_6810 ( .ZN(net_4941), .A(net_4940) );
NAND2_X2 inst_3728 ( .A1(net_8511), .ZN(net_5733), .A2(net_5732) );
CLKBUF_X2 inst_11576 ( .A(net_11494), .Z(net_11495) );
CLKBUF_X2 inst_13379 ( .A(net_12289), .Z(net_13298) );
INV_X2 inst_6843 ( .ZN(net_3580), .A(net_3438) );
NOR3_X2 inst_2416 ( .ZN(net_5369), .A1(net_5368), .A3(net_5367), .A2(net_2406) );
INV_X4 inst_6270 ( .A(net_9211), .ZN(net_769) );
INV_X4 inst_5453 ( .A(net_2617), .ZN(net_1078) );
NAND2_X2 inst_3812 ( .A1(net_10081), .A2(net_4534), .ZN(net_4526) );
INV_X4 inst_5405 ( .A(net_2298), .ZN(net_1163) );
DFF_X1 inst_8810 ( .QN(net_10279), .D(net_3608), .CK(net_10619) );
CLKBUF_X2 inst_13317 ( .A(net_13235), .Z(net_13236) );
DFF_X2 inst_7879 ( .Q(net_9847), .D(net_6151), .CK(net_11950) );
NAND2_X2 inst_3959 ( .ZN(net_3618), .A2(net_3457), .A1(net_3456) );
INV_X2 inst_7193 ( .A(net_9204), .ZN(net_491) );
NOR2_X2 inst_2503 ( .A2(net_9436), .A1(net_9067), .ZN(net_8509) );
AOI221_X2 inst_9839 ( .A(net_6889), .B2(net_6888), .C2(net_6887), .ZN(net_6879), .B1(net_5845), .C1(x4937) );
CLKBUF_X2 inst_15347 ( .A(net_15265), .Z(net_15266) );
INV_X4 inst_5420 ( .ZN(net_1138), .A(net_1137) );
INV_X4 inst_4877 ( .A(net_3591), .ZN(net_3348) );
INV_X8 inst_4518 ( .ZN(net_8921), .A(net_8920) );
CLKBUF_X2 inst_11185 ( .A(net_11103), .Z(net_11104) );
AOI221_X2 inst_9994 ( .B2(net_10084), .C2(net_10083), .B1(net_10066), .C1(net_10065), .ZN(net_2113), .A(net_1422) );
CLKBUF_X2 inst_15415 ( .A(net_15333), .Z(net_15334) );
AND4_X2 inst_10348 ( .A3(net_9278), .A2(net_9277), .A1(net_9276), .ZN(net_1469), .A4(net_592) );
XNOR2_X2 inst_94 ( .B(net_8925), .ZN(net_8494), .A(net_8388) );
AOI222_X1 inst_9726 ( .B1(net_7583), .C1(net_4723), .ZN(net_3992), .A2(net_3078), .A1(net_2887), .C2(net_2618), .B2(net_2614) );
CLKBUF_X2 inst_10946 ( .A(net_10652), .Z(net_10865) );
INV_X2 inst_6832 ( .A(net_4135), .ZN(net_3994) );
CLKBUF_X2 inst_14234 ( .A(net_14152), .Z(net_14153) );
CLKBUF_X2 inst_14615 ( .A(net_12417), .Z(net_14534) );
DFF_X2 inst_7958 ( .QN(net_10202), .D(net_5631), .CK(net_13248) );
CLKBUF_X2 inst_11858 ( .A(net_11439), .Z(net_11777) );
CLKBUF_X2 inst_13060 ( .A(net_12978), .Z(net_12979) );
CLKBUF_X2 inst_11237 ( .A(net_11155), .Z(net_11156) );
NAND2_X2 inst_4345 ( .A2(net_4177), .A1(net_1847), .ZN(net_1027) );
XNOR2_X2 inst_424 ( .B(net_9942), .A(net_1413), .ZN(net_1375) );
SDFF_X2 inst_591 ( .Q(net_9262), .SE(net_4589), .D(net_145), .SI(net_111), .CK(net_12550) );
CLKBUF_X2 inst_15504 ( .A(net_15422), .Z(net_15423) );
NAND3_X4 inst_3166 ( .A1(net_8929), .ZN(net_8698), .A3(net_8681), .A2(net_8531) );
CLKBUF_X2 inst_15338 ( .A(net_15256), .Z(net_15257) );
CLKBUF_X2 inst_14218 ( .A(net_14136), .Z(net_14137) );
DFF_X2 inst_7452 ( .QN(net_9645), .D(net_8160), .CK(net_15383) );
CLKBUF_X2 inst_13807 ( .A(net_13725), .Z(net_13726) );
AND2_X4 inst_10428 ( .A2(net_10540), .A1(net_6203), .ZN(net_4006) );
NAND2_X2 inst_3656 ( .ZN(net_6652), .A1(net_6651), .A2(net_6226) );
CLKBUF_X2 inst_12497 ( .A(net_12415), .Z(net_12416) );
OAI211_X2 inst_2237 ( .C1(net_7198), .C2(net_6480), .ZN(net_6467), .B(net_5620), .A(net_3527) );
NAND2_X2 inst_4417 ( .A2(net_10191), .A1(net_10178), .ZN(net_574) );
CLKBUF_X2 inst_10784 ( .A(net_10702), .Z(net_10703) );
AOI22_X2 inst_9155 ( .A1(net_9754), .A2(net_6382), .ZN(net_6327), .B2(net_5263), .B1(net_3528) );
CLKBUF_X2 inst_14905 ( .A(net_14823), .Z(net_14824) );
DFF_X2 inst_8320 ( .Q(net_10398), .D(net_3925), .CK(net_12325) );
CLKBUF_X2 inst_14570 ( .A(net_14488), .Z(net_14489) );
INV_X2 inst_6834 ( .ZN(net_3941), .A(net_3940) );
INV_X4 inst_5727 ( .ZN(net_808), .A(net_756) );
CLKBUF_X2 inst_14012 ( .A(net_11318), .Z(net_13931) );
CLKBUF_X2 inst_11861 ( .A(net_11779), .Z(net_11780) );
INV_X2 inst_6853 ( .A(net_3909), .ZN(net_3374) );
NOR2_X2 inst_2706 ( .A2(net_4411), .ZN(net_4272), .A1(net_2680) );
DFF_X1 inst_8640 ( .QN(net_9611), .D(net_7145), .CK(net_15401) );
SDFF_X2 inst_476 ( .SE(net_9540), .SI(net_8233), .Q(net_292), .D(net_292), .CK(net_13975) );
AOI211_X4 inst_10249 ( .A(net_8995), .C2(net_8984), .ZN(net_7083), .B(net_5997), .C1(net_2246) );
INV_X2 inst_6684 ( .ZN(net_8344), .A(net_8278) );
NAND2_X2 inst_3742 ( .A1(net_5930), .ZN(net_5709), .A2(net_5360) );
CLKBUF_X2 inst_10701 ( .A(net_10550), .Z(net_10620) );
NOR2_X2 inst_2499 ( .ZN(net_9021), .A1(net_8525), .A2(net_8524) );
NOR2_X2 inst_2827 ( .ZN(net_2500), .A1(net_2499), .A2(net_1952) );
CLKBUF_X2 inst_11542 ( .A(net_11460), .Z(net_11461) );
AOI22_X2 inst_9062 ( .B1(net_9682), .A2(net_6684), .B2(net_6683), .ZN(net_6604), .A1(net_251) );
XOR2_X2 inst_20 ( .B(net_9152), .Z(net_2727), .A(net_1479) );
NOR3_X2 inst_2448 ( .ZN(net_2948), .A2(net_2712), .A3(net_2711), .A1(net_1763) );
AOI21_X2 inst_10007 ( .B1(net_8929), .ZN(net_8706), .B2(net_8681), .A(net_8530) );
CLKBUF_X2 inst_13421 ( .A(net_13339), .Z(net_13340) );
INV_X4 inst_5549 ( .ZN(net_6673), .A(net_932) );
INV_X4 inst_4994 ( .ZN(net_4714), .A(net_2222) );
CLKBUF_X2 inst_15387 ( .A(net_15305), .Z(net_15306) );
NOR2_X2 inst_2541 ( .ZN(net_8309), .A2(net_8308), .A1(net_8082) );
CLKBUF_X2 inst_14477 ( .A(net_13413), .Z(net_14396) );
CLKBUF_X2 inst_13590 ( .A(net_11699), .Z(net_13509) );
SDFF_X2 inst_576 ( .D(net_9128), .SE(net_933), .CK(net_10930), .SI(x2707), .Q(x1282) );
OAI221_X2 inst_1693 ( .C1(net_7231), .ZN(net_5465), .B1(net_5464), .B2(net_4477), .C2(net_4455), .A(net_3731) );
CLKBUF_X2 inst_14398 ( .A(net_14316), .Z(net_14317) );
AOI21_X2 inst_10182 ( .B2(net_9035), .B1(net_7504), .ZN(net_3515), .A(net_3514) );
AOI21_X2 inst_10131 ( .B2(net_10129), .ZN(net_4423), .A(net_2008), .B1(net_2007) );
NAND3_X2 inst_3306 ( .ZN(net_3638), .A1(net_1000), .A3(net_907), .A2(net_772) );
OAI22_X2 inst_1020 ( .A2(net_8036), .ZN(net_8019), .B2(net_8018), .A1(net_1402), .B1(net_766) );
CLKBUF_X2 inst_11007 ( .A(net_10895), .Z(net_10926) );
AND3_X2 inst_10376 ( .A3(net_9164), .ZN(net_3542), .A1(net_3541), .A2(x589) );
DFF_X2 inst_7721 ( .Q(net_9907), .D(net_6507), .CK(net_15070) );
NOR2_X2 inst_2876 ( .A2(net_10456), .A1(net_10455), .ZN(net_2459) );
NAND4_X2 inst_3055 ( .ZN(net_5731), .A4(net_4775), .A3(net_4213), .A1(net_3859), .A2(net_3413) );
CLKBUF_X2 inst_11057 ( .A(net_10975), .Z(net_10976) );
CLKBUF_X2 inst_13886 ( .A(net_13804), .Z(net_13805) );
OAI22_X2 inst_976 ( .ZN(net_8800), .A2(net_8798), .B1(net_4635), .B2(net_4223), .A1(net_1314) );
NAND2_X2 inst_3952 ( .A1(net_10263), .ZN(net_3711), .A2(net_3425) );
AOI221_X2 inst_9919 ( .B2(net_6443), .C2(net_6442), .ZN(net_5884), .A(net_5197), .B1(net_2287), .C1(net_1816) );
CLKBUF_X2 inst_12084 ( .A(net_12002), .Z(net_12003) );
OAI22_X2 inst_1279 ( .B2(net_7671), .A1(net_7602), .ZN(net_4457), .B1(net_4456), .A2(net_3878) );
NAND2_X2 inst_3588 ( .A1(net_7721), .ZN(net_7560), .A2(net_7374) );
INV_X2 inst_7027 ( .ZN(net_1501), .A(net_1500) );
INV_X4 inst_6562 ( .A(net_10256), .ZN(net_7481) );
CLKBUF_X2 inst_15120 ( .A(net_15038), .Z(net_15039) );
INV_X4 inst_5559 ( .ZN(net_1105), .A(net_923) );
OAI22_X2 inst_1096 ( .A1(net_9188), .A2(net_6299), .B2(net_6298), .ZN(net_6297), .B1(net_1729) );
CLKBUF_X2 inst_13011 ( .A(net_12929), .Z(net_12930) );
DFF_X2 inst_7474 ( .D(net_8062), .Q(net_209), .CK(net_15173) );
CLKBUF_X2 inst_13280 ( .A(net_12436), .Z(net_13199) );
CLKBUF_X2 inst_13287 ( .A(net_13205), .Z(net_13206) );
INV_X4 inst_4552 ( .ZN(net_8552), .A(net_8540) );
CLKBUF_X2 inst_11036 ( .A(net_10954), .Z(net_10955) );
DFF_X2 inst_8025 ( .QN(net_10430), .D(net_5466), .CK(net_11467) );
AOI22_X2 inst_9260 ( .A2(net_8042), .B2(net_6120), .ZN(net_6045), .B1(net_6044), .A1(net_5983) );
INV_X4 inst_5637 ( .ZN(net_2216), .A(net_1732) );
OAI21_X2 inst_1839 ( .B1(net_7157), .ZN(net_6216), .A(net_5776), .B2(net_5775) );
CLKBUF_X2 inst_14708 ( .A(net_10663), .Z(net_14627) );
DFF_X2 inst_8041 ( .QN(net_9547), .D(net_9253), .CK(net_13867) );
DFF_X2 inst_7723 ( .Q(net_9703), .D(net_6284), .CK(net_15066) );
NAND2_X2 inst_3399 ( .A1(net_8953), .A2(net_8941), .ZN(net_8874) );
NAND2_X2 inst_3414 ( .ZN(net_9112), .A1(net_8478), .A2(net_8436) );
CLKBUF_X2 inst_13095 ( .A(net_12366), .Z(net_13014) );
INV_X8 inst_4495 ( .ZN(net_6778), .A(net_5445) );
OAI222_X2 inst_1432 ( .ZN(net_2733), .C2(net_2732), .A2(net_2732), .B1(net_2731), .B2(net_2330), .C1(net_982), .A1(net_745) );
OR2_X4 inst_725 ( .ZN(net_7906), .A2(net_7701), .A1(net_7655) );
INV_X4 inst_5667 ( .A(net_10229), .ZN(net_815) );
CLKBUF_X2 inst_12840 ( .A(net_10804), .Z(net_12759) );
CLKBUF_X2 inst_12159 ( .A(net_12077), .Z(net_12078) );
INV_X4 inst_6326 ( .A(net_10431), .ZN(net_1950) );
NAND4_X2 inst_3084 ( .A3(net_9568), .A4(net_9563), .ZN(net_5343), .A2(net_4297), .A1(net_2850) );
CLKBUF_X2 inst_15562 ( .A(net_14638), .Z(net_15481) );
CLKBUF_X2 inst_11739 ( .A(net_10729), .Z(net_11658) );
OAI222_X2 inst_1337 ( .ZN(net_7661), .A1(net_7660), .B2(net_7659), .C2(net_7658), .A2(net_7552), .B1(net_7030), .C1(net_635) );
AOI221_X2 inst_9790 ( .B1(net_9968), .A(net_7090), .B2(net_7089), .C1(net_7088), .ZN(net_7061), .C2(net_240) );
INV_X4 inst_5375 ( .A(net_2258), .ZN(net_1540) );
NOR2_X4 inst_2464 ( .ZN(net_9033), .A1(net_8529), .A2(net_8527) );
NAND4_X2 inst_3096 ( .ZN(net_4347), .A1(net_3865), .A2(net_3864), .A3(net_3758), .A4(net_3442) );
CLKBUF_X2 inst_15532 ( .A(net_15450), .Z(net_15451) );
DFF_X1 inst_8776 ( .Q(net_10274), .D(net_4954), .CK(net_11770) );
NOR2_X2 inst_3015 ( .A2(net_9240), .A1(net_9172), .ZN(net_821) );
CLKBUF_X2 inst_11197 ( .A(net_10829), .Z(net_11116) );
AOI22_X2 inst_9433 ( .A1(net_9855), .B1(net_6828), .ZN(net_4496), .A2(net_4495), .B2(net_4494) );
CLKBUF_X2 inst_14432 ( .A(net_11172), .Z(net_14351) );
CLKBUF_X2 inst_15373 ( .A(net_15291), .Z(net_15292) );
NAND2_X2 inst_4010 ( .A2(net_9037), .ZN(net_3092), .A1(net_564) );
CLKBUF_X2 inst_13254 ( .A(net_11968), .Z(net_13173) );
AOI222_X1 inst_9677 ( .B1(net_9504), .ZN(net_8313), .A2(net_8295), .B2(net_8294), .C2(net_8293), .C1(net_8231), .A1(x3249) );
NAND2_X4 inst_3328 ( .A2(net_8934), .ZN(net_8608), .A1(net_8578) );
CLKBUF_X2 inst_11618 ( .A(net_11536), .Z(net_11537) );
NOR3_X2 inst_2441 ( .ZN(net_2944), .A2(net_2943), .A3(net_2709), .A1(net_2687) );
DFF_X2 inst_8399 ( .Q(net_10199), .D(net_10198), .CK(net_12236) );
CLKBUF_X2 inst_14495 ( .A(net_14413), .Z(net_14414) );
OAI22_X2 inst_1111 ( .A1(net_6623), .A2(net_6190), .B2(net_6184), .ZN(net_5952), .B1(net_968) );
CLKBUF_X2 inst_11945 ( .A(net_11863), .Z(net_11864) );
AOI22_X2 inst_9122 ( .A1(net_9674), .A2(net_6420), .ZN(net_6367), .B2(net_5263), .B1(net_112) );
NOR2_X2 inst_2658 ( .ZN(net_5372), .A2(net_5190), .A1(net_552) );
AOI222_X1 inst_9714 ( .C2(net_10137), .B1(net_10136), .ZN(net_7795), .A2(net_7711), .B2(net_7548), .C1(net_7331), .A1(net_7305) );
DFF_X2 inst_7427 ( .QN(net_9406), .D(net_8358), .CK(net_13944) );
OR2_X2 inst_878 ( .ZN(net_6612), .A1(net_6344), .A2(net_5956) );
CLKBUF_X2 inst_11496 ( .A(net_11414), .Z(net_11415) );
INV_X4 inst_4959 ( .ZN(net_3701), .A(net_2924) );
CLKBUF_X2 inst_13442 ( .A(net_12848), .Z(net_13361) );
INV_X2 inst_6782 ( .ZN(net_6016), .A(net_5826) );
SDFF_X2 inst_480 ( .SE(net_9540), .SI(net_8229), .Q(net_295), .D(net_295), .CK(net_13918) );
OAI21_X2 inst_1926 ( .ZN(net_4511), .B2(net_4066), .A(net_3347), .B1(net_3289) );
INV_X4 inst_4631 ( .ZN(net_7306), .A(net_6335) );
NAND2_X2 inst_4351 ( .A2(net_10248), .ZN(net_2732), .A1(net_639) );
INV_X4 inst_6211 ( .ZN(net_7184), .A(x5003) );
CLKBUF_X2 inst_12761 ( .A(net_12679), .Z(net_12680) );
INV_X4 inst_6383 ( .A(net_9971), .ZN(net_395) );
SDFF_X2 inst_564 ( .SE(net_9210), .Q(net_9210), .SI(net_6436), .D(net_6154), .CK(net_11785) );
NOR2_X2 inst_2986 ( .A1(net_10325), .ZN(net_1173), .A2(net_931) );
DFF_X2 inst_8074 ( .Q(net_9559), .D(net_9265), .CK(net_12615) );
OAI211_X2 inst_2206 ( .C1(net_7184), .C2(net_6501), .ZN(net_6499), .B(net_5567), .A(net_3679) );
CLKBUF_X2 inst_13597 ( .A(net_12154), .Z(net_13516) );
NOR2_X2 inst_2792 ( .ZN(net_3012), .A2(net_3011), .A1(net_2643) );
CLKBUF_X2 inst_12795 ( .A(net_11329), .Z(net_12714) );
AOI211_X2 inst_10262 ( .C2(net_7932), .ZN(net_7929), .C1(net_7928), .B(net_7806), .A(net_5686) );
OR2_X4 inst_739 ( .A1(net_9099), .ZN(net_7293), .A2(net_4905) );
CLKBUF_X2 inst_11210 ( .A(net_10612), .Z(net_11129) );
INV_X4 inst_6637 ( .A(net_9060), .ZN(net_9059) );
INV_X4 inst_6500 ( .A(net_10034), .ZN(net_5103) );
XOR2_X2 inst_46 ( .A(net_7634), .B(net_7632), .Z(net_1191) );
OR2_X2 inst_934 ( .A1(net_9204), .ZN(net_2517), .A2(net_2516) );
NOR2_X2 inst_2537 ( .ZN(net_8294), .A2(net_8293), .A1(net_8082) );
CLKBUF_X2 inst_15530 ( .A(net_11533), .Z(net_15449) );
OAI22_X2 inst_1000 ( .ZN(net_8548), .A2(net_8546), .B2(net_8545), .A1(net_2004), .B1(net_864) );
CLKBUF_X2 inst_12361 ( .A(net_12279), .Z(net_12280) );
OAI22_X2 inst_1126 ( .B1(net_9941), .A1(net_7182), .ZN(net_5154), .A2(net_5139), .B2(net_5138) );
CLKBUF_X2 inst_13065 ( .A(net_12983), .Z(net_12984) );
NAND2_X2 inst_3470 ( .A1(net_9439), .A2(net_8952), .ZN(net_8886) );
OR2_X4 inst_796 ( .ZN(net_2143), .A2(net_1386), .A1(net_1362) );
NOR2_X2 inst_2585 ( .ZN(net_7058), .A1(net_7057), .A2(net_6622) );
CLKBUF_X2 inst_12044 ( .A(net_11962), .Z(net_11963) );
NOR3_X2 inst_2364 ( .ZN(net_8805), .A1(net_8802), .A3(net_8629), .A2(net_7908) );
CLKBUF_X2 inst_14135 ( .A(net_14053), .Z(net_14054) );
CLKBUF_X2 inst_11727 ( .A(net_10673), .Z(net_11646) );
NAND2_X2 inst_4299 ( .A2(net_10159), .ZN(net_1531), .A1(net_1233) );
CLKBUF_X2 inst_11281 ( .A(net_11199), .Z(net_11200) );
OAI21_X2 inst_1882 ( .ZN(net_5223), .B1(net_5217), .B2(net_5216), .A(net_4382) );
CLKBUF_X2 inst_14510 ( .A(net_14428), .Z(net_14429) );
CLKBUF_X2 inst_13787 ( .A(net_11400), .Z(net_13706) );
CLKBUF_X2 inst_14482 ( .A(net_12477), .Z(net_14401) );
DFF_X2 inst_7812 ( .Q(net_10015), .D(net_6470), .CK(net_14756) );
CLKBUF_X2 inst_15030 ( .A(net_11027), .Z(net_14949) );
DFF_X2 inst_7628 ( .D(net_6777), .QN(net_178), .CK(net_14329) );
INV_X2 inst_6699 ( .A(net_8381), .ZN(net_8204) );
DFF_X1 inst_8441 ( .D(net_8453), .CK(net_11163), .Q(x962) );
DFF_X2 inst_8218 ( .Q(net_10185), .D(net_4832), .CK(net_12968) );
INV_X4 inst_6578 ( .A(net_10113), .ZN(net_5845) );
OAI221_X2 inst_1499 ( .C2(net_9063), .B2(net_9056), .ZN(net_7362), .C1(net_7224), .A(net_6996), .B1(net_5457) );
NOR2_X2 inst_2972 ( .A2(net_9211), .ZN(net_1567), .A1(net_1535) );
CLKBUF_X2 inst_12849 ( .A(net_12767), .Z(net_12768) );
AOI22_X2 inst_9470 ( .A1(net_10393), .B1(net_9877), .A2(net_4062), .ZN(net_3857), .B2(net_2973) );
INV_X4 inst_5531 ( .A(net_9371), .ZN(net_7902) );
INV_X4 inst_5397 ( .A(net_4166), .ZN(net_1599) );
OR2_X4 inst_727 ( .A1(net_9163), .ZN(net_8812), .A2(net_7592) );
CLKBUF_X2 inst_11795 ( .A(net_10776), .Z(net_11714) );
CLKBUF_X2 inst_15554 ( .A(net_15472), .Z(net_15473) );
INV_X4 inst_4804 ( .A(net_7832), .ZN(net_7704) );
CLKBUF_X2 inst_11686 ( .A(net_10917), .Z(net_11605) );
AOI22_X2 inst_9293 ( .B1(net_9902), .A1(net_5759), .B2(net_5758), .ZN(net_5699), .A2(net_241) );
NOR2_X2 inst_2874 ( .ZN(net_2645), .A2(net_1948), .A1(net_1127) );
CLKBUF_X2 inst_12345 ( .A(net_12263), .Z(net_12264) );
INV_X4 inst_6485 ( .A(net_9843), .ZN(net_669) );
INV_X4 inst_4607 ( .A(net_9310), .ZN(net_7694) );
NOR3_X2 inst_2431 ( .A3(net_9610), .A2(net_9104), .ZN(net_3715), .A1(net_3714) );
NAND3_X2 inst_3297 ( .A1(net_9247), .ZN(net_3018), .A3(net_1644), .A2(net_1340) );
DFF_X1 inst_8861 ( .QN(net_8847), .D(net_872), .CK(net_12662) );
INV_X4 inst_5931 ( .ZN(net_5473), .A(net_2702) );
INV_X4 inst_5429 ( .A(net_6808), .ZN(net_1130) );
CLKBUF_X2 inst_12556 ( .A(net_12474), .Z(net_12475) );
CLKBUF_X2 inst_12052 ( .A(net_11970), .Z(net_11971) );
NAND2_X1 inst_4423 ( .ZN(net_4184), .A1(net_4183), .A2(net_4182) );
AND2_X4 inst_10438 ( .A1(net_3134), .ZN(net_2358), .A2(net_2357) );
CLKBUF_X2 inst_13384 ( .A(net_13302), .Z(net_13303) );
CLKBUF_X2 inst_11880 ( .A(net_11798), .Z(net_11799) );
DFF_X2 inst_8274 ( .Q(net_10051), .D(net_4748), .CK(net_13165) );
DFF_X2 inst_7607 ( .QN(net_10148), .D(net_7159), .CK(net_13518) );
OAI33_X1 inst_953 ( .B1(net_7449), .A1(net_7345), .A3(net_7343), .ZN(net_7342), .B3(net_7341), .B2(net_1749), .A2(net_1158) );
CLKBUF_X2 inst_13674 ( .A(net_13592), .Z(net_13593) );
CLKBUF_X2 inst_11524 ( .A(net_11442), .Z(net_11443) );
NAND2_X2 inst_4342 ( .ZN(net_2056), .A1(net_840), .A2(net_839) );
CLKBUF_X2 inst_15691 ( .A(net_15580), .Z(net_15610) );
INV_X4 inst_5483 ( .A(net_9638), .ZN(net_6158) );
DFF_X1 inst_8664 ( .D(net_6742), .Q(net_144), .CK(net_15112) );
CLKBUF_X2 inst_12887 ( .A(net_12805), .Z(net_12806) );
AND2_X4 inst_10398 ( .A2(net_9103), .ZN(net_6944), .A1(net_4798) );
INV_X4 inst_5060 ( .A(net_4723), .ZN(net_3207) );
NAND2_X2 inst_4339 ( .A2(net_2017), .ZN(net_1781), .A1(net_1073) );
CLKBUF_X2 inst_14187 ( .A(net_13627), .Z(net_14106) );
OAI222_X2 inst_1421 ( .B2(net_7665), .A2(net_7664), .C2(net_7663), .ZN(net_4923), .B1(net_4104), .A1(net_2815), .C1(net_1930) );
INV_X2 inst_6694 ( .ZN(net_8322), .A(net_8205) );
NAND2_X4 inst_3373 ( .A2(net_9421), .ZN(net_6625), .A1(net_705) );
CLKBUF_X2 inst_12819 ( .A(net_11482), .Z(net_12738) );
INV_X4 inst_4902 ( .ZN(net_4962), .A(net_2577) );
NAND2_X2 inst_4262 ( .ZN(net_4110), .A2(net_1093), .A1(net_996) );
CLKBUF_X2 inst_12607 ( .A(net_12525), .Z(net_12526) );
DFF_X2 inst_8298 ( .Q(net_9513), .D(net_4612), .CK(net_12480) );
AND2_X4 inst_10406 ( .ZN(net_4906), .A1(net_4905), .A2(net_4904) );
CLKBUF_X2 inst_13882 ( .A(net_10856), .Z(net_13801) );
AOI222_X1 inst_9688 ( .B1(net_9505), .ZN(net_8296), .A2(net_8295), .B2(net_8294), .C2(net_8293), .C1(net_8224), .A1(x3194) );
NAND2_X2 inst_3664 ( .A2(net_10170), .ZN(net_6259), .A1(net_1966) );
AOI221_X2 inst_9961 ( .C1(net_10493), .B1(net_10283), .C2(net_6415), .B2(net_4774), .ZN(net_4770), .A(net_4341) );
DFF_X2 inst_7613 ( .QN(net_9215), .D(net_7059), .CK(net_11847) );
CLKBUF_X2 inst_11464 ( .A(net_11229), .Z(net_11383) );
AND2_X2 inst_10536 ( .ZN(net_4158), .A2(net_3703), .A1(net_3678) );
INV_X4 inst_6011 ( .A(net_10015), .ZN(net_526) );
INV_X2 inst_6956 ( .ZN(net_2794), .A(net_668) );
INV_X4 inst_4720 ( .ZN(net_4725), .A(net_4547) );
NAND2_X2 inst_3486 ( .ZN(net_8392), .A2(net_8391), .A1(net_8368) );
CLKBUF_X2 inst_13246 ( .A(net_13164), .Z(net_13165) );
CLKBUF_X2 inst_11488 ( .A(net_10829), .Z(net_11407) );
DFF_X1 inst_8833 ( .Q(net_9613), .D(net_2387), .CK(net_14118) );
CLKBUF_X2 inst_13961 ( .A(net_13879), .Z(net_13880) );
INV_X4 inst_4986 ( .ZN(net_2988), .A(net_2230) );
AOI22_X2 inst_9636 ( .A1(net_10084), .B1(net_10010), .A2(net_5319), .ZN(net_3406), .B2(net_2468) );
INV_X4 inst_6378 ( .A(net_9301), .ZN(net_666) );
XNOR2_X2 inst_294 ( .ZN(net_3475), .A(net_2797), .B(net_2452) );
CLKBUF_X2 inst_13510 ( .A(net_11120), .Z(net_13429) );
CLKBUF_X2 inst_13358 ( .A(net_13276), .Z(net_13277) );
CLKBUF_X2 inst_12099 ( .A(net_12017), .Z(net_12018) );
DFF_X2 inst_8275 ( .Q(net_9755), .D(net_4740), .CK(net_15417) );
DFF_X2 inst_7842 ( .Q(net_9696), .D(net_6530), .CK(net_15421) );
CLKBUF_X2 inst_15428 ( .A(net_15346), .Z(net_15347) );
CLKBUF_X2 inst_13769 ( .A(net_13687), .Z(net_13688) );
NAND2_X2 inst_3384 ( .ZN(net_8774), .A2(net_8757), .A1(net_1677) );
CLKBUF_X2 inst_11202 ( .A(net_11100), .Z(net_11121) );
INV_X4 inst_6628 ( .A(net_8978), .ZN(net_8977) );
AOI21_X2 inst_10029 ( .B1(net_9369), .A(net_7916), .B2(net_7915), .ZN(net_7850) );
DFF_X2 inst_7621 ( .QN(net_10265), .D(net_6932), .CK(net_11666) );
OR2_X4 inst_810 ( .A1(net_10157), .ZN(net_2427), .A2(net_1225) );
CLKBUF_X2 inst_13877 ( .A(net_13795), .Z(net_13796) );
CLKBUF_X1 inst_8982 ( .A(x185142), .Z(x911) );
XNOR2_X2 inst_230 ( .ZN(net_4388), .A(net_3941), .B(net_2335) );
INV_X4 inst_5903 ( .A(net_1115), .ZN(net_971) );
AOI22_X2 inst_9511 ( .B1(net_10508), .A1(net_9698), .B2(net_6415), .ZN(net_3812), .A2(net_3039) );
AOI221_X2 inst_9767 ( .ZN(net_7587), .C2(net_7586), .B2(net_7584), .A(net_7436), .B1(net_2187), .C1(net_1826) );
NAND4_X2 inst_3035 ( .A4(net_9605), .A2(net_9604), .ZN(net_8796), .A3(net_7647), .A1(net_313) );
AOI21_X2 inst_10089 ( .B1(net_10490), .A(net_6680), .ZN(net_5768), .B2(net_5200) );
CLKBUF_X2 inst_14855 ( .A(net_14312), .Z(net_14774) );
OAI21_X2 inst_1893 ( .B1(net_7241), .B2(net_4862), .ZN(net_4859), .A(net_4531) );
CLKBUF_X2 inst_12063 ( .A(net_10807), .Z(net_11982) );
INV_X4 inst_4728 ( .ZN(net_8116), .A(net_7277) );
INV_X4 inst_5101 ( .ZN(net_6564), .A(net_5954) );
DFF_X2 inst_8325 ( .Q(net_9617), .D(net_3269), .CK(net_14066) );
INV_X4 inst_6480 ( .A(net_9929), .ZN(net_915) );
NAND2_X2 inst_4385 ( .A2(net_9345), .ZN(net_1390), .A1(net_554) );
DFF_X2 inst_7836 ( .Q(net_9896), .D(net_6483), .CK(net_15681) );
AOI21_X2 inst_10010 ( .B1(net_8902), .ZN(net_8643), .A(net_8437), .B2(net_8391) );
CLKBUF_X2 inst_14573 ( .A(net_14491), .Z(net_14492) );
CLKBUF_X2 inst_11984 ( .A(net_11902), .Z(net_11903) );
SDFF_X2 inst_481 ( .SE(net_9540), .SI(net_8228), .Q(net_297), .D(net_297), .CK(net_13967) );
INV_X4 inst_5992 ( .A(net_10005), .ZN(net_536) );
INV_X4 inst_4606 ( .ZN(net_8647), .A(net_7592) );
DFF_X1 inst_8633 ( .Q(net_9882), .D(net_7222), .CK(net_14390) );
CLKBUF_X2 inst_14375 ( .A(net_14293), .Z(net_14294) );
XNOR2_X1 inst_452 ( .A(net_3223), .ZN(net_2478), .B(net_1723) );
AND4_X4 inst_10338 ( .ZN(net_3212), .A1(net_2428), .A3(net_2185), .A4(net_1684), .A2(net_1236) );
AOI22_X2 inst_9392 ( .B1(net_9905), .A1(net_5759), .B2(net_5758), .ZN(net_5421), .A2(net_244) );
CLKBUF_X2 inst_13699 ( .A(net_11873), .Z(net_13618) );
DFF_X2 inst_8397 ( .D(net_10541), .Q(net_9659), .CK(net_10850) );
NAND4_X2 inst_3061 ( .ZN(net_5725), .A4(net_4770), .A3(net_4212), .A1(net_3830), .A2(net_3434) );
INV_X4 inst_6208 ( .A(net_10436), .ZN(net_1210) );
CLKBUF_X2 inst_13146 ( .A(net_13064), .Z(net_13065) );
CLKBUF_X2 inst_14000 ( .A(net_13763), .Z(net_13919) );
NAND2_X2 inst_4144 ( .ZN(net_2926), .A2(net_2368), .A1(net_2320) );
AOI211_X2 inst_10254 ( .A(net_8190), .ZN(net_8188), .C2(net_7896), .C1(net_4632), .B(net_3298) );
CLKBUF_X2 inst_14308 ( .A(net_12775), .Z(net_14227) );
CLKBUF_X2 inst_11180 ( .A(net_11076), .Z(net_11099) );
OR2_X4 inst_728 ( .ZN(net_7782), .A1(net_7749), .A2(net_7556) );
CLKBUF_X2 inst_13056 ( .A(net_12974), .Z(net_12975) );
AND3_X2 inst_10372 ( .ZN(net_4690), .A1(net_4689), .A3(net_4688), .A2(net_2355) );
NOR2_X2 inst_2780 ( .ZN(net_3867), .A1(net_3145), .A2(net_3042) );
NAND4_X2 inst_3121 ( .A1(net_4041), .A3(net_3891), .ZN(net_3391), .A4(net_3390), .A2(net_3089) );
NOR2_X2 inst_2485 ( .ZN(net_8767), .A1(net_8766), .A2(net_8765) );
CLKBUF_X2 inst_15034 ( .A(net_13594), .Z(net_14953) );
AOI22_X2 inst_9087 ( .A1(net_9665), .ZN(net_6407), .A2(net_6402), .B2(net_5263), .B1(net_103) );
AND2_X2 inst_10584 ( .A1(net_9204), .ZN(net_2518), .A2(net_2516) );
INV_X2 inst_6655 ( .ZN(net_8503), .A(net_8502) );
CLKBUF_X2 inst_13353 ( .A(net_11472), .Z(net_13272) );
NAND2_X2 inst_4152 ( .ZN(net_2048), .A2(net_2047), .A1(net_1161) );
OAI211_X2 inst_2217 ( .C1(net_7198), .C2(net_6501), .ZN(net_6488), .B(net_5556), .A(net_3679) );
CLKBUF_X2 inst_13707 ( .A(net_13625), .Z(net_13626) );
CLKBUF_X2 inst_11031 ( .A(net_10949), .Z(net_10950) );
OR2_X2 inst_850 ( .A2(net_9577), .A1(net_9576), .ZN(net_8575) );
NOR2_X2 inst_2844 ( .ZN(net_2266), .A1(net_2265), .A2(net_1501) );
DFF_X2 inst_7612 ( .Q(net_9216), .D(net_6982), .CK(net_11848) );
NOR2_X2 inst_2492 ( .A2(net_9581), .ZN(net_8680), .A1(net_2578) );
CLKBUF_X2 inst_11175 ( .A(net_11093), .Z(net_11094) );
CLKBUF_X2 inst_15571 ( .A(net_15150), .Z(net_15490) );
NAND2_X2 inst_3582 ( .A2(net_10242), .ZN(net_7404), .A1(net_1115) );
NAND2_X2 inst_3480 ( .A1(net_9459), .A2(net_8951), .ZN(net_8432) );
CLKBUF_X2 inst_14125 ( .A(net_13096), .Z(net_14044) );
CLKBUF_X2 inst_12642 ( .A(net_10831), .Z(net_12561) );
CLKBUF_X2 inst_11721 ( .A(net_11639), .Z(net_11640) );
CLKBUF_X2 inst_14485 ( .A(net_14403), .Z(net_14404) );
NOR3_X2 inst_2438 ( .A2(net_9544), .ZN(net_7573), .A1(net_7546), .A3(net_3088) );
INV_X4 inst_5705 ( .ZN(net_776), .A(net_775) );
CLKBUF_X2 inst_15577 ( .A(net_15495), .Z(net_15496) );
CLKBUF_X2 inst_10879 ( .A(net_10797), .Z(net_10798) );
AND2_X4 inst_10391 ( .ZN(net_7322), .A2(net_7321), .A1(net_1085) );
INV_X4 inst_5479 ( .ZN(net_6054), .A(net_1956) );
XNOR2_X2 inst_237 ( .ZN(net_4260), .A(net_4108), .B(net_1813) );
NOR2_X2 inst_2543 ( .ZN(net_8300), .A2(net_8299), .A1(net_8082) );
NOR2_X2 inst_2772 ( .ZN(net_3233), .A2(net_3232), .A1(net_2649) );
CLKBUF_X2 inst_15314 ( .A(net_15232), .Z(net_15233) );
CLKBUF_X2 inst_11449 ( .A(net_11367), .Z(net_11368) );
DFF_X1 inst_8836 ( .Q(net_9858), .D(net_2159), .CK(net_10805) );
CLKBUF_X2 inst_13178 ( .A(net_13096), .Z(net_13097) );
DFF_X2 inst_7638 ( .D(net_6735), .QN(net_151), .CK(net_13877) );
DFF_X2 inst_8056 ( .QN(net_10120), .D(net_5510), .CK(net_12335) );
CLKBUF_X2 inst_14776 ( .A(net_14694), .Z(net_14695) );
CLKBUF_X2 inst_11017 ( .A(net_10629), .Z(net_10936) );
INV_X2 inst_7093 ( .A(net_2622), .ZN(net_1100) );
INV_X4 inst_4818 ( .ZN(net_3540), .A(net_3059) );
XOR2_X1 inst_51 ( .Z(net_6942), .A(net_6012), .B(net_1937) );
OR2_X4 inst_813 ( .ZN(net_2074), .A2(net_1363), .A1(net_844) );
AND3_X2 inst_10379 ( .A3(net_10224), .A1(net_3196), .ZN(net_2734), .A2(net_1287) );
INV_X2 inst_6691 ( .ZN(net_8333), .A(net_8271) );
CLKBUF_X2 inst_14874 ( .A(net_10884), .Z(net_14793) );
CLKBUF_X2 inst_13373 ( .A(net_13291), .Z(net_13292) );
CLKBUF_X2 inst_11195 ( .A(net_11113), .Z(net_11114) );
AND3_X2 inst_10381 ( .ZN(net_2100), .A1(net_2099), .A3(net_2098), .A2(net_451) );
OAI21_X2 inst_1837 ( .ZN(net_7060), .A(net_6563), .B2(net_2508), .B1(net_1420) );
OAI22_X2 inst_974 ( .A1(net_8813), .B2(net_8812), .ZN(net_8807), .A2(net_8805), .B1(net_426) );
CLKBUF_X2 inst_13198 ( .A(net_13116), .Z(net_13117) );
AOI22_X2 inst_9100 ( .A1(net_9681), .A2(net_6420), .ZN(net_6392), .B2(net_5263), .B1(net_853) );
INV_X4 inst_5686 ( .ZN(net_1085), .A(net_801) );
CLKBUF_X2 inst_10944 ( .A(net_10862), .Z(net_10863) );
NAND3_X2 inst_3291 ( .A2(net_4714), .A3(net_3591), .ZN(net_2942), .A1(net_2941) );
XNOR2_X2 inst_64 ( .ZN(net_8729), .A(net_8707), .B(net_8133) );
OAI22_X2 inst_1001 ( .ZN(net_8547), .A2(net_8546), .B2(net_8545), .A1(net_2633), .B1(net_435) );
CLKBUF_X2 inst_13964 ( .A(net_13882), .Z(net_13883) );
OR2_X4 inst_743 ( .A1(net_10058), .ZN(net_5899), .A2(net_5898) );
OAI211_X2 inst_2106 ( .C2(net_6778), .ZN(net_6742), .A(net_6370), .B(net_6100), .C1(net_490) );
NAND2_X2 inst_4051 ( .A2(net_3142), .ZN(net_2809), .A1(net_2808) );
NOR2_X2 inst_2723 ( .A2(net_10385), .ZN(net_4322), .A1(net_3872) );
NOR2_X1 inst_3033 ( .A1(net_2972), .A2(net_2555), .ZN(net_2462) );
INV_X4 inst_5825 ( .A(net_2210), .ZN(net_917) );
NOR2_X2 inst_2925 ( .A2(net_10353), .A1(net_10352), .ZN(net_2006) );
DFF_X2 inst_7843 ( .Q(net_9920), .D(net_6487), .CK(net_14221) );
AOI22_X2 inst_9141 ( .A1(net_9724), .A2(net_6382), .ZN(net_6345), .B1(net_6344), .B2(net_5263) );
NAND2_X2 inst_4265 ( .A1(net_10261), .ZN(net_4114), .A2(net_1367) );
AND2_X2 inst_10537 ( .ZN(net_3999), .A2(net_3657), .A1(net_203) );
AOI22_X2 inst_9510 ( .B1(net_9895), .A1(net_9764), .B2(net_4969), .ZN(net_3813), .A2(net_2462) );
OAI21_X2 inst_1828 ( .B1(net_7157), .ZN(net_6454), .B2(net_5439), .A(net_5426) );
DFF_X1 inst_8628 ( .Q(net_9787), .D(net_7207), .CK(net_13360) );
OAI21_X2 inst_1809 ( .ZN(net_7390), .B2(net_7060), .A(net_5345), .B1(net_5344) );
NAND2_X2 inst_3388 ( .ZN(net_8765), .A2(net_8742), .A1(net_8737) );
NAND2_X2 inst_3735 ( .A1(net_10510), .ZN(net_5426), .A2(net_5425) );
INV_X2 inst_6664 ( .ZN(net_8364), .A(net_8307) );
CLKBUF_X2 inst_11238 ( .A(net_11156), .Z(net_11157) );
NOR2_X2 inst_2675 ( .ZN(net_5288), .A2(net_4781), .A1(net_3298) );
INV_X4 inst_5311 ( .ZN(net_1503), .A(net_1287) );
DFF_X2 inst_8272 ( .Q(net_10052), .D(net_4756), .CK(net_13167) );
CLKBUF_X2 inst_14602 ( .A(net_14520), .Z(net_14521) );
CLKBUF_X2 inst_12172 ( .A(net_11894), .Z(net_12091) );
CLKBUF_X2 inst_11866 ( .A(net_11784), .Z(net_11785) );
XNOR2_X2 inst_141 ( .ZN(net_7303), .A(net_6666), .B(net_2026) );
AND2_X2 inst_10578 ( .A1(net_9654), .ZN(net_3307), .A2(net_2829) );
NOR2_X2 inst_2520 ( .A1(net_8714), .ZN(net_8395), .A2(net_8249) );
NAND2_X2 inst_4344 ( .A2(net_4019), .A1(net_1970), .ZN(net_1032) );
DFF_X2 inst_8111 ( .Q(net_9936), .D(net_5120), .CK(net_14301) );
DFF_X1 inst_8541 ( .Q(net_9975), .D(net_7371), .CK(net_14630) );
CLKBUF_X2 inst_15404 ( .A(net_15322), .Z(net_15323) );
CLKBUF_X2 inst_14717 ( .A(net_11811), .Z(net_14636) );
SDFF_X2 inst_571 ( .D(net_9131), .SE(net_933), .CK(net_10596), .SI(x2531), .Q(x1248) );
NAND2_X2 inst_4011 ( .ZN(net_3091), .A1(net_3090), .A2(net_3089) );
OAI21_X2 inst_1974 ( .ZN(net_2990), .B1(net_2760), .B2(net_2100), .A(net_850) );
INV_X4 inst_6007 ( .A(net_9987), .ZN(net_529) );
CLKBUF_X2 inst_11478 ( .A(net_11396), .Z(net_11397) );
AND2_X4 inst_10432 ( .ZN(net_3486), .A2(net_3009), .A1(net_1102) );
OAI21_X2 inst_2017 ( .ZN(net_8857), .B1(net_2678), .B2(net_2677), .A(net_2676) );
OAI22_X2 inst_1154 ( .A1(net_7243), .A2(net_5139), .B2(net_5138), .ZN(net_5119), .B1(net_2636) );
CLKBUF_X2 inst_15556 ( .A(net_11687), .Z(net_15475) );
CLKBUF_X2 inst_14901 ( .A(net_12209), .Z(net_14820) );
CLKBUF_X2 inst_14609 ( .A(net_14527), .Z(net_14528) );
DFF_X2 inst_7728 ( .Q(net_10003), .D(net_6271), .CK(net_12563) );
CLKBUF_X2 inst_12413 ( .A(net_11865), .Z(net_12332) );
INV_X4 inst_6445 ( .A(net_10475), .ZN(net_1035) );
AOI22_X2 inst_9584 ( .A1(net_10067), .B1(net_10046), .A2(net_5320), .B2(net_5174), .ZN(net_3578) );
INV_X2 inst_7224 ( .A(net_9547), .ZN(net_424) );
DFF_X2 inst_8045 ( .QN(net_10117), .D(net_5498), .CK(net_12338) );
DFF_X2 inst_7436 ( .QN(net_9415), .D(net_8349), .CK(net_11690) );
SDFF_X2 inst_469 ( .SE(net_8747), .SI(net_8622), .Q(net_236), .D(net_105), .CK(net_11579) );
DFF_X1 inst_8598 ( .Q(net_9683), .D(net_7263), .CK(net_15737) );
DFF_X2 inst_7468 ( .QN(net_9519), .D(net_8100), .CK(net_12751) );
CLKBUF_X2 inst_11689 ( .A(net_11392), .Z(net_11608) );
NOR2_X2 inst_2980 ( .A1(net_10431), .ZN(net_2643), .A2(net_686) );
INV_X4 inst_5197 ( .ZN(net_7583), .A(net_2488) );
INV_X2 inst_7133 ( .ZN(net_849), .A(net_848) );
INV_X2 inst_6837 ( .ZN(net_3888), .A(net_3887) );
CLKBUF_X2 inst_15013 ( .A(net_13567), .Z(net_14932) );
AOI21_X2 inst_10184 ( .ZN(net_3426), .A(net_3425), .B2(net_3105), .B1(net_2628) );
OR2_X2 inst_915 ( .ZN(net_3470), .A2(net_3469), .A1(net_2731) );
AOI221_X2 inst_9869 ( .B1(net_9777), .B2(net_9098), .A(net_6940), .C2(net_6939), .ZN(net_6833), .C1(net_247) );
DFF_X1 inst_8866 ( .Q(net_95), .CK(net_11859), .D(x3327) );
INV_X4 inst_6507 ( .A(net_9171), .ZN(net_761) );
INV_X4 inst_6642 ( .A(net_9084), .ZN(net_9083) );
NAND2_X2 inst_4416 ( .A2(net_10191), .A1(net_10184), .ZN(net_575) );
AOI21_X2 inst_10008 ( .B1(net_8944), .ZN(net_8689), .A(net_8317), .B2(net_8186) );
NOR4_X2 inst_2339 ( .ZN(net_3392), .A2(net_3198), .A4(net_2694), .A3(net_2363), .A1(net_1711) );
CLKBUF_X2 inst_12300 ( .A(net_11793), .Z(net_12219) );
INV_X4 inst_5660 ( .ZN(net_2668), .A(net_821) );
CLKBUF_X2 inst_14017 ( .A(net_13935), .Z(net_13936) );
CLKBUF_X2 inst_11603 ( .A(net_11521), .Z(net_11522) );
DFF_X2 inst_8260 ( .Q(net_10286), .D(net_4821), .CK(net_14521) );
OAI22_X2 inst_1216 ( .A1(net_7190), .A2(net_5107), .B2(net_5105), .ZN(net_5033), .B1(net_5032) );
CLKBUF_X2 inst_15544 ( .A(net_15462), .Z(net_15463) );
INV_X2 inst_6697 ( .ZN(net_8389), .A(net_8340) );
AOI22_X2 inst_9552 ( .B1(net_9988), .A1(net_9754), .A2(net_6442), .ZN(net_3768), .B2(net_2541) );
CLKBUF_X2 inst_14703 ( .A(net_11558), .Z(net_14622) );
CLKBUF_X2 inst_12591 ( .A(net_12509), .Z(net_12510) );
OAI33_X1 inst_952 ( .B1(net_7449), .ZN(net_7346), .A1(net_7345), .A2(net_7344), .A3(net_7343), .B3(net_5889), .B2(net_3088) );
INV_X4 inst_4807 ( .ZN(net_4232), .A(net_3611) );
OAI221_X2 inst_1668 ( .C1(net_7219), .A(net_5637), .B2(net_5591), .ZN(net_5501), .C2(net_4902), .B1(net_938) );
INV_X4 inst_5972 ( .A(net_10115), .ZN(net_696) );
CLKBUF_X2 inst_11169 ( .A(net_11087), .Z(net_11088) );
AOI221_X2 inst_9987 ( .B1(net_3885), .ZN(net_3603), .B2(net_3602), .C2(net_2916), .A(net_2903), .C1(net_2115) );
INV_X2 inst_7254 ( .A(net_9404), .ZN(net_8194) );
CLKBUF_X2 inst_15425 ( .A(net_15343), .Z(net_15344) );
INV_X4 inst_4811 ( .ZN(net_4076), .A(net_3561) );
CLKBUF_X2 inst_11942 ( .A(net_11860), .Z(net_11861) );
INV_X2 inst_7068 ( .ZN(net_1253), .A(net_817) );
CLKBUF_X2 inst_14710 ( .A(net_14628), .Z(net_14629) );
OR3_X2 inst_721 ( .A2(net_9529), .A1(net_9526), .ZN(net_2575), .A3(net_1696) );
CLKBUF_X2 inst_11135 ( .A(net_10646), .Z(net_11054) );
CLKBUF_X2 inst_10838 ( .A(net_10756), .Z(net_10757) );
INV_X2 inst_7211 ( .A(net_9392), .ZN(net_8211) );
XNOR2_X2 inst_293 ( .ZN(net_3497), .B(net_3496), .A(net_3266) );
INV_X4 inst_4741 ( .ZN(net_5012), .A(net_4687) );
CLKBUF_X2 inst_11078 ( .A(net_10996), .Z(net_10997) );
CLKBUF_X2 inst_13667 ( .A(net_13585), .Z(net_13586) );
OAI222_X2 inst_1366 ( .B1(net_7728), .A2(net_7727), .C2(net_7726), .ZN(net_6285), .B2(net_5738), .A1(net_4134), .C1(net_1290) );
NOR2_X2 inst_3009 ( .ZN(net_1372), .A1(net_840), .A2(net_839) );
NAND2_X2 inst_3744 ( .A1(net_5881), .ZN(net_5588), .A2(net_5322) );
CLKBUF_X2 inst_15346 ( .A(net_15264), .Z(net_15265) );
CLKBUF_X2 inst_13079 ( .A(net_12973), .Z(net_12998) );
OAI21_X2 inst_1915 ( .ZN(net_4596), .A(net_4439), .B2(net_4296), .B1(net_1902) );
NOR2_X2 inst_2794 ( .A1(net_9289), .A2(net_7502), .ZN(net_2970) );
INV_X4 inst_5402 ( .ZN(net_1971), .A(net_1166) );
OAI22_X2 inst_1254 ( .B1(net_7184), .A2(net_4826), .B2(net_4825), .ZN(net_4820), .A1(net_474) );
NOR2_X2 inst_2953 ( .A1(net_10369), .ZN(net_2641), .A2(net_600) );
INV_X2 inst_7111 ( .ZN(net_1003), .A(net_1002) );
CLKBUF_X2 inst_14412 ( .A(net_14330), .Z(net_14331) );
CLKBUF_X2 inst_14031 ( .A(net_13949), .Z(net_13950) );
NAND2_X2 inst_3553 ( .A1(net_10404), .ZN(net_7871), .A2(net_7863) );
CLKBUF_X2 inst_13000 ( .A(net_12918), .Z(net_12919) );
DFF_X2 inst_8219 ( .Q(net_10080), .D(net_4855), .CK(net_10730) );
XNOR2_X2 inst_98 ( .B(net_9431), .ZN(net_8411), .A(net_6208) );
OAI21_X2 inst_1811 ( .ZN(net_7085), .B1(net_6937), .B2(net_6898), .A(net_6239) );
INV_X4 inst_4544 ( .ZN(net_8644), .A(net_8586) );
CLKBUF_X2 inst_11147 ( .A(net_11065), .Z(net_11066) );
CLKBUF_X2 inst_11351 ( .A(net_11269), .Z(net_11270) );
NAND4_X2 inst_3087 ( .ZN(net_4489), .A2(net_4054), .A1(net_3804), .A3(net_3775), .A4(net_3732) );
OAI33_X1 inst_959 ( .A1(net_7602), .ZN(net_4513), .A3(net_4512), .B1(net_4071), .B3(net_3887), .B2(net_1515), .A2(net_1515) );
CLKBUF_X2 inst_14479 ( .A(net_14397), .Z(net_14398) );
CLKBUF_X2 inst_10801 ( .A(net_10719), .Z(net_10720) );
AOI21_X2 inst_10102 ( .B2(net_5174), .ZN(net_4899), .A(net_4502), .B1(net_702) );
CLKBUF_X2 inst_14611 ( .A(net_11870), .Z(net_14530) );
INV_X2 inst_7054 ( .ZN(net_1317), .A(net_1316) );
CLKBUF_X2 inst_14834 ( .A(net_12475), .Z(net_14753) );
DFF_X1 inst_8826 ( .QN(net_9566), .D(net_3245), .CK(net_12080) );
AOI22_X2 inst_9156 ( .A1(net_9755), .A2(net_6418), .ZN(net_6325), .B2(net_5263), .B1(net_1403) );
XNOR2_X2 inst_163 ( .ZN(net_9019), .B(net_5972), .A(net_5250) );
DFF_X1 inst_8455 ( .QN(net_10383), .D(net_8060), .CK(net_10678) );
XNOR2_X2 inst_394 ( .ZN(net_1999), .B(net_666), .A(net_209) );
CLKBUF_X2 inst_13343 ( .A(net_13261), .Z(net_13262) );
CLKBUF_X2 inst_11619 ( .A(net_11537), .Z(net_11538) );
DFF_X2 inst_7626 ( .D(net_6688), .QN(net_174), .CK(net_15614) );
SDFF_X2 inst_605 ( .Q(net_10517), .D(net_10517), .SE(net_4560), .CK(net_10551), .SI(x6028) );
AOI21_X4 inst_9998 ( .B1(net_9015), .ZN(net_8180), .A(net_7380), .B2(net_6905) );
OAI21_X2 inst_1814 ( .B2(net_10240), .ZN(net_6920), .A(net_1702), .B1(net_622) );
DFF_X2 inst_7481 ( .D(net_8065), .Q(net_216), .CK(net_12533) );
NOR2_X2 inst_2799 ( .A2(net_3117), .ZN(net_2892), .A1(net_2262) );
MUX2_X1 inst_4470 ( .S(net_6041), .A(net_5798), .B(x6264), .Z(x355) );
CLKBUF_X2 inst_10988 ( .A(net_10906), .Z(net_10907) );
CLKBUF_X2 inst_10875 ( .A(net_10793), .Z(net_10794) );
OAI211_X2 inst_2048 ( .C2(net_10486), .B(net_8821), .ZN(net_7840), .A(net_7765), .C1(net_1134) );
XNOR2_X2 inst_361 ( .ZN(net_3724), .A(net_2728), .B(net_2448) );
NOR2_X2 inst_2948 ( .ZN(net_4409), .A1(net_796), .A2(net_754) );
DFF_X2 inst_7900 ( .QN(net_10112), .D(net_6027), .CK(net_15516) );
CLKBUF_X2 inst_11358 ( .A(net_11276), .Z(net_11277) );
AND2_X4 inst_10396 ( .ZN(net_7088), .A2(net_6164), .A1(net_4794) );
NAND2_X2 inst_3400 ( .A2(net_8935), .A1(net_8894), .ZN(net_8607) );
DFF_X2 inst_8127 ( .Q(net_9836), .D(net_5135), .CK(net_12023) );
CLKBUF_X2 inst_11643 ( .A(net_11561), .Z(net_11562) );
CLKBUF_X2 inst_13850 ( .A(net_10786), .Z(net_13769) );
CLKBUF_X2 inst_12134 ( .A(net_12052), .Z(net_12053) );
OAI21_X2 inst_1931 ( .ZN(net_4914), .B1(net_4103), .A(net_4099), .B2(net_4097) );
DFF_X2 inst_8082 ( .QN(net_9169), .D(net_5788), .CK(net_11309) );
CLKBUF_X2 inst_11008 ( .A(net_10926), .Z(net_10927) );
INV_X4 inst_4735 ( .ZN(net_4787), .A(net_4467) );
INV_X4 inst_6631 ( .A(net_9039), .ZN(net_9035) );
CLKBUF_X2 inst_11926 ( .A(net_11844), .Z(net_11845) );
DFF_X2 inst_8402 ( .QN(net_9040), .CK(net_12993), .D(x3653) );
NOR2_X2 inst_3002 ( .ZN(net_2487), .A2(net_755), .A1(net_664) );
CLKBUF_X2 inst_13007 ( .A(net_11349), .Z(net_12926) );
CLKBUF_X2 inst_14852 ( .A(net_14770), .Z(net_14771) );
NAND2_X2 inst_4389 ( .A2(net_4190), .A1(net_1976), .ZN(net_799) );
OR2_X4 inst_786 ( .A1(net_9239), .ZN(net_3347), .A2(net_2751) );
INV_X2 inst_6828 ( .ZN(net_4082), .A(net_4081) );
CLKBUF_X2 inst_15153 ( .A(net_15071), .Z(net_15072) );
NOR2_X2 inst_2940 ( .A1(net_10474), .ZN(net_2576), .A2(net_1210) );
CLKBUF_X2 inst_11855 ( .A(net_11773), .Z(net_11774) );
DFF_X2 inst_7533 ( .QN(net_9311), .D(net_7784), .CK(net_15328) );
AOI22_X2 inst_9383 ( .B1(net_9702), .A1(net_5755), .B2(net_5754), .ZN(net_5441), .A2(net_239) );
INV_X4 inst_6606 ( .A(net_10440), .ZN(net_703) );
XOR2_X2 inst_2 ( .B(net_9068), .Z(net_6627), .A(net_6626) );
CLKBUF_X2 inst_11267 ( .A(net_10775), .Z(net_11186) );
CLKBUF_X2 inst_15048 ( .A(net_14966), .Z(net_14967) );
CLKBUF_X2 inst_11003 ( .A(net_10921), .Z(net_10922) );
INV_X2 inst_7022 ( .A(net_1786), .ZN(net_1525) );
NAND2_X2 inst_3474 ( .A2(net_9443), .A1(net_8952), .ZN(net_8907) );
CLKBUF_X2 inst_12328 ( .A(net_11319), .Z(net_12247) );
SDFF_X2 inst_578 ( .SE(net_5386), .D(net_3367), .CK(net_13474), .SI(x526), .Q(x526) );
OR2_X2 inst_888 ( .A1(net_10167), .ZN(net_6634), .A2(net_5971) );
CLKBUF_X2 inst_12306 ( .A(net_12224), .Z(net_12225) );
OAI21_X2 inst_1769 ( .ZN(net_8013), .B1(net_8012), .A(net_7874), .B2(net_7870) );
NAND2_X2 inst_3625 ( .ZN(net_7101), .A1(net_6869), .A2(net_6671) );
INV_X4 inst_5999 ( .ZN(net_726), .A(net_176) );
CLKBUF_X2 inst_14197 ( .A(net_14115), .Z(net_14116) );
CLKBUF_X2 inst_13063 ( .A(net_11817), .Z(net_12982) );
INV_X4 inst_6598 ( .A(net_10004), .ZN(net_318) );
INV_X4 inst_5979 ( .A(net_9642), .ZN(net_1028) );
CLKBUF_X2 inst_15164 ( .A(net_15082), .Z(net_15083) );
INV_X2 inst_7317 ( .A(net_9103), .ZN(net_9101) );
DFF_X2 inst_7817 ( .Q(net_10022), .D(net_6455), .CK(net_15540) );
NOR2_X2 inst_2581 ( .ZN(net_7308), .A2(net_7077), .A1(net_4601) );
NAND2_X2 inst_4110 ( .ZN(net_2362), .A1(net_1973), .A2(net_1689) );
OAI211_X2 inst_2164 ( .C1(net_7184), .C2(net_6548), .ZN(net_6547), .A(net_6546), .B(net_5673) );
OAI221_X2 inst_1498 ( .C2(net_9063), .B2(net_9056), .ZN(net_7365), .C1(net_7229), .A(net_6998), .B1(net_5473) );
OAI222_X2 inst_1358 ( .B1(net_7732), .A2(net_7731), .C2(net_7730), .ZN(net_6931), .B2(net_5975), .A1(net_4434), .C1(net_3100) );
INV_X2 inst_7198 ( .A(net_9590), .ZN(net_483) );
CLKBUF_X2 inst_13208 ( .A(net_13126), .Z(net_13127) );
DFF_X2 inst_8343 ( .D(net_10542), .QN(net_10515), .CK(net_10872) );
CLKBUF_X2 inst_11696 ( .A(net_11614), .Z(net_11615) );
NAND2_X2 inst_4392 ( .A2(net_10296), .A1(net_10289), .ZN(net_765) );
CLKBUF_X2 inst_11093 ( .A(net_11011), .Z(net_11012) );
DFF_X1 inst_8590 ( .Q(net_9668), .D(net_7111), .CK(net_12097) );
INV_X4 inst_4915 ( .A(net_7095), .ZN(net_3298) );
CLKBUF_X2 inst_15758 ( .A(net_11813), .Z(net_15677) );
CLKBUF_X2 inst_14424 ( .A(net_14342), .Z(net_14343) );
CLKBUF_X2 inst_12456 ( .A(net_12374), .Z(net_12375) );
INV_X4 inst_4775 ( .ZN(net_4014), .A(net_4013) );
DFF_X1 inst_8530 ( .Q(net_9968), .D(net_7320), .CK(net_15649) );
AOI22_X2 inst_9655 ( .B1(net_9735), .ZN(net_2551), .A1(net_2209), .A2(net_2208), .B2(net_1669) );
CLKBUF_X2 inst_11245 ( .A(net_10597), .Z(net_11164) );
CLKBUF_X2 inst_10831 ( .A(net_10749), .Z(net_10750) );
MUX2_X1 inst_4450 ( .S(net_6041), .A(net_296), .B(x5143), .Z(x132) );
CLKBUF_X2 inst_12817 ( .A(net_12735), .Z(net_12736) );
CLKBUF_X2 inst_12460 ( .A(net_12378), .Z(net_12379) );
NAND3_X2 inst_3182 ( .ZN(net_8109), .A1(net_8108), .A2(net_8107), .A3(net_1584) );
NAND2_X2 inst_3385 ( .ZN(net_8768), .A1(net_8766), .A2(net_8765) );
CLKBUF_X2 inst_14557 ( .A(net_14475), .Z(net_14476) );
OAI221_X2 inst_1572 ( .C1(net_10316), .C2(net_9047), .B2(net_7287), .B1(net_7234), .ZN(net_7177), .A(net_6844) );
CLKBUF_X2 inst_11753 ( .A(net_11671), .Z(net_11672) );
NOR2_X2 inst_2866 ( .A2(net_2403), .ZN(net_2042), .A1(net_2041) );
INV_X2 inst_6805 ( .A(net_5360), .ZN(net_5143) );
INV_X4 inst_4906 ( .ZN(net_4774), .A(net_2461) );
CLKBUF_X2 inst_11528 ( .A(net_11050), .Z(net_11447) );
CLKBUF_X2 inst_11546 ( .A(net_11464), .Z(net_11465) );
CLKBUF_X2 inst_14932 ( .A(net_14850), .Z(net_14851) );
INV_X4 inst_5379 ( .ZN(net_1591), .A(net_1199) );
OR2_X4 inst_838 ( .A2(net_10361), .A1(net_10360), .ZN(net_2432) );
CLKBUF_X2 inst_14815 ( .A(net_13680), .Z(net_14734) );
CLKBUF_X2 inst_15634 ( .A(net_10788), .Z(net_15553) );
CLKBUF_X2 inst_14026 ( .A(net_13656), .Z(net_13945) );
AOI21_X2 inst_10221 ( .ZN(net_2803), .B1(net_2296), .B2(net_1852), .A(net_1170) );
CLKBUF_X2 inst_12905 ( .A(net_12823), .Z(net_12824) );
INV_X4 inst_4978 ( .ZN(net_2592), .A(net_1517) );
OAI222_X2 inst_1405 ( .B2(net_7728), .A2(net_7727), .C2(net_7726), .ZN(net_5325), .B1(net_4107), .A1(net_3252), .C1(net_1913) );
DFF_X2 inst_7875 ( .QN(net_10355), .D(net_6002), .CK(net_13658) );
INV_X2 inst_6811 ( .ZN(net_4932), .A(net_4931) );
NAND2_X2 inst_4058 ( .A2(net_8861), .ZN(net_4583), .A1(net_2766) );
INV_X2 inst_6786 ( .A(net_9258), .ZN(net_5804) );
AOI22_X2 inst_9172 ( .A1(net_9924), .B1(net_9825), .ZN(net_6146), .B2(net_6140), .A2(net_6109) );
NOR2_X2 inst_2749 ( .A1(net_3687), .ZN(net_3673), .A2(net_3672) );
INV_X4 inst_5584 ( .ZN(net_2938), .A(net_886) );
AOI222_X1 inst_9721 ( .C1(net_10494), .B1(net_10389), .C2(net_6415), .A2(net_6413), .B2(net_4062), .ZN(net_4061), .A1(net_619) );
INV_X2 inst_6963 ( .ZN(net_1838), .A(net_1126) );
CLKBUF_X2 inst_12048 ( .A(net_11966), .Z(net_11967) );
DFF_X1 inst_8823 ( .Q(net_9197), .D(net_3607), .CK(net_13603) );
CLKBUF_X2 inst_11118 ( .A(net_11036), .Z(net_11037) );
CLKBUF_X2 inst_14647 ( .A(net_14565), .Z(net_14566) );
INV_X4 inst_5567 ( .A(net_3448), .ZN(net_3172) );
AND4_X2 inst_10346 ( .ZN(net_4240), .A2(net_4239), .A3(net_3722), .A4(net_3629), .A1(net_2690) );
NAND2_X2 inst_4367 ( .A2(net_4026), .A1(net_1978), .ZN(net_920) );
OAI21_X2 inst_2013 ( .A(net_4033), .B2(net_4022), .ZN(net_1709), .B1(net_1708) );
INV_X8 inst_4506 ( .ZN(net_6402), .A(net_5295) );
NOR2_X2 inst_2756 ( .A1(net_7435), .A2(net_3919), .ZN(net_3605) );
DFF_X2 inst_7712 ( .QN(net_10145), .D(net_6273), .CK(net_13513) );
AOI21_X2 inst_10071 ( .ZN(net_6620), .A(net_6619), .B1(net_4677), .B2(net_4555) );
SDFF_X2 inst_492 ( .SE(net_9540), .SI(net_8217), .Q(net_308), .D(net_308), .CK(net_11653) );
OAI21_X2 inst_1731 ( .ZN(net_8758), .A(net_8756), .B1(net_8739), .B2(net_8734) );
DFF_X1 inst_8635 ( .Q(net_9884), .D(net_7230), .CK(net_12161) );
INV_X2 inst_7229 ( .A(net_9414), .ZN(net_8219) );
INV_X4 inst_5414 ( .A(net_1345), .ZN(net_1151) );
NOR2_X2 inst_2960 ( .ZN(net_1842), .A2(net_1057), .A1(net_826) );
DFF_X2 inst_7960 ( .QN(net_10204), .D(net_5628), .CK(net_14361) );
OAI21_X2 inst_1909 ( .B2(net_10131), .A(net_10130), .ZN(net_4676), .B1(net_4675) );
CLKBUF_X2 inst_12589 ( .A(net_12288), .Z(net_12508) );
NAND2_X2 inst_4318 ( .A2(net_10455), .ZN(net_1624), .A1(net_584) );
INV_X4 inst_6616 ( .A(net_8938), .ZN(net_8937) );
CLKBUF_X2 inst_12292 ( .A(net_12210), .Z(net_12211) );
CLKBUF_X2 inst_11080 ( .A(net_10998), .Z(net_10999) );
XNOR2_X2 inst_82 ( .A(net_8953), .ZN(net_8623), .B(net_2930) );
NAND2_X2 inst_4335 ( .ZN(net_1687), .A2(net_1363), .A1(net_594) );
NAND2_X2 inst_4187 ( .ZN(net_2118), .A2(net_1859), .A1(net_1239) );
NAND2_X2 inst_4239 ( .A1(net_2761), .ZN(net_1508), .A2(net_1507) );
CLKBUF_X2 inst_15586 ( .A(net_15504), .Z(net_15505) );
CLKBUF_X2 inst_11669 ( .A(net_11587), .Z(net_11588) );
HA_X1 inst_7335 ( .CO(net_7325), .S(net_6961), .A(net_6960), .B(net_5989) );
DFF_X2 inst_7991 ( .QN(net_10418), .D(net_5535), .CK(net_11747) );
AOI22_X2 inst_9063 ( .B1(net_9683), .A2(net_6684), .B2(net_6683), .ZN(net_6603), .A1(net_252) );
CLKBUF_X2 inst_12171 ( .A(net_12089), .Z(net_12090) );
DFF_X1 inst_8443 ( .Q(net_9436), .D(net_8404), .CK(net_14938) );
OAI22_X2 inst_1121 ( .A2(net_9087), .ZN(net_5419), .B1(net_2545), .A1(net_1326), .B2(net_876) );
DFF_X2 inst_7455 ( .QN(net_9646), .D(net_8187), .CK(net_13143) );
CLKBUF_X2 inst_12185 ( .A(net_12103), .Z(net_12104) );
NAND4_X2 inst_3161 ( .A4(net_2786), .A2(net_2785), .ZN(net_2150), .A3(net_2090), .A1(net_1729) );
NAND3_X2 inst_3187 ( .ZN(net_7725), .A3(net_7724), .A1(net_7721), .A2(net_7640) );
CLKBUF_X2 inst_14908 ( .A(net_14826), .Z(net_14827) );
CLKBUF_X2 inst_11053 ( .A(net_10971), .Z(net_10972) );
XNOR2_X2 inst_307 ( .ZN(net_3228), .B(net_2807), .A(net_2662) );
DFF_X1 inst_8411 ( .QN(net_9309), .D(net_8799), .CK(net_14200) );
DFF_X2 inst_8292 ( .Q(net_10397), .D(net_4814), .CK(net_15198) );
AOI21_X2 inst_10032 ( .B1(net_10490), .ZN(net_7869), .A(net_6680), .B2(net_263) );
CLKBUF_X2 inst_12663 ( .A(net_12581), .Z(net_12582) );
CLKBUF_X2 inst_11462 ( .A(net_11380), .Z(net_11381) );
NOR2_X2 inst_2816 ( .ZN(net_2609), .A1(net_2608), .A2(net_2607) );
OAI211_X2 inst_2034 ( .C2(net_8102), .ZN(net_8100), .B(net_8098), .A(net_7999), .C1(net_2819) );
XNOR2_X2 inst_276 ( .ZN(net_3947), .A(net_3239), .B(net_2638) );
OR3_X2 inst_717 ( .A2(net_3529), .ZN(net_3055), .A3(net_3054), .A1(net_2466) );
OAI221_X2 inst_1505 ( .B2(net_9063), .C2(net_9056), .ZN(net_7356), .B1(net_7226), .A(net_6997), .C1(net_5480) );
CLKBUF_X2 inst_15097 ( .A(net_15015), .Z(net_15016) );
CLKBUF_X2 inst_13380 ( .A(net_13136), .Z(net_13299) );
AND2_X4 inst_10439 ( .A1(net_2684), .ZN(net_2338), .A2(net_1793) );
NAND2_X4 inst_3339 ( .A2(net_8885), .A1(net_8884), .ZN(net_8527) );
DFF_X1 inst_8460 ( .QN(net_10173), .D(net_7979), .CK(net_10822) );
NAND2_X2 inst_3791 ( .ZN(net_6679), .A2(net_5915), .A1(net_4634) );
CLKBUF_X2 inst_11557 ( .A(net_11391), .Z(net_11476) );
INV_X2 inst_7166 ( .A(net_3496), .ZN(net_566) );
INV_X4 inst_5297 ( .A(net_7902), .ZN(net_1306) );
XNOR2_X2 inst_91 ( .ZN(net_8564), .A(net_8506), .B(net_8422) );
OAI21_X2 inst_1762 ( .ZN(net_8406), .B1(net_8405), .A(net_8341), .B2(net_8329) );
OAI211_X4 inst_2023 ( .C2(net_9628), .C1(net_8972), .ZN(net_8126), .B(net_7959), .A(net_3728) );
NOR2_X2 inst_2779 ( .A1(net_9614), .A2(net_9613), .ZN(net_3146) );
DFF_X2 inst_7944 ( .QN(net_10324), .D(net_5488), .CK(net_12140) );
NAND2_X2 inst_3686 ( .ZN(net_6660), .A2(net_5990), .A1(net_2512) );
NAND2_X2 inst_3842 ( .ZN(net_4440), .A2(net_4269), .A1(net_2426) );
INV_X4 inst_6508 ( .ZN(net_5953), .A(net_277) );
CLKBUF_X2 inst_12186 ( .A(net_12104), .Z(net_12105) );
OAI221_X2 inst_1703 ( .C2(net_7671), .B1(net_7602), .ZN(net_5270), .A(net_4718), .C1(net_4508), .B2(net_3879) );
INV_X4 inst_4919 ( .ZN(net_6413), .A(net_4661) );
CLKBUF_X2 inst_13250 ( .A(net_13168), .Z(net_13169) );
INV_X4 inst_5886 ( .ZN(net_838), .A(net_617) );
INV_X4 inst_6566 ( .A(net_9209), .ZN(net_2758) );
INV_X2 inst_7167 ( .A(net_8439), .ZN(net_559) );
INV_X4 inst_4715 ( .ZN(net_5322), .A(net_4710) );
DFF_X2 inst_7424 ( .QN(net_9395), .D(net_8335), .CK(net_14012) );
CLKBUF_X2 inst_14894 ( .A(net_14812), .Z(net_14813) );
CLKBUF_X2 inst_14139 ( .A(net_12191), .Z(net_14058) );
CLKBUF_X2 inst_13680 ( .A(net_13058), .Z(net_13599) );
DFF_X2 inst_7788 ( .Q(net_9795), .D(net_6508), .CK(net_13207) );
SDFF_X2 inst_614 ( .SI(net_10541), .Q(net_10541), .SE(net_3633), .D(net_3393), .CK(net_11231) );
CLKBUF_X2 inst_14079 ( .A(net_11101), .Z(net_13998) );
CLKBUF_X2 inst_11897 ( .A(net_11409), .Z(net_11816) );
INV_X4 inst_6648 ( .ZN(net_9110), .A(net_959) );
AOI22_X2 inst_9080 ( .A1(net_9726), .ZN(net_6422), .A2(net_6404), .B2(net_5263), .B1(net_3060) );
DFF_X1 inst_8851 ( .Q(net_10527), .D(net_99), .CK(net_11203) );
CLKBUF_X2 inst_12197 ( .A(net_11645), .Z(net_12116) );
OAI21_X2 inst_1896 ( .B1(net_7136), .B2(net_4862), .ZN(net_4856), .A(net_4528) );
OAI22_X2 inst_1031 ( .A1(net_9270), .A2(net_7906), .B2(net_7904), .ZN(net_7903), .B1(net_7902) );
DFF_X2 inst_8075 ( .QN(net_10471), .D(net_5310), .CK(net_11377) );
OAI33_X1 inst_945 ( .B3(net_8850), .ZN(net_8771), .A3(net_8769), .A1(net_8749), .B2(net_8745), .A2(net_8743), .B1(net_8680) );
CLKBUF_X2 inst_11187 ( .A(net_11105), .Z(net_11106) );
XNOR2_X2 inst_369 ( .ZN(net_2507), .A(net_1738), .B(net_223) );
INV_X4 inst_6415 ( .ZN(net_7234), .A(x5427) );
INV_X4 inst_5161 ( .A(net_2292), .ZN(net_1572) );
OAI21_X2 inst_1900 ( .B1(net_7182), .B2(net_4862), .ZN(net_4852), .A(net_4524) );
CLKBUF_X2 inst_15044 ( .A(net_10655), .Z(net_14963) );
CLKBUF_X2 inst_12899 ( .A(net_12624), .Z(net_12818) );
DFF_X2 inst_7984 ( .QN(net_10428), .D(net_5543), .CK(net_14593) );
CLKBUF_X2 inst_12850 ( .A(net_12768), .Z(net_12769) );
INV_X4 inst_6489 ( .A(net_9739), .ZN(net_358) );
INV_X4 inst_5695 ( .ZN(net_787), .A(net_786) );
NOR2_X2 inst_2916 ( .ZN(net_1475), .A2(net_1474), .A1(net_816) );
XNOR2_X2 inst_266 ( .B(net_9656), .ZN(net_3972), .A(net_3650) );
OAI22_X2 inst_1286 ( .B1(net_9239), .A2(net_4319), .ZN(net_4036), .B2(net_1509), .A1(net_1177) );
AOI22_X2 inst_9288 ( .B1(net_9706), .A1(net_5755), .B2(net_5754), .ZN(net_5712), .A2(net_243) );
OAI211_X2 inst_2051 ( .ZN(net_7824), .C1(net_7823), .B(net_7718), .A(net_5354), .C2(net_2053) );
DFF_X2 inst_8382 ( .D(net_9234), .Q(net_9233), .CK(net_13536) );
DFF_X1 inst_8812 ( .QN(net_10172), .D(net_3537), .CK(net_10818) );
OAI22_X2 inst_1198 ( .A1(net_7249), .A2(net_5139), .B2(net_5138), .ZN(net_5055), .B1(net_1079) );
XNOR2_X2 inst_171 ( .ZN(net_5739), .A(net_4818), .B(net_2039) );
XNOR2_X2 inst_77 ( .B(net_8760), .ZN(net_8646), .A(net_8609) );
INV_X4 inst_6399 ( .A(net_9183), .ZN(net_2091) );
DFF_X2 inst_8224 ( .D(net_4866), .Q(net_229), .CK(net_10831) );
CLKBUF_X2 inst_10950 ( .A(net_10868), .Z(net_10869) );
XNOR2_X2 inst_374 ( .ZN(net_2474), .A(net_1772), .B(net_1724) );
CLKBUF_X2 inst_12832 ( .A(net_11102), .Z(net_12751) );
XNOR2_X2 inst_103 ( .ZN(net_8255), .A(net_8114), .B(net_6247) );
CLKBUF_X2 inst_14864 ( .A(net_14044), .Z(net_14783) );
CLKBUF_X2 inst_13328 ( .A(net_13246), .Z(net_13247) );
NAND2_X2 inst_3690 ( .A2(net_9252), .A1(net_9096), .ZN(net_6239) );
CLKBUF_X2 inst_11710 ( .A(net_10843), .Z(net_11629) );
CLKBUF_X2 inst_10763 ( .A(net_10681), .Z(net_10682) );
INV_X2 inst_7086 ( .A(net_3270), .ZN(net_1147) );
AOI22_X2 inst_9642 ( .ZN(net_3647), .B2(net_3011), .A2(net_2128), .A1(net_2127), .B1(net_1759) );
CLKBUF_X2 inst_11716 ( .A(net_11634), .Z(net_11635) );
INV_X4 inst_6061 ( .A(net_10497), .ZN(net_506) );
INV_X4 inst_6353 ( .A(net_10155), .ZN(net_756) );
AOI221_X2 inst_9905 ( .B1(net_9862), .B2(net_9101), .A(net_6945), .C2(net_6944), .C1(net_6813), .ZN(net_6789) );
CLKBUF_X2 inst_15713 ( .A(net_15631), .Z(net_15632) );
NAND2_X2 inst_3738 ( .A1(net_9160), .A2(net_7530), .ZN(net_5955) );
CLKBUF_X2 inst_11881 ( .A(net_11472), .Z(net_11800) );
DFF_X2 inst_8247 ( .Q(net_10089), .D(net_4846), .CK(net_10718) );
NOR2_X2 inst_2855 ( .A1(net_9657), .ZN(net_2109), .A2(net_1405) );
AOI21_X2 inst_10097 ( .B2(net_10490), .A(net_6680), .ZN(net_5425), .B1(net_627) );
INV_X2 inst_6749 ( .A(net_6903), .ZN(net_6621) );
CLKBUF_X2 inst_13553 ( .A(net_13471), .Z(net_13472) );
OR2_X4 inst_809 ( .A1(net_10264), .ZN(net_2203), .A2(net_1334) );
OAI211_X2 inst_2058 ( .A(net_7783), .C2(net_7782), .ZN(net_7775), .B(net_7680), .C1(net_2477) );
CLKBUF_X2 inst_14691 ( .A(net_13082), .Z(net_14610) );
AOI22_X2 inst_9637 ( .A1(net_10081), .B1(net_10007), .A2(net_5319), .ZN(net_3405), .B2(net_2468) );
CLKBUF_X2 inst_15821 ( .A(net_15739), .Z(net_15740) );
NAND2_X2 inst_3675 ( .A1(net_9075), .ZN(net_6616), .A2(net_6233) );
DFF_X2 inst_7816 ( .Q(net_9993), .D(net_6464), .CK(net_14610) );
OAI22_X2 inst_1234 ( .B1(net_7184), .A2(net_4890), .B2(net_4889), .ZN(net_4883), .A1(net_523) );
NOR2_X2 inst_2562 ( .A2(net_8614), .ZN(net_8612), .A1(net_7719) );
AOI21_X2 inst_10040 ( .B1(net_9051), .ZN(net_7699), .B2(net_7638), .A(net_7501) );
CLKBUF_X2 inst_14245 ( .A(net_14163), .Z(net_14164) );
NOR3_X2 inst_2398 ( .ZN(net_7612), .A3(net_7528), .A1(net_3984), .A2(x3390) );
CLKBUF_X2 inst_13925 ( .A(net_13843), .Z(net_13844) );
OAI22_X2 inst_1022 ( .A2(net_8036), .B2(net_8018), .ZN(net_8016), .A1(net_2522), .B1(net_595) );
NOR2_X2 inst_2595 ( .ZN(net_6899), .A2(net_6898), .A1(net_6240) );
INV_X4 inst_5614 ( .ZN(net_1314), .A(net_644) );
CLKBUF_X2 inst_15054 ( .A(net_11374), .Z(net_14973) );
AOI22_X2 inst_9248 ( .A1(net_9954), .B1(net_9855), .B2(net_6133), .A2(net_6111), .ZN(net_6063) );
CLKBUF_X2 inst_11938 ( .A(net_11856), .Z(net_11857) );
AOI22_X2 inst_9400 ( .ZN(net_5980), .A2(net_4703), .B1(net_3710), .B2(net_2700), .A1(net_2388) );
NOR3_X2 inst_2371 ( .A1(net_8190), .ZN(net_8157), .A2(net_8122), .A3(net_7933) );
NOR2_X2 inst_2939 ( .A1(net_10159), .ZN(net_2325), .A2(net_1233) );
INV_X2 inst_6818 ( .ZN(net_4678), .A(net_4677) );
AND2_X4 inst_10416 ( .ZN(net_4287), .A2(x3645), .A1(x813) );
OAI22_X2 inst_1223 ( .A1(net_7108), .A2(net_5139), .B2(net_5138), .ZN(net_5024), .B1(net_1898) );
NOR2_X2 inst_2785 ( .ZN(net_3419), .A1(net_3102), .A2(net_3101) );
CLKBUF_X2 inst_13636 ( .A(net_13554), .Z(net_13555) );
NAND2_X2 inst_3906 ( .ZN(net_3898), .A1(net_3897), .A2(net_3059) );
INV_X4 inst_6241 ( .A(net_9538), .ZN(net_457) );
INV_X4 inst_6574 ( .A(net_9556), .ZN(net_8439) );
OR4_X4 inst_681 ( .ZN(net_5937), .A1(net_5867), .A2(net_5359), .A4(net_5358), .A3(net_1240) );
DFF_X1 inst_8657 ( .Q(net_9765), .D(net_7242), .CK(net_13457) );
INV_X4 inst_5432 ( .ZN(net_1977), .A(net_1664) );
CLKBUF_X2 inst_13785 ( .A(net_13703), .Z(net_13704) );
DFF_X2 inst_7665 ( .Q(net_9279), .D(net_6838), .CK(net_15358) );
INV_X4 inst_4886 ( .ZN(net_5173), .A(net_2843) );
CLKBUF_X2 inst_15376 ( .A(net_15294), .Z(net_15295) );
AOI22_X2 inst_9322 ( .B1(net_9697), .A1(net_6808), .A2(net_5755), .B2(net_5754), .ZN(net_5654) );
OAI21_X2 inst_2010 ( .B1(net_5464), .B2(net_2016), .ZN(net_2003), .A(net_2002) );
CLKBUF_X2 inst_13181 ( .A(net_13099), .Z(net_13100) );
CLKBUF_X2 inst_15604 ( .A(net_15522), .Z(net_15523) );
CLKBUF_X2 inst_15103 ( .A(net_15021), .Z(net_15022) );
CLKBUF_X2 inst_11575 ( .A(net_11493), .Z(net_11494) );
CLKBUF_X2 inst_10665 ( .A(net_10554), .Z(net_10584) );
INV_X4 inst_5547 ( .A(net_10335), .ZN(net_1069) );
NOR2_X2 inst_2915 ( .A1(net_2753), .A2(net_2406), .ZN(net_1480) );
NAND3_X2 inst_3296 ( .A1(net_3630), .A3(net_2744), .ZN(net_2742), .A2(net_221) );
CLKBUF_X2 inst_14792 ( .A(net_12780), .Z(net_14711) );
AOI22_X2 inst_9135 ( .A1(net_9719), .A2(net_6404), .ZN(net_6353), .B2(net_5263), .B1(net_4188) );
OR2_X2 inst_871 ( .A1(net_8412), .ZN(net_7039), .A2(net_7038) );
INV_X4 inst_6148 ( .ZN(net_605), .A(net_175) );
NOR2_X2 inst_2684 ( .A2(net_10376), .ZN(net_4575), .A1(net_2257) );
INV_X4 inst_6320 ( .A(net_9963), .ZN(net_420) );
INV_X4 inst_6379 ( .A(net_9730), .ZN(net_895) );
SDFF_X2 inst_532 ( .Q(net_9304), .D(net_9304), .SI(net_9155), .SE(net_7553), .CK(net_14051) );
INV_X2 inst_6842 ( .A(net_8122), .ZN(net_3713) );
OAI22_X2 inst_1171 ( .A1(net_7184), .A2(net_5107), .B2(net_5105), .ZN(net_5091), .B1(net_5090) );
NOR3_X2 inst_2382 ( .ZN(net_7829), .A1(net_7828), .A3(net_7698), .A2(x3390) );
NOR2_X2 inst_2965 ( .A1(net_10224), .ZN(net_2679), .A2(net_2628) );
NAND4_X2 inst_3164 ( .ZN(net_1049), .A1(net_149), .A4(net_141), .A3(net_140), .A2(net_139) );
CLKBUF_X2 inst_12228 ( .A(net_11877), .Z(net_12147) );
NOR2_X2 inst_2969 ( .ZN(net_1779), .A2(net_1090), .A1(x6351) );
INV_X4 inst_5274 ( .A(net_5886), .ZN(net_1569) );
INV_X4 inst_5493 ( .ZN(net_2255), .A(net_1378) );
NAND3_X2 inst_3314 ( .A1(net_7344), .A3(net_7146), .ZN(net_1159), .A2(net_1158) );
INV_X4 inst_5616 ( .A(net_1817), .ZN(net_868) );
DFF_X2 inst_8192 ( .Q(net_9727), .D(net_5153), .CK(net_15119) );
INV_X4 inst_5766 ( .ZN(net_1000), .A(net_723) );
CLKBUF_X2 inst_14854 ( .A(net_14772), .Z(net_14773) );
NOR2_X2 inst_2594 ( .ZN(net_6906), .A2(net_6905), .A1(net_6244) );
INV_X4 inst_5113 ( .ZN(net_4267), .A(net_1646) );
CLKBUF_X2 inst_15294 ( .A(net_12948), .Z(net_15213) );
CLKBUF_X2 inst_14052 ( .A(net_13970), .Z(net_13971) );
NAND2_X2 inst_4037 ( .ZN(net_3042), .A2(net_2926), .A1(net_2924) );
NAND2_X2 inst_3976 ( .A1(net_3591), .ZN(net_3290), .A2(net_3289) );
CLKBUF_X2 inst_13277 ( .A(net_13195), .Z(net_13196) );
CLKBUF_X2 inst_13566 ( .A(net_11881), .Z(net_13485) );
CLKBUF_X2 inst_12073 ( .A(net_11991), .Z(net_11992) );
OAI22_X2 inst_1327 ( .B2(net_9744), .ZN(net_1430), .A2(net_1429), .B1(net_1413), .A1(net_194) );
AND2_X2 inst_10598 ( .A1(net_9653), .ZN(net_2829), .A2(net_2166) );
CLKBUF_X2 inst_11715 ( .A(net_11633), .Z(net_11634) );
CLKBUF_X2 inst_11773 ( .A(net_11403), .Z(net_11692) );
AOI22_X2 inst_9444 ( .A1(net_10523), .B1(net_9796), .ZN(net_4057), .A2(net_4056), .B2(net_2556) );
OAI22_X2 inst_1119 ( .ZN(net_5990), .A2(net_4967), .B2(net_4966), .B1(net_3712), .A1(net_2231) );
CLKBUF_X2 inst_15430 ( .A(net_15348), .Z(net_15349) );
CLKBUF_X2 inst_14748 ( .A(net_14666), .Z(net_14667) );
NAND2_X2 inst_3699 ( .ZN(net_6560), .A1(net_5938), .A2(net_5764) );
INV_X4 inst_5082 ( .ZN(net_1805), .A(net_1804) );
AOI222_X1 inst_9684 ( .B1(net_9504), .ZN(net_8303), .A2(net_8301), .B2(net_8300), .C2(net_8299), .C1(net_8228), .A1(x2278) );
OAI22_X2 inst_1255 ( .B1(net_7182), .A2(net_4826), .B2(net_4825), .ZN(net_4819), .A1(net_324) );
INV_X4 inst_6066 ( .ZN(net_3032), .A(net_201) );
AOI221_X2 inst_9844 ( .A(net_6889), .B2(net_6888), .C2(net_6887), .ZN(net_6874), .B1(net_5835), .C1(x5850) );
INV_X4 inst_5050 ( .ZN(net_2225), .A(net_1891) );
CLKBUF_X2 inst_10947 ( .A(net_10865), .Z(net_10866) );
AOI22_X2 inst_9279 ( .B1(net_9898), .A1(net_5759), .B2(net_5758), .ZN(net_5741), .A2(net_237) );
OAI21_X2 inst_1791 ( .B2(net_7505), .ZN(net_7490), .A(net_7489), .B1(net_564) );
AOI22_X2 inst_9112 ( .A1(net_9672), .A2(net_6382), .ZN(net_6377), .B2(net_5263), .B1(net_110) );
NAND2_X2 inst_3420 ( .ZN(net_8514), .A2(net_8481), .A1(net_8480) );
INV_X4 inst_4925 ( .ZN(net_2957), .A(net_2688) );
DFF_X1 inst_8834 ( .QN(net_10056), .D(net_2162), .CK(net_11223) );
INV_X2 inst_7021 ( .A(net_10351), .ZN(net_1529) );
MUX2_X1 inst_4457 ( .S(net_6041), .A(net_289), .B(x5601), .Z(x223) );
INV_X4 inst_6133 ( .ZN(net_5972), .A(net_276) );
CLKBUF_X2 inst_12341 ( .A(net_12259), .Z(net_12260) );
INV_X4 inst_5064 ( .ZN(net_1868), .A(net_1867) );
CLKBUF_X2 inst_11827 ( .A(net_11745), .Z(net_11746) );
SDFF_X2 inst_528 ( .SI(net_9337), .Q(net_9282), .D(net_9282), .SE(net_7588), .CK(net_14673) );
AOI22_X2 inst_9360 ( .B1(net_9920), .A1(net_6816), .A2(net_5759), .B2(net_5758), .ZN(net_5562) );
OR2_X2 inst_903 ( .ZN(net_4909), .A2(net_4500), .A1(net_4243) );
CLKBUF_X2 inst_14806 ( .A(net_14724), .Z(net_14725) );
CLKBUF_X2 inst_13574 ( .A(net_10708), .Z(net_13493) );
AOI221_X2 inst_9782 ( .C1(net_9350), .B1(net_9159), .A(net_7157), .B2(net_7155), .C2(net_7154), .ZN(net_7152) );
OAI21_X4 inst_1725 ( .B1(net_8948), .ZN(net_8169), .A(net_7472), .B2(net_7253) );
INV_X4 inst_5391 ( .ZN(net_5073), .A(net_1183) );
CLKBUF_X2 inst_13173 ( .A(net_13091), .Z(net_13092) );
INV_X4 inst_4957 ( .ZN(net_5454), .A(net_2547) );
INV_X2 inst_7238 ( .A(net_9612), .ZN(net_833) );
DFF_X1 inst_8607 ( .Q(net_9762), .D(net_7244), .CK(net_15471) );
CLKBUF_X2 inst_11377 ( .A(net_11295), .Z(net_11296) );
DFF_X1 inst_8602 ( .Q(net_9692), .D(net_7254), .CK(net_12009) );
OR2_X2 inst_846 ( .A2(net_9581), .A1(net_9580), .ZN(net_8679) );
INV_X4 inst_5925 ( .A(net_1947), .ZN(net_896) );
AOI222_X1 inst_9700 ( .B1(net_9511), .A2(net_8286), .B2(net_8285), .C2(net_8284), .ZN(net_8278), .C1(net_8198), .A1(x1418) );
NAND2_X2 inst_3504 ( .ZN(net_8961), .A1(net_8177), .A2(net_8176) );
NAND2_X2 inst_3924 ( .A1(net_4723), .A2(net_4319), .ZN(net_3883) );
OAI21_X2 inst_1734 ( .A(net_8756), .ZN(net_8738), .B2(net_8716), .B1(net_8715) );
CLKBUF_X2 inst_14408 ( .A(net_14326), .Z(net_14327) );
INV_X8 inst_4510 ( .ZN(net_8117), .A(net_6319) );
INV_X2 inst_7036 ( .ZN(net_1400), .A(net_1399) );
INV_X4 inst_4646 ( .ZN(net_6012), .A(net_6011) );
AOI22_X2 inst_9548 ( .A1(net_9875), .B2(net_5174), .ZN(net_3773), .B1(net_3772), .A2(net_2973) );
INV_X4 inst_4572 ( .ZN(net_8127), .A(net_8126) );
INV_X4 inst_5189 ( .A(net_2276), .ZN(net_1867) );
CLKBUF_X2 inst_13053 ( .A(net_12971), .Z(net_12972) );
CLKBUF_X2 inst_11203 ( .A(net_11121), .Z(net_11122) );
NAND2_X2 inst_3464 ( .A1(net_9467), .A2(net_8475), .ZN(net_8459) );
OAI22_X2 inst_1044 ( .A1(net_9365), .B2(net_7638), .ZN(net_7636), .A2(net_7635), .B1(net_7634) );
AOI22_X2 inst_9233 ( .A1(net_9897), .B1(net_9798), .A2(net_6141), .B2(net_6133), .ZN(net_6078) );
NAND2_X4 inst_3354 ( .ZN(net_8419), .A2(net_8385), .A1(net_8380) );
INV_X4 inst_6187 ( .A(net_9355), .ZN(net_5938) );
AOI211_X2 inst_10309 ( .B(net_5954), .ZN(net_2985), .A(net_2984), .C1(net_2983), .C2(net_2982) );
INV_X4 inst_4993 ( .ZN(net_4192), .A(net_2222) );
DFF_X2 inst_7554 ( .QN(net_9326), .D(net_7691), .CK(net_15306) );
AOI22_X2 inst_9509 ( .B1(net_10297), .A1(net_10192), .B2(net_4774), .A2(net_4217), .ZN(net_3814) );
CLKBUF_X2 inst_14389 ( .A(net_10729), .Z(net_14308) );
AOI22_X2 inst_9500 ( .B1(net_9920), .A1(net_9722), .B2(net_4969), .ZN(net_3823), .A2(net_3039) );
DFF_X2 inst_8327 ( .QN(net_10062), .D(net_3257), .CK(net_10713) );
NOR2_X2 inst_3014 ( .A1(net_10115), .ZN(net_1170), .A2(net_793) );
DFF_X2 inst_8199 ( .QN(net_9929), .D(net_5024), .CK(net_13689) );
CLKBUF_X2 inst_15112 ( .A(net_13264), .Z(net_15031) );
INV_X4 inst_6256 ( .ZN(net_454), .A(net_279) );
XNOR2_X2 inst_227 ( .ZN(net_4405), .B(net_4403), .A(net_3475) );
OAI221_X2 inst_1532 ( .B1(net_10306), .B2(net_9047), .C2(net_7287), .C1(net_7243), .ZN(net_7239), .A(net_6800) );
NAND2_X2 inst_4303 ( .A2(net_10456), .ZN(net_1611), .A1(net_1209) );
INV_X4 inst_5861 ( .ZN(net_807), .A(net_641) );
OAI211_X2 inst_2136 ( .C2(net_6774), .ZN(net_6712), .A(net_6406), .B(net_6143), .C1(net_376) );
NOR2_X2 inst_2718 ( .A2(net_10480), .A1(net_5175), .ZN(net_4959) );
NOR2_X2 inst_2891 ( .A1(net_5272), .A2(net_2913), .ZN(net_1775) );
NAND2_X2 inst_3927 ( .A1(net_4717), .A2(net_4319), .ZN(net_3879) );
XOR2_X1 inst_58 ( .Z(net_1539), .B(net_1538), .A(net_1238) );
CLKBUF_X2 inst_11653 ( .A(net_11571), .Z(net_11572) );
AOI22_X2 inst_9574 ( .B2(net_6443), .A2(net_6442), .ZN(net_3732), .A1(net_1559), .B1(net_1518) );
NAND2_X2 inst_3633 ( .A1(net_10191), .ZN(net_6983), .A2(net_6974) );
DFF_X2 inst_7557 ( .QN(net_10465), .D(net_7729), .CK(net_11409) );
DFF_X1 inst_8642 ( .Q(net_9890), .D(net_7210), .CK(net_14376) );
INV_X4 inst_6036 ( .A(net_10000), .ZN(net_516) );
AOI221_X2 inst_9775 ( .C1(net_9525), .C2(net_8001), .ZN(net_7475), .B2(net_7474), .B1(net_5198), .A(net_3298) );
CLKBUF_X2 inst_13792 ( .A(net_12044), .Z(net_13711) );
OAI221_X2 inst_1469 ( .ZN(net_7835), .A(net_7756), .C2(net_7449), .B2(net_7345), .C1(net_3689), .B1(net_3304) );
CLKBUF_X2 inst_12056 ( .A(net_11974), .Z(net_11975) );
AOI211_X2 inst_10295 ( .B(net_4007), .ZN(net_3747), .A(net_3746), .C1(net_3338), .C2(net_3321) );
AOI221_X2 inst_9944 ( .ZN(net_5336), .C2(net_5335), .B2(net_5335), .A(net_4644), .B1(net_3097), .C1(net_3083) );
INV_X4 inst_5029 ( .ZN(net_7672), .A(net_7512) );
CLKBUF_X2 inst_12878 ( .A(net_11788), .Z(net_12797) );
INV_X4 inst_5690 ( .ZN(net_1269), .A(net_794) );
AOI21_X2 inst_10200 ( .ZN(net_2877), .B1(net_2876), .B2(net_2242), .A(net_1333) );
CLKBUF_X2 inst_15457 ( .A(net_15375), .Z(net_15376) );
AOI22_X2 inst_9592 ( .ZN(net_3530), .A1(net_3529), .B1(net_3528), .A2(net_3503), .B2(net_3285) );
SDFF_X2 inst_581 ( .D(net_9133), .SE(net_933), .CK(net_10945), .SI(x2400), .Q(x1231) );
NOR2_X2 inst_2551 ( .A2(net_9512), .A1(net_8913), .ZN(net_7990) );
INV_X4 inst_5288 ( .ZN(net_5462), .A(net_2943) );
XOR2_X2 inst_28 ( .Z(net_2155), .A(net_2154), .B(net_623) );
NAND2_X2 inst_4407 ( .A2(net_9229), .A1(net_9228), .ZN(net_1440) );
NOR3_X2 inst_2424 ( .A2(net_9243), .A1(net_7602), .A3(net_4512), .ZN(net_4316) );
INV_X8 inst_4517 ( .A(net_8924), .ZN(net_8919) );
AOI22_X2 inst_9410 ( .A1(net_9954), .B1(net_6828), .ZN(net_4744), .A2(net_4734), .B2(net_4733) );
CLKBUF_X2 inst_12656 ( .A(net_12574), .Z(net_12575) );
AOI22_X2 inst_9434 ( .A1(net_9852), .B1(net_6813), .ZN(net_4493), .A2(net_4491), .B2(net_4490) );
CLKBUF_X2 inst_13719 ( .A(net_12826), .Z(net_13638) );
AOI22_X2 inst_9401 ( .ZN(net_5978), .A2(net_4702), .B1(net_3708), .B2(net_2551), .A1(net_2371) );
DFF_X2 inst_7440 ( .QN(net_9391), .D(net_8345), .CK(net_14004) );
NAND4_X2 inst_3144 ( .ZN(net_2423), .A4(net_1125), .A2(net_1051), .A1(net_624), .A3(net_574) );
CLKBUF_X2 inst_13386 ( .A(net_13304), .Z(net_13305) );
SDFF_X2 inst_592 ( .QN(net_9258), .SE(net_4589), .D(net_141), .SI(net_107), .CK(net_13828) );
INV_X4 inst_6124 ( .A(net_9206), .ZN(net_487) );
INV_X2 inst_7289 ( .A(net_8986), .ZN(net_8983) );
CLKBUF_X2 inst_13841 ( .A(net_13069), .Z(net_13760) );
CLKBUF_X2 inst_11530 ( .A(net_11448), .Z(net_11449) );
OAI22_X2 inst_993 ( .B1(net_9266), .A2(net_8962), .B2(net_8659), .ZN(net_8639), .A1(net_7171) );
NAND2_X2 inst_3666 ( .A2(net_10170), .A1(net_10169), .ZN(net_7069) );
CLKBUF_X2 inst_14882 ( .A(net_10835), .Z(net_14801) );
INV_X4 inst_5143 ( .ZN(net_3960), .A(net_1756) );
INV_X4 inst_5177 ( .ZN(net_1849), .A(net_1558) );
CLKBUF_X2 inst_14590 ( .A(net_14508), .Z(net_14509) );
INV_X4 inst_6407 ( .A(net_10393), .ZN(net_388) );
CLKBUF_X2 inst_15118 ( .A(net_15036), .Z(net_15037) );
INV_X2 inst_7264 ( .A(net_9400), .ZN(net_8233) );
CLKBUF_X2 inst_13855 ( .A(net_11905), .Z(net_13774) );
CLKBUF_X2 inst_13504 ( .A(net_13422), .Z(net_13423) );
DFF_X2 inst_7858 ( .Q(net_9701), .D(net_6224), .CK(net_15054) );
CLKBUF_X2 inst_14755 ( .A(net_11155), .Z(net_14674) );
CLKBUF_X2 inst_12876 ( .A(net_12794), .Z(net_12795) );
INV_X4 inst_5096 ( .ZN(net_2598), .A(net_1722) );
SDFF_X2 inst_630 ( .Q(net_9445), .D(net_9445), .SE(net_3293), .CK(net_12448), .SI(x2826) );
NAND2_X2 inst_3948 ( .A1(net_9533), .ZN(net_4149), .A2(net_3508) );
INV_X4 inst_5535 ( .A(net_1691), .ZN(net_1234) );
CLKBUF_X2 inst_11413 ( .A(net_11331), .Z(net_11332) );
INV_X4 inst_5227 ( .A(net_2873), .ZN(net_1834) );
CLKBUF_X2 inst_14157 ( .A(net_14075), .Z(net_14076) );
INV_X4 inst_5268 ( .ZN(net_5017), .A(net_3016) );
CLKBUF_X2 inst_11796 ( .A(net_11714), .Z(net_11715) );
AOI22_X2 inst_9662 ( .B2(net_10194), .A2(net_10193), .B1(net_10180), .A1(net_10179), .ZN(net_1051) );
OAI22_X2 inst_1273 ( .ZN(net_4748), .A1(net_4747), .A2(net_4746), .B2(net_4745), .B1(net_1130) );
CLKBUF_X2 inst_12791 ( .A(net_12709), .Z(net_12710) );
CLKBUF_X2 inst_11337 ( .A(net_10664), .Z(net_11256) );
SDFF_X2 inst_512 ( .Q(net_9327), .D(net_9327), .SI(net_9152), .SE(net_7588), .CK(net_13100) );
CLKBUF_X2 inst_11808 ( .A(net_11726), .Z(net_11727) );
INV_X4 inst_4966 ( .ZN(net_2485), .A(net_2133) );
OAI22_X2 inst_1301 ( .ZN(net_3097), .A1(net_3095), .B2(net_2921), .A2(net_2920), .B1(net_943) );
CLKBUF_X2 inst_14307 ( .A(net_14225), .Z(net_14226) );
CLKBUF_X2 inst_15308 ( .A(net_15226), .Z(net_15227) );
CLKBUF_X2 inst_12278 ( .A(net_11832), .Z(net_12197) );
OAI211_X2 inst_2151 ( .C2(net_6774), .ZN(net_6697), .A(net_6412), .B(net_6059), .C1(net_5066) );
CLKBUF_X2 inst_14109 ( .A(net_14027), .Z(net_14028) );
SDFF_X2 inst_647 ( .Q(net_9464), .D(net_9464), .SE(net_3293), .CK(net_11882), .SI(x1660) );
NOR2_X2 inst_2830 ( .ZN(net_3457), .A2(net_2168), .A1(x6445) );
NAND4_X2 inst_3054 ( .ZN(net_5870), .A4(net_4980), .A1(net_3769), .A3(net_3764), .A2(net_3752) );
CLKBUF_X2 inst_15450 ( .A(net_15368), .Z(net_15369) );
CLKBUF_X2 inst_12871 ( .A(net_12789), .Z(net_12790) );
CLKBUF_X2 inst_11744 ( .A(net_10734), .Z(net_11663) );
INV_X4 inst_4764 ( .ZN(net_4474), .A(net_4366) );
INV_X4 inst_5137 ( .ZN(net_3761), .A(net_1594) );
CLKBUF_X2 inst_13271 ( .A(net_13189), .Z(net_13190) );
NOR2_X2 inst_2985 ( .A1(net_10249), .ZN(net_2344), .A2(net_778) );
AOI221_X2 inst_9821 ( .B1(net_9867), .B2(net_9101), .A(net_6945), .C1(net_6944), .ZN(net_6933), .C2(net_238) );
DFF_X2 inst_8156 ( .QN(net_9740), .D(net_5070), .CK(net_12876) );
CLKBUF_X2 inst_15755 ( .A(net_15673), .Z(net_15674) );
OR2_X4 inst_833 ( .A2(net_10151), .A1(net_10150), .ZN(net_2430) );
NAND2_X2 inst_3772 ( .A1(net_8866), .ZN(net_4818), .A2(net_4758) );
NAND2_X2 inst_4210 ( .A1(net_9388), .A2(net_8914), .ZN(net_1748) );
CLKBUF_X2 inst_11968 ( .A(net_11886), .Z(net_11887) );
OAI33_X1 inst_960 ( .B2(net_9622), .ZN(net_4500), .A2(net_4499), .A1(net_4357), .A3(net_4355), .B3(net_4077), .B1(net_3530) );
OAI211_X2 inst_2043 ( .ZN(net_7934), .B(net_7836), .C1(net_7823), .C2(net_7341), .A(net_5262) );
XNOR2_X2 inst_118 ( .ZN(net_7716), .A(net_7715), .B(net_7055) );
INV_X4 inst_4924 ( .ZN(net_2697), .A(net_2696) );
NOR3_X2 inst_2411 ( .ZN(net_5811), .A2(net_5809), .A3(net_5808), .A1(net_5271) );
CLKBUF_X2 inst_12709 ( .A(net_12627), .Z(net_12628) );
CLKBUF_X2 inst_14433 ( .A(net_14351), .Z(net_14352) );
CLKBUF_X2 inst_10781 ( .A(net_10674), .Z(net_10700) );
XOR2_X2 inst_38 ( .A(net_9154), .B(net_9153), .Z(net_1724) );
INV_X4 inst_6591 ( .A(net_9992), .ZN(net_322) );
XNOR2_X2 inst_381 ( .B(net_10040), .ZN(net_2290), .A(net_2281) );
OAI211_X2 inst_2037 ( .C2(net_8102), .ZN(net_8080), .A(net_7998), .C1(net_3566), .B(net_3507) );
NOR2_X2 inst_2601 ( .ZN(net_6661), .A2(net_6660), .A1(net_3199) );
DFF_X1 inst_8578 ( .Q(net_9676), .D(net_7264), .CK(net_14825) );
CLKBUF_X2 inst_14846 ( .A(net_10993), .Z(net_14765) );
CLKBUF_X2 inst_13532 ( .A(net_13450), .Z(net_13451) );
AOI22_X2 inst_9448 ( .A1(net_10521), .B1(net_9794), .A2(net_4056), .ZN(net_4048), .B2(net_2556) );
INV_X2 inst_6930 ( .ZN(net_1945), .A(net_1944) );
AOI22_X2 inst_9102 ( .A1(net_9682), .A2(net_6402), .ZN(net_6390), .B2(net_5263), .B1(net_4017) );
NAND2_X2 inst_3837 ( .A2(net_4448), .ZN(net_4310), .A1(net_4309) );
CLKBUF_X2 inst_15343 ( .A(net_15261), .Z(net_15262) );
CLKBUF_X2 inst_12276 ( .A(net_12194), .Z(net_12195) );
OR2_X2 inst_883 ( .A2(net_7038), .ZN(net_6288), .A1(net_6287) );
INV_X2 inst_6876 ( .A(net_3891), .ZN(net_3360) );
DFF_X2 inst_7577 ( .QN(net_10161), .D(net_7541), .CK(net_13521) );
CLKBUF_X2 inst_12536 ( .A(net_12454), .Z(net_12455) );
CLKBUF_X2 inst_13108 ( .A(net_10625), .Z(net_13027) );
CLKBUF_X2 inst_12710 ( .A(net_12628), .Z(net_12629) );
AND3_X4 inst_10355 ( .ZN(net_4949), .A1(net_4948), .A3(net_4947), .A2(net_2571) );
OR2_X4 inst_756 ( .ZN(net_4399), .A2(net_4398), .A1(net_1670) );
DFF_X2 inst_8068 ( .QN(net_10469), .D(net_5312), .CK(net_11454) );
INV_X4 inst_5496 ( .A(net_10158), .ZN(net_2623) );
CLKBUF_X2 inst_13880 ( .A(net_13798), .Z(net_13799) );
INV_X4 inst_6002 ( .A(net_10495), .ZN(net_532) );
CLKBUF_X2 inst_13423 ( .A(net_12253), .Z(net_13342) );
AOI21_X2 inst_10228 ( .B1(net_2298), .ZN(net_2013), .A(net_2012), .B2(net_1178) );
AOI22_X2 inst_9270 ( .B1(net_9906), .ZN(net_5761), .A1(net_5759), .B2(net_5758), .A2(net_245) );
CLKBUF_X2 inst_15628 ( .A(net_15546), .Z(net_15547) );
INV_X2 inst_7150 ( .A(net_3433), .ZN(net_3163) );
CLKBUF_X2 inst_15500 ( .A(net_15418), .Z(net_15419) );
CLKBUF_X2 inst_14599 ( .A(net_14517), .Z(net_14518) );
CLKBUF_X2 inst_15008 ( .A(net_14926), .Z(net_14927) );
OAI22_X2 inst_1188 ( .A1(net_7294), .A2(net_5107), .B2(net_5105), .ZN(net_5067), .B1(net_5066) );
INV_X4 inst_4597 ( .ZN(net_7915), .A(net_7741) );
INV_X4 inst_5503 ( .ZN(net_1393), .A(net_982) );
AOI221_X2 inst_9873 ( .B1(net_9762), .B2(net_9097), .A(net_6940), .C2(net_6939), .ZN(net_6829), .C1(net_6828) );
AOI222_X1 inst_9685 ( .B1(net_9506), .ZN(net_8302), .A2(net_8301), .B2(net_8300), .C2(net_8299), .C1(net_8226), .A1(x2165) );
OAI22_X2 inst_1165 ( .A1(net_7245), .ZN(net_5108), .A2(net_5107), .B1(net_5106), .B2(net_5105) );
CLKBUF_X2 inst_14579 ( .A(net_14497), .Z(net_14498) );
INV_X4 inst_5439 ( .A(net_1273), .ZN(net_1110) );
CLKBUF_X2 inst_11029 ( .A(net_10569), .Z(net_10948) );
NOR2_X2 inst_2644 ( .A2(net_5449), .ZN(net_5446), .A1(net_2156) );
INV_X2 inst_6922 ( .ZN(net_2084), .A(net_2083) );
NOR2_X2 inst_2626 ( .A2(net_9252), .A1(net_9096), .ZN(net_6898) );
CLKBUF_X2 inst_13462 ( .A(net_12459), .Z(net_13381) );
AOI221_X2 inst_9960 ( .C1(net_10492), .B1(net_10282), .C2(net_6415), .B2(net_4774), .ZN(net_4771), .A(net_4342) );
AOI22_X2 inst_9314 ( .B1(net_9719), .A2(net_5755), .B2(net_5754), .ZN(net_5663), .A1(net_256) );
INV_X4 inst_4629 ( .A(net_7783), .ZN(net_7749) );
INV_X2 inst_6957 ( .ZN(net_1877), .A(net_1876) );
INV_X2 inst_7184 ( .A(net_10262), .ZN(net_520) );
CLKBUF_X2 inst_14140 ( .A(net_14058), .Z(net_14059) );
INV_X4 inst_5983 ( .A(net_9962), .ZN(net_541) );
AOI22_X2 inst_9056 ( .B1(net_9662), .A1(net_6834), .A2(net_6684), .B2(net_6683), .ZN(net_6610) );
DFF_X2 inst_8363 ( .QN(net_10337), .D(net_2267), .CK(net_11055) );
NAND2_X2 inst_3873 ( .ZN(net_4629), .A2(net_4227), .A1(net_4080) );
INV_X2 inst_6883 ( .A(net_3080), .ZN(net_3052) );
OAI22_X2 inst_992 ( .A2(net_8962), .B2(net_8659), .ZN(net_8640), .A1(net_7039), .B1(net_6242) );
SDFF_X2 inst_488 ( .SE(net_9540), .SI(net_8221), .Q(net_304), .D(net_304), .CK(net_13906) );
CLKBUF_X2 inst_14085 ( .A(net_14003), .Z(net_14004) );
DFF_X2 inst_7809 ( .Q(net_9822), .D(net_6460), .CK(net_11964) );
XNOR2_X2 inst_387 ( .A(net_2630), .ZN(net_2273), .B(net_2272) );
INV_X4 inst_5196 ( .ZN(net_4037), .A(net_1540) );
DFF_X1 inst_8666 ( .D(net_6773), .Q(net_111), .CK(net_12605) );
INV_X2 inst_7308 ( .A(net_9082), .ZN(net_9081) );
XNOR2_X2 inst_254 ( .ZN(net_4106), .A(net_3468), .B(net_2877) );
INV_X4 inst_6053 ( .ZN(net_642), .A(net_172) );
CLKBUF_X2 inst_15416 ( .A(net_14680), .Z(net_15335) );
INV_X4 inst_4601 ( .A(net_8812), .ZN(net_7720) );
CLKBUF_X2 inst_14769 ( .A(net_14687), .Z(net_14688) );
AOI22_X2 inst_9543 ( .B1(net_9906), .A1(net_9874), .B2(net_4969), .ZN(net_3778), .A2(net_2973) );
CLKBUF_X2 inst_12784 ( .A(net_12702), .Z(net_12703) );
DFF_X1 inst_8801 ( .QN(net_10235), .D(net_3980), .CK(net_10938) );
OAI211_X2 inst_2129 ( .C2(net_6774), .ZN(net_6719), .A(net_6345), .B(net_6083), .C1(net_512) );
OAI222_X2 inst_1412 ( .B2(net_7728), .A2(net_7727), .C2(net_7726), .ZN(net_5307), .B1(net_3947), .A1(net_2535), .C1(net_2292) );
INV_X4 inst_5750 ( .ZN(net_912), .A(net_739) );
CLKBUF_X2 inst_11273 ( .A(net_11191), .Z(net_11192) );
AOI221_X2 inst_9862 ( .A(net_6889), .B2(net_6888), .C2(net_6887), .ZN(net_6856), .B1(net_1126), .C1(x4449) );
OAI22_X2 inst_1181 ( .A1(net_7224), .A2(net_5139), .B2(net_5138), .ZN(net_5078), .B1(net_3538) );
CLKBUF_X2 inst_10957 ( .A(net_10875), .Z(net_10876) );
CLKBUF_X1 inst_8986 ( .A(x185142), .Z(x931) );
INV_X4 inst_6165 ( .A(net_9606), .ZN(net_758) );
CLKBUF_X2 inst_15382 ( .A(net_15300), .Z(net_15301) );
CLKBUF_X2 inst_13364 ( .A(net_13282), .Z(net_13283) );
CLKBUF_X2 inst_12774 ( .A(net_12692), .Z(net_12693) );
INV_X4 inst_5045 ( .A(net_3037), .ZN(net_1911) );
SDFF_X2 inst_661 ( .SI(net_9498), .Q(net_9498), .SE(net_3073), .CK(net_11879), .D(x1547) );
INV_X4 inst_6265 ( .A(net_10097), .ZN(net_5841) );
DFF_X2 inst_7416 ( .QN(net_9416), .D(net_8348), .CK(net_11707) );
OAI221_X2 inst_1548 ( .C1(net_10213), .C2(net_7295), .B2(net_7293), .ZN(net_7212), .B1(net_7211), .A(net_6852) );
CLKBUF_X2 inst_10817 ( .A(net_10640), .Z(net_10736) );
OAI211_X2 inst_2073 ( .C2(net_6778), .ZN(net_6776), .A(net_6377), .B(net_6145), .C1(net_411) );
HA_X1 inst_7346 ( .S(net_4588), .CO(net_4587), .B(net_4126), .A(net_2091) );
AOI221_X2 inst_9913 ( .ZN(net_6445), .B2(net_6443), .C2(net_6442), .A(net_5723), .B1(net_1418), .C1(net_709) );
DFF_X1 inst_8661 ( .Q(net_9121), .D(net_6911), .CK(net_10591) );
CLKBUF_X2 inst_11418 ( .A(net_11336), .Z(net_11337) );
CLKBUF_X2 inst_14255 ( .A(net_14173), .Z(net_14174) );
AOI22_X2 inst_9457 ( .A2(net_10269), .B2(net_8844), .ZN(net_3935), .A1(net_1148), .B1(net_1014) );
NAND2_X2 inst_3984 ( .ZN(net_3239), .A2(net_3238), .A1(net_2782) );
INV_X4 inst_4682 ( .ZN(net_5000), .A(net_4735) );
INV_X2 inst_7013 ( .A(net_2198), .ZN(net_1588) );
CLKBUF_X2 inst_11310 ( .A(net_10854), .Z(net_11229) );
XNOR2_X2 inst_419 ( .A(net_9654), .B(net_2928), .ZN(net_1405) );
CLKBUF_X2 inst_10899 ( .A(net_10817), .Z(net_10818) );
DFF_X2 inst_7488 ( .D(net_7992), .Q(net_207), .CK(net_12526) );
CLKBUF_X2 inst_12546 ( .A(net_12464), .Z(net_12465) );
CLKBUF_X2 inst_12098 ( .A(net_12016), .Z(net_12017) );
INV_X4 inst_5715 ( .ZN(net_999), .A(net_767) );
INV_X4 inst_6495 ( .ZN(net_864), .A(net_221) );
CLKBUF_X2 inst_15763 ( .A(net_13536), .Z(net_15682) );
DFF_X1 inst_8470 ( .Q(net_9271), .D(net_7981), .CK(net_15189) );
INV_X2 inst_6941 ( .A(net_4929), .ZN(net_1914) );
AND2_X4 inst_10462 ( .A1(net_10264), .ZN(net_1656), .A2(net_1334) );
DFF_X2 inst_7799 ( .Q(net_9914), .D(net_6493), .CK(net_13413) );
CLKBUF_X2 inst_10629 ( .A(net_10545), .Z(net_10548) );
CLKBUF_X2 inst_14298 ( .A(net_14216), .Z(net_14217) );
CLKBUF_X2 inst_14283 ( .A(net_14201), .Z(net_14202) );
CLKBUF_X2 inst_12018 ( .A(net_10870), .Z(net_11937) );
CLKBUF_X2 inst_12377 ( .A(net_11536), .Z(net_12296) );
DFF_X2 inst_7898 ( .QN(net_10460), .D(net_6004), .CK(net_11397) );
INV_X4 inst_5130 ( .ZN(net_1598), .A(net_1597) );
CLKBUF_X2 inst_12749 ( .A(net_12140), .Z(net_12668) );
CLKBUF_X2 inst_11160 ( .A(net_10793), .Z(net_11079) );
XOR2_X2 inst_34 ( .Z(net_2930), .A(net_700), .B(net_405) );
NAND2_X2 inst_3717 ( .A1(net_6289), .ZN(net_6011), .A2(net_5823) );
CLKBUF_X2 inst_15447 ( .A(net_15365), .Z(net_15366) );
CLKBUF_X2 inst_14629 ( .A(net_14547), .Z(net_14548) );
AOI22_X2 inst_9120 ( .A1(net_9705), .A2(net_6418), .ZN(net_6369), .B2(net_5263), .B1(net_145) );
XOR2_X2 inst_12 ( .Z(net_2874), .A(net_2873), .B(net_2291) );
CLKBUF_X2 inst_12690 ( .A(net_10821), .Z(net_12609) );
AOI221_X2 inst_9823 ( .B1(net_9865), .B2(net_9101), .A(net_6945), .C1(net_6944), .ZN(net_6928), .C2(net_236) );
INV_X4 inst_5489 ( .ZN(net_2622), .A(net_996) );
CLKBUF_X2 inst_13946 ( .A(net_11776), .Z(net_13865) );
DFF_X2 inst_7765 ( .Q(net_9714), .D(net_6540), .CK(net_13434) );
CLKBUF_X2 inst_14662 ( .A(net_11666), .Z(net_14581) );
AOI221_X2 inst_9856 ( .A(net_6889), .B2(net_6888), .C2(net_6887), .ZN(net_6862), .B1(net_1866), .C1(x4041) );
AOI221_X2 inst_9760 ( .B2(net_7770), .ZN(net_7698), .C1(net_7697), .A(net_7604), .B1(net_7514), .C2(net_2596) );
DFF_X1 inst_8682 ( .D(net_6736), .Q(net_150), .CK(net_13273) );
OAI222_X2 inst_1424 ( .ZN(net_3911), .A2(net_3910), .B2(net_3909), .C1(net_3908), .A1(net_3908), .C2(net_3907), .B1(net_2559) );
INV_X4 inst_5290 ( .A(net_2129), .ZN(net_1315) );
AOI21_X2 inst_10239 ( .ZN(net_8851), .B1(net_8320), .B2(net_8319), .A(net_8318) );
OAI222_X2 inst_1425 ( .A1(net_4509), .B2(net_3910), .C2(net_3907), .ZN(net_3906), .A2(net_3612), .C1(net_1515), .B1(net_1515) );
DFF_X1 inst_8585 ( .Q(net_9768), .D(net_7137), .CK(net_15620) );
NOR4_X2 inst_2307 ( .A2(net_9381), .ZN(net_7630), .A4(net_7629), .A1(net_7502), .A3(net_5370) );
OAI211_X2 inst_2198 ( .C1(net_7216), .C2(net_6542), .ZN(net_6509), .B(net_5607), .A(net_3679) );
CLKBUF_X2 inst_11611 ( .A(net_11529), .Z(net_11530) );
XNOR2_X2 inst_258 ( .ZN(net_4060), .A(net_3852), .B(net_1919) );
NOR2_X2 inst_2611 ( .A2(net_6846), .ZN(net_6245), .A1(net_1311) );
CLKBUF_X2 inst_13469 ( .A(net_11189), .Z(net_13388) );
INV_X4 inst_5004 ( .ZN(net_3095), .A(net_2182) );
AOI221_X2 inst_9926 ( .B2(net_5867), .A(net_5859), .ZN(net_5852), .C1(net_5851), .C2(net_4725), .B1(x5143) );
NOR3_X2 inst_2405 ( .A1(net_7345), .A3(net_7343), .ZN(net_7148), .A2(net_1305) );
CLKBUF_X2 inst_13126 ( .A(net_13044), .Z(net_13045) );
NOR2_X2 inst_2994 ( .A1(net_10253), .ZN(net_1474), .A2(net_1062) );
NOR2_X2 inst_3023 ( .A2(net_9206), .A1(net_9205), .ZN(net_1504) );
OAI22_X2 inst_1243 ( .A1(net_7241), .A2(net_4871), .B2(net_4870), .ZN(net_4867), .B1(net_372) );
CLKBUF_X2 inst_13155 ( .A(net_13073), .Z(net_13074) );
CLKBUF_X2 inst_14970 ( .A(net_14888), .Z(net_14889) );
CLKBUF_X2 inst_13074 ( .A(net_11235), .Z(net_12993) );
AOI22_X2 inst_9512 ( .B1(net_10298), .A1(net_9666), .A2(net_5966), .B2(net_4774), .ZN(net_3811) );
NAND4_X2 inst_3076 ( .A1(net_5168), .A2(net_5167), .A4(net_5166), .ZN(net_5165), .A3(net_5164) );
CLKBUF_X2 inst_10964 ( .A(net_10811), .Z(net_10883) );
SDFF_X2 inst_482 ( .SE(net_9540), .SI(net_8227), .Q(net_298), .D(net_298), .CK(net_13917) );
AND2_X2 inst_10514 ( .ZN(net_4976), .A2(net_4686), .A1(net_206) );
CLKBUF_X2 inst_14639 ( .A(net_10825), .Z(net_14558) );
AOI221_X2 inst_9804 ( .B1(net_9983), .A(net_7090), .B2(net_7089), .C2(net_7088), .ZN(net_6998), .C1(net_6821) );
NAND2_X2 inst_3534 ( .A2(net_9632), .A1(net_8973), .ZN(net_8052) );
NAND3_X2 inst_3276 ( .ZN(net_4069), .A2(net_4068), .A3(net_4067), .A1(net_3870) );
INV_X4 inst_5958 ( .A(net_5953), .ZN(net_552) );
AOI21_X2 inst_10230 ( .B2(net_10117), .ZN(net_2316), .A(net_2008), .B1(net_2007) );
OAI22_X2 inst_1093 ( .A1(net_9204), .A2(net_9064), .B2(net_6639), .ZN(net_6554), .B1(net_2814) );
NAND2_X2 inst_3996 ( .A2(net_3390), .ZN(net_3373), .A1(net_1681) );
INV_X2 inst_7059 ( .A(net_5314), .ZN(net_1279) );
SDFF_X2 inst_539 ( .D(net_9125), .SE(net_933), .CK(net_10907), .SI(x2890), .Q(x1313) );
DFF_X2 inst_7646 ( .D(net_6723), .QN(net_162), .CK(net_14247) );
CLKBUF_X2 inst_12915 ( .A(net_11355), .Z(net_12834) );
CLKBUF_X2 inst_11066 ( .A(net_10984), .Z(net_10985) );
CLKBUF_X2 inst_14728 ( .A(net_11743), .Z(net_14647) );
OR2_X2 inst_895 ( .A1(net_10188), .ZN(net_5775), .A2(net_5774) );
CLKBUF_X2 inst_11042 ( .A(net_10960), .Z(net_10961) );
AOI21_X2 inst_10054 ( .ZN(net_7144), .B2(net_6682), .B1(net_6254), .A(net_5427) );
CLKBUF_X2 inst_14516 ( .A(net_14434), .Z(net_14435) );
CLKBUF_X2 inst_10707 ( .A(net_10625), .Z(net_10626) );
OAI222_X2 inst_1430 ( .ZN(net_3152), .C2(net_3151), .B2(net_3151), .A2(net_2314), .A1(net_2303), .C1(net_1473), .B1(net_978) );
NAND3_X2 inst_3271 ( .A3(net_10453), .ZN(net_4146), .A1(net_4145), .A2(net_866) );
NAND3_X2 inst_3257 ( .ZN(net_4498), .A1(net_4234), .A2(net_3357), .A3(net_3356) );
CLKBUF_X2 inst_10759 ( .A(net_10677), .Z(net_10678) );
INV_X4 inst_6583 ( .A(net_9833), .ZN(net_690) );
CLKBUF_X2 inst_14081 ( .A(net_13999), .Z(net_14000) );
CLKBUF_X2 inst_11498 ( .A(net_11416), .Z(net_11417) );
AOI21_X2 inst_10034 ( .B1(net_10280), .ZN(net_7865), .A(net_6678), .B2(net_263) );
NOR4_X2 inst_2341 ( .ZN(net_3094), .A4(net_2704), .A1(net_2547), .A2(net_2410), .A3(net_1219) );
INV_X4 inst_5526 ( .ZN(net_1247), .A(net_956) );
CLKBUF_X2 inst_10685 ( .A(net_10603), .Z(net_10604) );
AND2_X2 inst_10616 ( .ZN(net_2509), .A2(net_1740), .A1(net_829) );
AOI221_X2 inst_9979 ( .C1(net_10182), .B1(net_9741), .B2(net_6442), .ZN(net_4219), .C2(net_4217), .A(net_3590) );
NAND2_X2 inst_4122 ( .ZN(net_2335), .A1(net_2334), .A2(net_1620) );
CLKBUF_X2 inst_12557 ( .A(net_11664), .Z(net_12476) );
OR2_X4 inst_763 ( .ZN(net_4742), .A1(net_4324), .A2(net_4322) );
NOR4_X2 inst_2330 ( .ZN(net_5218), .A2(net_5217), .A4(net_5216), .A3(net_4549), .A1(net_3534) );
DFF_X2 inst_7377 ( .Q(net_9369), .D(net_8673), .CK(net_14186) );
NAND2_X2 inst_3636 ( .A2(net_7557), .ZN(net_7441), .A1(net_564) );
CLKBUF_X2 inst_13184 ( .A(net_13102), .Z(net_13103) );
CLKBUF_X2 inst_11069 ( .A(net_10987), .Z(net_10988) );
CLKBUF_X2 inst_14018 ( .A(net_13019), .Z(net_13937) );
AOI221_X2 inst_9901 ( .B1(net_9886), .B2(net_9101), .A(net_6945), .C2(net_6944), .ZN(net_6793), .C1(net_257) );
AND4_X4 inst_10324 ( .ZN(net_3535), .A2(net_3534), .A3(net_3533), .A4(net_3532), .A1(net_2947) );
CLKBUF_X2 inst_13754 ( .A(net_12503), .Z(net_13673) );
AOI22_X2 inst_9189 ( .A1(net_9861), .B1(net_9762), .A2(net_8042), .ZN(net_6125), .B2(net_6120) );
SDFF_X2 inst_537 ( .D(net_9139), .SE(net_933), .CK(net_10982), .SI(x2027), .Q(x1187) );
INV_X4 inst_4797 ( .A(net_3727), .ZN(net_3662) );
INV_X4 inst_6082 ( .ZN(net_928), .A(net_189) );
DFF_X1 inst_8482 ( .QN(net_9628), .D(net_7948), .CK(net_15022) );
OR2_X4 inst_826 ( .A2(net_10458), .ZN(net_1675), .A1(net_1094) );
AOI22_X2 inst_9343 ( .B1(net_9819), .A2(net_5766), .B2(net_5765), .ZN(net_5609), .A1(net_257) );
NAND2_X2 inst_4002 ( .ZN(net_4456), .A2(net_3390), .A1(net_2221) );
INV_X4 inst_5069 ( .A(net_2906), .ZN(net_2871) );
CLKBUF_X2 inst_14009 ( .A(net_13927), .Z(net_13928) );
AND3_X4 inst_10362 ( .A1(net_6203), .ZN(net_4655), .A2(net_4233), .A3(net_4226) );
XNOR2_X2 inst_159 ( .ZN(net_5981), .A(net_5980), .B(net_1744) );
INV_X2 inst_7042 ( .ZN(net_1369), .A(net_1368) );
CLKBUF_X2 inst_13220 ( .A(net_12548), .Z(net_13139) );
AOI22_X2 inst_9572 ( .B2(net_6443), .A2(net_6442), .ZN(net_3735), .A1(net_989), .B1(net_893) );
CLKBUF_X2 inst_14977 ( .A(net_14895), .Z(net_14896) );
INV_X2 inst_7141 ( .A(net_858), .ZN(net_819) );
CLKBUF_X2 inst_15281 ( .A(net_15199), .Z(net_15200) );
CLKBUF_X2 inst_15232 ( .A(net_13901), .Z(net_15151) );
CLKBUF_X2 inst_14341 ( .A(net_14259), .Z(net_14260) );
INV_X4 inst_5759 ( .A(net_1354), .ZN(net_938) );
CLKBUF_X2 inst_13657 ( .A(net_13575), .Z(net_13576) );
CLKBUF_X2 inst_11005 ( .A(net_10923), .Z(net_10924) );
CLKBUF_X2 inst_10786 ( .A(net_10704), .Z(net_10705) );
DFF_X1 inst_8431 ( .D(net_8641), .QN(net_277), .CK(net_14950) );
INV_X4 inst_6318 ( .A(net_10286), .ZN(net_422) );
DFF_X2 inst_7379 ( .D(net_8642), .QN(net_276), .CK(net_14929) );
DFF_X1 inst_8863 ( .Q(net_96), .CK(net_11864), .D(x3320) );
NAND2_X2 inst_3950 ( .ZN(net_3666), .A2(net_3488), .A1(net_917) );
NAND2_X2 inst_4288 ( .A2(net_9735), .ZN(net_1793), .A1(net_898) );
CLKBUF_X2 inst_15491 ( .A(net_15409), .Z(net_15410) );
OR2_X2 inst_869 ( .ZN(net_7712), .A1(net_7547), .A2(net_7416) );
CLKBUF_X2 inst_10671 ( .A(net_10589), .Z(net_10590) );
DFF_X2 inst_8339 ( .D(net_3099), .QN(net_132), .CK(net_14271) );
XOR2_X2 inst_19 ( .Z(net_2770), .B(net_2563), .A(net_1248) );
NOR2_X2 inst_2646 ( .A1(net_9354), .ZN(net_7015), .A2(net_5402) );
CLKBUF_X2 inst_13623 ( .A(net_13541), .Z(net_13542) );
CLKBUF_X2 inst_11509 ( .A(net_11427), .Z(net_11428) );
AND3_X2 inst_10378 ( .A1(net_3131), .ZN(net_2735), .A2(net_1153), .A3(net_841) );
CLKBUF_X2 inst_13599 ( .A(net_13517), .Z(net_13518) );
INV_X4 inst_6543 ( .A(net_9928), .ZN(net_902) );
CLKBUF_X2 inst_13229 ( .A(net_13147), .Z(net_13148) );
AOI221_X2 inst_9753 ( .ZN(net_7773), .B2(net_7770), .A(net_7675), .C2(net_4464), .B1(net_3371), .C1(net_2857) );
NAND2_X2 inst_4268 ( .A2(net_9246), .A1(net_9245), .ZN(net_2934) );
CLKBUF_X2 inst_14170 ( .A(net_14088), .Z(net_14089) );
NAND2_X2 inst_3830 ( .ZN(net_7726), .A2(net_4442), .A1(net_691) );
CLKBUF_X2 inst_13649 ( .A(net_13567), .Z(net_13568) );
AOI221_X2 inst_9849 ( .A(net_6889), .B2(net_6888), .C2(net_6887), .ZN(net_6869), .B1(net_5825), .C1(x5548) );
NAND3_X2 inst_3267 ( .A1(net_6203), .ZN(net_4841), .A2(net_4233), .A3(net_4227) );
CLKBUF_X2 inst_12287 ( .A(net_12205), .Z(net_12206) );
OAI221_X2 inst_1686 ( .B1(net_7198), .C2(net_5642), .ZN(net_5476), .C1(net_5475), .B2(net_4905), .A(net_3731) );
NAND3_X2 inst_3205 ( .ZN(net_6935), .A1(net_6416), .A3(net_3803), .A2(net_3751) );
CLKBUF_X2 inst_14315 ( .A(net_13883), .Z(net_14234) );
AND2_X2 inst_10541 ( .A1(net_9206), .ZN(net_3966), .A2(net_3513) );
INV_X4 inst_6048 ( .A(net_9982), .ZN(net_510) );
CLKBUF_X2 inst_15732 ( .A(net_15650), .Z(net_15651) );
SDFF_X2 inst_612 ( .QN(net_10197), .D(net_4413), .SE(net_3684), .SI(net_661), .CK(net_10847) );
CLKBUF_X2 inst_12505 ( .A(net_12423), .Z(net_12424) );
OAI21_X2 inst_1789 ( .ZN(net_7593), .A(net_7509), .B2(net_1259), .B1(net_1001) );
OAI221_X2 inst_1692 ( .C1(net_7203), .ZN(net_5466), .B2(net_4477), .C2(net_4455), .A(net_3507), .B1(net_978) );
INV_X4 inst_6185 ( .A(net_10372), .ZN(net_473) );
CLKBUF_X2 inst_14664 ( .A(net_10979), .Z(net_14583) );
INV_X2 inst_7192 ( .ZN(net_914), .A(net_178) );
CLKBUF_X2 inst_14832 ( .A(net_14750), .Z(net_14751) );
CLKBUF_X2 inst_15803 ( .A(net_15721), .Z(net_15722) );
NAND2_X2 inst_3986 ( .A1(net_9853), .A2(net_6413), .ZN(net_3190) );
DFF_X2 inst_7627 ( .D(net_6696), .QN(net_175), .CK(net_14957) );
AOI22_X2 inst_9437 ( .A1(net_6892), .B2(net_6625), .ZN(net_6251), .B1(net_4304), .A2(net_3971) );
NAND2_X2 inst_3441 ( .A1(net_9447), .ZN(net_8887), .A2(net_8479) );
INV_X2 inst_6955 ( .A(net_3712), .ZN(net_1879) );
CLKBUF_X2 inst_13137 ( .A(net_13055), .Z(net_13056) );
CLKBUF_X2 inst_14328 ( .A(net_14246), .Z(net_14247) );
INV_X2 inst_7275 ( .A(net_8948), .ZN(net_8947) );
CLKBUF_X2 inst_10819 ( .A(net_10737), .Z(net_10738) );
CLKBUF_X2 inst_12332 ( .A(net_12250), .Z(net_12251) );
CLKBUF_X2 inst_14535 ( .A(net_14453), .Z(net_14454) );
AOI22_X2 inst_9413 ( .A1(net_10182), .ZN(net_4658), .A2(net_4656), .B2(net_4655), .B1(x5077) );
NOR3_X2 inst_2455 ( .A1(net_3529), .A3(net_2984), .A2(net_2564), .ZN(net_2009) );
DFF_X2 inst_8000 ( .QN(net_10124), .D(net_5512), .CK(net_12361) );
CLKBUF_X2 inst_12923 ( .A(net_12841), .Z(net_12842) );
CLKBUF_X2 inst_11535 ( .A(net_11453), .Z(net_11454) );
AND2_X2 inst_10575 ( .ZN(net_3312), .A1(net_3032), .A2(net_2834) );
CLKBUF_X2 inst_15690 ( .A(net_15608), .Z(net_15609) );
CLKBUF_X2 inst_15250 ( .A(net_15168), .Z(net_15169) );
INV_X2 inst_6724 ( .ZN(net_7778), .A(net_7744) );
CLKBUF_X2 inst_11581 ( .A(net_11092), .Z(net_11500) );
INV_X4 inst_4828 ( .A(net_7157), .ZN(net_5575) );
INV_X4 inst_5218 ( .A(net_1515), .ZN(net_1514) );
INV_X4 inst_5389 ( .A(net_2294), .ZN(net_1188) );
CLKBUF_X2 inst_12516 ( .A(net_11456), .Z(net_12435) );
INV_X4 inst_4860 ( .ZN(net_6443), .A(net_4274) );
CLKBUF_X2 inst_14923 ( .A(net_14841), .Z(net_14842) );
CLKBUF_X2 inst_12226 ( .A(net_11667), .Z(net_12145) );
INV_X2 inst_6770 ( .ZN(net_6032), .A(net_5857) );
OAI222_X2 inst_1344 ( .B1(net_7660), .A2(net_7659), .C2(net_7658), .ZN(net_7578), .B2(net_7419), .A1(net_6173), .C1(net_1825) );
OAI221_X2 inst_1460 ( .C1(net_8981), .B2(net_7974), .C2(net_7973), .ZN(net_7964), .A(net_7963), .B1(net_3108) );
OAI211_X2 inst_2287 ( .C1(net_7297), .C2(net_6548), .ZN(net_6180), .B(net_5404), .A(net_3679) );
OR2_X2 inst_885 ( .A2(net_7038), .ZN(net_6220), .A1(net_6219) );
NOR2_X2 inst_2630 ( .A2(net_7721), .ZN(net_6186), .A1(net_5954) );
CLKBUF_X2 inst_15422 ( .A(net_15340), .Z(net_15341) );
INV_X4 inst_5803 ( .ZN(net_2865), .A(net_1733) );
CLKBUF_X2 inst_10748 ( .A(net_10666), .Z(net_10667) );
OAI221_X2 inst_1443 ( .B2(net_9602), .ZN(net_8567), .B1(net_8566), .C1(net_8565), .C2(net_8494), .A(net_3902) );
OAI22_X2 inst_1028 ( .A2(net_8036), .B2(net_8018), .ZN(net_7984), .A1(net_4953), .B1(net_331) );
INV_X4 inst_5891 ( .ZN(net_1378), .A(net_842) );
AOI21_X2 inst_10107 ( .B2(net_10236), .ZN(net_5187), .B1(net_3270), .A(net_3024) );
NAND2_X2 inst_3935 ( .A2(net_3698), .ZN(net_3691), .A1(net_564) );
NAND2_X2 inst_3610 ( .ZN(net_7256), .A2(net_6876), .A1(net_6592) );
CLKBUF_X2 inst_13097 ( .A(net_10971), .Z(net_13016) );
NOR2_X2 inst_2999 ( .A1(net_10465), .ZN(net_1700), .A2(net_703) );
AOI22_X2 inst_9645 ( .A2(net_2783), .B2(net_2782), .ZN(net_2781), .A1(net_2780), .B1(net_1189) );
OAI22_X2 inst_1271 ( .ZN(net_4754), .A1(net_4753), .A2(net_4752), .B2(net_4751), .B1(net_1300) );
CLKBUF_X2 inst_12822 ( .A(net_12740), .Z(net_12741) );
DFF_X2 inst_8351 ( .QN(net_10164), .D(net_2813), .CK(net_12242) );
CLKBUF_X2 inst_12110 ( .A(net_12028), .Z(net_12029) );
NOR4_X2 inst_2321 ( .A2(net_9949), .ZN(net_6636), .A3(net_6060), .A4(net_5791), .A1(net_3744) );
DFF_X2 inst_8188 ( .QN(net_10245), .D(net_5194), .CK(net_12196) );
INV_X4 inst_5956 ( .ZN(net_1363), .A(net_554) );
CLKBUF_X2 inst_13927 ( .A(net_13845), .Z(net_13846) );
NAND2_X2 inst_4156 ( .A1(net_2950), .A2(net_2034), .ZN(net_2030) );
INV_X4 inst_5305 ( .ZN(net_2198), .A(net_1295) );
AOI221_X2 inst_9875 ( .B1(net_9782), .B2(net_9097), .A(net_6940), .C2(net_6939), .ZN(net_6826), .C1(net_252) );
AOI221_X2 inst_9928 ( .B2(net_5867), .A(net_5859), .ZN(net_5848), .C1(net_5847), .C2(net_4725), .B1(x5003) );
XNOR2_X2 inst_200 ( .ZN(net_4987), .B(net_4986), .A(net_4709) );
NAND2_X1 inst_4425 ( .ZN(net_2616), .A1(net_1959), .A2(net_1078) );
CLKBUF_X2 inst_11986 ( .A(net_11571), .Z(net_11905) );
AOI222_X1 inst_9727 ( .C1(net_9963), .A2(net_5173), .B2(net_4694), .ZN(net_3913), .A1(net_3032), .C2(net_2541), .B1(net_228) );
MUX2_X1 inst_4461 ( .S(net_6041), .A(net_285), .B(x5850), .Z(x268) );
INV_X4 inst_6626 ( .ZN(net_8974), .A(net_8972) );
CLKBUF_X2 inst_14332 ( .A(net_12946), .Z(net_14251) );
NAND2_X2 inst_4373 ( .A2(net_10265), .ZN(net_2513), .A1(net_1063) );
AOI221_X2 inst_9939 ( .B2(net_5867), .A(net_5859), .ZN(net_5826), .C1(net_5825), .C2(net_4725), .B1(x5548) );
AOI22_X2 inst_9198 ( .A1(net_9888), .B1(net_9789), .A2(net_8042), .B2(net_8041), .ZN(net_6115) );
DFF_X2 inst_7407 ( .QN(net_9399), .D(net_8366), .CK(net_11762) );
CLKBUF_X2 inst_12343 ( .A(net_11394), .Z(net_12262) );
OAI21_X2 inst_1750 ( .ZN(net_8650), .A(net_8648), .B1(net_8647), .B2(net_8616) );
CLKBUF_X2 inst_10807 ( .A(net_10725), .Z(net_10726) );
INV_X4 inst_5242 ( .ZN(net_6514), .A(net_1467) );
OAI211_X2 inst_2236 ( .C1(net_7224), .C2(net_6480), .ZN(net_6468), .B(net_5679), .A(net_3679) );
NAND2_X4 inst_3368 ( .ZN(net_9096), .A1(net_4034), .A2(net_3895) );
INV_X2 inst_7307 ( .A(net_9078), .ZN(net_9077) );
OAI221_X2 inst_1553 ( .C2(net_7295), .B2(net_7293), .B1(net_7231), .ZN(net_7205), .A(net_6830), .C1(net_1492) );
CLKBUF_X2 inst_13038 ( .A(net_12956), .Z(net_12957) );
CLKBUF_X2 inst_13937 ( .A(net_13855), .Z(net_13856) );
CLKBUF_X2 inst_15322 ( .A(net_15240), .Z(net_15241) );
AND2_X4 inst_10458 ( .ZN(net_1649), .A2(net_1386), .A1(net_1362) );
AOI21_X2 inst_10155 ( .ZN(net_4130), .A(net_3661), .B2(net_3279), .B1(net_2627) );
DFF_X2 inst_7758 ( .QN(net_9209), .D(net_6441), .CK(net_11315) );
DFF_X2 inst_7593 ( .QN(net_10463), .D(net_7433), .CK(net_13666) );
OAI221_X2 inst_1635 ( .C1(net_10312), .B1(net_7136), .A(net_5637), .C2(net_5591), .ZN(net_5571), .B2(net_4902) );
NAND2_X2 inst_4130 ( .ZN(net_2602), .A1(net_2247), .A2(net_940) );
CLKBUF_X2 inst_12121 ( .A(net_12039), .Z(net_12040) );
AOI22_X2 inst_9569 ( .B1(net_9801), .A2(net_6443), .A1(net_6054), .ZN(net_3750), .B2(net_2556) );
CLKBUF_X2 inst_13102 ( .A(net_13020), .Z(net_13021) );
OAI221_X2 inst_1500 ( .C2(net_9063), .B2(net_9056), .ZN(net_7361), .C1(net_7219), .A(net_6999), .B1(net_843) );
CLKBUF_X2 inst_14737 ( .A(net_14655), .Z(net_14656) );
CLKBUF_X2 inst_11731 ( .A(net_11649), .Z(net_11650) );
CLKBUF_X2 inst_12294 ( .A(net_10764), .Z(net_12213) );
NOR2_X2 inst_2805 ( .ZN(net_4103), .A2(net_2982), .A1(net_2711) );
INV_X4 inst_6438 ( .A(net_9217), .ZN(net_2496) );
NAND2_X2 inst_3499 ( .ZN(net_8695), .A1(net_8186), .A2(net_8185) );
NOR2_X2 inst_2932 ( .A2(net_6960), .ZN(net_2400), .A1(net_730) );
OR2_X2 inst_893 ( .A1(net_10482), .ZN(net_6256), .A2(net_5806) );
INV_X2 inst_6917 ( .ZN(net_2585), .A(net_1977) );
AOI22_X2 inst_9483 ( .B1(net_9914), .A1(net_9882), .B2(net_4969), .ZN(net_3840), .A2(net_2973) );
NAND4_X2 inst_3048 ( .ZN(net_7405), .A2(net_7068), .A4(net_7067), .A3(net_6258), .A1(net_2946) );
CLKBUF_X2 inst_10911 ( .A(net_10829), .Z(net_10830) );
INV_X4 inst_4854 ( .ZN(net_3268), .A(net_3267) );
DFF_X2 inst_8128 ( .Q(net_9837), .D(net_5132), .CK(net_14289) );
CLKBUF_X2 inst_15711 ( .A(net_11476), .Z(net_15630) );
CLKBUF_X2 inst_15435 ( .A(net_13738), .Z(net_15354) );
CLKBUF_X2 inst_13862 ( .A(net_10782), .Z(net_13781) );
SDFF_X2 inst_569 ( .D(net_9144), .SE(net_933), .CK(net_11024), .SI(x1743), .Q(x1142) );
NAND2_X4 inst_3346 ( .ZN(net_8519), .A1(net_8465), .A2(net_8464) );
NOR2_X2 inst_2992 ( .A1(net_10434), .ZN(net_2402), .A2(net_530) );
AOI22_X2 inst_9209 ( .A1(net_9869), .B1(net_9770), .B2(net_6120), .A2(net_6109), .ZN(net_6102) );
CLKBUF_X2 inst_12763 ( .A(net_12026), .Z(net_12682) );
OAI22_X2 inst_1080 ( .A1(net_7157), .ZN(net_6579), .A2(net_5919), .B2(net_5917), .B1(net_410) );
INV_X4 inst_6405 ( .A(net_10392), .ZN(net_389) );
CLKBUF_X2 inst_15440 ( .A(net_14628), .Z(net_15359) );
CLKBUF_X2 inst_14730 ( .A(net_14648), .Z(net_14649) );
NOR3_X2 inst_2374 ( .A1(net_8190), .ZN(net_8123), .A2(net_8122), .A3(net_7936) );
CLKBUF_X2 inst_14451 ( .A(net_11187), .Z(net_14370) );
DFF_X2 inst_7473 ( .Q(net_10063), .D(net_8038), .CK(net_11185) );
CLKBUF_X2 inst_15723 ( .A(net_15641), .Z(net_15642) );
CLKBUF_X2 inst_12554 ( .A(net_12472), .Z(net_12473) );
OAI22_X2 inst_1103 ( .A1(net_9190), .A2(net_6299), .B2(net_6298), .ZN(net_6204), .B1(net_5100) );
INV_X4 inst_6535 ( .A(net_10051), .ZN(net_4747) );
DFF_X1 inst_8620 ( .Q(net_9666), .D(net_7104), .CK(net_14257) );
CLKBUF_X2 inst_10678 ( .A(net_10556), .Z(net_10597) );
AOI22_X2 inst_9256 ( .B2(net_6140), .A2(net_6109), .ZN(net_6050), .A1(net_3807), .B1(net_1932) );
DFF_X2 inst_7494 ( .D(net_8005), .Q(net_204), .CK(net_12517) );
SDFF_X2 inst_549 ( .SI(net_9358), .Q(net_9358), .D(net_9156), .SE(net_7248), .CK(net_15351) );
NAND2_X2 inst_4329 ( .ZN(net_1631), .A2(net_870), .A1(net_699) );
CLKBUF_X2 inst_12566 ( .A(net_12484), .Z(net_12485) );
NAND2_X2 inst_4220 ( .ZN(net_2711), .A2(net_1263), .A1(net_929) );
INV_X4 inst_4708 ( .ZN(net_4739), .A(net_4623) );
SDFF_X2 inst_522 ( .Q(net_9339), .D(net_9339), .SI(net_9331), .SE(net_7588), .CK(net_14688) );
INV_X4 inst_5202 ( .ZN(net_1938), .A(net_1597) );
CLKBUF_X2 inst_13617 ( .A(net_13535), .Z(net_13536) );
INV_X4 inst_5040 ( .ZN(net_5515), .A(net_1925) );
CLKBUF_X2 inst_14458 ( .A(net_14161), .Z(net_14377) );
CLKBUF_X2 inst_12408 ( .A(net_12326), .Z(net_12327) );
AOI22_X2 inst_9037 ( .ZN(net_7429), .A2(net_6961), .B1(net_6960), .B2(net_5255), .A1(net_5251) );
AOI221_X2 inst_9842 ( .A(net_6889), .B2(net_6888), .C2(net_6887), .ZN(net_6876), .B1(net_5839), .C1(x3889) );
INV_X4 inst_6231 ( .A(net_9294), .ZN(net_2545) );
NOR2_X2 inst_2809 ( .A2(net_2680), .ZN(net_2658), .A1(net_2657) );
CLKBUF_X2 inst_15147 ( .A(net_15065), .Z(net_15066) );
CLKBUF_X2 inst_14011 ( .A(net_13929), .Z(net_13930) );
AOI22_X2 inst_9654 ( .B1(net_3194), .A1(net_2355), .B2(net_2325), .ZN(net_2229), .A2(net_1531) );
CLKBUF_X2 inst_13776 ( .A(net_13459), .Z(net_13695) );
CLKBUF_X2 inst_12478 ( .A(net_12396), .Z(net_12397) );
CLKBUF_X2 inst_13141 ( .A(net_13059), .Z(net_13060) );
INV_X4 inst_6331 ( .A(net_9273), .ZN(net_7875) );
CLKBUF_X2 inst_12797 ( .A(net_12367), .Z(net_12716) );
AOI222_X1 inst_9737 ( .B2(net_10507), .C2(net_10505), .A2(net_10504), .B1(net_10494), .C1(net_10492), .A1(net_10491), .ZN(net_1251) );
NOR2_X2 inst_2673 ( .ZN(net_5286), .A2(net_4783), .A1(net_3298) );
CLKBUF_X2 inst_13592 ( .A(net_13510), .Z(net_13511) );
OAI221_X2 inst_1618 ( .B1(net_10315), .C1(net_7127), .A(net_6546), .ZN(net_5592), .B2(net_5591), .C2(net_4902) );
INV_X4 inst_5062 ( .ZN(net_2222), .A(net_1871) );
INV_X2 inst_6936 ( .ZN(net_1924), .A(net_1923) );
CLKBUF_X2 inst_14166 ( .A(net_13899), .Z(net_14085) );
OAI211_X2 inst_2126 ( .C2(net_6778), .ZN(net_6722), .A(net_6369), .B(net_6142), .C1(net_319) );
AND2_X2 inst_10484 ( .ZN(net_8437), .A2(net_8407), .A1(net_8182) );
INV_X2 inst_6911 ( .A(net_2619), .ZN(net_2228) );
AOI22_X2 inst_9144 ( .A1(net_9697), .A2(net_6402), .ZN(net_6341), .B2(net_5263), .B1(net_137) );
DFF_X2 inst_7776 ( .Q(net_9793), .D(net_6525), .CK(net_15236) );
CLKBUF_X2 inst_11131 ( .A(net_11049), .Z(net_11050) );
AOI22_X2 inst_8997 ( .B1(net_9501), .A1(net_9493), .ZN(net_8501), .A2(net_8476), .B2(net_8473) );
NOR2_X2 inst_2765 ( .A2(net_9036), .ZN(net_3301), .A1(net_1575) );
NAND2_X2 inst_3600 ( .ZN(net_7266), .A2(net_6878), .A1(net_6605) );
CLKBUF_X2 inst_14779 ( .A(net_14697), .Z(net_14698) );
INV_X4 inst_6493 ( .A(net_9548), .ZN(net_356) );
XNOR2_X2 inst_219 ( .ZN(net_4604), .B(net_4603), .A(net_4451) );
CLKBUF_X2 inst_15699 ( .A(net_15617), .Z(net_15618) );
OR3_X2 inst_719 ( .ZN(net_3634), .A2(net_2935), .A3(net_2934), .A1(net_2441) );
AOI21_X2 inst_10195 ( .B1(net_3875), .ZN(net_3162), .A(net_3161), .B2(net_3160) );
NAND2_X2 inst_4166 ( .A1(net_3885), .ZN(net_2901), .A2(net_1384) );
INV_X4 inst_4881 ( .ZN(net_2986), .A(net_2781) );
CLKBUF_X2 inst_15320 ( .A(net_14158), .Z(net_15239) );
CLKBUF_X1 inst_8980 ( .A(x185142), .Z(x898) );
DFF_X1 inst_8695 ( .D(net_6709), .QN(net_182), .CK(net_12084) );
NAND2_X2 inst_3868 ( .ZN(net_4364), .A2(net_4227), .A1(net_4083) );
OAI22_X2 inst_1134 ( .A1(net_7203), .A2(net_5151), .B2(net_5150), .ZN(net_5144), .B1(net_710) );
INV_X4 inst_5501 ( .ZN(net_1815), .A(net_984) );
OAI211_X2 inst_2204 ( .C1(net_7245), .ZN(net_6502), .C2(net_6501), .B(net_5644), .A(net_3507) );
OAI221_X2 inst_1609 ( .B1(net_10205), .C1(net_7108), .A(net_6546), .B2(net_5642), .ZN(net_5627), .C2(net_4905) );
NAND2_X2 inst_4105 ( .ZN(net_2377), .A1(net_2149), .A2(net_1680) );
NAND2_X2 inst_3546 ( .ZN(net_8949), .A2(net_7822), .A1(net_7279) );
XNOR2_X2 inst_408 ( .A(net_9371), .B(net_7848), .ZN(net_2725) );
INV_X4 inst_5748 ( .A(net_1429), .ZN(net_740) );
OAI22_X2 inst_1144 ( .A1(net_7186), .A2(net_5134), .B2(net_5133), .ZN(net_5129), .B1(net_417) );
INV_X4 inst_4701 ( .ZN(net_4794), .A(net_4793) );
INV_X4 inst_5165 ( .ZN(net_1880), .A(net_1568) );
INV_X4 inst_5644 ( .ZN(net_1984), .A(net_844) );
CLKBUF_X2 inst_12419 ( .A(net_12337), .Z(net_12338) );
CLKBUF_X2 inst_11212 ( .A(net_10565), .Z(net_11131) );
INV_X4 inst_5366 ( .ZN(net_1216), .A(net_1215) );
INV_X4 inst_6426 ( .A(net_9837), .ZN(net_381) );
INV_X4 inst_5551 ( .A(net_4997), .ZN(net_2183) );
NOR2_X2 inst_2568 ( .ZN(net_7493), .A2(net_7319), .A1(net_6232) );
INV_X4 inst_5596 ( .A(net_5794), .ZN(net_1202) );
OAI211_X2 inst_2295 ( .ZN(net_4385), .A(net_4094), .B(net_3451), .C2(net_1297), .C1(net_1132) );
CLKBUF_X2 inst_13021 ( .A(net_12939), .Z(net_12940) );
CLKBUF_X2 inst_11591 ( .A(net_11509), .Z(net_11510) );
CLKBUF_X2 inst_10719 ( .A(net_10637), .Z(net_10638) );
NAND2_X2 inst_3814 ( .A1(net_10083), .A2(net_4534), .ZN(net_4524) );
CLKBUF_X2 inst_12968 ( .A(net_12886), .Z(net_12887) );
DFF_X1 inst_8498 ( .Q(net_9857), .D(net_7838), .CK(net_15655) );
CLKBUF_X2 inst_15605 ( .A(net_15523), .Z(net_15524) );
NOR2_X1 inst_3028 ( .ZN(net_3039), .A1(net_2964), .A2(net_2955) );
NAND2_X2 inst_3532 ( .A2(net_9624), .A1(net_8975), .ZN(net_8054) );
AOI22_X2 inst_9190 ( .A1(net_9880), .B1(net_9781), .A2(net_8042), .B2(net_6129), .ZN(net_6124) );
AOI22_X2 inst_9432 ( .A1(net_9854), .B1(net_6834), .ZN(net_4497), .A2(net_4495), .B2(net_4494) );
NAND2_X2 inst_3854 ( .A1(net_6349), .ZN(net_4185), .A2(net_4182) );
DFF_X2 inst_7871 ( .QN(net_10141), .D(net_6035), .CK(net_13492) );
CLKBUF_X2 inst_10881 ( .A(net_10641), .Z(net_10800) );
NAND2_X2 inst_3514 ( .A2(net_8136), .ZN(net_8134), .A1(net_8057) );
CLKBUF_X2 inst_10826 ( .A(net_10744), .Z(net_10745) );
OAI221_X2 inst_1530 ( .B1(net_10204), .B2(net_7295), .C2(net_7293), .ZN(net_7242), .C1(net_7241), .A(net_6807) );
INV_X2 inst_7089 ( .A(net_4007), .ZN(net_1122) );
OAI221_X2 inst_1510 ( .C1(net_10411), .B2(net_9063), .C2(net_9056), .ZN(net_7350), .B1(net_7243), .A(net_7005) );
XNOR2_X2 inst_121 ( .B(net_9423), .ZN(net_7616), .A(net_6316) );
INV_X4 inst_5421 ( .ZN(net_6289), .A(net_1135) );
CLKBUF_X2 inst_12449 ( .A(net_10712), .Z(net_12368) );
OAI22_X2 inst_1065 ( .A2(net_7036), .B2(net_7035), .ZN(net_6964), .A1(net_1751), .B1(net_1750) );
DFF_X2 inst_7635 ( .D(net_6757), .QN(net_126), .CK(net_13453) );
CLKBUF_X2 inst_12002 ( .A(net_11879), .Z(net_11921) );
INV_X4 inst_6308 ( .A(net_10500), .ZN(net_425) );
CLKBUF_X2 inst_11599 ( .A(net_11517), .Z(net_11518) );
NAND2_X2 inst_4119 ( .A1(net_4558), .ZN(net_2339), .A2(net_1609) );
INV_X4 inst_5948 ( .A(net_693), .ZN(net_560) );
NAND2_X2 inst_4332 ( .A1(net_10368), .ZN(net_2768), .A2(net_1956) );
CLKBUF_X2 inst_13766 ( .A(net_12747), .Z(net_13685) );
AOI22_X2 inst_9340 ( .B1(net_9816), .A1(net_6823), .A2(net_5766), .B2(net_5765), .ZN(net_5612) );
CLKBUF_X2 inst_13318 ( .A(net_11244), .Z(net_13237) );
CLKBUF_X2 inst_10955 ( .A(net_10873), .Z(net_10874) );
AOI21_X2 inst_10076 ( .B2(net_10238), .A(net_10237), .ZN(net_5944), .B1(net_1506) );
INV_X4 inst_6282 ( .A(net_10432), .ZN(net_2302) );
CLKBUF_X2 inst_12111 ( .A(net_12029), .Z(net_12030) );
CLKBUF_X2 inst_14348 ( .A(net_11037), .Z(net_14267) );
AOI22_X2 inst_9495 ( .B1(net_10388), .A1(net_9886), .B2(net_4062), .ZN(net_3828), .A2(net_2973) );
INV_X4 inst_5353 ( .ZN(net_5513), .A(net_1234) );
CLKBUF_X2 inst_14189 ( .A(net_14107), .Z(net_14108) );
CLKBUF_X2 inst_13876 ( .A(net_13794), .Z(net_13795) );
AOI221_X2 inst_9981 ( .C1(net_10185), .B2(net_6442), .C2(net_4217), .ZN(net_4216), .A(net_3585), .B1(net_1429) );
CLKBUF_X2 inst_12586 ( .A(net_12504), .Z(net_12505) );
INV_X4 inst_4671 ( .A(net_9539), .ZN(net_5818) );
INV_X4 inst_6244 ( .A(net_9210), .ZN(net_1535) );
DFF_X1 inst_8753 ( .Q(net_10537), .D(net_10536), .CK(net_10966) );
NAND2_X2 inst_4174 ( .ZN(net_2946), .A2(net_2202), .A1(net_1960) );
SDFF_X2 inst_530 ( .SI(net_9340), .Q(net_9285), .D(net_9285), .SE(net_7588), .CK(net_14668) );
AOI22_X2 inst_9009 ( .B1(net_9304), .A2(net_8030), .B2(net_8029), .ZN(net_8027), .A1(net_212) );
DFF_X2 inst_8004 ( .QN(net_10119), .D(net_5504), .CK(net_12347) );
CLKBUF_X2 inst_15133 ( .A(net_15051), .Z(net_15052) );
OAI222_X2 inst_1353 ( .B1(net_9256), .C1(net_9090), .ZN(net_7376), .A2(net_7275), .C2(net_7274), .B2(net_7274), .A1(net_7050) );
INV_X4 inst_6369 ( .A(net_8834), .ZN(net_2706) );
DFF_X2 inst_7370 ( .Q(net_9365), .D(net_8692), .CK(net_10547) );
NOR2_X2 inst_2502 ( .A2(net_9575), .A1(net_9574), .ZN(net_8534) );
CLKBUF_X2 inst_15483 ( .A(net_12033), .Z(net_15402) );
OR2_X4 inst_769 ( .A1(net_9237), .A2(net_4070), .ZN(net_3543) );
CLKBUF_X2 inst_13334 ( .A(net_13252), .Z(net_13253) );
CLKBUF_X2 inst_12429 ( .A(net_11046), .Z(net_12348) );
OAI22_X2 inst_1200 ( .A1(net_7249), .A2(net_5107), .B2(net_5105), .ZN(net_5052), .B1(net_5051) );
CLKBUF_X2 inst_15593 ( .A(net_15511), .Z(net_15512) );
CLKBUF_X2 inst_10888 ( .A(net_10806), .Z(net_10807) );
AOI21_X2 inst_10120 ( .B2(net_9739), .ZN(net_4783), .A(net_4472), .B1(net_627) );
AOI22_X2 inst_9114 ( .A1(net_9667), .A2(net_6418), .ZN(net_6375), .B2(net_5263), .B1(net_105) );
CLKBUF_X2 inst_15473 ( .A(net_15391), .Z(net_15392) );
CLKBUF_X2 inst_11233 ( .A(net_11151), .Z(net_11152) );
CLKBUF_X2 inst_10918 ( .A(net_10836), .Z(net_10837) );
DFF_X1 inst_8523 ( .Q(net_8820), .D(net_7402), .CK(net_11415) );
NOR2_X2 inst_3021 ( .ZN(net_647), .A2(net_266), .A1(net_265) );
NAND2_X2 inst_3974 ( .ZN(net_3300), .A1(net_3299), .A2(net_3050) );
INV_X4 inst_6349 ( .A(net_9830), .ZN(net_639) );
CLKBUF_X2 inst_13290 ( .A(net_13208), .Z(net_13209) );
HA_X1 inst_7365 ( .B(net_9275), .A(net_9274), .S(net_1067), .CO(net_1066) );
INV_X4 inst_6474 ( .A(net_10016), .ZN(net_368) );
CLKBUF_X2 inst_12601 ( .A(net_12519), .Z(net_12520) );
CLKBUF_X2 inst_12232 ( .A(net_12150), .Z(net_12151) );
CLKBUF_X2 inst_11664 ( .A(net_10589), .Z(net_11583) );
CLKBUF_X2 inst_15084 ( .A(net_15002), .Z(net_15003) );
CLKBUF_X2 inst_11501 ( .A(net_11419), .Z(net_11420) );
XNOR2_X2 inst_213 ( .ZN(net_4933), .A(net_4397), .B(net_2373) );
CLKBUF_X2 inst_12618 ( .A(net_12536), .Z(net_12537) );
XNOR2_X2 inst_205 ( .ZN(net_4953), .A(net_4686), .B(net_206) );
OAI221_X2 inst_1645 ( .C1(net_10428), .B1(net_7182), .ZN(net_5543), .C2(net_4477), .B2(net_4455), .A(net_3507) );
CLKBUF_X2 inst_13045 ( .A(net_12963), .Z(net_12964) );
DFF_X2 inst_7904 ( .QN(net_10159), .D(net_6003), .CK(net_13477) );
NAND2_X2 inst_3722 ( .A2(net_10274), .ZN(net_7068), .A1(net_2202) );
INV_X4 inst_5410 ( .ZN(net_1949), .A(net_1155) );
DFF_X2 inst_8043 ( .Q(net_9549), .D(net_9255), .CK(net_13760) );
NAND2_X2 inst_4311 ( .A2(net_9243), .ZN(net_2935), .A1(net_858) );
CLKBUF_X2 inst_11922 ( .A(net_11197), .Z(net_11841) );
CLKBUF_X2 inst_15618 ( .A(net_15536), .Z(net_15537) );
CLKBUF_X2 inst_14790 ( .A(net_14708), .Z(net_14709) );
NAND2_X2 inst_3911 ( .ZN(net_4013), .A2(net_3896), .A1(net_3891) );
CLKBUF_X2 inst_14469 ( .A(net_14387), .Z(net_14388) );
OAI221_X2 inst_1515 ( .C1(net_10417), .B2(net_9063), .C2(net_9056), .ZN(net_7328), .B1(net_7136), .A(net_7081) );
INV_X2 inst_6777 ( .ZN(net_6021), .A(net_5836) );
AOI221_X2 inst_9743 ( .B2(net_9647), .A(net_9571), .ZN(net_8205), .C2(net_8190), .B1(net_5283), .C1(net_3125) );
DFF_X2 inst_7546 ( .QN(net_10360), .D(net_7733), .CK(net_12233) );
CLKBUF_X2 inst_14916 ( .A(net_14834), .Z(net_14835) );
CLKBUF_X2 inst_13088 ( .A(net_13006), .Z(net_13007) );
CLKBUF_X2 inst_15388 ( .A(net_15076), .Z(net_15307) );
CLKBUF_X2 inst_14117 ( .A(net_14035), .Z(net_14036) );
OAI21_X2 inst_1782 ( .B2(net_7757), .ZN(net_7702), .A(net_7643), .B1(net_1229) );
INV_X4 inst_5173 ( .A(net_7435), .ZN(net_1871) );
CLKBUF_X2 inst_15274 ( .A(net_11902), .Z(net_15193) );
NOR2_X2 inst_2951 ( .A1(net_10250), .ZN(net_2343), .A2(net_1214) );
INV_X4 inst_6464 ( .A(net_9214), .ZN(net_2497) );
AOI22_X2 inst_9176 ( .A1(net_9903), .B1(net_9804), .ZN(net_6142), .A2(net_6141), .B2(net_6140) );
NAND2_X2 inst_3890 ( .ZN(net_4414), .A2(net_4003), .A1(net_1222) );
MUX2_X1 inst_4472 ( .S(net_6041), .A(net_4910), .B(x6303), .Z(x374) );
DFF_X2 inst_7513 ( .QN(net_9588), .D(net_7977), .CK(net_11604) );
OAI22_X2 inst_1015 ( .A2(net_8247), .B2(net_8246), .ZN(net_8202), .A1(net_6197), .B1(net_1198) );
CLKBUF_X2 inst_15776 ( .A(net_15694), .Z(net_15695) );
INV_X2 inst_7003 ( .A(net_2398), .ZN(net_1620) );
CLKBUF_X2 inst_14390 ( .A(net_14308), .Z(net_14309) );
NAND2_X2 inst_3899 ( .ZN(net_4074), .A2(net_3606), .A1(x6599) );
CLKBUF_X2 inst_13526 ( .A(net_12229), .Z(net_13445) );
CLKBUF_X2 inst_14226 ( .A(net_12573), .Z(net_14145) );
NAND3_X2 inst_3213 ( .A2(net_10092), .A3(net_8511), .A1(net_7832), .ZN(net_6430) );
AOI21_X2 inst_10209 ( .ZN(net_2529), .A(net_2528), .B1(net_2527), .B2(net_1782) );
NOR2_X2 inst_2535 ( .A2(net_9597), .ZN(net_8316), .A1(net_8117) );
CLKBUF_X2 inst_15771 ( .A(net_15689), .Z(net_15690) );
INV_X4 inst_4569 ( .A(net_8385), .ZN(net_8381) );
OAI221_X2 inst_1661 ( .C1(net_7198), .A(net_5637), .C2(net_5520), .ZN(net_5508), .B2(net_4547), .B1(net_1807) );
CLKBUF_X2 inst_12393 ( .A(net_11106), .Z(net_12312) );
MUX2_X1 inst_4480 ( .S(net_6041), .A(net_279), .B(x6186), .Z(x304) );
CLKBUF_X2 inst_13583 ( .A(net_13501), .Z(net_13502) );
XNOR2_X2 inst_283 ( .ZN(net_3646), .A(net_3012), .B(net_2293) );
CLKBUF_X2 inst_15193 ( .A(net_15111), .Z(net_15112) );
CLKBUF_X2 inst_10723 ( .A(net_10641), .Z(net_10642) );
INV_X2 inst_6676 ( .ZN(net_8352), .A(net_8289) );
NOR2_X2 inst_2519 ( .A1(net_9554), .ZN(net_8405), .A2(net_8250) );
NAND2_X2 inst_3406 ( .ZN(net_8542), .A2(net_8491), .A1(net_7040) );
AOI22_X2 inst_9378 ( .B1(net_10019), .A1(net_6816), .A2(net_5743), .B2(net_5742), .ZN(net_5527) );
OAI221_X2 inst_1597 ( .C1(net_10212), .B1(net_7139), .C2(net_5642), .ZN(net_5640), .A(net_5637), .B2(net_4905) );
INV_X4 inst_5639 ( .ZN(net_1189), .A(net_805) );
NAND2_X2 inst_3502 ( .ZN(net_8251), .A2(net_8126), .A1(net_603) );
DFF_X2 inst_7574 ( .D(net_9387), .QN(net_8869), .CK(net_14710) );
NAND2_X2 inst_3473 ( .A1(net_9442), .ZN(net_9022), .A2(net_8952) );
CLKBUF_X2 inst_14584 ( .A(net_14502), .Z(net_14503) );
INV_X4 inst_6018 ( .A(net_10119), .ZN(net_754) );
CLKBUF_X2 inst_14644 ( .A(net_13653), .Z(net_14563) );
AOI221_X2 inst_9942 ( .B1(net_9899), .C1(net_9867), .ZN(net_5339), .B2(net_4969), .A(net_4664), .C2(net_2973) );
DFF_X1 inst_8502 ( .QN(net_9268), .D(net_7792), .CK(net_12540) );
DFF_X2 inst_7705 ( .Q(net_9705), .D(net_6440), .CK(net_13875) );
INV_X4 inst_5822 ( .ZN(net_670), .A(net_669) );
XNOR2_X2 inst_431 ( .A(net_9655), .B(net_2928), .ZN(net_1072) );
INV_X4 inst_6063 ( .A(net_10123), .ZN(net_729) );
INV_X4 inst_6448 ( .A(net_9999), .ZN(net_376) );
XNOR2_X2 inst_348 ( .B(net_9223), .ZN(net_2840), .A(net_2543) );
CLKBUF_X2 inst_11331 ( .A(net_11249), .Z(net_11250) );
DFF_X2 inst_7676 ( .QN(net_10370), .D(net_6931), .CK(net_12213) );
INV_X2 inst_6906 ( .ZN(net_2251), .A(net_2250) );
DFF_X2 inst_7429 ( .QN(net_9407), .D(net_8359), .CK(net_13941) );
DFF_X1 inst_8737 ( .Q(net_9136), .D(net_5731), .CK(net_10633) );
NOR2_X2 inst_2686 ( .A2(net_10271), .A1(net_10270), .ZN(net_5216) );
INV_X4 inst_5123 ( .ZN(net_1603), .A(net_1602) );
CLKBUF_X2 inst_14911 ( .A(net_14829), .Z(net_14830) );
CLKBUF_X2 inst_10774 ( .A(net_10692), .Z(net_10693) );
CLKBUF_X2 inst_15657 ( .A(net_15575), .Z(net_15576) );
NAND2_X2 inst_3740 ( .ZN(net_5950), .A2(net_5393), .A1(net_5392) );
AOI22_X2 inst_9600 ( .ZN(net_3958), .B2(net_3230), .B1(net_2878), .A2(net_2486), .A1(net_2483) );
OAI211_X2 inst_2293 ( .C2(net_4661), .ZN(net_4660), .C1(net_4659), .B(net_4235), .A(net_3505) );
OAI222_X2 inst_1364 ( .A2(net_7660), .C2(net_7659), .B2(net_7658), .ZN(net_6318), .A1(net_2503), .B1(net_1881), .C1(net_1565) );
CLKBUF_X2 inst_11299 ( .A(net_11217), .Z(net_11218) );
CLKBUF_X2 inst_11514 ( .A(net_11432), .Z(net_11433) );
SDFF_X2 inst_645 ( .Q(net_9448), .D(net_9448), .SE(net_3293), .CK(net_14144), .SI(x2648) );
CLKBUF_X2 inst_13299 ( .A(net_13136), .Z(net_13218) );
CLKBUF_X2 inst_15615 ( .A(net_15522), .Z(net_15534) );
CLKBUF_X2 inst_14460 ( .A(net_14378), .Z(net_14379) );
NAND4_X2 inst_3041 ( .A4(net_9310), .ZN(net_7617), .A1(net_862), .A2(net_856), .A3(net_404) );
CLKBUF_X2 inst_14967 ( .A(net_14885), .Z(net_14886) );
NOR4_X2 inst_2352 ( .A4(net_3706), .ZN(net_3322), .A2(net_3102), .A1(net_2622), .A3(net_2621) );
NOR2_X2 inst_2719 ( .ZN(net_4552), .A2(net_4108), .A1(net_1812) );
XNOR2_X2 inst_269 ( .B(net_9159), .ZN(net_4403), .A(net_3953) );
INV_X2 inst_6847 ( .A(net_10269), .ZN(net_3460) );
INV_X2 inst_6864 ( .ZN(net_4893), .A(net_3263) );
CLKBUF_X2 inst_14563 ( .A(net_14481), .Z(net_14482) );
CLKBUF_X2 inst_14801 ( .A(net_14719), .Z(net_14720) );
CLKBUF_X2 inst_12534 ( .A(net_12452), .Z(net_12453) );
CLKBUF_X2 inst_14278 ( .A(net_12432), .Z(net_14197) );
CLKBUF_X2 inst_11278 ( .A(net_10934), .Z(net_11197) );
AOI22_X2 inst_9560 ( .B1(net_9860), .A1(net_9694), .ZN(net_3759), .A2(net_3039), .B2(net_2973) );
NOR2_X2 inst_2544 ( .ZN(net_8301), .A2(net_8299), .A1(net_8081) );
AOI221_X2 inst_9796 ( .B1(net_9976), .A(net_7090), .B2(net_7089), .C2(net_7088), .ZN(net_7008), .C1(net_248) );
CLKBUF_X2 inst_15329 ( .A(net_15247), .Z(net_15248) );
SDFF_X2 inst_514 ( .Q(net_9329), .D(net_9329), .SI(net_9154), .SE(net_7588), .CK(net_14692) );
CLKBUF_X2 inst_14364 ( .A(net_12832), .Z(net_14283) );
CLKBUF_X2 inst_12707 ( .A(net_10732), .Z(net_12626) );
OAI221_X2 inst_1541 ( .B2(net_7295), .C2(net_7293), .C1(net_7226), .ZN(net_7223), .A(net_6820), .B1(net_986) );
NAND2_X2 inst_4236 ( .A2(net_10369), .ZN(net_1944), .A1(net_1116) );
OR4_X2 inst_685 ( .ZN(net_8603), .A1(net_8602), .A4(net_8601), .A2(net_8574), .A3(net_5433) );
CLKBUF_X2 inst_13281 ( .A(net_13199), .Z(net_13200) );
AOI22_X2 inst_9586 ( .B1(net_9984), .A2(net_5173), .ZN(net_3574), .B2(net_2541), .A1(net_218) );
CLKBUF_X2 inst_12952 ( .A(net_12870), .Z(net_12871) );
CLKBUF_X2 inst_15478 ( .A(net_15396), .Z(net_15397) );
CLKBUF_X2 inst_15236 ( .A(net_15154), .Z(net_15155) );
CLKBUF_X2 inst_13829 ( .A(net_12947), .Z(net_13748) );
CLKBUF_X2 inst_14061 ( .A(net_13979), .Z(net_13980) );
INV_X4 inst_4656 ( .A(net_9262), .ZN(net_6241) );
CLKBUF_X2 inst_10658 ( .A(net_10576), .Z(net_10577) );
AOI22_X2 inst_9150 ( .A1(net_9747), .A2(net_6402), .ZN(net_6334), .B2(net_5263), .B1(net_353) );
INV_X4 inst_6338 ( .A(net_9537), .ZN(net_610) );
CLKBUF_X2 inst_14358 ( .A(net_14276), .Z(net_14277) );
INV_X4 inst_5621 ( .A(net_10199), .ZN(net_4221) );
CLKBUF_X2 inst_11585 ( .A(net_11503), .Z(net_11504) );
CLKBUF_X2 inst_10636 ( .A(net_10554), .Z(net_10555) );
NAND2_X2 inst_3432 ( .A1(net_9473), .A2(net_8487), .ZN(net_8484) );
CLKBUF_X2 inst_14047 ( .A(net_10814), .Z(net_13966) );
DFF_X2 inst_7693 ( .Q(net_10402), .D(net_6572), .CK(net_15147) );
CLKBUF_X2 inst_15760 ( .A(net_15678), .Z(net_15679) );
INV_X4 inst_6561 ( .ZN(net_3380), .A(net_168) );
CLKBUF_X2 inst_12700 ( .A(net_12618), .Z(net_12619) );
CLKBUF_X2 inst_12678 ( .A(net_11783), .Z(net_12597) );
CLKBUF_X2 inst_13984 ( .A(net_11153), .Z(net_13903) );
INV_X2 inst_6886 ( .ZN(net_3000), .A(net_2826) );
CLKBUF_X2 inst_15211 ( .A(net_15129), .Z(net_15130) );
XNOR2_X2 inst_427 ( .B(net_7499), .ZN(net_1133), .A(net_210) );
NAND2_X2 inst_3840 ( .ZN(net_7859), .A1(net_4299), .A2(net_4298) );
INV_X2 inst_6881 ( .ZN(net_2991), .A(net_2225) );
CLKBUF_X2 inst_13113 ( .A(net_13031), .Z(net_13032) );
CLKBUF_X2 inst_13852 ( .A(net_13770), .Z(net_13771) );
AOI22_X2 inst_9477 ( .B1(net_10400), .A1(net_9826), .A2(net_6413), .B2(net_4062), .ZN(net_3846) );
CLKBUF_X2 inst_11952 ( .A(net_11870), .Z(net_11871) );
OAI211_X2 inst_2144 ( .C2(net_6778), .ZN(net_6704), .A(net_6330), .B(net_6067), .C1(net_5094) );
CLKBUF_X2 inst_15327 ( .A(net_15245), .Z(net_15246) );
INV_X4 inst_5721 ( .ZN(net_1004), .A(net_761) );
INV_X4 inst_6121 ( .A(net_9235), .ZN(net_681) );
XNOR2_X2 inst_138 ( .ZN(net_7398), .B(net_6937), .A(net_6899) );
INV_X2 inst_6793 ( .A(net_5888), .ZN(net_5707) );
INV_X2 inst_6973 ( .A(net_2682), .ZN(net_1697) );
NOR2_X2 inst_2810 ( .A1(net_4409), .ZN(net_2653), .A2(net_1954) );
INV_X4 inst_5333 ( .ZN(net_1574), .A(net_1259) );
CLKBUF_X2 inst_13971 ( .A(net_13889), .Z(net_13890) );
OR2_X2 inst_899 ( .A1(net_10188), .ZN(net_5657), .A2(net_5431) );
INV_X4 inst_4944 ( .A(net_4714), .ZN(net_4509) );
INV_X2 inst_7170 ( .A(net_9194), .ZN(net_547) );
CLKBUF_X2 inst_10975 ( .A(net_10893), .Z(net_10894) );
AOI211_X2 inst_10259 ( .ZN(net_7988), .A(net_7987), .B(net_7986), .C2(net_7487), .C1(net_7344) );
CLKBUF_X2 inst_12304 ( .A(net_12222), .Z(net_12223) );
XNOR2_X2 inst_312 ( .ZN(net_3224), .B(net_3223), .A(net_2482) );
CLKBUF_X2 inst_13346 ( .A(net_13264), .Z(net_13265) );
CLKBUF_X2 inst_13256 ( .A(net_10840), .Z(net_13175) );
CLKBUF_X2 inst_13429 ( .A(net_13347), .Z(net_13348) );
AOI22_X2 inst_9554 ( .B1(net_9727), .B2(net_6442), .A2(net_5173), .ZN(net_3766), .A1(net_1401) );
XNOR2_X2 inst_309 ( .ZN(net_3953), .B(net_2558), .A(net_2471) );
AOI221_X2 inst_9889 ( .B1(net_9860), .B2(net_9101), .A(net_6945), .C2(net_6944), .C1(net_6834), .ZN(net_6805) );
NAND2_X2 inst_3416 ( .ZN(net_9025), .A1(net_8463), .A2(net_8433) );
OAI211_X2 inst_2149 ( .C2(net_6778), .ZN(net_6699), .A(net_6304), .B(net_6046), .C1(net_5027) );
CLKBUF_X2 inst_13765 ( .A(net_13683), .Z(net_13684) );
DFF_X2 inst_8356 ( .QN(net_10338), .D(net_2493), .CK(net_11031) );
INV_X2 inst_6980 ( .ZN(net_1676), .A(net_1675) );
INV_X4 inst_5001 ( .ZN(net_4719), .A(net_2605) );
AOI22_X2 inst_9365 ( .B1(net_9921), .A2(net_5759), .B2(net_5758), .ZN(net_5557), .A1(net_260) );
CLKBUF_X2 inst_11875 ( .A(net_11793), .Z(net_11794) );
INV_X2 inst_7265 ( .A(net_8914), .ZN(net_8913) );
CLKBUF_X2 inst_14470 ( .A(net_14388), .Z(net_14389) );
AOI221_X2 inst_9833 ( .A(net_6889), .B2(net_6888), .C2(net_6887), .ZN(net_6885), .B1(net_5858), .C1(x5364) );
NOR2_X2 inst_2694 ( .A2(net_10481), .A1(net_10480), .ZN(net_4958) );
DFF_X2 inst_7386 ( .D(net_8654), .QN(net_272), .CK(net_14921) );
DFF_X2 inst_8038 ( .QN(net_9558), .D(net_9264), .CK(net_12625) );
CLKBUF_X2 inst_15207 ( .A(net_13447), .Z(net_15126) );
AOI221_X2 inst_9950 ( .ZN(net_5176), .B1(net_5175), .B2(net_5174), .C2(net_5173), .A(net_4489), .C1(net_3332) );
AOI22_X2 inst_9319 ( .B1(net_9696), .A1(net_6813), .A2(net_5755), .B2(net_5754), .ZN(net_5658) );
DFF_X2 inst_8172 ( .QN(net_9728), .D(net_5040), .CK(net_14533) );
CLKBUF_X2 inst_13899 ( .A(net_11818), .Z(net_13818) );
DFF_X1 inst_8876 ( .Q(net_94), .CK(net_11852), .D(x3338) );
OAI21_X2 inst_1968 ( .A(net_3266), .ZN(net_3256), .B1(net_3255), .B2(net_2812) );
CLKBUF_X2 inst_12983 ( .A(net_12901), .Z(net_12902) );
NAND2_X2 inst_4078 ( .A1(net_9533), .ZN(net_7644), .A2(net_2615) );
CLKBUF_X2 inst_12168 ( .A(net_12086), .Z(net_12087) );
NAND2_X2 inst_4067 ( .ZN(net_3165), .A1(net_2719), .A2(net_2099) );
CLKBUF_X2 inst_12038 ( .A(net_11956), .Z(net_11957) );
OAI222_X2 inst_1330 ( .B1(net_9600), .A1(net_8963), .ZN(net_8540), .B2(net_8539), .A2(net_8539), .C2(net_8538), .C1(net_8138) );
CLKBUF_X2 inst_13963 ( .A(net_13881), .Z(net_13882) );
CLKBUF_X2 inst_13728 ( .A(net_11487), .Z(net_13647) );
CLKBUF_X2 inst_12410 ( .A(net_12146), .Z(net_12329) );
AOI22_X2 inst_9109 ( .A1(net_9690), .ZN(net_6383), .A2(net_6382), .B1(net_6381), .B2(net_5263) );
OAI21_X2 inst_1898 ( .B1(net_7186), .B2(net_4862), .ZN(net_4854), .A(net_4526) );
AOI21_X2 inst_10175 ( .ZN(net_3614), .A(net_3613), .B2(net_3122), .B1(net_1980) );
CLKBUF_X2 inst_14972 ( .A(net_13411), .Z(net_14891) );
CLKBUF_X2 inst_15644 ( .A(net_15562), .Z(net_15563) );
CLKBUF_X2 inst_14180 ( .A(net_11789), .Z(net_14099) );
DFF_X1 inst_8885 ( .Q(net_9508), .D(net_9284), .CK(net_13724) );
NAND2_X2 inst_3883 ( .A2(net_4028), .ZN(net_4020), .A1(net_4019) );
AOI21_X2 inst_10020 ( .ZN(net_8308), .A(net_8082), .B2(net_7986), .B1(net_1690) );
DFF_X1 inst_8551 ( .Q(net_9989), .D(net_7359), .CK(net_14405) );
OAI221_X2 inst_1714 ( .ZN(net_3623), .A(net_3154), .C2(net_2316), .B1(net_2198), .B2(net_2129), .C1(net_668) );
INV_X4 inst_6275 ( .A(net_9345), .ZN(net_594) );
CLKBUF_X2 inst_11811 ( .A(net_11256), .Z(net_11730) );
CLKBUF_X2 inst_13451 ( .A(net_13369), .Z(net_13370) );
AOI22_X2 inst_9164 ( .A2(net_6382), .ZN(net_6308), .B2(net_5263), .B1(net_2583), .A1(net_1867) );
CLKBUF_X2 inst_14630 ( .A(net_14548), .Z(net_14549) );
AOI22_X2 inst_9096 ( .A1(net_9677), .A2(net_6420), .ZN(net_6396), .B2(net_5263), .B1(net_115) );
AOI22_X2 inst_9428 ( .A1(net_9754), .B1(net_6808), .ZN(net_4619), .A2(net_4618), .B2(net_4617) );
INV_X4 inst_4777 ( .ZN(net_4306), .A(net_4000) );
CLKBUF_X2 inst_15789 ( .A(net_15707), .Z(net_15708) );
CLKBUF_X2 inst_10851 ( .A(net_10769), .Z(net_10770) );
CLKBUF_X2 inst_10762 ( .A(net_10616), .Z(net_10681) );
CLKBUF_X2 inst_15333 ( .A(net_15251), .Z(net_15252) );
INV_X4 inst_5818 ( .ZN(net_1365), .A(net_674) );
CLKBUF_X2 inst_11292 ( .A(net_11210), .Z(net_11211) );
OAI221_X2 inst_1496 ( .C2(net_9063), .B2(net_9056), .ZN(net_7367), .C1(net_7231), .A(net_7006), .B1(net_5464) );
INV_X4 inst_5510 ( .A(net_10125), .ZN(net_1431) );
AOI22_X2 inst_9091 ( .A1(net_9662), .A2(net_6420), .ZN(net_6401), .B2(net_5263), .B1(net_100) );
INV_X2 inst_7041 ( .ZN(net_1373), .A(net_1372) );
CLKBUF_X2 inst_13005 ( .A(net_12923), .Z(net_12924) );
AOI22_X2 inst_9381 ( .B1(net_10022), .A2(net_5743), .B2(net_5742), .ZN(net_5524), .A1(net_262) );
NAND2_X2 inst_4297 ( .A2(net_10229), .A1(net_7481), .ZN(net_1236) );
OR2_X2 inst_924 ( .ZN(net_3313), .A2(net_3058), .A1(net_2254) );
OAI221_X2 inst_1565 ( .C1(net_10308), .C2(net_9047), .B2(net_7287), .B1(net_7190), .ZN(net_7188), .A(net_6786) );
DFF_X1 inst_8415 ( .Q(net_9569), .D(net_8791), .CK(net_11636) );
CLKBUF_X2 inst_12632 ( .A(net_11328), .Z(net_12551) );
AOI211_X2 inst_10308 ( .B(net_9182), .C1(net_9180), .ZN(net_3017), .A(net_3016), .C2(net_2196) );
XNOR2_X2 inst_287 ( .ZN(net_6655), .A(net_6625), .B(net_1143) );
AND2_X2 inst_10614 ( .A1(net_9175), .ZN(net_1746), .A2(net_1064) );
NOR2_X2 inst_2577 ( .ZN(net_7993), .A1(net_7253), .A2(net_7252) );
DFF_X2 inst_7929 ( .QN(net_10305), .D(net_5593), .CK(net_12036) );
CLKBUF_X2 inst_15319 ( .A(net_15237), .Z(net_15238) );
CLKBUF_X2 inst_12030 ( .A(net_11948), .Z(net_11949) );
DFF_X2 inst_7565 ( .Q(net_9289), .D(net_7650), .CK(net_13120) );
NAND4_X2 inst_3094 ( .ZN(net_4351), .A2(net_3791), .A3(net_3548), .A1(net_3186), .A4(net_2745) );
CLKBUF_X2 inst_13267 ( .A(net_12409), .Z(net_13186) );
CLKBUF_X2 inst_13830 ( .A(net_13748), .Z(net_13749) );
NOR2_X2 inst_2903 ( .ZN(net_2680), .A2(net_1169), .A1(net_917) );
NAND2_X2 inst_4045 ( .A2(net_8868), .ZN(net_4580), .A1(net_2827) );
INV_X4 inst_6431 ( .A(net_10494), .ZN(net_380) );
CLKBUF_X2 inst_12623 ( .A(net_12541), .Z(net_12542) );
INV_X4 inst_4890 ( .ZN(net_2937), .A(net_2733) );
INV_X2 inst_7131 ( .ZN(net_853), .A(net_852) );
OAI22_X2 inst_984 ( .B1(net_9258), .A2(net_8962), .B2(net_8659), .ZN(net_8656), .A1(net_6428) );
NAND2_X2 inst_3804 ( .A1(net_10073), .ZN(net_4535), .A2(net_4534) );
INV_X2 inst_6734 ( .A(net_7605), .ZN(net_7516) );
OAI211_X2 inst_2064 ( .A(net_9534), .ZN(net_7713), .B(net_7620), .C2(net_7619), .C1(net_7618) );
CLKBUF_X2 inst_14604 ( .A(net_14522), .Z(net_14523) );
OAI211_X2 inst_2266 ( .C1(net_7129), .C2(net_6542), .ZN(net_6279), .B(net_5705), .A(net_3679) );
CLKBUF_X2 inst_15057 ( .A(net_13671), .Z(net_14976) );
CLKBUF_X2 inst_14331 ( .A(net_14249), .Z(net_14250) );
OAI22_X2 inst_1292 ( .B1(net_5092), .A2(net_4274), .ZN(net_3590), .A1(net_3589), .B2(net_3588) );
INV_X2 inst_7148 ( .A(net_4211), .ZN(net_3536) );
CLKBUF_X2 inst_15769 ( .A(net_15687), .Z(net_15688) );
CLKBUF_X2 inst_13206 ( .A(net_13124), .Z(net_13125) );
INV_X4 inst_5014 ( .ZN(net_2811), .A(net_2117) );
OAI21_X2 inst_1963 ( .ZN(net_3499), .A(net_3267), .B2(net_3027), .B1(net_843) );
OAI22_X2 inst_1056 ( .ZN(net_7450), .B2(net_7449), .A1(net_7343), .A2(net_6969), .B1(net_3510) );
CLKBUF_X2 inst_11818 ( .A(net_11736), .Z(net_11737) );
CLKBUF_X2 inst_13440 ( .A(net_13358), .Z(net_13359) );
NAND2_X2 inst_3648 ( .ZN(net_6783), .A2(net_6448), .A1(net_3827) );
NAND2_X2 inst_4247 ( .ZN(net_1438), .A1(net_1437), .A2(net_1436) );
CLKBUF_X2 inst_14434 ( .A(net_11986), .Z(net_14353) );
DFF_X1 inst_8744 ( .Q(net_9150), .D(net_5680), .CK(net_11064) );
CLKBUF_X2 inst_12023 ( .A(net_11941), .Z(net_11942) );
CLKBUF_X2 inst_13437 ( .A(net_13262), .Z(net_13356) );
NOR2_X2 inst_2514 ( .A1(net_9057), .ZN(net_8270), .A2(net_8154) );
DFF_X2 inst_7869 ( .QN(net_10263), .D(net_5959), .CK(net_11665) );
CLKBUF_X2 inst_14359 ( .A(net_14277), .Z(net_14278) );
OAI22_X2 inst_1128 ( .A1(net_7245), .ZN(net_5152), .A2(net_5151), .B2(net_5150), .B1(net_482) );
INV_X4 inst_4988 ( .ZN(net_2567), .A(net_2227) );
INV_X4 inst_6524 ( .A(net_9839), .ZN(net_601) );
DFF_X2 inst_8009 ( .QN(net_10438), .D(net_5500), .CK(net_13717) );
CLKBUF_X2 inst_11325 ( .A(net_11243), .Z(net_11244) );
NAND3_X2 inst_3222 ( .A2(net_9533), .A1(net_5353), .ZN(net_5352), .A3(net_5351) );
NAND2_X2 inst_3759 ( .A2(net_5383), .ZN(net_5230), .A1(net_440) );
CLKBUF_X2 inst_15074 ( .A(net_14992), .Z(net_14993) );
CLKBUF_X2 inst_10928 ( .A(net_10712), .Z(net_10847) );
DFF_X2 inst_7422 ( .QN(net_9393), .D(net_8339), .CK(net_14017) );
CLKBUF_X2 inst_14216 ( .A(net_10744), .Z(net_14135) );
CLKBUF_X2 inst_14996 ( .A(net_14914), .Z(net_14915) );
CLKBUF_X2 inst_11677 ( .A(net_11595), .Z(net_11596) );
CLKBUF_X2 inst_11559 ( .A(net_11186), .Z(net_11478) );
AOI21_X2 inst_10064 ( .ZN(net_7024), .A(net_7023), .B1(net_5185), .B2(net_4928) );
CLKBUF_X2 inst_10999 ( .A(net_10732), .Z(net_10918) );
NAND2_X2 inst_4070 ( .ZN(net_7615), .A1(net_2845), .A2(net_2368) );
AOI22_X2 inst_9077 ( .B1(net_9676), .A1(net_6684), .B2(net_6683), .ZN(net_6559), .A2(net_245) );
OAI21_X2 inst_1924 ( .B2(net_10489), .ZN(net_4515), .B1(net_3748), .A(x3698) );
AOI22_X2 inst_9023 ( .B1(net_9523), .A1(net_8002), .B2(net_8001), .ZN(net_7996), .A2(net_7949) );
CLKBUF_X2 inst_12714 ( .A(net_12632), .Z(net_12633) );
AND2_X2 inst_10502 ( .ZN(net_6619), .A1(net_5961), .A2(net_5782) );
AOI21_X2 inst_10244 ( .ZN(net_8864), .B1(net_2399), .B2(net_2398), .A(net_2397) );
CLKBUF_X2 inst_14750 ( .A(net_13369), .Z(net_14669) );
DFF_X2 inst_7650 ( .D(net_6697), .QN(net_180), .CK(net_15243) );
INV_X4 inst_4748 ( .ZN(net_5642), .A(net_4517) );
DFF_X2 inst_8296 ( .Q(net_9854), .D(net_4616), .CK(net_15412) );
NAND2_X2 inst_4160 ( .A1(net_4183), .ZN(net_1979), .A2(net_1396) );
INV_X4 inst_5685 ( .ZN(net_1112), .A(net_992) );
CLKBUF_X2 inst_12160 ( .A(net_12078), .Z(net_12079) );
OAI33_X1 inst_961 ( .B3(net_9649), .A2(net_9640), .ZN(net_5200), .A1(net_1792), .B1(net_1769), .B2(net_1028), .A3(net_1024) );
NAND3_X2 inst_3255 ( .ZN(net_4505), .A3(net_4065), .A2(net_3552), .A1(net_3440) );
CLKBUF_X2 inst_12246 ( .A(net_10991), .Z(net_12165) );
CLKBUF_X2 inst_13119 ( .A(net_13037), .Z(net_13038) );
OAI221_X2 inst_1590 ( .B2(net_10376), .ZN(net_5984), .B1(net_5983), .A(net_5225), .C2(net_5215), .C1(net_4248) );
CLKBUF_X2 inst_11082 ( .A(net_11000), .Z(net_11001) );
DFF_X2 inst_7591 ( .D(net_7496), .QN(net_193), .CK(net_15363) );
CLKBUF_X2 inst_12800 ( .A(net_12718), .Z(net_12719) );
DFF_X2 inst_8077 ( .QN(net_10354), .D(net_5326), .CK(net_13617) );
CLKBUF_X2 inst_10931 ( .A(net_10849), .Z(net_10850) );
CLKBUF_X2 inst_10648 ( .A(net_10550), .Z(net_10567) );
DFF_X2 inst_8332 ( .Q(net_9615), .D(net_3144), .CK(net_14062) );
INV_X4 inst_6229 ( .A(net_9944), .ZN(net_2287) );
XNOR2_X2 inst_399 ( .B(net_9616), .ZN(net_1754), .A(net_1545) );
NOR4_X2 inst_2318 ( .ZN(net_7173), .A1(net_6612), .A3(net_6349), .A4(net_6347), .A2(net_3616) );
INV_X4 inst_5347 ( .A(net_1247), .ZN(net_1241) );
CLKBUF_X2 inst_12433 ( .A(net_12351), .Z(net_12352) );
INV_X4 inst_5103 ( .ZN(net_4233), .A(net_2963) );
NAND2_X2 inst_3957 ( .ZN(net_3474), .A2(net_3473), .A1(net_2032) );
CLKBUF_X2 inst_11364 ( .A(net_10792), .Z(net_11283) );
AOI221_X2 inst_9953 ( .C2(net_10444), .B1(net_10443), .ZN(net_4799), .A(net_4300), .B2(net_4137), .C1(net_3985) );
NAND2_X2 inst_4020 ( .A1(net_9538), .ZN(net_5180), .A2(net_3072) );
CLKBUF_X2 inst_13404 ( .A(net_11368), .Z(net_13323) );
DFF_X1 inst_8489 ( .QN(net_9627), .D(net_7921), .CK(net_15007) );
NOR4_X2 inst_2316 ( .ZN(net_7178), .A4(net_7175), .A2(net_5270), .A3(net_4510), .A1(net_3359) );
NOR2_X2 inst_2737 ( .ZN(net_4154), .A1(net_3298), .A2(net_3145) );
INV_X2 inst_6654 ( .ZN(net_8551), .A(net_8533) );
CLKBUF_X2 inst_14266 ( .A(net_14184), .Z(net_14185) );
SDFF_X2 inst_499 ( .SE(net_9540), .SI(net_8210), .Q(net_288), .D(net_288), .CK(net_12694) );
OAI22_X2 inst_1299 ( .A2(net_10127), .B2(net_8845), .ZN(net_3395), .A1(net_3173), .B1(net_1243) );
DFF_X2 inst_8404 ( .Q(net_9153), .CK(net_11292), .D(x3613) );
INV_X4 inst_6450 ( .ZN(net_1972), .A(net_153) );
CLKBUF_X2 inst_13487 ( .A(net_11555), .Z(net_13406) );
AND2_X4 inst_10404 ( .ZN(net_5159), .A2(net_5158), .A1(net_4327) );
INV_X4 inst_6175 ( .ZN(net_7201), .A(x4694) );
AOI22_X2 inst_9468 ( .B1(net_9909), .A1(net_9711), .B2(net_4969), .ZN(net_3859), .A2(net_3039) );
CLKBUF_X2 inst_14683 ( .A(net_14601), .Z(net_14602) );
SDFF_X2 inst_674 ( .SI(net_9485), .Q(net_9485), .SE(net_3073), .CK(net_12385), .D(x2333) );
NOR3_X2 inst_2400 ( .A2(net_9544), .A3(net_9542), .ZN(net_7619), .A1(net_7546) );
INV_X4 inst_5259 ( .A(net_6673), .ZN(net_1846) );
OAI221_X2 inst_1451 ( .ZN(net_8061), .C2(net_7881), .A(net_7879), .B2(net_7834), .B1(net_7794), .C1(net_6837) );
NAND2_X2 inst_4082 ( .ZN(net_3344), .A2(net_1977), .A1(net_593) );
INV_X4 inst_4781 ( .A(net_8122), .ZN(x813) );
INV_X4 inst_5518 ( .ZN(net_970), .A(net_969) );
CLKBUF_X2 inst_14151 ( .A(net_14069), .Z(net_14070) );
CLKBUF_X2 inst_14207 ( .A(net_11592), .Z(net_14126) );
CLKBUF_X2 inst_10859 ( .A(net_10673), .Z(net_10778) );
OAI211_X2 inst_2253 ( .C1(net_7249), .C2(net_6548), .ZN(net_6438), .B(net_5441), .A(net_3679) );
CLKBUF_X2 inst_13670 ( .A(net_13588), .Z(net_13589) );
OAI21_X2 inst_2009 ( .ZN(net_2004), .A(net_1329), .B2(net_221), .B1(net_220) );
AOI21_X2 inst_10115 ( .ZN(net_4556), .B1(net_4553), .B2(net_4552), .A(net_2951) );
AOI222_X2 inst_9674 ( .ZN(net_3116), .A1(net_3115), .C2(net_3114), .B2(net_3114), .A2(net_2252), .B1(net_1449), .C1(net_908) );
SDFF_X2 inst_501 ( .SE(net_9540), .SI(net_8208), .Q(net_290), .D(net_290), .CK(net_13965) );
NOR2_X2 inst_2868 ( .ZN(net_2029), .A2(net_2028), .A1(net_1341) );
CLKBUF_X2 inst_12254 ( .A(net_12172), .Z(net_12173) );
OAI211_X2 inst_2093 ( .C2(net_6778), .ZN(net_6755), .A(net_6383), .B(net_6115), .C1(net_529) );
INV_X4 inst_6522 ( .A(net_9938), .ZN(net_587) );
OAI22_X2 inst_1081 ( .A1(net_7157), .ZN(net_6578), .A2(net_5911), .B2(net_5910), .B1(net_540) );
NAND3_X2 inst_3195 ( .ZN(net_8993), .A3(net_7144), .A2(net_7087), .A1(net_4730) );
DFF_X1 inst_8873 ( .Q(net_98), .CK(net_11855), .D(x3307) );
CLKBUF_X2 inst_14549 ( .A(net_14467), .Z(net_14468) );
CLKBUF_X2 inst_10731 ( .A(net_10580), .Z(net_10650) );
CLKBUF_X2 inst_12261 ( .A(net_12179), .Z(net_12180) );
CLKBUF_X2 inst_15828 ( .A(net_10616), .Z(net_15747) );
OAI21_X2 inst_1832 ( .B2(net_10450), .ZN(net_6335), .A(net_1172), .B1(net_679) );
NOR2_X2 inst_2905 ( .ZN(net_2744), .A1(net_1199), .A2(net_1101) );
CLKBUF_X2 inst_13241 ( .A(net_13159), .Z(net_13160) );
NOR2_X2 inst_2819 ( .A1(net_7672), .A2(net_3065), .ZN(net_2597) );
CLKBUF_X2 inst_15740 ( .A(net_15658), .Z(net_15659) );
CLKBUF_X2 inst_12263 ( .A(net_11835), .Z(net_12182) );
SDFF_X2 inst_640 ( .Q(net_9449), .D(net_9449), .SE(net_3293), .CK(net_14150), .SI(x2589) );
INV_X4 inst_4562 ( .ZN(net_8424), .A(net_8242) );
AOI221_X2 inst_9893 ( .B1(net_9879), .B2(net_9101), .A(net_6945), .C2(net_6944), .ZN(net_6801), .C1(net_250) );
DFF_X2 inst_7500 ( .Q(net_9278), .D(net_8034), .CK(net_13127) );
INV_X4 inst_6293 ( .A(net_9939), .ZN(net_3589) );
OAI221_X2 inst_1478 ( .ZN(net_7645), .B1(net_7644), .B2(net_7426), .C1(net_5180), .C2(net_4894), .A(net_3264) );
INV_X4 inst_6098 ( .A(net_9985), .ZN(net_494) );
CLKBUF_X2 inst_15016 ( .A(net_14934), .Z(net_14935) );
AOI221_X2 inst_9963 ( .C1(net_9967), .B2(net_5173), .ZN(net_4768), .A(net_4339), .C2(net_2541), .B1(net_205) );
OAI22_X2 inst_1114 ( .B2(net_7525), .ZN(net_5686), .A1(net_5685), .B1(net_5684), .A2(net_4759) );
DFF_X2 inst_7982 ( .QN(net_10425), .D(net_5546), .CK(net_11751) );
AOI22_X2 inst_9327 ( .B1(net_9994), .A1(net_6808), .A2(net_5743), .B2(net_5742), .ZN(net_5648) );
AOI22_X2 inst_9535 ( .B1(net_9705), .A2(net_5173), .ZN(net_3786), .B2(net_3039), .A1(net_208) );
NAND2_X2 inst_4163 ( .ZN(net_2918), .A1(net_1976), .A2(net_1975) );
CLKBUF_X2 inst_15391 ( .A(net_15309), .Z(net_15310) );
AOI22_X2 inst_9020 ( .A1(net_8002), .B2(net_8001), .ZN(net_7999), .A2(net_7952), .B1(net_2818) );
CLKBUF_X2 inst_12957 ( .A(net_12875), .Z(net_12876) );
AOI22_X2 inst_9085 ( .A1(net_9738), .A2(net_6418), .ZN(net_6410), .B2(net_5263), .B1(net_951) );
CLKBUF_X2 inst_13739 ( .A(net_13657), .Z(net_13658) );
OAI21_X2 inst_1982 ( .B2(net_9045), .ZN(net_8565), .A(net_2850), .B1(net_2849) );
INV_X4 inst_6075 ( .A(net_9306), .ZN(net_502) );
OAI211_X2 inst_2089 ( .C2(net_6774), .ZN(net_6759), .A(net_6386), .B(net_6119), .C1(net_336) );
CLKBUF_X2 inst_15128 ( .A(net_13844), .Z(net_15047) );
CLKBUF_X2 inst_11805 ( .A(net_11723), .Z(net_11724) );
CLKBUF_X2 inst_11378 ( .A(net_10733), .Z(net_11297) );
OAI21_X2 inst_1849 ( .ZN(net_5883), .A(net_5597), .B1(net_5511), .B2(net_5323) );
OAI221_X2 inst_1679 ( .B1(net_10324), .C1(net_7231), .B2(net_5591), .ZN(net_5488), .C2(net_4902), .A(net_3507) );
INV_X4 inst_5540 ( .ZN(net_942), .A(net_187) );
CLKBUF_X2 inst_11123 ( .A(net_10944), .Z(net_11042) );
OAI21_X2 inst_1976 ( .ZN(net_2883), .B2(net_2882), .A(net_2773), .B1(net_1492) );
INV_X4 inst_4932 ( .ZN(net_3628), .A(net_2602) );
NOR2_X2 inst_2744 ( .A1(net_3687), .ZN(net_3684), .A2(net_3683) );
NAND2_X2 inst_3681 ( .ZN(net_6166), .A1(net_6165), .A2(net_6164) );
INV_X2 inst_6909 ( .A(net_2871), .ZN(net_2583) );
CLKBUF_X2 inst_13238 ( .A(net_13156), .Z(net_13157) );
OAI211_X2 inst_2215 ( .C1(net_7226), .C2(net_6501), .ZN(net_6490), .B(net_5553), .A(net_3679) );
XNOR2_X2 inst_337 ( .ZN(net_2977), .A(net_2383), .B(net_2144) );
OAI21_X2 inst_1855 ( .ZN(net_6846), .A(net_6190), .B2(net_5802), .B1(net_4975) );
INV_X4 inst_5277 ( .ZN(net_2051), .A(net_916) );
NOR3_X2 inst_2384 ( .A3(net_9612), .ZN(net_7809), .A1(net_7808), .A2(net_2889) );
INV_X4 inst_4614 ( .ZN(net_7338), .A(net_7153) );
CLKBUF_X2 inst_11564 ( .A(net_11482), .Z(net_11483) );
AOI22_X2 inst_9606 ( .B1(net_9803), .A2(net_5174), .ZN(net_3447), .B2(net_2556), .A1(net_1036) );
OAI22_X2 inst_1212 ( .A1(net_7192), .A2(net_5139), .B2(net_5138), .ZN(net_5037), .B1(net_2593) );
CLKBUF_X2 inst_11193 ( .A(net_11111), .Z(net_11112) );
SDFF_X2 inst_670 ( .SI(net_9499), .Q(net_9499), .SE(net_3073), .CK(net_12391), .D(x1503) );
CLKBUF_X2 inst_15355 ( .A(net_13699), .Z(net_15274) );
INV_X4 inst_6220 ( .A(net_10371), .ZN(net_699) );
CLKBUF_X2 inst_13355 ( .A(net_11796), .Z(net_13274) );
NAND2_X2 inst_4180 ( .ZN(net_2659), .A2(net_1561), .A1(net_1195) );
INV_X4 inst_5789 ( .A(net_3380), .ZN(net_1732) );
CLKBUF_X2 inst_11105 ( .A(net_11023), .Z(net_11024) );
CLKBUF_X2 inst_13775 ( .A(net_13693), .Z(net_13694) );
AOI22_X2 inst_9612 ( .A1(net_10085), .B1(net_10011), .A2(net_5319), .ZN(net_3441), .B2(net_2468) );
NAND2_X2 inst_3901 ( .ZN(net_3905), .A2(net_3903), .A1(net_101) );
AOI22_X2 inst_9262 ( .B2(net_10236), .A1(net_10235), .ZN(net_5933), .A2(net_5188), .B1(net_4929) );
INV_X2 inst_6679 ( .ZN(net_8349), .A(net_8283) );
DFF_X2 inst_7738 ( .Q(net_10014), .D(net_6472), .CK(net_12801) );
CLKBUF_X2 inst_15200 ( .A(net_15118), .Z(net_15119) );
NOR3_X2 inst_2396 ( .A1(net_9163), .ZN(net_7637), .A3(net_7593), .A2(net_3542) );
CLKBUF_X2 inst_15704 ( .A(net_15622), .Z(net_15623) );
AOI21_X2 inst_10232 ( .ZN(net_1952), .A(net_1951), .B1(net_1299), .B2(net_886) );
AOI211_X2 inst_10281 ( .C2(net_9072), .ZN(net_5995), .A(net_5994), .C1(net_5993), .B(net_5812) );
CLKBUF_X2 inst_14295 ( .A(net_14213), .Z(net_14214) );
CLKBUF_X2 inst_14093 ( .A(net_14011), .Z(net_14012) );
INV_X4 inst_5898 ( .ZN(net_1817), .A(net_602) );
DFF_X1 inst_8647 ( .Q(net_9876), .D(net_7181), .CK(net_15459) );
CLKBUF_X2 inst_14628 ( .A(net_10684), .Z(net_14547) );
CLKBUF_X2 inst_10845 ( .A(net_10763), .Z(net_10764) );
XNOR2_X2 inst_246 ( .ZN(net_4134), .A(net_3979), .B(net_1289) );
INV_X4 inst_5908 ( .A(net_1211), .ZN(net_992) );
CLKBUF_X2 inst_12384 ( .A(net_12302), .Z(net_12303) );
SDFF_X2 inst_635 ( .Q(net_9469), .D(net_9469), .SE(net_3293), .CK(net_11365), .SI(x1418) );
MUX2_X1 inst_4443 ( .S(net_6041), .A(net_303), .B(x4587), .Z(x91) );
AOI221_X2 inst_9814 ( .B1(net_9963), .A(net_7090), .B2(net_7089), .C2(net_7088), .ZN(net_6988), .C1(net_235) );
INV_X4 inst_5787 ( .ZN(net_697), .A(net_696) );
CLKBUF_X2 inst_14502 ( .A(net_14420), .Z(net_14421) );
OR2_X4 inst_807 ( .ZN(net_3118), .A1(net_1387), .A2(net_1371) );
OR3_X2 inst_705 ( .ZN(net_8636), .A2(net_8635), .A1(net_8613), .A3(net_7720) );
AND2_X2 inst_10569 ( .A1(net_3270), .A2(net_3023), .ZN(net_3020) );
DFF_X1 inst_8510 ( .QN(net_9661), .D(net_7695), .CK(net_11209) );
OR2_X2 inst_911 ( .ZN(net_4408), .A2(net_3958), .A1(net_2214) );
CLKBUF_X2 inst_15140 ( .A(net_15058), .Z(net_15059) );
SDFF_X2 inst_519 ( .Q(net_9335), .D(net_9335), .SI(net_9327), .SE(net_7588), .CK(net_13076) );
CLKBUF_X2 inst_10921 ( .A(net_10839), .Z(net_10840) );
DFF_X2 inst_7641 ( .D(net_6729), .QN(net_156), .CK(net_12822) );
NAND2_X2 inst_3796 ( .ZN(net_4711), .A2(net_4599), .A1(net_1349) );
CLKBUF_X2 inst_15746 ( .A(net_15664), .Z(net_15665) );
AOI22_X2 inst_9359 ( .B1(net_9916), .A1(net_6821), .A2(net_5759), .B2(net_5758), .ZN(net_5563) );
OAI22_X2 inst_1003 ( .A2(net_8546), .B2(net_8545), .ZN(net_8543), .A1(net_2507), .B1(net_550) );
CLKBUF_X2 inst_14893 ( .A(net_14494), .Z(net_14812) );
CLKBUF_X2 inst_13804 ( .A(net_13722), .Z(net_13723) );
CLKBUF_X2 inst_12758 ( .A(net_12676), .Z(net_12677) );
CLKBUF_X2 inst_12174 ( .A(net_12092), .Z(net_12093) );
OAI22_X2 inst_1053 ( .ZN(net_7523), .A1(net_7522), .B1(net_7521), .A2(net_6855), .B2(net_5401) );
INV_X4 inst_5158 ( .ZN(net_4050), .A(net_2202) );
CLKBUF_X2 inst_14889 ( .A(net_13215), .Z(net_14808) );
AOI211_X2 inst_10284 ( .ZN(net_5887), .C1(net_5886), .C2(net_5885), .B(net_5162), .A(net_2850) );
NAND2_X2 inst_3469 ( .A2(net_9438), .A1(net_8952), .ZN(net_8890) );
INV_X2 inst_7231 ( .A(net_9541), .ZN(net_392) );
CLKBUF_X2 inst_14673 ( .A(net_14591), .Z(net_14592) );
NOR2_X2 inst_2774 ( .ZN(net_4468), .A1(net_3298), .A2(net_3192) );
INV_X4 inst_6026 ( .A(net_9311), .ZN(net_2524) );
INV_X2 inst_6871 ( .ZN(net_3043), .A(net_3042) );
CLKBUF_X2 inst_12202 ( .A(net_11318), .Z(net_12121) );
INV_X4 inst_5456 ( .ZN(net_1595), .A(net_1069) );
XNOR2_X2 inst_239 ( .ZN(net_4257), .A(net_4111), .B(net_1810) );
INV_X4 inst_4577 ( .ZN(net_8136), .A(net_8119) );
OAI22_X2 inst_1193 ( .A1(net_7249), .A2(net_5151), .B2(net_5150), .ZN(net_5060), .B1(net_1164) );
OAI211_X2 inst_2080 ( .C2(net_6778), .ZN(net_6768), .A(net_6395), .B(net_6128), .C1(net_340) );
CLKBUF_X2 inst_14770 ( .A(net_12655), .Z(net_14689) );
OAI221_X2 inst_1625 ( .C1(net_10322), .B1(net_7184), .A(net_5637), .C2(net_5591), .ZN(net_5582), .B2(net_4902) );
DFF_X2 inst_7710 ( .Q(net_10018), .D(net_6467), .CK(net_13439) );
SDFF_X2 inst_593 ( .Q(net_9257), .SE(net_4589), .D(net_140), .SI(net_106), .CK(net_13825) );
INV_X4 inst_5707 ( .ZN(net_891), .A(net_773) );
CLKBUF_X2 inst_15664 ( .A(net_15582), .Z(net_15583) );
OAI211_X2 inst_2223 ( .C1(net_7245), .ZN(net_6482), .C2(net_6480), .B(net_5649), .A(net_3527) );
CLKBUF_X2 inst_15228 ( .A(net_15146), .Z(net_15147) );
AND2_X2 inst_10582 ( .ZN(net_3009), .A2(net_2563), .A1(net_960) );
INV_X8 inst_4522 ( .ZN(net_8933), .A(net_8605) );
INV_X4 inst_6137 ( .A(net_9845), .ZN(net_2021) );
CLKBUF_X2 inst_12426 ( .A(net_12344), .Z(net_12345) );
AOI21_X2 inst_10099 ( .A(net_5101), .ZN(net_5018), .B1(net_5017), .B2(net_2153) );
CLKBUF_X2 inst_12395 ( .A(net_11444), .Z(net_12314) );
SDFF_X2 inst_601 ( .QN(net_9173), .D(net_4802), .SI(net_4801), .SE(net_1033), .CK(net_11232) );
INV_X4 inst_5738 ( .A(net_3967), .ZN(net_854) );
INV_X4 inst_6091 ( .A(net_10014), .ZN(net_495) );
CLKBUF_X2 inst_13709 ( .A(net_13627), .Z(net_13628) );
DFF_X2 inst_7391 ( .D(net_8585), .QN(net_234), .CK(net_12076) );
DFF_X2 inst_7952 ( .QN(net_10212), .D(net_5640), .CK(net_14793) );
DFF_X2 inst_7845 ( .Q(net_9713), .D(net_6544), .CK(net_12787) );
DFF_X2 inst_8097 ( .QN(net_9166), .D(net_5018), .CK(net_13552) );
AOI22_X2 inst_9065 ( .B1(net_9685), .A1(net_6823), .A2(net_6684), .B2(net_6683), .ZN(net_6601) );
AOI21_X2 inst_10045 ( .ZN(net_7443), .A(net_7122), .B2(net_3313), .B1(net_2713) );
SDFF_X2 inst_479 ( .SE(net_9540), .SI(net_8230), .Q(net_294), .D(net_294), .CK(net_13972) );
OAI21_X2 inst_1773 ( .ZN(net_7925), .B1(net_7924), .B2(net_7861), .A(net_7511) );
AND2_X4 inst_10448 ( .A2(net_9344), .ZN(net_2235), .A1(net_1383) );
NOR4_X2 inst_2344 ( .A4(net_9826), .ZN(net_2947), .A1(net_2946), .A3(net_2945), .A2(net_2194) );
AOI211_X2 inst_10278 ( .A(net_7343), .ZN(net_7122), .B(net_6968), .C2(net_6967), .C1(net_980) );
AOI21_X2 inst_10133 ( .B2(net_10339), .ZN(net_4419), .A(net_2006), .B1(net_2005) );
NAND2_X4 inst_3326 ( .ZN(net_9084), .A1(net_8606), .A2(net_8604) );
INV_X2 inst_7288 ( .A(net_8982), .ZN(net_8981) );
DFF_X2 inst_7683 ( .Q(net_10066), .D(net_6570), .CK(net_11181) );
OR2_X4 inst_771 ( .A2(net_4333), .ZN(net_3336), .A1(net_3142) );
OAI221_X2 inst_1583 ( .B1(net_10317), .B2(net_9047), .C2(net_7287), .C1(net_7139), .ZN(net_7123), .A(net_6917) );
CLKBUF_X2 inst_12892 ( .A(net_12810), .Z(net_12811) );
NAND2_X2 inst_4387 ( .A2(net_10458), .ZN(net_806), .A1(net_805) );
AOI22_X2 inst_9420 ( .A1(net_10184), .A2(net_4656), .B2(net_4655), .ZN(net_4649), .B1(x4937) );
INV_X4 inst_6325 ( .A(net_10163), .ZN(net_7029) );
CLKBUF_X2 inst_11552 ( .A(net_10900), .Z(net_11471) );
CLKBUF_X2 inst_15068 ( .A(net_14986), .Z(net_14987) );
INV_X2 inst_7113 ( .A(net_9949), .ZN(net_1228) );
CLKBUF_X2 inst_15654 ( .A(net_15572), .Z(net_15573) );
INV_X4 inst_5780 ( .ZN(net_987), .A(net_705) );
INV_X16 inst_7324 ( .ZN(net_5867), .A(net_5520) );
AOI22_X2 inst_9334 ( .B1(net_9810), .A2(net_5766), .B2(net_5765), .ZN(net_5618), .A1(net_248) );
DFF_X2 inst_7402 ( .QN(net_8955), .D(net_8414), .CK(net_11766) );
INV_X2 inst_7138 ( .A(net_10247), .ZN(net_829) );
DFF_X2 inst_8169 ( .QN(net_9928), .D(net_5046), .CK(net_12120) );
CLKBUF_X2 inst_12945 ( .A(net_12863), .Z(net_12864) );
AND2_X2 inst_10523 ( .ZN(net_4451), .A1(net_4157), .A2(net_4156) );
CLKBUF_X2 inst_13873 ( .A(net_13791), .Z(net_13792) );
INV_X4 inst_5782 ( .A(net_1031), .ZN(net_985) );
AND2_X2 inst_10520 ( .ZN(net_4449), .A1(net_4172), .A2(net_4171) );
INV_X8 inst_4497 ( .ZN(net_8041), .A(net_5298) );
OAI22_X2 inst_1319 ( .B2(net_9845), .ZN(net_2022), .A2(net_2021), .A1(net_1817), .B1(net_868) );
NOR2_X2 inst_2651 ( .ZN(net_5896), .A2(net_5329), .A1(net_2180) );
INV_X4 inst_4756 ( .ZN(net_4330), .A(net_4329) );
NAND2_X2 inst_4201 ( .A1(net_9519), .ZN(net_2546), .A2(net_1786) );
INV_X4 inst_5658 ( .A(net_10124), .ZN(net_1543) );
XOR2_X2 inst_48 ( .B(net_7595), .Z(net_2929), .A(net_623) );
XNOR2_X2 inst_358 ( .ZN(net_2774), .B(net_2773), .A(net_2048) );
MUX2_X1 inst_4462 ( .S(net_6041), .A(net_284), .B(x5901), .Z(x277) );
OAI21_X2 inst_1756 ( .ZN(net_8508), .A(net_8450), .B2(net_8449), .B1(net_7157) );
OAI211_X2 inst_2246 ( .A(net_8098), .C1(net_7213), .C2(net_6501), .ZN(net_6458), .B(net_5557) );
DFF_X2 inst_7507 ( .QN(net_9374), .D(net_7939), .CK(net_14181) );
CLKBUF_X2 inst_14037 ( .A(net_13955), .Z(net_13956) );
DFF_X1 inst_8794 ( .Q(net_10237), .D(net_4286), .CK(net_10910) );
INV_X2 inst_6766 ( .A(net_6560), .ZN(net_6167) );
CLKBUF_X2 inst_15215 ( .A(net_15133), .Z(net_15134) );
AOI22_X2 inst_9309 ( .B1(net_9714), .A2(net_5755), .B2(net_5754), .ZN(net_5669), .A1(net_251) );
INV_X2 inst_7108 ( .ZN(net_1014), .A(net_1013) );
XNOR2_X2 inst_443 ( .A(net_9651), .ZN(net_877), .B(net_313) );
CLKBUF_X2 inst_14177 ( .A(net_11232), .Z(net_14096) );
CLKBUF_X2 inst_11022 ( .A(net_10940), .Z(net_10941) );
DFF_X1 inst_8766 ( .Q(net_10379), .D(net_5202), .CK(net_14374) );
SDFF_X2 inst_655 ( .SI(net_9480), .Q(net_9480), .SE(net_3073), .CK(net_12419), .D(x2648) );
NAND2_X2 inst_4259 ( .A1(net_10156), .ZN(net_4109), .A2(net_1374) );
INV_X4 inst_5914 ( .ZN(net_1127), .A(net_589) );
CLKBUF_X2 inst_12152 ( .A(net_12070), .Z(net_12071) );
INV_X4 inst_5817 ( .A(net_3032), .ZN(net_675) );
AOI22_X2 inst_9060 ( .B1(net_9681), .A2(net_6684), .B2(net_6683), .ZN(net_6606), .A1(net_250) );
DFF_X1 inst_8422 ( .D(net_8752), .Q(net_242), .CK(net_13891) );
INV_X4 inst_5934 ( .ZN(net_983), .A(net_973) );
AOI22_X2 inst_9373 ( .B1(net_10007), .A2(net_5743), .B2(net_5742), .ZN(net_5532), .A1(net_247) );
OAI221_X2 inst_1700 ( .C1(net_7221), .ZN(net_5453), .B1(net_5452), .B2(net_4477), .C2(net_4455), .A(net_3507) );
CLKBUF_X2 inst_15814 ( .A(net_15732), .Z(net_15733) );
CLKBUF_X2 inst_11316 ( .A(net_11234), .Z(net_11235) );
NOR2_X2 inst_2571 ( .A1(net_9648), .A2(net_9647), .ZN(net_7605) );
MUX2_X1 inst_4438 ( .S(net_6041), .A(net_308), .B(x4209), .Z(x57) );
CLKBUF_X2 inst_12481 ( .A(net_12399), .Z(net_12400) );
INV_X2 inst_6662 ( .ZN(net_8366), .A(net_8312) );
DFF_X1 inst_8800 ( .QN(net_10377), .D(net_4118), .CK(net_12148) );
OR2_X4 inst_730 ( .ZN(net_7171), .A1(net_7170), .A2(net_7038) );
CLKBUF_X2 inst_11430 ( .A(net_10615), .Z(net_11349) );
AOI21_X2 inst_10116 ( .B2(net_10446), .ZN(net_4677), .B1(net_3670), .A(net_3490) );
INV_X4 inst_6303 ( .A(net_9960), .ZN(net_428) );
INV_X2 inst_6754 ( .A(net_7083), .ZN(net_6264) );
XNOR2_X2 inst_321 ( .ZN(net_3033), .B(net_3032), .A(net_2834) );
INV_X4 inst_5623 ( .A(net_873), .ZN(net_863) );
CLKBUF_X2 inst_10977 ( .A(net_10841), .Z(net_10896) );
AOI22_X2 inst_9669 ( .B2(net_10299), .A2(net_10298), .B1(net_10291), .A1(net_10290), .ZN(net_953) );
CLKBUF_X2 inst_11996 ( .A(net_11914), .Z(net_11915) );
CLKBUF_X2 inst_11516 ( .A(net_11434), .Z(net_11435) );
XOR2_X2 inst_41 ( .Z(net_2479), .B(net_2450), .A(net_941) );
CLKBUF_X2 inst_12569 ( .A(net_12487), .Z(net_12488) );
CLKBUF_X2 inst_11743 ( .A(net_11661), .Z(net_11662) );
NAND4_X2 inst_3131 ( .ZN(net_4481), .A3(net_2001), .A2(net_1818), .A4(net_1430), .A1(net_1412) );
CLKBUF_X2 inst_12684 ( .A(net_12602), .Z(net_12603) );
CLKBUF_X2 inst_14788 ( .A(net_13802), .Z(net_14707) );
CLKBUF_X2 inst_13308 ( .A(net_13226), .Z(net_13227) );
CLKBUF_X2 inst_11868 ( .A(net_11786), .Z(net_11787) );
OAI21_X2 inst_1989 ( .B1(net_9735), .ZN(net_2896), .B2(net_2684), .A(net_1794) );
CLKBUF_X2 inst_13260 ( .A(net_13178), .Z(net_13179) );
AOI222_X1 inst_9694 ( .B1(net_9505), .ZN(net_8287), .A2(net_8286), .B2(net_8285), .C2(net_8284), .C1(net_8219), .A1(x1743) );
DFF_X2 inst_8264 ( .Q(net_10386), .D(net_4812), .CK(net_12937) );
XNOR2_X2 inst_152 ( .ZN(net_6645), .A(net_6261), .B(net_2660) );
INV_X4 inst_5609 ( .ZN(net_1134), .A(net_873) );
CLKBUF_X2 inst_11111 ( .A(net_10818), .Z(net_11030) );
INV_X2 inst_6944 ( .ZN(net_1907), .A(net_1906) );
CLKBUF_X2 inst_12314 ( .A(net_12232), .Z(net_12233) );
OAI22_X2 inst_1152 ( .A1(net_7234), .A2(net_5139), .B2(net_5138), .ZN(net_5121), .B1(net_338) );
INV_X2 inst_6878 ( .A(net_3558), .ZN(net_2853) );
INV_X4 inst_6388 ( .A(net_10161), .ZN(net_6960) );
CLKBUF_X2 inst_15255 ( .A(net_10720), .Z(net_15174) );
OAI222_X2 inst_1400 ( .B2(net_7732), .A2(net_7731), .C2(net_7730), .ZN(net_5333), .B1(net_2979), .A1(net_2859), .C1(net_1965) );
CLKBUF_X2 inst_14374 ( .A(net_14292), .Z(net_14293) );
INV_X4 inst_6517 ( .ZN(net_346), .A(net_204) );
XNOR2_X2 inst_89 ( .A(net_8941), .B(net_8935), .ZN(net_8609) );
INV_X4 inst_5233 ( .ZN(net_4204), .A(net_1963) );
OAI221_X2 inst_1520 ( .B2(net_9081), .ZN(net_7300), .C2(net_6265), .A(net_5999), .C1(net_5996), .B1(net_1548) );
INV_X2 inst_6823 ( .ZN(net_4420), .A(net_4419) );
OAI221_X2 inst_1535 ( .C1(net_10211), .C2(net_7295), .B2(net_7293), .ZN(net_7235), .B1(net_7234), .A(net_6866) );
CLKBUF_X2 inst_14112 ( .A(net_10630), .Z(net_14031) );
CLKBUF_X2 inst_13609 ( .A(net_13527), .Z(net_13528) );
DFF_X1 inst_8670 ( .D(net_6752), .Q(net_102), .CK(net_14343) );
XNOR2_X2 inst_182 ( .ZN(net_5245), .A(net_4699), .B(net_2328) );
OR2_X4 inst_788 ( .ZN(net_2261), .A2(net_1756), .A1(net_808) );
CLKBUF_X2 inst_15525 ( .A(net_15443), .Z(net_15444) );
OR2_X2 inst_931 ( .A2(net_8863), .ZN(net_4691), .A1(net_2754) );
AOI22_X2 inst_9205 ( .A1(net_9865), .B1(net_9766), .B2(net_6120), .A2(net_6111), .ZN(net_6106) );
NAND3_X2 inst_3174 ( .A3(net_10090), .ZN(net_8554), .A2(net_8511), .A1(net_7832) );
DFF_X2 inst_7526 ( .QN(net_9537), .D(net_7812), .CK(net_12748) );
CLKBUF_X2 inst_13391 ( .A(net_13309), .Z(net_13310) );
OAI221_X2 inst_1674 ( .B1(net_7213), .C1(net_6289), .C2(net_5591), .ZN(net_5495), .B2(net_4902), .A(net_3527) );
NAND2_X2 inst_3824 ( .A1(net_10530), .ZN(net_4478), .A2(net_4469) );
INV_X4 inst_5990 ( .A(net_10283), .ZN(net_537) );
INV_X2 inst_6895 ( .ZN(net_2588), .A(net_2587) );
CLKBUF_X2 inst_12807 ( .A(net_12583), .Z(net_12726) );
DFF_X1 inst_8438 ( .D(net_8508), .CK(net_10709), .Q(x1010) );
OAI221_X2 inst_1579 ( .B1(net_10209), .B2(net_7295), .C2(net_7293), .ZN(net_7130), .C1(net_7129), .A(net_6923) );
INV_X4 inst_5407 ( .ZN(net_1515), .A(net_664) );
CLKBUF_X2 inst_13482 ( .A(net_13400), .Z(net_13401) );
DFF_X2 inst_8315 ( .QN(net_10166), .D(net_3949), .CK(net_12251) );
XNOR2_X2 inst_193 ( .ZN(net_5202), .A(net_4447), .B(net_2359) );
CLKBUF_X2 inst_14568 ( .A(net_14486), .Z(net_14487) );
NAND2_X2 inst_4089 ( .A1(net_10261), .ZN(net_3105), .A2(net_2532) );
CLKBUF_X2 inst_14320 ( .A(net_13981), .Z(net_14239) );
CLKBUF_X2 inst_11704 ( .A(net_11432), .Z(net_11623) );
OAI222_X2 inst_1415 ( .A2(net_7665), .C2(net_7664), .B2(net_7663), .ZN(net_5195), .C1(net_2882), .A1(net_2273), .B1(net_1291) );
OAI221_X2 inst_1709 ( .B2(net_7437), .ZN(net_4001), .B1(net_3290), .A(net_2888), .C2(net_2635), .C1(net_2240) );
CLKBUF_X2 inst_15358 ( .A(net_15276), .Z(net_15277) );
CLKBUF_X2 inst_12089 ( .A(net_12007), .Z(net_12008) );
CLKBUF_X2 inst_13631 ( .A(net_13549), .Z(net_13550) );
NAND3_X2 inst_3301 ( .ZN(net_3492), .A2(net_2419), .A1(net_1701), .A3(net_1647) );
INV_X4 inst_5997 ( .A(net_9974), .ZN(net_533) );
INV_X4 inst_6469 ( .A(net_9850), .ZN(net_3433) );
OAI211_X2 inst_2202 ( .C1(net_7190), .C2(net_6542), .ZN(net_6505), .B(net_5602), .A(net_3527) );
DFF_X2 inst_7531 ( .QN(net_9324), .D(net_7778), .CK(net_13053) );
CLKBUF_X2 inst_11673 ( .A(net_11591), .Z(net_11592) );
NAND3_X2 inst_3180 ( .ZN(net_8129), .A1(net_8056), .A3(net_7969), .A2(net_3379) );
DFF_X2 inst_7969 ( .QN(net_10320), .D(net_5584), .CK(net_15585) );
INV_X4 inst_4737 ( .ZN(net_4789), .A(net_4462) );
AOI221_X2 inst_9965 ( .C1(net_9704), .B2(net_5173), .ZN(net_4766), .A(net_4337), .C2(net_3039), .B1(net_207) );
AND2_X2 inst_10618 ( .A1(net_9212), .ZN(net_2164), .A2(net_1567) );
NOR2_X2 inst_2987 ( .A1(net_10148), .ZN(net_1717), .A2(net_501) );
CLKBUF_X2 inst_12571 ( .A(net_12489), .Z(net_12490) );
CLKBUF_X2 inst_15162 ( .A(net_15080), .Z(net_15081) );
CLKBUF_X2 inst_11645 ( .A(net_11563), .Z(net_11564) );
CLKBUF_X2 inst_13433 ( .A(net_10705), .Z(net_13352) );
INV_X4 inst_5578 ( .ZN(net_1273), .A(net_1094) );
CLKBUF_X2 inst_11853 ( .A(net_10603), .Z(net_11772) );
INV_X4 inst_5884 ( .A(net_2302), .ZN(net_867) );
CLKBUF_X2 inst_13396 ( .A(net_13314), .Z(net_13315) );
CLKBUF_X2 inst_11170 ( .A(net_11088), .Z(net_11089) );
DFF_X1 inst_8655 ( .Q(net_9764), .D(net_7191), .CK(net_15447) );
CLKBUF_X2 inst_11459 ( .A(net_11360), .Z(net_11378) );
INV_X4 inst_4599 ( .ZN(net_7805), .A(net_7709) );
DFF_X2 inst_8147 ( .QN(net_10042), .D(net_5087), .CK(net_12485) );
INV_X4 inst_5906 ( .A(net_1210), .ZN(net_828) );
INV_X4 inst_4677 ( .A(net_5393), .ZN(net_5391) );
CLKBUF_X2 inst_12874 ( .A(net_12424), .Z(net_12793) );
CLKBUF_X2 inst_14796 ( .A(net_14714), .Z(net_14715) );
NOR2_X4 inst_2473 ( .ZN(net_9026), .A1(net_8517), .A2(net_8516) );
INV_X4 inst_5516 ( .A(net_4978), .ZN(net_1262) );
OAI221_X2 inst_1698 ( .B1(net_7224), .A(net_6546), .C2(net_5642), .ZN(net_5456), .B2(net_4905), .C1(net_2232) );
CLKBUF_X2 inst_11698 ( .A(net_11213), .Z(net_11617) );
OR2_X2 inst_944 ( .A2(net_10430), .A1(net_10429), .ZN(net_1197) );
INV_X4 inst_5248 ( .ZN(net_5331), .A(net_1476) );
INV_X2 inst_7125 ( .ZN(net_1217), .A(net_174) );
CLKBUF_X2 inst_12442 ( .A(net_12360), .Z(net_12361) );
INV_X8 inst_4516 ( .A(net_8924), .ZN(net_8918) );
CLKBUF_X2 inst_15488 ( .A(net_15406), .Z(net_15407) );
DFF_X2 inst_7992 ( .QN(net_10419), .D(net_5534), .CK(net_15576) );
CLKBUF_X2 inst_13952 ( .A(net_13870), .Z(net_13871) );
SDFF_X2 inst_459 ( .SE(net_8747), .SI(net_8722), .Q(net_240), .D(net_109), .CK(net_13861) );
DFF_X2 inst_8259 ( .Q(net_10285), .D(net_4822), .CK(net_12940) );
CLKBUF_X2 inst_11737 ( .A(net_11655), .Z(net_11656) );
DFF_X1 inst_8532 ( .Q(net_9966), .D(net_7328), .CK(net_12837) );
NOR2_X2 inst_2864 ( .ZN(net_2713), .A2(net_2053), .A1(net_558) );
CLKBUF_X2 inst_14645 ( .A(net_13861), .Z(net_14564) );
NAND2_X2 inst_3476 ( .A1(net_9455), .A2(net_8951), .ZN(net_8909) );
AOI21_X2 inst_10084 ( .B2(net_10133), .A(net_10132), .ZN(net_5395), .B1(net_1579) );
DFF_X2 inst_7461 ( .QN(net_9638), .D(net_8123), .CK(net_15378) );
CLKBUF_X2 inst_12861 ( .A(net_11673), .Z(net_12780) );
NAND2_X2 inst_3789 ( .ZN(net_6680), .A2(net_5918), .A1(net_4634) );
CLKBUF_X2 inst_15001 ( .A(net_14919), .Z(net_14920) );
INV_X2 inst_7096 ( .A(net_5317), .ZN(net_1084) );
CLKBUF_X2 inst_13723 ( .A(net_13641), .Z(net_13642) );
NAND2_X2 inst_3393 ( .ZN(net_9003), .A1(net_8878), .A2(net_8701) );
DFF_X1 inst_8613 ( .Q(net_9877), .D(net_7180), .CK(net_13290) );
XNOR2_X2 inst_367 ( .B(net_9617), .ZN(net_2520), .A(net_2197) );
DFF_X2 inst_8148 ( .Q(net_10046), .D(net_5085), .CK(net_14725) );
CLKBUF_X2 inst_11589 ( .A(net_11030), .Z(net_11508) );
OAI33_X1 inst_957 ( .B1(net_6041), .A1(net_5442), .A3(net_4638), .A2(net_4608), .B3(net_4326), .B2(net_314), .ZN(x0) );
INV_X4 inst_4976 ( .ZN(net_4642), .A(net_2291) );
AOI22_X2 inst_9657 ( .ZN(net_2698), .A1(net_2204), .A2(net_2203), .B1(net_2202), .B2(net_1656) );
NAND2_X2 inst_3409 ( .ZN(net_9006), .A1(net_8474), .A2(net_8472) );
OAI21_X2 inst_1871 ( .ZN(net_5293), .A(net_5292), .B2(net_4367), .B1(x4587) );
CLKBUF_X2 inst_13252 ( .A(net_13170), .Z(net_13171) );
NAND2_X2 inst_3591 ( .ZN(net_9067), .A2(net_7033), .A1(net_3384) );
OAI211_X2 inst_2300 ( .ZN(net_4039), .B(net_3598), .C2(net_3165), .A(net_2721), .C1(net_1959) );
INV_X4 inst_5970 ( .A(net_10221), .ZN(net_1947) );
INV_X4 inst_6460 ( .A(net_9940), .ZN(net_3644) );
DFF_X2 inst_7552 ( .QN(net_9355), .D(net_7708), .CK(net_15311) );
CLKBUF_X2 inst_10800 ( .A(net_10620), .Z(net_10719) );
XNOR2_X1 inst_450 ( .ZN(net_7053), .A(net_7052), .B(net_2353) );
AOI222_X1 inst_9723 ( .C1(net_9870), .B1(net_9771), .A2(net_6413), .A1(net_6056), .ZN(net_4055), .C2(net_2973), .B2(net_2462) );
CLKBUF_X2 inst_11694 ( .A(net_11612), .Z(net_11613) );
OR2_X4 inst_745 ( .A1(net_9356), .ZN(net_7721), .A2(net_6190) );
SDFF_X2 inst_520 ( .Q(net_9336), .D(net_9336), .SI(net_9328), .SE(net_7588), .CK(net_14691) );
INV_X4 inst_5717 ( .A(net_767), .ZN(net_764) );
NAND2_X2 inst_3658 ( .A2(net_10380), .ZN(net_6644), .A1(net_1956) );
INV_X2 inst_7024 ( .ZN(net_2380), .A(net_1516) );
AOI21_X2 inst_10019 ( .ZN(net_8293), .A(net_8082), .B1(net_7987), .B2(net_7986) );
CLKBUF_X2 inst_11622 ( .A(net_11540), .Z(net_11541) );
CLKBUF_X2 inst_11667 ( .A(net_10780), .Z(net_11586) );
OAI211_X2 inst_2032 ( .ZN(net_8103), .C2(net_8102), .A(net_8003), .B(net_3507), .C1(net_1705) );
INV_X4 inst_4554 ( .ZN(net_8550), .A(net_8515) );
CLKBUF_X2 inst_14850 ( .A(net_14768), .Z(net_14769) );
INV_X4 inst_5977 ( .A(net_9247), .ZN(net_664) );
NAND2_X2 inst_4113 ( .ZN(net_2356), .A2(net_2355), .A1(net_1640) );
OAI211_X2 inst_2026 ( .ZN(net_8448), .B(net_8447), .C2(net_8256), .C1(net_4763), .A(x987) );
XNOR2_X2 inst_80 ( .ZN(net_8633), .A(net_8592), .B(net_8392) );
NAND2_X2 inst_3623 ( .ZN(net_7103), .A1(net_6890), .A2(net_6675) );
OR2_X4 inst_836 ( .A2(net_10466), .A1(net_10465), .ZN(net_2419) );
DFF_X2 inst_7698 ( .QN(net_9503), .D(net_6985), .CK(net_12733) );
OAI221_X2 inst_1556 ( .C2(net_7295), .B2(net_7293), .B1(net_7219), .ZN(net_7200), .A(net_6824), .C1(net_917) );
AOI22_X2 inst_9228 ( .A1(net_9922), .B1(net_9823), .A2(net_8042), .B2(net_8041), .ZN(net_6083) );
CLKBUF_X2 inst_14820 ( .A(net_10969), .Z(net_14739) );
AOI22_X2 inst_9521 ( .B1(net_9701), .A1(net_9669), .A2(net_5966), .ZN(net_3801), .B2(net_3039) );
DFF_X1 inst_8821 ( .QN(net_10277), .D(net_3164), .CK(net_10618) );
INV_X2 inst_6796 ( .ZN(net_5414), .A(net_5413) );
CLKBUF_X2 inst_15636 ( .A(net_15554), .Z(net_15555) );
CLKBUF_X2 inst_10771 ( .A(net_10689), .Z(net_10690) );
INV_X4 inst_6564 ( .A(net_10036), .ZN(net_328) );
CLKBUF_X2 inst_11243 ( .A(net_11161), .Z(net_11162) );
AOI22_X2 inst_9562 ( .A1(net_10392), .B1(net_9876), .A2(net_4062), .ZN(net_3757), .B2(net_2973) );
CLKBUF_X2 inst_12075 ( .A(net_11993), .Z(net_11994) );
XNOR2_X2 inst_241 ( .ZN(net_4254), .A(net_4253), .B(net_2065) );
NAND2_X2 inst_4409 ( .A2(net_10195), .A1(net_10187), .ZN(net_607) );
INV_X4 inst_5120 ( .ZN(net_1614), .A(net_1613) );
CLKBUF_X2 inst_14705 ( .A(net_14623), .Z(net_14624) );
INV_X4 inst_4934 ( .ZN(net_2593), .A(net_2592) );
CLKBUF_X2 inst_15384 ( .A(net_15302), .Z(net_15303) );
CLKBUF_X2 inst_14410 ( .A(net_14328), .Z(net_14329) );
OR2_X2 inst_862 ( .A1(net_10293), .ZN(net_7866), .A2(net_7865) );
NAND2_X2 inst_4358 ( .A2(net_10226), .ZN(net_2094), .A1(net_962) );
NAND2_X2 inst_4390 ( .A2(net_10432), .ZN(net_1759), .A1(net_364) );
INV_X2 inst_6690 ( .ZN(net_8334), .A(net_8272) );
CLKBUF_X2 inst_15534 ( .A(net_15452), .Z(net_15453) );
CLKBUF_X2 inst_14142 ( .A(net_14060), .Z(net_14061) );
CLKBUF_X2 inst_13491 ( .A(net_13409), .Z(net_13410) );
NAND2_X2 inst_3918 ( .A2(net_9053), .ZN(net_7963), .A1(net_680) );
CLKBUF_X2 inst_14618 ( .A(net_14536), .Z(net_14537) );
NOR2_X2 inst_2758 ( .A2(net_10280), .ZN(net_4073), .A1(net_3872) );
OAI22_X2 inst_1116 ( .A1(net_8985), .ZN(net_5427), .B2(net_4993), .A2(net_4991), .B1(net_1435) );
INV_X8 inst_4504 ( .ZN(net_6109), .A(net_5296) );
DFF_X2 inst_7947 ( .QN(net_10350), .D(net_5702), .CK(net_13647) );
AND2_X2 inst_10620 ( .A1(net_9616), .ZN(net_2197), .A2(net_1545) );
NAND2_X2 inst_3753 ( .ZN(net_5294), .A2(net_4778), .A1(net_3755) );
INV_X4 inst_5545 ( .ZN(net_939), .A(net_938) );
OAI21_X2 inst_1764 ( .ZN(net_8370), .B2(net_8369), .B1(net_8338), .A(net_8095) );
CLKBUF_X2 inst_14024 ( .A(net_13942), .Z(net_13943) );
INV_X4 inst_5271 ( .A(net_5407), .ZN(net_2192) );
CLKBUF_X2 inst_12050 ( .A(net_11968), .Z(net_11969) );
CLKBUF_X2 inst_14799 ( .A(net_14717), .Z(net_14718) );
INV_X4 inst_5323 ( .ZN(net_3920), .A(net_3172) );
CLKBUF_X2 inst_15366 ( .A(net_11613), .Z(net_15285) );
DFF_X2 inst_7472 ( .QN(net_9520), .D(net_8039), .CK(net_14962) );
CLKBUF_X2 inst_11555 ( .A(net_11473), .Z(net_11474) );
OAI22_X2 inst_1159 ( .A1(net_7203), .A2(net_5139), .B2(net_5138), .ZN(net_5114), .B1(net_556) );
DFF_X1 inst_8740 ( .Q(net_9144), .D(net_5728), .CK(net_11040) );
AOI22_X2 inst_9550 ( .A1(net_9936), .B1(net_9805), .A2(net_6443), .ZN(net_3770), .B2(net_2556) );
DFF_X1 inst_8659 ( .Q(net_9868), .D(net_7250), .CK(net_13342) );
XNOR2_X2 inst_402 ( .A(net_9158), .B(net_9157), .ZN(net_2469) );
NAND4_X2 inst_3136 ( .ZN(net_5337), .A4(net_5272), .A2(net_2912), .A3(net_2911), .A1(net_920) );
INV_X4 inst_6394 ( .A(net_10049), .ZN(net_702) );
CLKBUF_X2 inst_10962 ( .A(net_10880), .Z(net_10881) );
CLKBUF_X2 inst_11259 ( .A(net_11177), .Z(net_11178) );
AOI221_X2 inst_9835 ( .A(net_6889), .B2(net_6888), .C2(net_6887), .ZN(net_6883), .B1(net_5854), .C1(x5225) );
CLKBUF_X2 inst_13025 ( .A(net_12943), .Z(net_12944) );
OR2_X2 inst_938 ( .A1(net_9179), .ZN(net_2196), .A2(net_2195) );
CLKBUF_X2 inst_14521 ( .A(net_14439), .Z(net_14440) );
INV_X4 inst_5832 ( .A(net_2091), .ZN(net_660) );
CLKBUF_X2 inst_12815 ( .A(net_11086), .Z(net_12734) );
CLKBUF_X2 inst_11189 ( .A(net_10783), .Z(net_11108) );
HA_X1 inst_7350 ( .S(net_4428), .CO(net_4427), .B(net_4268), .A(net_539) );
CLKBUF_X2 inst_12552 ( .A(net_12470), .Z(net_12471) );
OAI22_X2 inst_1288 ( .A1(net_4509), .A2(net_4085), .ZN(net_3915), .B2(net_3914), .B1(net_1953) );
NAND2_X2 inst_3844 ( .ZN(net_4862), .A2(net_4238), .A1(net_3072) );
CLKBUF_X2 inst_12742 ( .A(net_12660), .Z(net_12661) );
INV_X4 inst_6646 ( .A(net_9109), .ZN(net_9108) );
AOI222_X1 inst_9698 ( .B1(net_9509), .A2(net_8286), .B2(net_8285), .C2(net_8284), .ZN(net_8280), .C1(net_8216), .A1(x1503) );
DFF_X2 inst_7610 ( .QN(net_9345), .D(net_7133), .CK(net_15284) );
NAND2_X2 inst_3638 ( .A2(net_9378), .ZN(net_7700), .A1(net_7505) );
NAND2_X2 inst_4365 ( .A2(net_10141), .ZN(net_1200), .A1(net_707) );
CLKBUF_X2 inst_11329 ( .A(net_10987), .Z(net_11248) );
AOI22_X2 inst_9399 ( .A1(net_6892), .B2(net_6625), .ZN(net_6182), .B1(net_5374), .A2(net_4666) );
CLKBUF_X2 inst_11845 ( .A(net_11763), .Z(net_11764) );
OAI22_X2 inst_1033 ( .A1(net_9092), .B1(net_8919), .A2(net_8915), .ZN(net_7951), .B2(net_1573) );
CLKBUF_X2 inst_11320 ( .A(net_11238), .Z(net_11239) );
INV_X4 inst_4673 ( .ZN(net_5823), .A(net_5259) );
CLKBUF_X2 inst_14253 ( .A(net_14171), .Z(net_14172) );
CLKBUF_X2 inst_14201 ( .A(net_14119), .Z(net_14120) );
INV_X4 inst_5582 ( .A(net_10325), .ZN(net_1285) );
OAI222_X2 inst_1348 ( .B1(net_7728), .A2(net_7727), .C2(net_7726), .ZN(net_7433), .B2(net_7053), .A1(net_4682), .C1(net_695) );
DFF_X2 inst_7426 ( .QN(net_9398), .D(net_8332), .CK(net_14008) );
OAI211_X2 inst_2102 ( .C2(net_6778), .ZN(net_6746), .A(net_6374), .B(net_6104), .C1(net_504) );
INV_X4 inst_5427 ( .A(net_6255), .ZN(net_5041) );
CLKBUF_X2 inst_14070 ( .A(net_12000), .Z(net_13989) );
AOI221_X2 inst_9762 ( .ZN(net_7657), .B1(net_7642), .C2(net_7641), .A(net_7533), .B2(net_5951), .C1(net_5411) );
OAI21_X2 inst_1748 ( .B2(net_8812), .ZN(net_8666), .A(net_8636), .B1(net_370) );
INV_X4 inst_4908 ( .A(net_3105), .ZN(net_2839) );
INV_X2 inst_7160 ( .A(net_7029), .ZN(net_635) );
CLKBUF_X2 inst_15686 ( .A(net_15604), .Z(net_15605) );
DFF_X2 inst_7619 ( .D(net_9543), .Q(net_9542), .CK(net_13980) );
CLKBUF_X2 inst_11423 ( .A(net_11341), .Z(net_11342) );
HA_X1 inst_7356 ( .CO(net_3161), .S(net_2736), .A(net_1875), .B(net_875) );
AND4_X2 inst_10343 ( .A1(net_5168), .A2(net_5167), .A4(net_5166), .ZN(net_5162), .A3(net_625) );
INV_X4 inst_6168 ( .A(net_9849), .ZN(net_476) );
DFF_X1 inst_8445 ( .Q(net_9432), .D(net_8170), .CK(net_14931) );
INV_X4 inst_5565 ( .ZN(net_6658), .A(net_913) );
CLKBUF_X2 inst_14781 ( .A(net_10892), .Z(net_14700) );
CLKBUF_X2 inst_11684 ( .A(net_11602), .Z(net_11603) );
CLKBUF_X2 inst_11864 ( .A(net_11782), .Z(net_11783) );
CLKBUF_X2 inst_14058 ( .A(net_13976), .Z(net_13977) );
CLKBUF_X2 inst_11182 ( .A(net_11100), .Z(net_11101) );
AOI21_X2 inst_10145 ( .B1(net_7583), .A(net_4512), .ZN(net_4208), .B2(net_4016) );
AOI222_X1 inst_9712 ( .C2(net_10347), .B1(net_10346), .ZN(net_7876), .A2(net_7793), .B2(net_7610), .C1(net_7479), .A1(net_7458) );
DFF_X1 inst_8637 ( .Q(net_9887), .D(net_7195), .CK(net_14384) );
AOI22_X2 inst_9216 ( .A1(net_9909), .B1(net_9810), .B2(net_6133), .A2(net_6111), .ZN(net_6095) );
OR2_X4 inst_784 ( .A2(net_2400), .ZN(net_2323), .A1(net_2322) );
NAND3_X2 inst_3237 ( .A1(net_7142), .ZN(net_4720), .A3(net_4719), .A2(net_4041) );
CLKBUF_X2 inst_11088 ( .A(net_11006), .Z(net_11007) );
OAI22_X2 inst_1264 ( .B1(net_7186), .A2(net_4842), .B2(net_4841), .ZN(net_4809), .A1(net_389) );
CLKBUF_X2 inst_12046 ( .A(net_10576), .Z(net_11965) );
OR3_X4 inst_690 ( .ZN(net_7659), .A3(net_4979), .A2(net_4978), .A1(net_4221) );
INV_X4 inst_6397 ( .A(net_10461), .ZN(net_963) );
CLKBUF_X2 inst_11895 ( .A(net_11813), .Z(net_11814) );
OAI211_X2 inst_2025 ( .ZN(net_8450), .B(net_8449), .C2(net_8260), .C1(net_4514), .A(x1010) );
HA_X1 inst_7337 ( .CO(net_7323), .S(net_6957), .A(net_6956), .B(net_5987) );
NOR2_X4 inst_2461 ( .A1(net_8872), .ZN(net_8785), .A2(net_3932) );
DFF_X2 inst_7819 ( .QN(net_9178), .D(net_6301), .CK(net_11314) );
AND2_X2 inst_10607 ( .A1(net_2685), .ZN(net_2024), .A2(net_2023) );
DFF_X1 inst_8814 ( .QN(net_10130), .D(net_3497), .CK(net_10764) );
OR2_X4 inst_732 ( .A2(net_7038), .ZN(net_6586), .A1(net_6585) );
INV_X4 inst_4717 ( .ZN(net_7846), .A(net_5973) );
CLKBUF_X2 inst_12722 ( .A(net_11403), .Z(net_12641) );
CLKBUF_X2 inst_13044 ( .A(net_11184), .Z(net_12963) );
CLKBUF_X2 inst_12183 ( .A(net_11506), .Z(net_12102) );
CLKBUF_X2 inst_10969 ( .A(net_10596), .Z(net_10888) );
AOI22_X2 inst_9666 ( .B2(net_10404), .A2(net_10403), .B1(net_10396), .A1(net_10395), .ZN(net_964) );
DFF_X2 inst_8023 ( .QN(net_10221), .D(net_5470), .CK(net_14457) );
XNOR2_X2 inst_75 ( .ZN(net_8664), .A(net_8621), .B(net_2725) );
INV_X4 inst_5968 ( .A(net_9993), .ZN(net_548) );
DFF_X2 inst_7714 ( .Q(net_9707), .D(net_6471), .CK(net_12577) );
CLKBUF_X2 inst_15656 ( .A(net_15574), .Z(net_15575) );
INV_X4 inst_6386 ( .A(net_9241), .ZN(net_723) );
XNOR2_X2 inst_79 ( .ZN(net_8634), .A(net_8594), .B(net_8337) );
CLKBUF_X2 inst_11250 ( .A(net_11168), .Z(net_11169) );
DFF_X2 inst_7986 ( .QN(net_10412), .D(net_5599), .CK(net_14586) );
NOR2_X2 inst_2654 ( .A1(net_9528), .ZN(net_5800), .A2(net_5258) );
INV_X2 inst_7088 ( .ZN(net_1140), .A(net_1139) );
AOI22_X2 inst_9286 ( .B1(net_9704), .A1(net_5755), .B2(net_5754), .ZN(net_5714), .A2(net_241) );
DFF_X2 inst_7600 ( .Q(net_9980), .D(net_7366), .CK(net_14758) );
CLKBUF_X2 inst_11662 ( .A(net_11345), .Z(net_11581) );
DFF_X2 inst_7891 ( .QN(net_10097), .D(net_6024), .CK(net_15530) );
CLKBUF_X2 inst_12082 ( .A(net_10815), .Z(net_12001) );
CLKBUF_X2 inst_11962 ( .A(net_11880), .Z(net_11881) );
DFF_X1 inst_8838 ( .QN(net_9957), .D(net_2160), .CK(net_11221) );
DFF_X2 inst_7895 ( .QN(net_10102), .D(net_6018), .CK(net_14906) );
CLKBUF_X2 inst_13938 ( .A(net_12897), .Z(net_13857) );
CLKBUF_X2 inst_10890 ( .A(net_10808), .Z(net_10809) );
NAND2_X2 inst_4413 ( .A2(net_10300), .A1(net_10292), .ZN(net_579) );
OAI21_X2 inst_1741 ( .B1(net_8945), .A(net_8852), .ZN(net_8717), .B2(net_8695) );
NOR2_X2 inst_2975 ( .A2(net_9212), .ZN(net_1638), .A1(net_769) );
AND4_X4 inst_10339 ( .ZN(net_3210), .A3(net_2430), .A1(net_2181), .A4(net_2068), .A2(net_1302) );
OAI22_X2 inst_1024 ( .A2(net_8036), .B2(net_8018), .ZN(net_8014), .A1(net_3333), .B1(net_651) );
INV_X4 inst_5827 ( .ZN(net_949), .A(net_667) );
INV_X4 inst_5594 ( .A(net_1225), .ZN(net_1168) );
CLKBUF_X2 inst_12144 ( .A(net_12062), .Z(net_12063) );
OAI211_X2 inst_2232 ( .C1(net_7219), .C2(net_6480), .ZN(net_6472), .B(net_5622), .A(net_3679) );
INV_X4 inst_4546 ( .ZN(net_8586), .A(net_8581) );
CLKBUF_X2 inst_13218 ( .A(net_13136), .Z(net_13137) );
OAI221_X2 inst_1658 ( .C1(net_7209), .ZN(net_5514), .B1(net_5513), .B2(net_4477), .C2(net_4455), .A(net_3731) );
CLKBUF_X2 inst_14991 ( .A(net_14909), .Z(net_14910) );
INV_X4 inst_6515 ( .A(net_9947), .ZN(net_348) );
CLKBUF_X2 inst_12061 ( .A(net_11979), .Z(net_11980) );
OAI221_X2 inst_1689 ( .C1(net_7203), .B2(net_5642), .ZN(net_5471), .C2(net_4905), .A(net_3731), .B1(net_1580) );
AOI22_X2 inst_9003 ( .A2(net_9956), .B2(net_9857), .ZN(net_8079), .A1(net_8042), .B1(net_8041) );
DFF_X2 inst_8279 ( .QN(net_10261), .D(net_4913), .CK(net_12182) );
NOR2_X2 inst_2846 ( .A2(net_6956), .ZN(net_2259), .A1(net_1520) );
NAND2_X2 inst_3965 ( .A2(net_6625), .ZN(net_3384), .A1(net_279) );
NAND2_X2 inst_4267 ( .A2(net_10436), .A1(net_10435), .ZN(net_2709) );
NAND2_X2 inst_3584 ( .ZN(net_7397), .A2(net_7396), .A1(net_5915) );
CLKBUF_X2 inst_11408 ( .A(net_11273), .Z(net_11327) );
AOI22_X2 inst_9472 ( .B1(net_9811), .A1(net_9680), .A2(net_5966), .ZN(net_3851), .B2(net_2556) );
OAI221_X2 inst_1448 ( .B2(net_9633), .B1(net_8980), .ZN(net_8178), .A(net_7971), .C2(net_3526), .C1(net_177) );
CLKBUF_X2 inst_12829 ( .A(net_12198), .Z(net_12748) );
DFF_X2 inst_8395 ( .Q(net_9152), .CK(net_11796), .D(x3621) );
OAI21_X2 inst_1816 ( .B2(net_7846), .ZN(net_6670), .A(net_6009), .B1(net_5261) );
XNOR2_X2 inst_440 ( .B(net_9220), .A(net_9219), .ZN(net_961) );
CLKBUF_X2 inst_11892 ( .A(net_11256), .Z(net_11811) );
CLKBUF_X2 inst_11723 ( .A(net_11641), .Z(net_11642) );
CLKBUF_X2 inst_14829 ( .A(net_14747), .Z(net_14748) );
CLKBUF_X2 inst_14386 ( .A(net_14304), .Z(net_14305) );
INV_X4 inst_5012 ( .ZN(net_2127), .A(net_1758) );
INV_X4 inst_4927 ( .ZN(net_5745), .A(net_2407) );
NAND2_X2 inst_3381 ( .ZN(net_8788), .A2(net_8784), .A1(net_7857) );
CLKBUF_X2 inst_14123 ( .A(net_14041), .Z(net_14042) );
CLKBUF_X2 inst_15423 ( .A(net_12177), .Z(net_15342) );
CLKBUF_X2 inst_15287 ( .A(net_15205), .Z(net_15206) );
OAI21_X2 inst_1887 ( .B2(net_10341), .A(net_10340), .ZN(net_4928), .B1(net_4927) );
OAI22_X2 inst_1091 ( .A2(net_9064), .B2(net_6639), .ZN(net_6556), .B1(net_3274), .A1(net_334) );
CLKBUF_X2 inst_11708 ( .A(net_10706), .Z(net_11627) );
CLKBUF_X2 inst_15108 ( .A(net_15026), .Z(net_15027) );
AOI221_X2 inst_9915 ( .B1(net_10509), .ZN(net_6417), .B2(net_6415), .C2(net_6413), .C1(net_6044), .A(net_5689) );
INV_X4 inst_4837 ( .ZN(net_4784), .A(net_3298) );
INV_X4 inst_5059 ( .A(net_3960), .ZN(net_2242) );
DFF_X2 inst_8206 ( .Q(net_10083), .D(net_4852), .CK(net_10691) );
AND2_X4 inst_10450 ( .A1(net_9345), .ZN(net_2368), .A2(net_1363) );
NAND2_X2 inst_3579 ( .A1(net_9065), .A2(net_8659), .ZN(net_7510) );
CLKBUF_X2 inst_13800 ( .A(net_13718), .Z(net_13719) );
NAND2_X2 inst_4154 ( .ZN(net_2040), .A2(net_1765), .A1(net_1360) );
AND3_X2 inst_10374 ( .ZN(net_4231), .A2(net_4230), .A3(net_4229), .A1(x6599) );
INV_X4 inst_5688 ( .A(net_2780), .ZN(net_798) );
INV_X4 inst_5398 ( .ZN(net_1590), .A(net_1168) );
OAI221_X2 inst_1672 ( .C1(net_7219), .ZN(net_5497), .B2(net_4477), .C2(net_4455), .A(net_3507), .B1(net_843) );
INV_X4 inst_4816 ( .ZN(net_4028), .A(net_3059) );
CLKBUF_X2 inst_13705 ( .A(net_12974), .Z(net_13624) );
CLKBUF_X2 inst_12120 ( .A(net_11198), .Z(net_12039) );
DFF_X1 inst_8625 ( .Q(net_9783), .D(net_7218), .CK(net_13365) );
OAI21_X2 inst_2015 ( .B1(net_10463), .ZN(net_2435), .A(net_1172), .B2(net_1118) );
CLKBUF_X2 inst_12108 ( .A(net_12026), .Z(net_12027) );
NAND3_X2 inst_3179 ( .ZN(net_8130), .A1(net_8055), .A3(net_7967), .A2(net_3377) );
NAND4_X2 inst_3059 ( .ZN(net_5727), .A4(net_4769), .A3(net_4214), .A2(net_3823), .A1(net_3432) );
NAND2_X2 inst_3937 ( .ZN(net_5685), .A2(net_3553), .A1(net_1476) );
NOR2_X2 inst_2970 ( .A1(net_10140), .ZN(net_1741), .A2(net_1071) );
CLKBUF_X2 inst_15297 ( .A(net_12225), .Z(net_15216) );
CLKBUF_X2 inst_14488 ( .A(net_14406), .Z(net_14407) );
CLKBUF_X2 inst_11357 ( .A(net_11275), .Z(net_11276) );
CLKBUF_X2 inst_11950 ( .A(net_11868), .Z(net_11869) );
CLKBUF_X2 inst_15660 ( .A(net_15578), .Z(net_15579) );
CLKBUF_X2 inst_10942 ( .A(net_10566), .Z(net_10861) );
AOI22_X2 inst_9281 ( .B1(net_9997), .A1(net_5743), .B2(net_5742), .ZN(net_5737), .A2(net_237) );
DFF_X2 inst_8278 ( .QN(net_10260), .D(net_4912), .CK(net_12186) );
NAND2_X2 inst_4085 ( .ZN(net_3875), .A2(net_2601), .A1(net_1593) );
CLKBUF_X2 inst_14719 ( .A(net_14598), .Z(net_14638) );
AOI22_X2 inst_9390 ( .B1(net_9806), .A1(net_5766), .B2(net_5765), .ZN(net_5430), .A2(net_244) );
CLKBUF_X2 inst_13183 ( .A(net_13101), .Z(net_13102) );
NOR2_X2 inst_2587 ( .A1(net_7274), .ZN(net_7055), .A2(net_7054) );
INV_X4 inst_4990 ( .ZN(net_2547), .A(net_2224) );
INV_X4 inst_5664 ( .ZN(net_1293), .A(net_896) );
AND4_X4 inst_10317 ( .ZN(net_8962), .A1(net_8577), .A4(net_8572), .A2(net_8553), .A3(net_8413) );
CLKBUF_X2 inst_12285 ( .A(net_12203), .Z(net_12204) );
INV_X2 inst_6680 ( .ZN(net_8348), .A(net_8282) );
DFF_X1 inst_8868 ( .Q(net_9507), .D(net_9283), .CK(net_13732) );
AOI22_X2 inst_9442 ( .ZN(net_4207), .B2(net_4206), .A2(net_2969), .A1(net_2792), .B1(net_746) );
CLKBUF_X2 inst_11090 ( .A(net_11008), .Z(net_11009) );
CLKBUF_X2 inst_13072 ( .A(net_12990), .Z(net_12991) );
OR2_X4 inst_815 ( .ZN(net_2144), .A2(net_883), .A1(net_560) );
DFF_X1 inst_8883 ( .Q(net_9506), .D(net_9282), .CK(net_14484) );
NOR2_X1 inst_3031 ( .ZN(net_2606), .A2(net_2605), .A1(net_1949) );
CLKBUF_X2 inst_15433 ( .A(net_13289), .Z(net_15352) );
OAI211_X2 inst_2165 ( .C1(net_7182), .C2(net_6548), .ZN(net_6545), .B(net_5672), .A(net_3679) );
OAI22_X2 inst_1257 ( .B1(net_7203), .A2(net_4826), .B2(net_4825), .ZN(net_4816), .A1(net_347) );
OR2_X2 inst_875 ( .A1(net_10293), .ZN(net_6973), .A2(net_6972) );
NAND3_X2 inst_3298 ( .ZN(net_2637), .A2(net_2636), .A1(net_1517), .A3(net_945) );
NAND4_X2 inst_3081 ( .A3(net_10385), .ZN(net_4797), .A4(net_4641), .A1(net_4516), .A2(net_4180) );
NAND2_X2 inst_3482 ( .A1(net_9548), .ZN(net_8425), .A2(net_8424) );
CLKBUF_X2 inst_12096 ( .A(net_12014), .Z(net_12015) );
INV_X4 inst_5075 ( .A(net_1832), .ZN(net_1830) );
INV_X4 inst_5187 ( .ZN(net_1553), .A(net_1552) );
OAI211_X2 inst_2069 ( .ZN(net_7401), .A(net_7300), .B(net_6264), .C1(net_5419), .C2(net_5267) );
DFF_X2 inst_8227 ( .D(net_4865), .Q(net_230), .CK(net_11124) );
INV_X2 inst_7006 ( .A(net_2395), .ZN(net_1610) );
CLKBUF_X2 inst_15032 ( .A(net_12746), .Z(net_14951) );
OAI211_X2 inst_2108 ( .C2(net_6778), .ZN(net_6740), .A(net_6366), .B(net_6098), .C1(net_318) );
NAND2_X2 inst_3572 ( .A1(net_8801), .A2(net_7753), .ZN(net_7701) );
NAND2_X2 inst_4098 ( .ZN(net_4067), .A2(net_2464), .A1(x6157) );
CLKBUF_X2 inst_12178 ( .A(net_12096), .Z(net_12097) );
CLKBUF_X2 inst_11220 ( .A(net_11138), .Z(net_11139) );
INV_X4 inst_5703 ( .ZN(net_1367), .A(net_778) );
DFF_X2 inst_7761 ( .Q(net_9711), .D(net_6547), .CK(net_12056) );
CLKBUF_X2 inst_11177 ( .A(net_11002), .Z(net_11096) );
NOR2_X2 inst_2978 ( .A1(net_10220), .ZN(net_1160), .A2(net_1021) );
XNOR2_X2 inst_413 ( .B(net_7499), .ZN(net_1416), .A(net_1415) );
CLKBUF_X2 inst_14817 ( .A(net_14735), .Z(net_14736) );
CLKBUF_X2 inst_14239 ( .A(net_14157), .Z(net_14158) );
CLKBUF_X2 inst_11033 ( .A(net_10738), .Z(net_10952) );
INV_X4 inst_5094 ( .A(net_2598), .ZN(net_1737) );
CLKBUF_X2 inst_11393 ( .A(net_11273), .Z(net_11312) );
OR2_X2 inst_859 ( .A1(net_9544), .ZN(net_7991), .A2(net_7990) );
INV_X4 inst_6623 ( .A(net_8960), .ZN(net_8957) );
DFF_X2 inst_8118 ( .Q(net_9726), .D(net_5152), .CK(net_15121) );
AOI211_X2 inst_10269 ( .A(net_7704), .ZN(net_7614), .C2(net_7518), .C1(net_5005), .B(x3390) );
CLKBUF_X2 inst_13446 ( .A(net_11333), .Z(net_13365) );
CLKBUF_X2 inst_14352 ( .A(net_14270), .Z(net_14271) );
CLKBUF_X2 inst_12634 ( .A(net_12552), .Z(net_12553) );
NAND2_X4 inst_3323 ( .ZN(net_8900), .A1(net_8883), .A2(net_8581) );
CLKBUF_X2 inst_13013 ( .A(net_12931), .Z(net_12932) );
OAI21_X2 inst_2019 ( .ZN(net_8859), .A(net_2427), .B2(net_1770), .B1(net_1686) );
CLKBUF_X2 inst_13679 ( .A(net_12288), .Z(net_13598) );
DFF_X2 inst_8323 ( .QN(net_10481), .D(net_3646), .CK(net_11437) );
INV_X4 inst_5186 ( .ZN(net_2821), .A(net_1554) );
INV_X4 inst_5938 ( .ZN(net_1334), .A(net_581) );
CLKBUF_X2 inst_13061 ( .A(net_12330), .Z(net_12980) );
CLKBUF_X2 inst_15061 ( .A(net_14979), .Z(net_14980) );
XNOR2_X2 inst_69 ( .ZN(net_8710), .A(net_8689), .B(net_8262) );
INV_X4 inst_5736 ( .ZN(net_1383), .A(net_747) );
CLKBUF_X2 inst_15542 ( .A(net_15460), .Z(net_15461) );
CLKBUF_X2 inst_14448 ( .A(net_14366), .Z(net_14367) );
CLKBUF_X2 inst_15626 ( .A(net_12246), .Z(net_15545) );
OAI221_X2 inst_1691 ( .C1(net_7229), .B2(net_5642), .A(net_5637), .ZN(net_5468), .B1(net_5467), .C2(net_4905) );
NOR2_X2 inst_2669 ( .ZN(net_4980), .A2(net_4704), .A1(net_4484) );
CLKBUF_X2 inst_15396 ( .A(net_15314), .Z(net_15315) );
AOI22_X2 inst_9019 ( .A1(net_8002), .B2(net_8001), .ZN(net_8000), .A2(net_7946), .B1(net_2139) );
CLKBUF_X2 inst_12844 ( .A(net_11103), .Z(net_12763) );
CLKBUF_X2 inst_11156 ( .A(net_11074), .Z(net_11075) );
OR2_X4 inst_844 ( .A2(net_10464), .A1(net_10463), .ZN(net_1172) );
NOR2_X2 inst_2489 ( .ZN(net_8716), .A1(net_8714), .A2(net_8713) );
CLKBUF_X2 inst_14712 ( .A(net_13294), .Z(net_14631) );
INV_X2 inst_6968 ( .A(net_4573), .ZN(net_1807) );
CLKBUF_X2 inst_15413 ( .A(net_15331), .Z(net_15332) );
NAND2_X2 inst_3619 ( .ZN(net_7111), .A1(net_6872), .A2(net_6686) );
NAND2_X2 inst_3688 ( .A2(net_9263), .A1(net_8965), .ZN(net_7379) );
INV_X2 inst_6709 ( .A(net_8181), .ZN(net_8128) );
INV_X4 inst_5805 ( .A(net_1028), .ZN(net_865) );
DFF_X2 inst_7716 ( .Q(net_9806), .D(net_6425), .CK(net_12576) );
INV_X2 inst_6939 ( .A(net_3670), .ZN(net_1918) );
INV_X4 inst_4641 ( .ZN(net_6037), .A(net_5868) );
INV_X2 inst_7056 ( .A(net_6658), .ZN(net_1304) );
CLKBUF_X2 inst_11038 ( .A(net_10956), .Z(net_10957) );
INV_X4 inst_5476 ( .ZN(net_1196), .A(net_1005) );
SDFF_X2 inst_460 ( .D(net_8712), .SE(net_758), .Q(net_241), .SI(net_110), .CK(net_13856) );
CLKBUF_X2 inst_10877 ( .A(net_10795), .Z(net_10796) );
OAI221_X2 inst_1455 ( .C1(net_9071), .ZN(net_7976), .A(net_7975), .B2(net_7974), .C2(net_7973), .B1(net_2586) );
INV_X4 inst_5776 ( .ZN(net_794), .A(net_711) );
INV_X2 inst_7135 ( .A(net_9243), .ZN(net_834) );
CLKBUF_X2 inst_12149 ( .A(net_12067), .Z(net_12068) );
NOR2_X2 inst_2497 ( .ZN(net_8568), .A1(net_8541), .A2(net_8509) );
CLKBUF_X2 inst_13124 ( .A(net_11696), .Z(net_13043) );
AOI21_X2 inst_10186 ( .ZN(net_3420), .A(net_3419), .B1(net_3102), .B2(net_3101) );
NAND2_X2 inst_3660 ( .A1(net_8511), .ZN(net_6431), .A2(net_6430) );
CLKBUF_X2 inst_11167 ( .A(net_11017), .Z(net_11086) );
SDFF_X2 inst_560 ( .D(net_9138), .SE(net_933), .CK(net_10980), .SI(x2098), .Q(x1192) );
CLKBUF_X2 inst_15678 ( .A(net_15596), .Z(net_15597) );
INV_X4 inst_5393 ( .A(net_2101), .ZN(net_1180) );
AOI222_X1 inst_9729 ( .ZN(net_3205), .A1(net_3204), .B2(net_3203), .A2(net_3203), .C2(net_3202), .C1(net_2538), .B1(net_656) );
NAND2_X2 inst_4230 ( .A2(net_10330), .A1(net_4166), .ZN(net_1621) );
INV_X4 inst_5199 ( .A(net_2935), .ZN(net_2692) );
CLKBUF_X2 inst_15316 ( .A(net_14670), .Z(net_15235) );
CLKBUF_X2 inst_12953 ( .A(net_12871), .Z(net_12872) );
DFF_X2 inst_7479 ( .D(net_8069), .Q(net_212), .CK(net_12902) );
INV_X4 inst_4809 ( .ZN(net_3563), .A(net_3401) );
INV_X4 inst_5571 ( .ZN(net_4986), .A(net_909) );
CLKBUF_X2 inst_13455 ( .A(net_13373), .Z(net_13374) );
OAI21_X2 inst_1802 ( .B2(net_10137), .A(net_10136), .ZN(net_7332), .B1(net_7331) );
OAI33_X1 inst_950 ( .B1(net_7557), .ZN(net_7508), .A1(net_7506), .A3(net_7505), .B3(net_7503), .A2(net_1574), .B2(net_910) );
AOI211_X2 inst_10260 ( .ZN(net_7936), .A(net_7837), .B(net_7561), .C1(net_6158), .C2(net_5885) );
INV_X2 inst_6851 ( .ZN(net_3387), .A(net_3386) );
CLKBUF_X2 inst_15444 ( .A(net_15362), .Z(net_15363) );
NOR2_X2 inst_2982 ( .A1(net_10358), .ZN(net_1720), .A2(net_321) );
NAND2_X2 inst_3955 ( .A1(net_10368), .ZN(net_3705), .A2(net_3419) );
CLKBUF_X2 inst_11837 ( .A(net_11755), .Z(net_11756) );
AOI21_X2 inst_10100 ( .B2(net_8117), .ZN(net_5994), .B1(net_1150), .A(net_593) );
OAI22_X2 inst_1218 ( .A1(net_7129), .A2(net_5134), .B2(net_5133), .ZN(net_5030), .B1(net_1889) );
NAND2_X4 inst_3359 ( .A2(net_9002), .A1(net_9001), .ZN(net_8106) );
DFF_X1 inst_8458 ( .Q(net_9571), .D(net_7983), .CK(net_11545) );
INV_X4 inst_6414 ( .A(net_10388), .ZN(net_385) );
DFF_X2 inst_7491 ( .Q(net_10509), .D(net_8013), .CK(net_12992) );
CLKBUF_X2 inst_14338 ( .A(net_13407), .Z(net_14257) );
NAND2_X2 inst_4418 ( .A2(net_9517), .A1(net_9516), .ZN(net_959) );
AOI22_X2 inst_9541 ( .B1(net_9923), .A1(net_9693), .A2(net_5966), .B2(net_4969), .ZN(net_3780) );
XNOR2_X2 inst_96 ( .B(net_9435), .ZN(net_8451), .A(net_7170) );
XNOR2_X2 inst_101 ( .ZN(net_8402), .A(net_8172), .B(net_7058) );
NAND2_X2 inst_4346 ( .A2(net_10115), .ZN(net_1852), .A1(net_793) );
DFF_X1 inst_8564 ( .Q(net_9772), .D(net_7235), .CK(net_15573) );
CLKBUF_X2 inst_14033 ( .A(net_12050), .Z(net_13952) );
NAND2_X2 inst_3555 ( .ZN(net_8626), .A2(net_7790), .A1(net_7638) );
CLKBUF_X2 inst_11205 ( .A(net_11123), .Z(net_11124) );
AOI21_X2 inst_10234 ( .ZN(net_2504), .B1(net_2002), .B2(net_1765), .A(net_1359) );
CLKBUF_X2 inst_14377 ( .A(net_14295), .Z(net_14296) );
AOI22_X2 inst_9330 ( .B1(net_10014), .A1(net_6823), .A2(net_5743), .B2(net_5742), .ZN(net_5622) );
CLKBUF_X2 inst_11388 ( .A(net_11306), .Z(net_11307) );
INV_X4 inst_4722 ( .ZN(net_4616), .A(net_4497) );
SDFF_X2 inst_510 ( .Q(net_9334), .D(net_9334), .SI(net_9159), .SE(net_7588), .CK(net_13105) );
CLKBUF_X2 inst_10912 ( .A(net_10830), .Z(net_10831) );
CLKBUF_X2 inst_15558 ( .A(net_15476), .Z(net_15477) );
CLKBUF_X2 inst_12194 ( .A(net_12112), .Z(net_12113) );
CLKBUF_X2 inst_14575 ( .A(net_12640), .Z(net_14494) );
NOR3_X2 inst_2436 ( .A2(net_5075), .ZN(net_3346), .A1(net_2944), .A3(net_1183) );
INV_X4 inst_6505 ( .ZN(net_1847), .A(net_155) );
OAI221_X2 inst_1677 ( .B1(net_7213), .C2(net_5642), .ZN(net_5490), .B2(net_4905), .A(net_3731), .C1(net_1589) );
NOR2_X2 inst_2832 ( .A1(net_4723), .A2(net_2751), .ZN(net_2439) );
OR2_X4 inst_830 ( .A2(net_9289), .ZN(net_8803), .A1(net_957) );
SDFF_X2 inst_603 ( .Q(net_10516), .D(net_10516), .SE(net_4560), .CK(net_10558), .SI(x6102) );
DFF_X1 inst_8433 ( .D(net_8638), .Q(net_279), .CK(net_14947) );
CLKBUF_X2 inst_15646 ( .A(net_13532), .Z(net_15565) );
XNOR2_X2 inst_291 ( .B(net_4273), .ZN(net_3519), .A(net_3041) );
NOR2_X2 inst_2878 ( .A2(net_10538), .ZN(net_2464), .A1(x3867) );
NOR2_X2 inst_2494 ( .A1(net_8714), .ZN(net_8599), .A2(net_8598) );
OR2_X4 inst_776 ( .ZN(net_4274), .A2(net_2971), .A1(net_2956) );
AOI22_X2 inst_9488 ( .A1(net_10176), .B1(net_9817), .A2(net_4217), .ZN(net_3835), .B2(net_2556) );
NOR2_X2 inst_2526 ( .A2(net_9114), .ZN(net_8166), .A1(net_392) );
CLKBUF_X2 inst_15521 ( .A(net_15439), .Z(net_15440) );
INV_X4 inst_5047 ( .ZN(net_8206), .A(net_1902) );
CLKBUF_X2 inst_12213 ( .A(net_12131), .Z(net_12132) );
CLKBUF_X2 inst_10787 ( .A(net_10705), .Z(net_10706) );
INV_X4 inst_5313 ( .ZN(net_5486), .A(net_1285) );
OAI21_X2 inst_1972 ( .ZN(net_3157), .B2(net_2958), .B1(net_2957), .A(net_2940) );
SDFF_X2 inst_558 ( .D(net_9119), .SE(net_933), .CK(net_10562), .SI(x3249), .Q(x1402) );
INV_X4 inst_6167 ( .A(net_9740), .ZN(net_596) );
CLKBUF_X2 inst_12704 ( .A(net_12622), .Z(net_12623) );
AOI211_X2 inst_10310 ( .B(net_5954), .A(net_2984), .ZN(net_2796), .C1(net_2712), .C2(net_2067) );
INV_X2 inst_6849 ( .A(net_10164), .ZN(net_3458) );
AOI22_X2 inst_9110 ( .A1(net_9691), .A2(net_6404), .ZN(net_6380), .B1(net_6379), .B2(net_5263) );
AND2_X2 inst_10591 ( .A2(net_4266), .A1(net_2427), .ZN(net_2384) );
XNOR2_X2 inst_389 ( .ZN(net_2270), .B(net_1467), .A(net_626) );
INV_X4 inst_5179 ( .A(net_1962), .ZN(net_1848) );
INV_X4 inst_6512 ( .ZN(net_6039), .A(net_275) );
CLKBUF_X2 inst_14301 ( .A(net_14219), .Z(net_14220) );
CLKBUF_X2 inst_13460 ( .A(net_13378), .Z(net_13379) );
NOR2_X2 inst_2712 ( .A2(net_5341), .ZN(net_4733), .A1(net_4170) );
AOI211_X2 inst_10252 ( .ZN(net_8191), .A(net_8190), .C2(net_7982), .C1(net_3978), .B(net_3298) );
INV_X4 inst_6152 ( .A(net_10037), .ZN(net_691) );
INV_X2 inst_6925 ( .ZN(net_1968), .A(net_1967) );
DFF_X1 inst_8650 ( .Q(net_8837), .D(net_7301), .CK(net_11776) );
DFF_X2 inst_7745 ( .QN(net_10140), .D(net_6318), .CK(net_14546) );
OAI222_X2 inst_1382 ( .B2(net_7660), .A2(net_7659), .C2(net_7658), .ZN(net_6003), .B1(net_5208), .A1(net_4201), .C1(net_1890) );
DFF_X1 inst_8841 ( .QN(net_10057), .D(net_2137), .CK(net_10739) );
DFF_X1 inst_8600 ( .Q(net_9689), .D(net_7258), .CK(net_15246) );
OAI21_X2 inst_1807 ( .ZN(net_7392), .B2(net_7060), .A(net_5342), .B1(net_5341) );
NOR2_X2 inst_2795 ( .ZN(net_4333), .A1(net_2928), .A2(net_2927) );
INV_X2 inst_7236 ( .A(net_10349), .ZN(net_857) );
AOI221_X2 inst_9989 ( .B1(net_4166), .ZN(net_3557), .C2(net_3129), .A(net_3124), .C1(net_2411), .B2(net_845) );
CLKBUF_X2 inst_12274 ( .A(net_12192), .Z(net_12193) );
OR2_X2 inst_913 ( .A1(net_9044), .A2(net_8566), .ZN(net_8441) );
INV_X4 inst_5266 ( .ZN(net_2869), .A(net_2600) );
CLKBUF_X2 inst_12712 ( .A(net_11477), .Z(net_12631) );
INV_X4 inst_4766 ( .ZN(net_4472), .A(net_4363) );
MUX2_X1 inst_4445 ( .S(net_6041), .A(net_301), .B(x4781), .Z(x106) );
INV_X4 inst_5895 ( .ZN(net_967), .A(net_606) );
CLKBUF_X2 inst_11785 ( .A(net_11703), .Z(net_11704) );
AOI221_X2 inst_9977 ( .C1(net_9800), .B2(net_5174), .ZN(net_4381), .B1(net_4380), .A(net_3943), .C2(net_2556) );
CLKBUF_X2 inst_12866 ( .A(net_12784), .Z(net_12785) );
CLKBUF_X2 inst_12766 ( .A(net_12684), .Z(net_12685) );
DFF_X2 inst_8365 ( .Q(net_9163), .D(net_1968), .CK(net_14056) );
CLKBUF_X2 inst_14195 ( .A(net_14113), .Z(net_14114) );
INV_X2 inst_7105 ( .ZN(net_1024), .A(net_1023) );
CLKBUF_X2 inst_15502 ( .A(net_15420), .Z(net_15421) );
CLKBUF_X2 inst_15188 ( .A(net_15106), .Z(net_15107) );
CLKBUF_X2 inst_10843 ( .A(net_10761), .Z(net_10762) );
CLKBUF_X2 inst_11613 ( .A(net_11531), .Z(net_11532) );
DFF_X2 inst_7687 ( .QN(net_9203), .D(net_6555), .CK(net_11333) );
INV_X4 inst_6633 ( .A(net_9039), .ZN(net_9038) );
CLKBUF_X2 inst_12004 ( .A(net_11922), .Z(net_11923) );
CLKBUF_X2 inst_11133 ( .A(net_11051), .Z(net_11052) );
AND4_X4 inst_10322 ( .ZN(net_4486), .A4(net_4057), .A1(net_3813), .A2(net_3737), .A3(net_3430) );
CLKBUF_X2 inst_11724 ( .A(net_11642), .Z(net_11643) );
CLKBUF_X2 inst_11214 ( .A(net_11132), .Z(net_11133) );
AOI22_X2 inst_9298 ( .B1(net_10001), .A1(net_5743), .B2(net_5742), .ZN(net_5687), .A2(net_241) );
NOR2_X2 inst_2483 ( .A2(net_9309), .ZN(net_8802), .A1(net_8801) );
CLKBUF_X2 inst_13321 ( .A(net_13239), .Z(net_13240) );
AOI22_X2 inst_9446 ( .A1(net_10526), .B1(net_9799), .A2(net_4056), .ZN(net_4053), .B2(net_2556) );
OAI222_X2 inst_1414 ( .A2(net_7665), .C2(net_7664), .B2(net_7663), .ZN(net_5196), .A1(net_3006), .C1(net_2138), .B1(net_860) );
DFF_X2 inst_7624 ( .QN(net_10462), .D(net_6922), .CK(net_13664) );
DFF_X1 inst_8451 ( .Q(net_9526), .D(net_8078), .CK(net_15042) );
XNOR2_X1 inst_449 ( .ZN(net_8671), .A(net_8662), .B(net_2446) );
NAND2_X2 inst_3994 ( .A1(net_4723), .A2(net_3390), .ZN(net_3375) );
CLKBUF_X2 inst_13467 ( .A(net_13385), .Z(net_13386) );
NAND2_X2 inst_4212 ( .ZN(net_1744), .A1(net_1743), .A2(net_1389) );
CLKBUF_X2 inst_10797 ( .A(net_10715), .Z(net_10716) );
AND3_X4 inst_10354 ( .ZN(net_5285), .A1(net_5284), .A2(net_5283), .A3(net_4600) );
NOR2_X2 inst_2790 ( .A1(net_3917), .A2(net_3065), .ZN(net_3064) );
OAI211_X2 inst_2138 ( .C2(net_6778), .ZN(net_6710), .A(net_6422), .B(net_6146), .C1(net_5106) );
INV_X4 inst_5599 ( .ZN(net_1154), .A(net_882) );
INV_X2 inst_7152 ( .A(net_809), .ZN(net_718) );
CLKBUF_X2 inst_11417 ( .A(net_11335), .Z(net_11336) );
INV_X4 inst_6593 ( .A(net_10333), .ZN(net_321) );
INV_X4 inst_6055 ( .ZN(net_4015), .A(net_132) );
CLKBUF_X2 inst_13362 ( .A(net_13280), .Z(net_13281) );
CLKBUF_X2 inst_15257 ( .A(net_14747), .Z(net_15176) );
CLKBUF_X2 inst_15716 ( .A(net_15634), .Z(net_15635) );
CLKBUF_X2 inst_11231 ( .A(net_10987), .Z(net_11150) );
NAND3_X2 inst_3249 ( .ZN(net_4585), .A1(net_4584), .A3(net_4583), .A2(net_2207) );
INV_X4 inst_4935 ( .A(net_4717), .ZN(net_2589) );
CLKBUF_X2 inst_12912 ( .A(net_11427), .Z(net_12831) );
CLKBUF_X2 inst_11759 ( .A(net_11677), .Z(net_11678) );
AOI22_X2 inst_9594 ( .A1(net_10044), .B1(net_9815), .A2(net_5174), .ZN(net_3505), .B2(net_2556) );
DFF_X2 inst_7498 ( .D(net_8015), .QN(net_201), .CK(net_12899) );
NOR4_X2 inst_2309 ( .A4(net_9611), .ZN(net_7594), .A2(net_7519), .A1(net_6187), .A3(net_2506) );
AOI221_X2 inst_9860 ( .A(net_6889), .B2(net_6888), .C2(net_6887), .ZN(net_6858), .B1(net_1193), .C1(x4781) );
CLKBUF_X2 inst_13369 ( .A(net_11267), .Z(net_13288) );
CLKBUF_X2 inst_12420 ( .A(net_11459), .Z(net_12339) );
CLKBUF_X2 inst_15011 ( .A(net_10811), .Z(net_14930) );
CLKBUF_X2 inst_11044 ( .A(net_10619), .Z(net_10963) );
CLKBUF_X2 inst_12973 ( .A(net_12891), .Z(net_12892) );
DFF_X2 inst_7644 ( .D(net_6725), .QN(net_160), .CK(net_15722) );
INV_X2 inst_7196 ( .A(net_9551), .ZN(net_8177) );
DFF_X2 inst_8201 ( .QN(net_9833), .D(net_5057), .CK(net_11727) );
CLKBUF_X2 inst_11283 ( .A(net_11201), .Z(net_11202) );
NOR2_X2 inst_2603 ( .ZN(net_6552), .A1(net_5764), .A2(net_3028) );
NAND2_X2 inst_3614 ( .A2(net_10452), .ZN(net_7119), .A1(net_571) );
CLKBUF_X2 inst_15792 ( .A(net_13701), .Z(net_15711) );
CLKBUF_X2 inst_11335 ( .A(net_11253), .Z(net_11254) );
INV_X4 inst_4603 ( .ZN(net_7748), .A(net_7690) );
AOI22_X2 inst_9339 ( .B1(net_9815), .A2(net_5766), .B2(net_5765), .ZN(net_5613), .A1(net_253) );
OAI211_X2 inst_2153 ( .C2(net_6778), .ZN(net_6695), .A(net_6323), .B(net_6062), .C1(net_5075) );
CLKBUF_X2 inst_12776 ( .A(net_11984), .Z(net_12695) );
CLKBUF_X2 inst_10752 ( .A(net_10670), .Z(net_10671) );
SDFF_X2 inst_588 ( .Q(net_9251), .SE(net_4589), .D(net_134), .SI(net_100), .CK(net_13832) );
AND2_X4 inst_10394 ( .A2(net_7572), .A1(net_7379), .ZN(net_6900) );
CLKBUF_X2 inst_11411 ( .A(net_11329), .Z(net_11330) );
CLKBUF_X2 inst_11271 ( .A(net_11189), .Z(net_11190) );
CLKBUF_X2 inst_11904 ( .A(net_11822), .Z(net_11823) );
CLKBUF_X2 inst_11798 ( .A(net_11716), .Z(net_11717) );
CLKBUF_X2 inst_14015 ( .A(net_13933), .Z(net_13934) );
AND4_X4 inst_10329 ( .ZN(net_3318), .A4(net_2961), .A3(net_2272), .A1(net_994), .A2(net_860) );
AOI22_X2 inst_9405 ( .A2(net_9095), .B2(net_9068), .ZN(net_4999), .A1(net_3380), .B1(net_708) );
INV_X4 inst_5494 ( .ZN(net_1292), .A(net_1249) );
CLKBUF_X2 inst_11060 ( .A(net_10978), .Z(net_10979) );
AND2_X2 inst_10586 ( .ZN(net_3182), .A2(net_2464), .A1(net_725) );
INV_X4 inst_4752 ( .ZN(net_5591), .A(net_4516) );
DFF_X2 inst_7674 ( .D(net_6699), .QN(net_176), .CK(net_12737) );
CLKBUF_X2 inst_12913 ( .A(net_12831), .Z(net_12832) );
OAI222_X2 inst_1356 ( .B1(net_7728), .A2(net_7727), .C2(net_7726), .ZN(net_6953), .B2(net_5981), .A1(net_4432), .C1(net_2715) );
INV_X4 inst_5441 ( .ZN(net_2306), .A(net_1102) );
AOI221_X2 inst_9906 ( .B1(net_9890), .B2(net_9101), .A(net_6945), .C2(net_6944), .C1(net_6811), .ZN(net_6788) );
NOR2_X2 inst_2628 ( .A2(net_9258), .A1(net_8116), .ZN(net_6228) );
INV_X4 inst_6447 ( .A(net_9291), .ZN(net_377) );
INV_X2 inst_6874 ( .ZN(net_2992), .A(net_2991) );
OAI211_X2 inst_2196 ( .C1(net_7224), .C2(net_6542), .ZN(net_6511), .B(net_5609), .A(net_3679) );
NAND2_X2 inst_3485 ( .A2(net_8968), .ZN(net_8393), .A1(net_8251) );
CLKBUF_X2 inst_14159 ( .A(net_14077), .Z(net_14078) );
INV_X4 inst_5854 ( .ZN(net_843), .A(net_643) );
INV_X2 inst_7145 ( .ZN(net_1075), .A(net_796) );
DFF_X2 inst_7754 ( .Q(net_10510), .D(net_6454), .CK(net_12981) );
CLKBUF_X2 inst_14083 ( .A(net_14001), .Z(net_14002) );
OAI22_X2 inst_1045 ( .A1(net_9364), .B2(net_7638), .A2(net_7635), .ZN(net_7633), .B1(net_7632) );
OR2_X2 inst_865 ( .ZN(net_7709), .A2(net_7694), .A1(net_7615) );
XNOR2_X2 inst_252 ( .ZN(net_4116), .A(net_3961), .B(net_2658) );
OAI33_X1 inst_956 ( .A2(net_9270), .A3(net_9269), .ZN(net_6583), .B2(net_6582), .B3(net_6581), .B1(net_5376), .A1(net_2669) );
DFF_X1 inst_8587 ( .Q(net_9866), .D(net_7121), .CK(net_14264) );
CLKBUF_X2 inst_10959 ( .A(net_10877), .Z(net_10878) );
DFF_X1 inst_8680 ( .D(net_6740), .Q(net_147), .CK(net_12596) );
AOI21_X2 inst_10177 ( .A(net_3741), .ZN(net_3608), .B2(net_2962), .B1(net_860) );
INV_X4 inst_4684 ( .ZN(net_4994), .A(net_4993) );
CLKBUF_X2 inst_12757 ( .A(net_12675), .Z(net_12676) );
SDFF_X2 inst_484 ( .SE(net_9540), .SI(net_8225), .Q(net_300), .D(net_300), .CK(net_13912) );
AOI22_X2 inst_9272 ( .B1(net_9700), .ZN(net_5757), .A1(net_5755), .B2(net_5754), .A2(net_237) );
MUX2_X1 inst_4474 ( .S(net_6041), .A(net_4273), .B(x6351), .Z(x389) );
INV_X2 inst_6678 ( .ZN(net_8350), .A(net_8287) );
AOI22_X2 inst_9129 ( .A1(net_9695), .A2(net_6418), .ZN(net_6359), .B2(net_5263), .B1(net_135) );
XOR2_X2 inst_32 ( .A(net_7856), .Z(net_1992), .B(net_623) );
OAI21_X2 inst_1821 ( .ZN(net_6630), .A(net_6629), .B1(net_6628), .B2(net_5970) );
AOI22_X2 inst_9616 ( .A1(net_10089), .B1(net_10015), .A2(net_5319), .ZN(net_3437), .B2(net_2468) );
CLKBUF_X2 inst_12798 ( .A(net_12716), .Z(net_12717) );
INV_X2 inst_7011 ( .ZN(net_7910), .A(net_1314) );
INV_X2 inst_7271 ( .A(net_8938), .ZN(net_8936) );
CLKBUF_X2 inst_10683 ( .A(net_10601), .Z(net_10602) );
SDFF_X2 inst_616 ( .Q(net_9462), .D(net_9462), .SE(net_3293), .CK(net_11904), .SI(x1792) );
INV_X2 inst_7201 ( .A(net_9380), .ZN(net_957) );
INV_X4 inst_5381 ( .ZN(net_1597), .A(net_1196) );
CLKBUF_X2 inst_11049 ( .A(net_10967), .Z(net_10968) );
AOI22_X2 inst_9649 ( .ZN(net_2696), .A1(net_2415), .A2(net_2381), .B2(net_1516), .B1(net_1365) );
AOI22_X2 inst_9320 ( .B1(net_9724), .A1(net_6811), .A2(net_5755), .B2(net_5754), .ZN(net_5656) );
SDFF_X2 inst_620 ( .Q(net_9467), .D(net_9467), .SE(net_3293), .CK(net_11373), .SI(x1503) );
OAI21_X2 inst_1784 ( .B1(net_9544), .ZN(net_7621), .A(net_7620), .B2(net_7488) );
INV_X4 inst_6496 ( .ZN(net_7245), .A(x6102) );
NAND4_X2 inst_3118 ( .ZN(net_4035), .A4(net_3343), .A1(net_3296), .A2(net_2872), .A3(net_1734) );
INV_X4 inst_6401 ( .A(net_9534), .ZN(net_7344) );
DFF_X2 inst_8040 ( .QN(net_9546), .D(net_9252), .CK(net_13868) );
INV_X2 inst_6869 ( .ZN(net_3053), .A(net_3052) );
CLKBUF_X2 inst_14921 ( .A(net_10993), .Z(net_14840) );
OAI211_X2 inst_2071 ( .ZN(net_6779), .C2(net_6778), .A(net_6337), .B(net_6073), .C1(net_5092) );
CLKBUF_X2 inst_14597 ( .A(net_14515), .Z(net_14516) );
CLKBUF_X2 inst_14514 ( .A(net_12955), .Z(net_14433) );
OAI222_X2 inst_1427 ( .B2(net_8858), .A2(net_8858), .ZN(net_3398), .C2(net_3397), .C1(net_2340), .B1(net_1585), .A1(net_1135) );
AND2_X4 inst_10421 ( .ZN(net_4398), .A2(net_4258), .A1(net_4109) );
OAI222_X2 inst_1409 ( .B2(net_7728), .A2(net_7727), .C2(net_7726), .ZN(net_5310), .B1(net_4262), .A1(net_3278), .C1(net_1192) );
CLKBUF_X2 inst_10757 ( .A(net_10675), .Z(net_10676) );
CLKBUF_X2 inst_11570 ( .A(net_11488), .Z(net_11489) );
AOI22_X2 inst_9183 ( .A1(net_9873), .B1(net_9774), .A2(net_8042), .B2(net_6140), .ZN(net_6132) );
CLKBUF_X2 inst_13752 ( .A(net_13670), .Z(net_13671) );
AOI21_X2 inst_10056 ( .A(net_7114), .ZN(net_7113), .B2(net_6948), .B1(net_3699) );
INV_X2 inst_7259 ( .A(net_10029), .ZN(net_325) );
CLKBUF_X2 inst_15613 ( .A(net_15531), .Z(net_15532) );
CLKBUF_X2 inst_14296 ( .A(net_14214), .Z(net_14215) );
INV_X4 inst_4662 ( .ZN(net_5710), .A(net_5709) );
XNOR2_X2 inst_87 ( .A(net_8937), .ZN(net_8611), .B(net_2154) );
CLKBUF_X2 inst_13509 ( .A(net_13427), .Z(net_13428) );
NOR2_X2 inst_2996 ( .ZN(net_1376), .A2(net_901), .A1(net_823) );
INV_X4 inst_5037 ( .ZN(net_3916), .A(net_3085) );
AND2_X2 inst_10601 ( .A2(net_4110), .ZN(net_2065), .A1(net_2064) );
NOR2_X2 inst_2918 ( .A2(net_4183), .ZN(net_3615), .A1(net_1396) );
AOI21_X2 inst_10036 ( .ZN(net_7772), .B2(net_7766), .A(net_7377), .B1(net_7275) );
CLKBUF_X2 inst_11946 ( .A(net_10978), .Z(net_11865) );
NOR2_X2 inst_2721 ( .A2(net_4512), .ZN(net_4320), .A1(net_4016) );
AOI22_X2 inst_9576 ( .B1(net_9985), .A2(net_5173), .ZN(net_3680), .B2(net_2541), .A1(net_219) );
AOI22_X2 inst_9517 ( .B1(net_9766), .A1(net_9667), .A2(net_5966), .ZN(net_3805), .B2(net_2462) );
OR2_X4 inst_800 ( .A1(net_10368), .ZN(net_2415), .A2(net_1956) );
NAND4_X2 inst_3074 ( .ZN(net_5170), .A1(net_5168), .A2(net_5167), .A4(net_5166), .A3(net_644) );
INV_X4 inst_5281 ( .ZN(net_2131), .A(net_1448) );
AOI221_X2 inst_9925 ( .B2(net_5867), .A(net_5862), .ZN(net_5855), .C1(net_5854), .C2(net_5853), .B1(x5225) );
XOR2_X2 inst_10 ( .Z(net_3702), .A(net_3265), .B(net_1126) );
CLKBUF_X2 inst_14002 ( .A(net_13920), .Z(net_13921) );
DFF_X1 inst_8763 ( .Q(net_9131), .D(net_5294), .CK(net_10578) );
XOR2_X2 inst_4 ( .Z(net_6503), .A(net_5589), .B(net_1234) );
NAND2_X2 inst_3795 ( .A2(net_9082), .ZN(net_4726), .A1(net_4687) );
DFF_X2 inst_7770 ( .Q(net_9721), .D(net_6533), .CK(net_13425) );
CLKBUF_X2 inst_15550 ( .A(net_13023), .Z(net_15469) );
NAND2_X2 inst_4337 ( .A1(net_9061), .A2(net_8955), .ZN(net_1689) );
AND2_X4 inst_10475 ( .A2(net_10153), .A1(net_10152), .ZN(net_2010) );
DFF_X2 inst_7981 ( .QN(net_10424), .D(net_5596), .CK(net_14902) );
NAND3_X2 inst_3272 ( .A3(net_10348), .ZN(net_4144), .A1(net_4143), .A2(net_857) );
CLKBUF_X2 inst_13555 ( .A(net_13473), .Z(net_13474) );
CLKBUF_X2 inst_13186 ( .A(net_13104), .Z(net_13105) );
AOI221_X2 inst_9846 ( .A(net_6889), .B2(net_6888), .C2(net_6887), .ZN(net_6872), .B1(net_5831), .C1(x5722) );
AOI22_X2 inst_9455 ( .A2(net_10479), .B2(net_8840), .ZN(net_3937), .A1(net_3429), .B1(net_3409) );
INV_X4 inst_5459 ( .ZN(net_1462), .A(net_647) );
AND2_X2 inst_10494 ( .ZN(net_6895), .A2(net_6894), .A1(net_6651) );
CLKBUF_X2 inst_14232 ( .A(net_12759), .Z(net_14151) );
AOI221_X2 inst_9867 ( .B1(net_9873), .B2(net_9101), .A(net_6945), .C1(net_6944), .ZN(net_6843), .C2(net_244) );
AOI21_X2 inst_10090 ( .B1(net_10385), .A(net_6677), .ZN(net_5777), .B2(net_5200) );
OAI21_X2 inst_1866 ( .ZN(net_5912), .A(net_5348), .B1(net_5347), .B2(net_5346) );
CLKBUF_X2 inst_15230 ( .A(net_15148), .Z(net_15149) );
DFF_X1 inst_8795 ( .Q(net_10342), .D(net_4285), .CK(net_10669) );
CLKBUF_X2 inst_11961 ( .A(net_10955), .Z(net_11880) );
OAI21_X2 inst_1878 ( .B2(net_10448), .ZN(net_5247), .A(net_2710), .B1(net_884) );
INV_X4 inst_5136 ( .ZN(net_2906), .A(net_1384) );
INV_X4 inst_6016 ( .A(net_10019), .ZN(net_524) );
INV_X2 inst_6700 ( .A(net_8249), .ZN(net_8167) );
CLKBUF_X2 inst_14462 ( .A(net_14380), .Z(net_14381) );
AOI211_X2 inst_10290 ( .ZN(net_4670), .C2(net_4250), .C1(net_3557), .A(net_3215), .B(net_2421) );
INV_X4 inst_4731 ( .ZN(net_4982), .A(net_4297) );
OAI22_X2 inst_1276 ( .B2(net_7671), .A1(net_7602), .ZN(net_4463), .A2(net_3883), .B1(net_3375) );
OR2_X4 inst_765 ( .ZN(net_4622), .A1(net_4323), .A2(net_4220) );
XNOR2_X2 inst_256 ( .ZN(net_4104), .A(net_3470), .B(net_2331) );
INV_X4 inst_6205 ( .A(net_9825), .ZN(net_2193) );
CLKBUF_X2 inst_10790 ( .A(net_10708), .Z(net_10709) );
AOI221_X2 inst_9870 ( .B1(net_9778), .B2(net_9098), .A(net_6940), .C2(net_6939), .ZN(net_6832), .C1(net_248) );
CLKBUF_X2 inst_10664 ( .A(net_10582), .Z(net_10583) );
AOI22_X2 inst_9180 ( .A1(net_9910), .B1(net_9811), .A2(net_6141), .ZN(net_6136), .B2(net_6129) );
OAI21_X2 inst_1902 ( .B1(net_7203), .B2(net_4862), .ZN(net_4850), .A(net_4522) );
DFF_X1 inst_8626 ( .Q(net_9784), .D(net_7200), .CK(net_13364) );
CLKBUF_X2 inst_14247 ( .A(net_14165), .Z(net_14166) );
AOI22_X2 inst_9635 ( .B1(net_9807), .A1(net_9775), .ZN(net_3407), .B2(net_2556), .A2(net_2462) );
INV_X4 inst_5052 ( .ZN(net_1888), .A(net_1887) );
INV_X4 inst_6038 ( .A(net_10192), .ZN(net_515) );
NAND2_X2 inst_3422 ( .A2(net_9014), .A1(net_9013), .ZN(net_8512) );
CLKBUF_X2 inst_13791 ( .A(net_13709), .Z(net_13710) );
CLKBUF_X2 inst_13266 ( .A(net_13184), .Z(net_13185) );
NAND2_X2 inst_3832 ( .ZN(net_4870), .A2(net_4370), .A1(net_3297) );
NAND2_X2 inst_3978 ( .A1(net_10020), .ZN(net_3282), .A2(net_2468) );
INV_X4 inst_6618 ( .ZN(net_9034), .A(net_8941) );
NAND2_X2 inst_4039 ( .A1(net_3090), .A2(net_3056), .ZN(net_2852) );
INV_X4 inst_6106 ( .ZN(net_3933), .A(net_267) );
CLKBUF_X2 inst_11264 ( .A(net_11182), .Z(net_11183) );
NOR2_X2 inst_2967 ( .A2(net_4446), .ZN(net_1632), .A1(net_1109) );
AOI22_X2 inst_9354 ( .B1(net_9794), .A1(net_6828), .A2(net_5766), .B2(net_5765), .ZN(net_5568) );
CLKBUF_X2 inst_13279 ( .A(net_13197), .Z(net_13198) );
AOI21_X2 inst_10214 ( .ZN(net_2429), .B1(net_2428), .B2(net_2185), .A(net_815) );
AOI21_X2 inst_10042 ( .A(net_9544), .B1(net_9535), .ZN(net_7577), .B2(net_7575) );
AOI22_X2 inst_9161 ( .A2(net_6404), .ZN(net_6313), .B2(net_5263), .B1(net_2590), .A1(net_1849) );
OAI211_X2 inst_2078 ( .C2(net_6778), .ZN(net_6770), .A(net_6397), .B(net_6131), .C1(net_387) );
INV_X4 inst_6555 ( .ZN(net_8455), .A(net_220) );
INV_X4 inst_5674 ( .ZN(net_4603), .A(net_3209) );
AOI22_X2 inst_9029 ( .A1(net_9757), .ZN(net_7935), .A2(net_6418), .B2(net_5263), .B1(net_2707) );
CLKBUF_X2 inst_14873 ( .A(net_13596), .Z(net_14792) );
OR3_X4 inst_699 ( .A3(net_10514), .A2(net_10037), .ZN(net_7728), .A1(net_4442) );
DFF_X1 inst_8509 ( .Q(net_9425), .D(net_7622), .CK(net_13783) );
OAI221_X2 inst_1462 ( .C1(net_9087), .B2(net_7974), .C2(net_7973), .ZN(net_7960), .A(net_7959), .B1(net_2992) );
DFF_X2 inst_8377 ( .Q(net_9200), .D(net_2751), .CK(net_11239) );
OAI211_X2 inst_2273 ( .C1(net_7211), .C2(net_6480), .ZN(net_6263), .B(net_5412), .A(net_3679) );
AOI22_X2 inst_9138 ( .A1(net_9722), .A2(net_6382), .ZN(net_6350), .B1(net_6349), .B2(net_5263) );
AOI221_X2 inst_9921 ( .B2(net_5867), .ZN(net_5865), .C1(net_5864), .A(net_5859), .C2(net_4725), .B1(x5498) );
CLKBUF_X2 inst_13944 ( .A(net_13862), .Z(net_13863) );
INV_X4 inst_6391 ( .A(net_10047), .ZN(net_5094) );
OAI21_X2 inst_2003 ( .ZN(net_2805), .A(net_2147), .B1(net_2146), .B2(net_1682) );
AOI22_X2 inst_9514 ( .B1(net_9892), .A1(net_9761), .B2(net_4969), .ZN(net_3809), .A2(net_2462) );
INV_X4 inst_5430 ( .ZN(net_1537), .A(net_1129) );
INV_X4 inst_6084 ( .A(net_10065), .ZN(net_500) );
INV_X4 inst_6100 ( .A(net_10332), .ZN(net_692) );
CLKBUF_X2 inst_13823 ( .A(net_13741), .Z(net_13742) );
INV_X4 inst_5119 ( .ZN(net_1617), .A(net_1549) );
INV_X4 inst_4963 ( .A(net_6165), .ZN(net_3071) );
NOR2_X2 inst_2787 ( .A1(net_4376), .ZN(net_3078), .A2(net_3074) );
CLKBUF_X2 inst_14880 ( .A(net_14798), .Z(net_14799) );
INV_X4 inst_5612 ( .ZN(net_3772), .A(net_871) );
CLKBUF_X2 inst_13638 ( .A(net_13556), .Z(net_13557) );
CLKBUF_X2 inst_13144 ( .A(net_13062), .Z(net_13063) );
CLKBUF_X2 inst_12455 ( .A(net_12373), .Z(net_12374) );
CLKBUF_X2 inst_11074 ( .A(net_10987), .Z(net_10993) );
AOI22_X2 inst_9386 ( .B1(net_9801), .A1(net_5766), .B2(net_5765), .ZN(net_5437), .A2(net_239) );
NOR3_X2 inst_2426 ( .A2(net_7648), .A1(net_4631), .ZN(net_4611), .A3(net_3336) );
NOR2_X2 inst_2599 ( .ZN(net_7079), .A2(net_6665), .A1(net_2678) );
INV_X4 inst_6254 ( .A(net_10287), .ZN(net_455) );
CLKBUF_X2 inst_14211 ( .A(net_14129), .Z(net_14130) );
NAND2_X2 inst_3971 ( .ZN(net_3516), .A1(net_3311), .A2(net_3310) );
INV_X4 inst_6377 ( .ZN(net_3528), .A(net_190) );
CLKBUF_X2 inst_14528 ( .A(net_11423), .Z(net_14447) );
OAI221_X2 inst_1485 ( .ZN(net_7455), .C1(net_7454), .B1(net_7454), .A(net_7176), .B2(net_3910), .C2(net_3907) );
CLKBUF_X2 inst_11573 ( .A(net_11491), .Z(net_11492) );
AOI221_X2 inst_9858 ( .A(net_6889), .B2(net_6888), .C2(net_6887), .ZN(net_6860), .B1(net_4573), .C1(x4209) );
CLKBUF_X2 inst_13596 ( .A(net_13514), .Z(net_13515) );
CLKBUF_X2 inst_12259 ( .A(net_11121), .Z(net_12178) );
OR2_X4 inst_750 ( .ZN(net_5295), .A2(net_5178), .A1(net_4481) );
XNOR2_X2 inst_317 ( .ZN(net_3218), .A(net_2801), .B(net_2647) );
AND2_X2 inst_10561 ( .A1(net_9224), .ZN(net_3480), .A2(net_3098) );
OAI22_X2 inst_1123 ( .B1(net_7602), .ZN(net_5172), .A2(net_4465), .B2(net_3880), .A1(net_2769) );
DFF_X1 inst_8747 ( .Q(net_10345), .D(net_5423), .CK(net_10627) );
CLKBUF_X2 inst_13383 ( .A(net_13301), .Z(net_13302) );
XNOR2_X2 inst_278 ( .ZN(net_3675), .A(net_3502), .B(net_1906) );
MUX2_X2 inst_4429 ( .B(net_9152), .S(net_7553), .Z(net_7498), .A(net_666) );
SDFF_X2 inst_467 ( .SE(net_8747), .SI(net_8633), .Q(net_238), .D(net_107), .CK(net_11580) );
CLKBUF_X2 inst_11763 ( .A(net_11681), .Z(net_11682) );
NAND2_X2 inst_3677 ( .A1(net_9087), .ZN(net_7275), .A2(net_6230) );
INV_X2 inst_7169 ( .A(net_10367), .ZN(net_549) );
NAND2_X2 inst_3456 ( .A1(net_9497), .A2(net_8473), .ZN(net_8468) );
DFF_X2 inst_8061 ( .QN(net_10456), .D(net_5340), .CK(net_14703) );
OAI221_X2 inst_1628 ( .C1(net_10307), .B1(net_7192), .C2(net_5591), .ZN(net_5579), .B2(net_4902), .A(net_3507) );
NOR2_X2 inst_2963 ( .ZN(net_2425), .A1(net_938), .A2(net_753) );
DFF_X2 inst_7923 ( .QN(net_10367), .D(net_5820), .CK(net_13652) );
INV_X2 inst_6844 ( .ZN(net_3545), .A(net_3544) );
AND2_X2 inst_10535 ( .ZN(net_3726), .A1(net_3725), .A2(net_3724) );
AOI22_X2 inst_9640 ( .B1(net_9960), .A2(net_4694), .ZN(net_3402), .B2(net_2541), .A1(net_225) );
OAI222_X2 inst_1329 ( .C2(net_9603), .ZN(net_8585), .C1(net_8566), .A1(net_8565), .A2(net_8564), .B2(net_3372), .B1(net_498) );
OAI22_X2 inst_1204 ( .A1(net_7124), .A2(net_5134), .B2(net_5133), .ZN(net_5047), .B1(net_3532) );
DFF_X1 inst_8687 ( .D(net_6715), .Q(net_139), .CK(net_14252) );
NAND2_X2 inst_4066 ( .ZN(net_2971), .A2(net_2536), .A1(x6445) );
XNOR2_X2 inst_225 ( .ZN(net_4417), .B(net_4157), .A(net_4156) );
INV_X4 inst_4840 ( .ZN(net_4175), .A(net_3336) );
DFF_X2 inst_7669 ( .D(net_6703), .QN(net_189), .CK(net_12281) );
CLKBUF_X2 inst_14261 ( .A(net_14179), .Z(net_14180) );
CLKBUF_X2 inst_13568 ( .A(net_11569), .Z(net_13487) );
CLKBUF_X2 inst_12530 ( .A(net_10732), .Z(net_12449) );
AOI22_X2 inst_9030 ( .B2(net_10381), .ZN(net_7667), .A2(net_7545), .A1(net_7477), .B1(net_903) );
INV_X4 inst_5020 ( .ZN(net_3719), .A(net_1983) );
CLKBUF_X2 inst_14808 ( .A(net_14726), .Z(net_14727) );
CLKBUF_X2 inst_13158 ( .A(net_12407), .Z(net_13077) );
AOI21_X2 inst_10162 ( .A(net_10304), .B1(net_10280), .ZN(net_4169), .B2(net_2828) );
HA_X1 inst_7349 ( .S(net_4430), .CO(net_4429), .B(net_4200), .A(net_979) );
SDFF_X2 inst_508 ( .SI(net_9342), .Q(net_9287), .D(net_9287), .SE(net_7588), .CK(net_14700) );
CLKBUF_X2 inst_11015 ( .A(net_10807), .Z(net_10934) );
INV_X4 inst_4888 ( .ZN(net_4070), .A(net_3390) );
DFF_X2 inst_8150 ( .QN(net_9752), .D(net_5081), .CK(net_12977) );
CLKBUF_X2 inst_11718 ( .A(net_10723), .Z(net_11637) );
CLKBUF_X2 inst_12611 ( .A(net_12529), .Z(net_12530) );
NOR2_X2 inst_2618 ( .ZN(net_6206), .A1(net_5764), .A2(net_1752) );
CLKBUF_X2 inst_15065 ( .A(net_14983), .Z(net_14984) );
CLKBUF_X2 inst_10952 ( .A(net_10870), .Z(net_10871) );
INV_X4 inst_4950 ( .ZN(net_3084), .A(net_2854) );
CLKBUF_X2 inst_14726 ( .A(net_14644), .Z(net_14645) );
DFF_X1 inst_8853 ( .Q(net_10525), .D(net_97), .CK(net_11202) );
CLKBUF_X2 inst_11443 ( .A(net_11361), .Z(net_11362) );
AOI22_X2 inst_9241 ( .A1(net_9945), .B1(net_9846), .A2(net_6141), .B2(net_6133), .ZN(net_6070) );
SDFF_X2 inst_590 ( .Q(net_9261), .SE(net_4589), .D(net_144), .SI(net_110), .CK(net_13829) );
NOR2_X2 inst_2553 ( .ZN(net_7862), .A2(net_7861), .A1(net_7859) );
CLKBUF_X2 inst_12209 ( .A(net_12127), .Z(net_12128) );
CLKBUF_X2 inst_13051 ( .A(net_12280), .Z(net_12970) );
CLKBUF_X2 inst_12671 ( .A(net_12589), .Z(net_12590) );
CLKBUF_X2 inst_14428 ( .A(net_11216), .Z(net_14347) );
CLKBUF_X2 inst_13897 ( .A(net_13815), .Z(net_13816) );
OAI21_X2 inst_1729 ( .ZN(net_8784), .A(net_8783), .B1(net_8773), .B2(net_8767) );
DFF_X2 inst_8346 ( .QN(net_10444), .D(net_2820), .CK(net_11115) );
OAI22_X2 inst_1105 ( .A1(net_7535), .ZN(net_6199), .A2(net_5733), .B2(net_5732), .B1(net_383) );
INV_X8 inst_4531 ( .A(net_9100), .ZN(net_9098) );
CLKBUF_X2 inst_14746 ( .A(net_14664), .Z(net_14665) );
CLKBUF_X2 inst_13175 ( .A(net_13093), .Z(net_13094) );
NOR2_X2 inst_2746 ( .A1(net_3687), .ZN(net_3682), .A2(net_3681) );
INV_X4 inst_6126 ( .A(net_9117), .ZN(net_627) );
CLKBUF_X2 inst_14387 ( .A(net_14305), .Z(net_14306) );
INV_X2 inst_6996 ( .ZN(net_1633), .A(net_1632) );
CLKBUF_X2 inst_13576 ( .A(net_13494), .Z(net_13495) );
CLKBUF_X2 inst_15202 ( .A(net_15120), .Z(net_15121) );
INV_X4 inst_4648 ( .ZN(net_6848), .A(net_6846) );
AND2_X4 inst_10469 ( .A2(net_9640), .A1(net_9637), .ZN(net_781) );
DFF_X2 inst_8200 ( .QN(net_9734), .D(net_5060), .CK(net_12254) );
INV_X2 inst_6961 ( .ZN(net_5511), .A(net_1866) );
XNOR2_X2 inst_330 ( .ZN(net_2997), .B(net_2728), .A(net_2449) );
CLKBUF_X2 inst_13345 ( .A(net_13263), .Z(net_13264) );
AOI211_X2 inst_10297 ( .ZN(net_3743), .A(net_3742), .B(net_3741), .C2(net_3318), .C1(net_2960) );
CLKBUF_X2 inst_13558 ( .A(net_13476), .Z(net_13477) );
CLKBUF_X2 inst_11460 ( .A(net_11378), .Z(net_11379) );
DFF_X2 inst_7595 ( .Q(net_10191), .D(net_7447), .CK(net_12286) );
XNOR2_X2 inst_165 ( .ZN(net_5946), .A(net_5369), .B(net_2329) );
NAND2_X2 inst_3733 ( .ZN(net_6299), .A2(net_5447), .A1(net_1397) );
NAND2_X2 inst_4305 ( .A2(net_10474), .ZN(net_1615), .A1(net_1210) );
CLKBUF_X2 inst_12101 ( .A(net_12019), .Z(net_12020) );
CLKBUF_X2 inst_13546 ( .A(net_13464), .Z(net_13465) );
INV_X4 inst_5376 ( .A(net_2761), .ZN(net_1959) );
DFF_X1 inst_8786 ( .Q(net_10134), .D(net_4574), .CK(net_10777) );
OAI22_X2 inst_1176 ( .A1(net_7229), .A2(net_5107), .B2(net_5105), .ZN(net_5085), .B1(net_5084) );
NAND2_X2 inst_3566 ( .A2(net_7748), .ZN(net_7682), .A1(net_7681) );
CLKBUF_X2 inst_13864 ( .A(net_13782), .Z(net_13783) );
CLKBUF_X2 inst_12537 ( .A(net_12455), .Z(net_12456) );
CLKBUF_X2 inst_11803 ( .A(net_11721), .Z(net_11722) );
DFF_X2 inst_8159 ( .QN(net_9934), .D(net_5063), .CK(net_13303) );
CLKBUF_X2 inst_15455 ( .A(net_15373), .Z(net_15374) );
CLKBUF_X2 inst_12696 ( .A(net_11268), .Z(net_12615) );
OAI22_X2 inst_1232 ( .B1(net_7213), .A2(net_4890), .B2(net_4889), .ZN(net_4885), .A1(net_508) );
INV_X4 inst_5450 ( .ZN(net_5053), .A(net_4380) );
CLKBUF_X2 inst_15706 ( .A(net_15624), .Z(net_15625) );
CLKBUF_X2 inst_14431 ( .A(net_14349), .Z(net_14350) );
CLKBUF_X2 inst_11340 ( .A(net_11258), .Z(net_11259) );
NAND2_X2 inst_4172 ( .A2(net_4788), .ZN(net_3695), .A1(net_610) );
CLKBUF_X2 inst_13388 ( .A(net_13306), .Z(net_13307) );
NOR2_X2 inst_2605 ( .ZN(net_6270), .A1(net_5764), .A2(net_2523) );
OR2_X4 inst_758 ( .ZN(net_4871), .A1(net_4371), .A2(net_4370) );
CLKBUF_X2 inst_14423 ( .A(net_13560), .Z(net_14342) );
CLKBUF_X2 inst_14147 ( .A(net_14065), .Z(net_14066) );
OAI211_X2 inst_2146 ( .C2(net_6774), .ZN(net_6702), .A(net_6327), .B(net_6065), .C1(net_4747) );
CLKBUF_X2 inst_13759 ( .A(net_13677), .Z(net_13678) );
CLKBUF_X2 inst_13332 ( .A(net_13250), .Z(net_13251) );
INV_X2 inst_7252 ( .A(net_8825), .ZN(net_345) );
DFF_X1 inst_8543 ( .Q(net_9977), .D(net_7348), .CK(net_14627) );
CLKBUF_X2 inst_13717 ( .A(net_13635), .Z(net_13636) );
NOR2_X2 inst_2703 ( .ZN(net_4826), .A1(net_4391), .A2(net_4082) );
NAND2_X2 inst_3437 ( .A2(net_9475), .ZN(net_8892), .A1(net_8482) );
CLKBUF_X2 inst_13425 ( .A(net_13343), .Z(net_13344) );
INV_X2 inst_6813 ( .ZN(net_4732), .A(net_4731) );
CLKBUF_X2 inst_13857 ( .A(net_13775), .Z(net_13776) );
AOI221_X2 inst_9784 ( .B1(net_9974), .ZN(net_7091), .A(net_7090), .B2(net_7089), .C1(net_7088), .C2(net_246) );
INV_X4 inst_5764 ( .ZN(net_1756), .A(net_724) );
XNOR2_X2 inst_143 ( .ZN(net_7301), .A(net_6659), .B(net_2179) );
DFF_X2 inst_7442 ( .QN(net_9299), .D(net_8196), .CK(net_11500) );
OAI21_X2 inst_1953 ( .B1(net_4071), .ZN(net_3921), .A(net_3920), .B2(net_3919) );
INV_X4 inst_4570 ( .ZN(net_9012), .A(net_8385) );
INV_X4 inst_5286 ( .ZN(net_5467), .A(net_1321) );
NOR2_X2 inst_3016 ( .A2(net_10408), .A1(net_10407), .ZN(net_750) );
INV_X4 inst_6260 ( .A(net_10281), .ZN(net_450) );
OAI21_X2 inst_1958 ( .ZN(net_3940), .B2(net_3471), .A(net_3109), .B1(net_2049) );
NAND2_X2 inst_4272 ( .A2(net_10142), .ZN(net_1500), .A1(net_895) );
CLKBUF_X2 inst_14050 ( .A(net_13968), .Z(net_13969) );
NOR4_X2 inst_2337 ( .ZN(net_3343), .A1(net_2874), .A2(net_2870), .A4(net_2800), .A3(net_2289) );
NAND3_X2 inst_3250 ( .ZN(net_4582), .A1(net_4581), .A3(net_4580), .A2(net_2204) );
CLKBUF_X2 inst_15052 ( .A(net_14970), .Z(net_14971) );
AOI22_X2 inst_9403 ( .ZN(net_5974), .A2(net_4700), .B1(net_3706), .B2(net_2696), .A1(net_2380) );
AOI22_X2 inst_9357 ( .B1(net_9912), .A2(net_5759), .B2(net_5758), .ZN(net_5565), .A1(net_251) );
OAI21_X2 inst_1778 ( .ZN(net_7787), .B1(net_7785), .A(net_7723), .B2(net_7722) );
NAND3_X2 inst_3240 ( .A1(net_7142), .ZN(net_4715), .A2(net_4714), .A3(net_4713) );
INV_X2 inst_6885 ( .A(net_4376), .ZN(net_2841) );
CLKBUF_X2 inst_12132 ( .A(net_12050), .Z(net_12051) );
DFF_X2 inst_8091 ( .QN(net_10037), .D(net_5067), .CK(net_11446) );
OAI21_X2 inst_1736 ( .B2(net_9049), .ZN(net_8987), .B1(net_8711), .A(net_8141) );
OAI22_X2 inst_1040 ( .A2(net_8921), .B1(net_8918), .A1(net_8116), .ZN(net_7949), .B2(net_3080) );
NAND2_X2 inst_4027 ( .ZN(net_3294), .A2(net_3084), .A1(net_610) );
CLKBUF_X2 inst_15218 ( .A(net_15136), .Z(net_15137) );
AOI22_X2 inst_9158 ( .A2(net_6418), .ZN(net_6323), .B2(net_5263), .A1(net_4211), .B1(net_2984) );
INV_X4 inst_6009 ( .A(net_10045), .ZN(net_6148) );
INV_X4 inst_5042 ( .A(net_5175), .ZN(net_5021) );
CLKBUF_X2 inst_13196 ( .A(net_13114), .Z(net_13115) );
XNOR2_X2 inst_111 ( .A(net_8946), .ZN(net_8084), .B(net_7056) );
OAI21_X4 inst_1723 ( .ZN(net_8778), .A(net_8761), .B1(net_8760), .B2(net_8759) );
NAND4_X2 inst_3146 ( .ZN(net_2161), .A4(net_1343), .A2(net_1053), .A1(net_607), .A3(net_575) );
NAND3_X2 inst_3278 ( .ZN(net_4049), .A1(net_4047), .A3(net_4046), .A2(net_3316) );
AOI21_X2 inst_10246 ( .ZN(net_8866), .B1(net_2394), .B2(net_2393), .A(net_2392) );
INV_X2 inst_7303 ( .A(net_9072), .ZN(net_9071) );
CLKBUF_X2 inst_11651 ( .A(net_11569), .Z(net_11570) );
CLKBUF_X2 inst_11425 ( .A(net_11343), .Z(net_11344) );
OAI211_X2 inst_2056 ( .ZN(net_7784), .A(net_7783), .C1(net_7782), .B(net_7688), .C2(net_4405) );
INV_X4 inst_5145 ( .A(net_3400), .ZN(net_1923) );
OAI211_X2 inst_2116 ( .C2(net_6778), .ZN(net_6732), .A(net_6359), .B(net_6093), .C1(net_322) );
CLKBUF_X2 inst_11296 ( .A(net_10607), .Z(net_11215) );
NOR2_X2 inst_2825 ( .A1(net_3207), .A2(net_3065), .ZN(net_2526) );
INV_X4 inst_5071 ( .ZN(net_3353), .A(net_1849) );
CLKBUF_X2 inst_13407 ( .A(net_13325), .Z(net_13326) );
NAND2_X2 inst_4031 ( .ZN(net_3473), .A2(net_3002), .A1(net_2031) );
CLKBUF_X2 inst_15370 ( .A(net_15288), .Z(net_15289) );
DFF_X2 inst_8135 ( .Q(net_9838), .D(net_5122), .CK(net_14287) );
XNOR2_X2 inst_346 ( .ZN(net_2861), .B(net_2860), .A(net_1517) );
DFF_X1 inst_8755 ( .Q(net_10170), .D(net_5246), .CK(net_12306) );
CLKBUF_X2 inst_14757 ( .A(net_14675), .Z(net_14676) );
OAI22_X2 inst_978 ( .A2(net_9581), .ZN(net_8688), .A1(net_8687), .B2(net_8677), .B1(net_8206) );
CLKBUF_X2 inst_13506 ( .A(net_13424), .Z(net_13425) );
CLKBUF_X2 inst_10711 ( .A(net_10594), .Z(net_10630) );
NOR2_X2 inst_2955 ( .ZN(net_2396), .A1(net_678), .A2(net_555) );
CLKBUF_X2 inst_12058 ( .A(net_11976), .Z(net_11977) );
NAND2_X2 inst_3926 ( .A2(net_4319), .ZN(net_3881), .A1(net_1936) );
INV_X2 inst_7293 ( .A(net_9046), .ZN(net_9043) );
INV_X4 inst_6195 ( .A(net_10117), .ZN(net_2129) );
AOI221_X2 inst_9777 ( .B1(net_8957), .ZN(net_7380), .C2(net_7379), .B2(net_7379), .C1(net_7378), .A(net_6906) );
CLKBUF_X2 inst_11347 ( .A(net_11265), .Z(net_11266) );
CLKBUF_X2 inst_13160 ( .A(net_13018), .Z(net_13079) );
CLKBUF_X2 inst_12972 ( .A(net_12890), .Z(net_12891) );
NAND2_X2 inst_3929 ( .A2(net_4319), .ZN(net_3877), .A1(net_2886) );
DFF_X1 inst_8856 ( .Q(net_10524), .D(net_96), .CK(net_11198) );
CLKBUF_X2 inst_12312 ( .A(net_12230), .Z(net_12231) );
AND2_X2 inst_10506 ( .A2(net_10273), .ZN(net_5969), .A1(net_5407) );
AOI221_X2 inst_9745 ( .ZN(net_7937), .A(net_7818), .C2(net_3106), .C1(net_2928), .B1(net_2846), .B2(net_2845) );
NAND2_X2 inst_3852 ( .A1(net_10530), .A2(net_4361), .ZN(net_4329) );
CLKBUF_X2 inst_15131 ( .A(net_11319), .Z(net_15050) );
CLKBUF_X2 inst_14168 ( .A(net_11351), .Z(net_14087) );
CLKBUF_X2 inst_14366 ( .A(net_14284), .Z(net_14285) );
OAI22_X2 inst_1051 ( .ZN(net_7533), .A1(net_7531), .B2(net_7530), .A2(net_7387), .B1(net_3093) );
SDFF_X2 inst_495 ( .SE(net_9540), .SI(net_8214), .Q(net_283), .D(net_283), .CK(net_12708) );
NOR2_X2 inst_2566 ( .ZN(net_7715), .A2(net_7517), .A1(net_7431) );
CLKBUF_X2 inst_15041 ( .A(net_14959), .Z(net_14960) );
INV_X4 inst_6102 ( .A(net_10026), .ZN(net_1209) );
INV_X4 inst_6437 ( .A(net_9552), .ZN(net_8182) );
OAI21_X2 inst_1864 ( .ZN(net_5910), .A(net_5363), .B1(net_5362), .B2(net_5346) );
CLKBUF_X2 inst_12901 ( .A(net_12819), .Z(net_12820) );
AOI22_X2 inst_9632 ( .A1(net_10053), .B1(net_9824), .A2(net_5174), .ZN(net_3411), .B2(net_2556) );
NAND2_X2 inst_3603 ( .ZN(net_7263), .A2(net_6857), .A1(net_6603) );
CLKBUF_X2 inst_11076 ( .A(net_10994), .Z(net_10995) );
NAND3_X2 inst_3224 ( .ZN(net_5282), .A1(net_4768), .A2(net_3800), .A3(net_3798) );
CLKBUF_X2 inst_10887 ( .A(net_10606), .Z(net_10806) );
NAND4_X2 inst_3043 ( .A1(net_8966), .A3(net_8959), .A2(net_8057), .ZN(net_7427), .A4(net_7093) );
DFF_X2 inst_8063 ( .QN(net_10457), .D(net_5330), .CK(net_12463) );
CLKBUF_X2 inst_13665 ( .A(net_12314), .Z(net_13584) );
DFF_X2 inst_7917 ( .Q(net_10044), .D(net_5874), .CK(net_11938) );
CLKBUF_X2 inst_15826 ( .A(net_15744), .Z(net_15745) );
CLKBUF_X2 inst_12616 ( .A(net_12534), .Z(net_12535) );
INV_X4 inst_5752 ( .A(net_2497), .ZN(net_736) );
CLKBUF_X2 inst_13305 ( .A(net_13223), .Z(net_13224) );
CLKBUF_X2 inst_12644 ( .A(net_12562), .Z(net_12563) );
INV_X2 inst_7286 ( .A(net_8980), .ZN(net_8979) );
CLKBUF_X2 inst_14969 ( .A(net_14887), .Z(net_14888) );
AND2_X2 inst_10548 ( .A1(net_3670), .A2(net_3489), .ZN(net_3484) );
CLKBUF_X2 inst_13781 ( .A(net_13699), .Z(net_13700) );
NOR2_X2 inst_2893 ( .ZN(net_1721), .A2(net_1720), .A1(net_811) );
CLKBUF_X2 inst_11360 ( .A(net_10925), .Z(net_11279) );
AOI22_X2 inst_9497 ( .A1(net_9887), .B1(net_9788), .ZN(net_3826), .A2(net_2973), .B2(net_2462) );
SDFF_X2 inst_573 ( .D(net_9129), .SE(net_933), .CK(net_10934), .SI(x2648), .Q(x1274) );
DFF_X2 inst_7736 ( .Q(net_9699), .D(net_6196), .CK(net_14236) );
CLKBUF_X2 inst_12447 ( .A(net_12365), .Z(net_12366) );
INV_X2 inst_6727 ( .A(net_7795), .ZN(net_7761) );
DFF_X2 inst_7937 ( .QN(net_10416), .D(net_5539), .CK(net_11597) );
AOI22_X2 inst_9041 ( .A1(net_9153), .A2(net_7155), .B2(net_7154), .ZN(net_7014), .B1(net_1988) );
INV_X4 inst_6347 ( .A(net_10251), .ZN(net_962) );
DFF_X2 inst_8088 ( .QN(net_10026), .D(net_5033), .CK(net_13712) );
INV_X4 inst_5364 ( .ZN(net_2308), .A(net_1218) );
OAI221_X2 inst_1453 ( .ZN(net_7980), .C2(net_7800), .A(net_7798), .B2(net_7762), .B1(net_7712), .C1(net_6211) );
NAND2_X2 inst_4245 ( .A1(net_10259), .A2(net_2014), .ZN(net_1785) );
CLKBUF_X2 inst_12466 ( .A(net_10957), .Z(net_12385) );
CLKBUF_X2 inst_12391 ( .A(net_12309), .Z(net_12310) );
DFF_X1 inst_8871 ( .Q(net_93), .CK(net_14114), .D(x3349) );
NOR2_X2 inst_3007 ( .A1(net_10457), .ZN(net_1185), .A2(net_842) );
CLKBUF_X1 inst_8978 ( .A(x185142), .Z(x19) );
CLKBUF_X2 inst_15081 ( .A(net_14999), .Z(net_15000) );
NAND2_X2 inst_4185 ( .ZN(net_2116), .A2(net_1864), .A1(net_969) );
CLKBUF_X2 inst_11018 ( .A(net_10936), .Z(net_10937) );
NAND2_X2 inst_3512 ( .A2(net_8238), .ZN(net_8168), .A1(net_8140) );
NAND2_X2 inst_3544 ( .ZN(net_9001), .A2(net_7989), .A1(net_2362) );
INV_X4 inst_6358 ( .ZN(net_708), .A(net_167) );
CLKBUF_X2 inst_11485 ( .A(net_11403), .Z(net_11404) );
CLKBUF_X2 inst_10738 ( .A(net_10656), .Z(net_10657) );
CLKBUF_X2 inst_10973 ( .A(net_10891), .Z(net_10892) );
INV_X4 inst_5632 ( .A(net_7562), .ZN(net_859) );
CLKBUF_X2 inst_14839 ( .A(net_10811), .Z(net_14758) );
OAI22_X2 inst_1206 ( .A1(net_7124), .A2(net_5139), .B2(net_5138), .ZN(net_5045), .B1(net_3718) );
DFF_X2 inst_7970 ( .QN(net_10321), .D(net_5583), .CK(net_14600) );
CLKBUF_X2 inst_15778 ( .A(net_12385), .Z(net_15697) );
CLKBUF_X2 inst_13607 ( .A(net_12466), .Z(net_13526) );
AOI22_X2 inst_9362 ( .B1(net_9922), .A1(net_6811), .A2(net_5759), .B2(net_5758), .ZN(net_5560) );
CLKBUF_X2 inst_15270 ( .A(net_15188), .Z(net_15189) );
INV_X4 inst_6367 ( .A(net_10406), .ZN(net_3672) );
INV_X2 inst_6773 ( .ZN(net_6028), .A(net_5850) );
CLKBUF_X2 inst_15485 ( .A(net_15403), .Z(net_15404) );
AND4_X4 inst_10328 ( .ZN(net_3321), .A4(net_3320), .A3(net_2275), .A2(net_1387), .A1(net_1385) );
INV_X2 inst_7075 ( .A(net_4921), .ZN(net_1224) );
NAND2_X2 inst_3466 ( .A1(net_9492), .A2(net_8476), .ZN(net_8457) );
DFF_X2 inst_8106 ( .QN(net_9944), .D(net_5113), .CK(net_12500) );
CLKBUF_X2 inst_13907 ( .A(net_11056), .Z(net_13826) );
DFF_X2 inst_8358 ( .QN(net_10442), .D(net_2268), .CK(net_11145) );
INV_X4 inst_4800 ( .A(net_3707), .ZN(net_3659) );
CLKBUF_X2 inst_15684 ( .A(net_10545), .Z(net_15603) );
NAND2_X2 inst_4394 ( .A2(net_10506), .A1(net_10493), .ZN(net_735) );
CLKBUF_X2 inst_11303 ( .A(net_10963), .Z(net_11222) );
INV_X4 inst_5553 ( .A(net_10220), .ZN(net_1245) );
CLKBUF_X2 inst_13086 ( .A(net_13004), .Z(net_13005) );
CLKBUF_X2 inst_12631 ( .A(net_12549), .Z(net_12550) );
CLKBUF_X2 inst_11518 ( .A(net_11436), .Z(net_11437) );
OAI221_X2 inst_1487 ( .B2(net_7671), .ZN(net_7438), .C2(net_7437), .A(net_7141), .B1(net_4085), .C1(net_3288) );
INV_X4 inst_6111 ( .A(net_10260), .ZN(net_1211) );
DFF_X2 inst_7807 ( .Q(net_9991), .D(net_6482), .CK(net_15235) );
CLKBUF_X2 inst_13169 ( .A(net_13087), .Z(net_13088) );
OAI21_X2 inst_1933 ( .B1(net_5457), .A(net_4414), .ZN(net_4372), .B2(net_4003) );
NAND2_X2 inst_3522 ( .A2(net_9595), .ZN(net_8314), .A1(net_8116) );
INV_X2 inst_7246 ( .ZN(net_363), .A(net_202) );
CLKBUF_X2 inst_15795 ( .A(net_15713), .Z(net_15714) );
INV_X4 inst_6306 ( .ZN(net_426), .A(x769) );
CLKBUF_X2 inst_14119 ( .A(net_14037), .Z(net_14038) );
DFF_X2 inst_7511 ( .Q(net_9535), .D(net_7934), .CK(net_13997) );
OAI21_X2 inst_1758 ( .ZN(net_8502), .B1(net_8443), .A(net_5787), .B2(net_5383) );
OAI22_X2 inst_1142 ( .A1(net_7243), .A2(net_5134), .B2(net_5133), .ZN(net_5131), .B1(net_390) );
INV_X4 inst_6280 ( .A(net_10400), .ZN(net_442) );
CLKBUF_X2 inst_12025 ( .A(net_11943), .Z(net_11944) );
NAND2_X2 inst_4320 ( .A1(net_4446), .ZN(net_2349), .A2(net_1109) );
NAND2_X2 inst_3816 ( .A1(net_10085), .A2(net_4534), .ZN(net_4522) );
CLKBUF_X2 inst_11138 ( .A(net_10696), .Z(net_11057) );
CLKBUF_X2 inst_14914 ( .A(net_14832), .Z(net_14833) );
CLKBUF_X2 inst_14772 ( .A(net_13690), .Z(net_14691) );
INV_X4 inst_5418 ( .A(net_8687), .ZN(net_8677) );
OAI222_X2 inst_1381 ( .B1(net_7728), .A2(net_7727), .C2(net_7726), .ZN(net_6004), .B2(net_5192), .A1(net_3995), .C1(net_1284) );
CLKBUF_X2 inst_15527 ( .A(net_15445), .Z(net_15446) );
SDFF_X2 inst_643 ( .Q(net_9442), .D(net_9442), .SE(net_3293), .CK(net_14146), .SI(x3022) );
DFF_X2 inst_7572 ( .QN(net_9239), .D(net_7570), .CK(net_11260) );
INV_X4 inst_6313 ( .A(net_9752), .ZN(net_6321) );
DFF_X2 inst_7680 ( .QN(net_9422), .D(net_6627), .CK(net_13876) );
CLKBUF_X2 inst_12471 ( .A(net_12389), .Z(net_12390) );
CLKBUF_X2 inst_15516 ( .A(net_15209), .Z(net_15435) );
CLKBUF_X2 inst_13726 ( .A(net_13644), .Z(net_13645) );
CLKBUF_X2 inst_14316 ( .A(net_13683), .Z(net_14235) );
CLKBUF_X2 inst_14228 ( .A(net_10655), .Z(net_14147) );
AOI22_X2 inst_9430 ( .ZN(net_4592), .A1(net_4419), .A2(net_4282), .B2(net_3394), .B1(net_3178) );
CLKBUF_X2 inst_14182 ( .A(net_11959), .Z(net_14101) );
CLKBUF_X2 inst_10745 ( .A(net_10663), .Z(net_10664) );
DFF_X2 inst_7763 ( .Q(net_9716), .D(net_6538), .CK(net_12799) );
INV_X4 inst_4771 ( .ZN(net_7785), .A(net_3507) );
CLKBUF_X2 inst_12117 ( .A(net_12035), .Z(net_12036) );
CLKBUF_X2 inst_12220 ( .A(net_11791), .Z(net_12139) );
INV_X4 inst_4961 ( .A(net_5171), .ZN(net_3072) );
INV_X4 inst_4669 ( .ZN(net_5764), .A(net_5391) );
DFF_X2 inst_7695 ( .Q(net_10403), .D(net_6571), .CK(net_15144) );
CLKBUF_X2 inst_15091 ( .A(net_15009), .Z(net_15010) );
CLKBUF_X2 inst_15476 ( .A(net_15394), .Z(net_15395) );
DFF_X1 inst_8588 ( .Q(net_9766), .D(net_7109), .CK(net_14262) );
DFF_X2 inst_8016 ( .QN(net_10325), .D(net_5487), .CK(net_12133) );
DFF_X1 inst_8707 ( .Q(net_8827), .D(net_6952), .CK(net_13069) );
INV_X4 inst_6466 ( .A(net_9181), .ZN(net_5100) );
CLKBUF_X2 inst_12165 ( .A(net_12083), .Z(net_12084) );
CLKBUF_X2 inst_15191 ( .A(net_13797), .Z(net_15110) );
CLKBUF_X2 inst_13204 ( .A(net_13122), .Z(net_13123) );
DFF_X1 inst_8581 ( .Q(net_9674), .D(net_7106), .CK(net_14824) );
INV_X4 inst_5447 ( .ZN(net_1541), .A(net_1085) );
INV_X4 inst_6371 ( .A(net_10258), .ZN(net_1021) );
NAND2_X2 inst_4146 ( .A2(net_2766), .A1(net_2207), .ZN(net_2080) );
CLKBUF_X2 inst_12526 ( .A(net_11256), .Z(net_12445) );
CLKBUF_X2 inst_12230 ( .A(net_10758), .Z(net_12149) );
CLKBUF_X2 inst_12959 ( .A(net_12877), .Z(net_12878) );
CLKBUF_X2 inst_15650 ( .A(net_13008), .Z(net_15569) );
OAI21_X2 inst_1997 ( .ZN(net_3003), .B1(net_2490), .A(net_1617), .B2(net_1612) );
INV_X2 inst_6971 ( .ZN(net_1716), .A(net_1715) );
OAI22_X2 inst_1017 ( .A2(net_8247), .B2(net_8246), .ZN(net_8196), .A1(net_5931), .B1(net_1934) );
CLKBUF_X2 inst_12669 ( .A(net_12587), .Z(net_12588) );
OAI211_X2 inst_2297 ( .ZN(net_4631), .A(net_3366), .B(net_3147), .C2(net_2926), .C1(net_2374) );
NAND2_X2 inst_3736 ( .A1(net_6040), .ZN(net_5796), .A2(net_5372) );
CLKBUF_X2 inst_13802 ( .A(net_13720), .Z(net_13721) );
XNOR2_X2 inst_281 ( .ZN(net_3669), .B(net_3668), .A(net_3486) );
NAND2_X4 inst_3341 ( .ZN(net_9030), .A2(net_8887), .A1(net_8886) );
AOI211_X2 inst_10306 ( .B(net_5813), .C1(net_4188), .C2(net_3897), .ZN(net_3305), .A(net_2672) );
DFF_X1 inst_8500 ( .Q(net_9757), .D(net_7752), .CK(net_12911) );
INV_X4 inst_6336 ( .A(net_10096), .ZN(net_5843) );
CLKBUF_X2 inst_13411 ( .A(net_13329), .Z(net_13330) );
INV_X2 inst_7062 ( .A(net_3272), .ZN(net_1268) );
OAI21_X2 inst_1836 ( .ZN(net_6257), .A(net_6256), .B1(net_6255), .B2(net_5806) );
INV_X4 inst_6374 ( .A(net_9990), .ZN(net_399) );
CLKBUF_X2 inst_15296 ( .A(net_15214), .Z(net_15215) );
CLKBUF_X2 inst_14913 ( .A(net_14831), .Z(net_14832) );
INV_X2 inst_7005 ( .ZN(net_1616), .A(net_1615) );
NOR2_X2 inst_2508 ( .ZN(net_8401), .A2(net_8389), .A1(net_362) );
AOI21_X2 inst_10207 ( .ZN(net_2533), .A(net_2532), .B2(net_1785), .B1(net_1112) );
OAI211_X2 inst_2170 ( .C1(net_7201), .C2(net_6548), .A(net_6546), .ZN(net_6539), .B(net_5667) );
NAND2_X2 inst_4250 ( .ZN(net_2053), .A2(net_987), .A1(net_382) );
NAND2_X2 inst_4274 ( .A2(net_10219), .ZN(net_2773), .A1(net_743) );
CLKBUF_X2 inst_14642 ( .A(net_12076), .Z(net_14561) );
CLKBUF_X2 inst_15490 ( .A(net_15408), .Z(net_15409) );
CLKBUF_X2 inst_13322 ( .A(net_10897), .Z(net_13241) );
OR2_X4 inst_773 ( .ZN(net_4460), .A1(net_3140), .A2(net_3139) );
DFF_X2 inst_7414 ( .QN(net_9413), .D(net_8351), .CK(net_11710) );
CLKBUF_X2 inst_14149 ( .A(net_14067), .Z(net_14068) );
AOI221_X2 inst_9940 ( .ZN(net_5720), .B1(net_5719), .C1(net_5718), .A(net_5361), .B2(net_2498), .C2(net_837) );
NOR2_X2 inst_2946 ( .A1(net_10156), .A2(net_3496), .ZN(net_2214) );
CLKBUF_X2 inst_10776 ( .A(net_10694), .Z(net_10695) );
CLKBUF_X2 inst_15642 ( .A(net_15560), .Z(net_15561) );
CLKBUF_X2 inst_15234 ( .A(net_15152), .Z(net_15153) );
CLKBUF_X2 inst_13091 ( .A(net_10764), .Z(net_13010) );
AOI21_X2 inst_10074 ( .B2(net_9094), .ZN(net_5996), .A(net_5418), .B1(net_2865) );
NAND2_X2 inst_3620 ( .ZN(net_7106), .A1(net_6885), .A2(net_6672) );
CLKBUF_X2 inst_13827 ( .A(net_13745), .Z(net_13746) );
CLKBUF_X2 inst_10828 ( .A(net_10677), .Z(net_10747) );
CLKBUF_X2 inst_14134 ( .A(net_14052), .Z(net_14053) );
CLKBUF_X2 inst_14763 ( .A(net_14681), .Z(net_14682) );
AOI221_X2 inst_9798 ( .B1(net_9978), .A(net_7090), .B2(net_7089), .C2(net_7088), .ZN(net_7006), .C1(net_250) );
XNOR2_X2 inst_260 ( .B(net_4554), .ZN(net_3995), .A(net_3484) );
CLKBUF_X2 inst_11277 ( .A(net_11060), .Z(net_11196) );
AOI22_X2 inst_9371 ( .B1(net_9915), .A1(net_6823), .A2(net_5759), .B2(net_5758), .ZN(net_5551) );
CLKBUF_X2 inst_11597 ( .A(net_11515), .Z(net_11516) );
NAND3_X2 inst_3211 ( .ZN(net_6449), .A1(net_5884), .A2(net_3843), .A3(net_3842) );
INV_X4 inst_4973 ( .ZN(net_2317), .A(net_2316) );
AND3_X4 inst_10364 ( .ZN(net_5280), .A1(net_1505), .A3(net_1504), .A2(net_854) );
CLKBUF_X2 inst_12702 ( .A(net_11798), .Z(net_12621) );
INV_X2 inst_7270 ( .A(net_8929), .ZN(net_8928) );
NAND2_X2 inst_4139 ( .ZN(net_2515), .A2(net_2184), .A1(net_867) );
INV_X2 inst_6762 ( .A(net_7018), .ZN(net_6189) );
INV_X4 inst_4611 ( .A(net_9542), .ZN(net_7575) );
CLKBUF_X2 inst_13839 ( .A(net_13757), .Z(net_13758) );
CLKBUF_X2 inst_14803 ( .A(net_14721), .Z(net_14722) );
CLKBUF_X2 inst_10906 ( .A(net_10693), .Z(net_10825) );
CLKBUF_X2 inst_10725 ( .A(net_10562), .Z(net_10644) );
INV_X4 inst_4567 ( .ZN(net_9009), .A(net_8168) );
NAND2_X2 inst_3889 ( .ZN(net_4415), .A2(net_4005), .A1(net_3194) );
NOR3_X2 inst_2386 ( .A1(net_7884), .A3(net_7805), .ZN(net_7804), .A2(net_1592) );
AOI221_X2 inst_9880 ( .B1(net_9787), .B2(net_9098), .A(net_6940), .C2(net_6939), .ZN(net_6819), .C1(net_257) );
DFF_X1 inst_8739 ( .Q(net_9138), .D(net_5729), .CK(net_10676) );
SDFF_X2 inst_516 ( .Q(net_9331), .D(net_9331), .SI(net_9156), .SE(net_7588), .CK(net_13085) );
CLKBUF_X2 inst_12243 ( .A(net_11156), .Z(net_12162) );
OAI211_X2 inst_2258 ( .C1(net_7211), .C2(net_6542), .ZN(net_6425), .B(net_5430), .A(net_3679) );
CLKBUF_X2 inst_13986 ( .A(net_13904), .Z(net_13905) );
CLKBUF_X2 inst_13846 ( .A(net_11994), .Z(net_13765) );
XNOR2_X2 inst_190 ( .ZN(net_5205), .A(net_4582), .B(net_2365) );
AOI22_X2 inst_9602 ( .B1(net_9780), .A2(net_6413), .ZN(net_3466), .B2(net_2462), .A1(net_669) );
OAI22_X2 inst_1267 ( .B1(net_7216), .A2(net_4842), .B2(net_4841), .ZN(net_4806), .A1(net_391) );
NAND2_X2 inst_4103 ( .ZN(net_2385), .A1(net_2143), .A2(net_1650) );
OAI221_X2 inst_1507 ( .B2(net_9063), .C2(net_9056), .ZN(net_7354), .B1(net_7216), .A(net_6994), .C1(net_950) );
CLKBUF_X2 inst_15276 ( .A(net_15194), .Z(net_15195) );
INV_X4 inst_4873 ( .A(net_6192), .ZN(net_3286) );
CLKBUF_X2 inst_13484 ( .A(net_13402), .Z(net_13403) );
AOI221_X2 inst_9932 ( .B2(net_5867), .A(net_5862), .ZN(net_5840), .C1(net_5839), .C2(net_4725), .B1(x3889) );
INV_X2 inst_7301 ( .A(net_9069), .ZN(net_9068) );
INV_X4 inst_6424 ( .ZN(net_1976), .A(net_157) );
OAI211_X2 inst_2062 ( .B(net_7783), .C2(net_7782), .ZN(net_7740), .A(net_7684), .C1(net_2778) );
CLKBUF_X2 inst_15442 ( .A(net_15360), .Z(net_15361) );
NOR4_X2 inst_2350 ( .A4(net_3710), .A2(net_3104), .ZN(net_2967), .A1(net_2626), .A3(net_2625) );
NAND2_X2 inst_3786 ( .ZN(net_4668), .A2(net_4385), .A1(net_3492) );
INV_X2 inst_7260 ( .A(net_9403), .ZN(net_8229) );
CLKBUF_X2 inst_15168 ( .A(net_15086), .Z(net_15087) );
CLKBUF_X2 inst_14960 ( .A(net_14878), .Z(net_14879) );
NAND2_X2 inst_3404 ( .ZN(net_9049), .A2(net_8532), .A1(net_8440) );
DFF_X2 inst_7367 ( .D(net_8754), .QN(net_261), .CK(net_11616) );
SDFF_X2 inst_542 ( .Q(net_9306), .D(net_9306), .SI(net_9157), .SE(net_7553), .CK(net_14043) );
INV_X4 inst_5351 ( .A(net_2257), .ZN(net_1546) );
DFF_X2 inst_7878 ( .Q(net_9946), .D(net_6150), .CK(net_11951) );
XNOR2_X2 inst_128 ( .ZN(net_7483), .A(net_7097), .B(net_2271) );
CLKBUF_X2 inst_13589 ( .A(net_13507), .Z(net_13508) );
CLKBUF_X2 inst_14322 ( .A(net_14240), .Z(net_14241) );
CLKBUF_X2 inst_14172 ( .A(net_13372), .Z(net_14091) );
CLKBUF_X2 inst_13100 ( .A(net_13018), .Z(net_13019) );
CLKBUF_X2 inst_13222 ( .A(net_13140), .Z(net_13141) );
CLKBUF_X2 inst_15363 ( .A(net_15281), .Z(net_15282) );
CLKBUF_X2 inst_15252 ( .A(net_15170), .Z(net_15171) );
CLKBUF_X2 inst_11911 ( .A(net_11829), .Z(net_11830) );
NAND2_X2 inst_4000 ( .ZN(net_3612), .A2(net_3390), .A1(net_664) );
CLKBUF_X2 inst_13625 ( .A(net_12556), .Z(net_13544) );
NAND2_X2 inst_3435 ( .A1(net_9474), .ZN(net_9018), .A2(net_8487) );
INV_X2 inst_6934 ( .A(net_4283), .ZN(net_1930) );
NAND3_X2 inst_3218 ( .A2(net_9218), .ZN(net_6639), .A1(net_5694), .A3(net_3261) );
AOI22_X2 inst_9345 ( .B1(net_9821), .A1(net_6816), .A2(net_5766), .B2(net_5765), .ZN(net_5607) );
OR2_X4 inst_829 ( .A2(net_3914), .ZN(net_1714), .A1(net_648) );
INV_X2 inst_6904 ( .ZN(net_2262), .A(net_2261) );
CLKBUF_X2 inst_15697 ( .A(net_12879), .Z(net_15616) );
DFF_X2 inst_8137 ( .Q(net_9935), .D(net_5121), .CK(net_14282) );
XNOR2_X2 inst_197 ( .ZN(net_5183), .B(net_4921), .A(net_4920) );
INV_X2 inst_7277 ( .ZN(net_9016), .A(net_8378) );
NOR2_X2 inst_2958 ( .A1(net_10459), .ZN(net_2398), .A2(net_612) );
INV_X4 inst_4702 ( .ZN(net_8999), .A(net_4782) );
INV_X4 inst_5723 ( .A(net_963), .ZN(net_884) );
XOR2_X2 inst_24 ( .Z(net_2269), .A(net_1216), .B(net_1194) );
AOI21_X2 inst_10129 ( .A(net_10514), .B1(net_10490), .ZN(net_4442), .B2(net_2825) );
CLKBUF_X2 inst_14866 ( .A(net_14784), .Z(net_14785) );
OAI22_X2 inst_1209 ( .A1(net_7192), .A2(net_5151), .B2(net_5150), .ZN(net_5040), .B1(net_1868) );
CLKBUF_X2 inst_12830 ( .A(net_12530), .Z(net_12749) );
DFF_X2 inst_8190 ( .QN(net_10259), .D(net_5196), .CK(net_12191) );
CLKBUF_X2 inst_11155 ( .A(net_10705), .Z(net_11074) );
DFF_X1 inst_8558 ( .QN(net_9423), .D(net_7398), .CK(net_12664) );
OAI221_X2 inst_1611 ( .B1(net_10207), .C1(net_7136), .B2(net_5642), .ZN(net_5625), .C2(net_4905), .A(net_3507) );
XNOR2_X2 inst_150 ( .ZN(net_6649), .A(net_6648), .B(net_2346) );
INV_X2 inst_6743 ( .ZN(net_6952), .A(net_6951) );
INV_X4 inst_5358 ( .A(net_3546), .ZN(net_1227) );
MUX2_X1 inst_4469 ( .S(net_6041), .A(net_6039), .B(x6252), .Z(x348) );
CLKBUF_X2 inst_12764 ( .A(net_12682), .Z(net_12683) );
INV_X2 inst_6779 ( .ZN(net_6019), .A(net_5832) );
INV_X4 inst_4540 ( .ZN(net_8702), .A(net_8701) );
OR2_X2 inst_887 ( .A2(net_8192), .ZN(net_6161), .A1(net_6160) );
DFF_X1 inst_8730 ( .Q(net_9126), .D(net_6157), .CK(net_10610) );
DFF_X1 inst_8466 ( .Q(net_9596), .D(net_7976), .CK(net_13808) );
INV_X4 inst_5849 ( .ZN(net_1109), .A(net_901) );
INV_X4 inst_5175 ( .ZN(net_3289), .A(net_2279) );
DFF_X2 inst_8036 ( .QN(net_9556), .D(net_9262), .CK(net_12635) );
OAI221_X2 inst_1663 ( .C1(net_7203), .C2(net_5520), .ZN(net_5506), .B2(net_4547), .A(net_3507), .B1(net_1089) );
NOR2_X2 inst_2714 ( .ZN(net_4123), .A2(net_4122), .A1(net_2403) );
CLKBUF_X2 inst_13223 ( .A(net_13141), .Z(net_13142) );
CLKBUF_X2 inst_15630 ( .A(net_14315), .Z(net_15549) );
DFF_X1 inst_8547 ( .Q(net_9982), .D(net_7361), .CK(net_14407) );
INV_X2 inst_7099 ( .ZN(net_1076), .A(net_1075) );
CLKBUF_X2 inst_13647 ( .A(net_13565), .Z(net_13566) );
NAND2_X2 inst_4316 ( .ZN(net_1884), .A1(net_1177), .A2(net_1074) );
NOR4_X2 inst_2357 ( .A3(net_7681), .A4(net_7679), .A1(net_7677), .A2(net_2481), .ZN(net_1421) );
CLKBUF_X2 inst_13036 ( .A(net_12420), .Z(net_12955) );
CLKBUF_X2 inst_13911 ( .A(net_12042), .Z(net_13830) );
INV_X4 inst_6541 ( .A(net_9983), .ZN(net_336) );
DFF_X2 inst_7962 ( .QN(net_10207), .D(net_5625), .CK(net_15590) );
CLKBUF_X2 inst_15730 ( .A(net_15648), .Z(net_15649) );
CLKBUF_X2 inst_12248 ( .A(net_12166), .Z(net_12167) );
OAI21_X2 inst_1961 ( .B1(net_5265), .ZN(net_3568), .A(net_3516), .B2(net_3310) );
CLKBUF_X2 inst_15420 ( .A(net_15338), .Z(net_15339) );
CLKBUF_X2 inst_14343 ( .A(net_14261), .Z(net_14262) );
INV_X4 inst_5799 ( .ZN(net_689), .A(net_688) );
CLKBUF_X2 inst_11285 ( .A(net_10854), .Z(net_11204) );
INV_X4 inst_5954 ( .A(net_1418), .ZN(net_556) );
OAI22_X2 inst_1010 ( .A2(net_8247), .B2(net_8246), .ZN(net_8245), .A1(net_2599), .B1(net_1737) );
CLKBUF_X2 inst_15088 ( .A(net_15006), .Z(net_15007) );
CLKBUF_X2 inst_14928 ( .A(net_14846), .Z(net_14847) );
CLKBUF_X2 inst_10713 ( .A(net_10631), .Z(net_10632) );
DFF_X2 inst_7934 ( .QN(net_10427), .D(net_5544), .CK(net_14605) );
CLKBUF_X2 inst_14939 ( .A(net_12675), .Z(net_14858) );
CLKBUF_X2 inst_14979 ( .A(net_14752), .Z(net_14898) );
OR2_X2 inst_867 ( .ZN(net_7793), .A1(net_7610), .A2(net_7542) );
OR2_X4 inst_820 ( .A1(net_10257), .ZN(net_2146), .A2(net_1013) );
INV_X4 inst_6021 ( .A(net_10028), .ZN(net_805) );
CLKBUF_X2 inst_14179 ( .A(net_14097), .Z(net_14098) );
OAI221_X2 inst_1441 ( .C1(net_9580), .ZN(net_8745), .A(net_8731), .B2(net_8705), .C2(net_8704), .B1(net_2604) );
XNOR2_X2 inst_157 ( .ZN(net_6163), .A(net_5318), .B(net_1105) );
NOR2_X2 inst_2929 ( .ZN(net_2041), .A1(net_645), .A2(net_643) );
CLKBUF_X2 inst_12154 ( .A(net_12072), .Z(net_12073) );
NAND2_X2 inst_3443 ( .A2(net_9449), .ZN(net_8880), .A1(net_8479) );
NAND2_X2 inst_3568 ( .A2(net_7748), .ZN(net_7678), .A1(net_7677) );
INV_X4 inst_6202 ( .ZN(net_3704), .A(net_269) );
INV_X4 inst_6159 ( .A(net_10387), .ZN(net_480) );
NAND2_X2 inst_4287 ( .A2(net_10459), .ZN(net_2334), .A1(net_325) );
CLKBUF_X2 inst_10986 ( .A(net_10707), .Z(net_10905) );
CLKBUF_X2 inst_10760 ( .A(net_10565), .Z(net_10679) );
OAI211_X2 inst_2177 ( .C1(net_7216), .C2(net_6548), .ZN(net_6532), .B(net_5660), .A(net_3527) );
INV_X4 inst_5491 ( .ZN(net_4921), .A(net_995) );
CLKBUF_X2 inst_15449 ( .A(net_11441), .Z(net_15368) );
CLKBUF_X2 inst_12364 ( .A(net_12282), .Z(net_12283) );
AOI22_X2 inst_9342 ( .B1(net_9818), .A2(net_5766), .B2(net_5765), .ZN(net_5610), .A1(net_256) );
AOI22_X2 inst_9588 ( .A1(net_10071), .B1(net_10019), .A2(net_5320), .ZN(net_3572), .B2(net_2468) );
NAND2_X2 inst_4158 ( .ZN(net_2020), .A1(net_2019), .A2(net_1205) );
CLKBUF_X2 inst_11481 ( .A(net_11045), .Z(net_11400) );
DFF_X2 inst_8348 ( .QN(net_10128), .D(net_2795), .CK(net_10799) );
OAI221_X2 inst_1643 ( .C1(net_10426), .B1(net_7186), .ZN(net_5545), .C2(net_4477), .B2(net_4455), .A(net_3731) );
DFF_X2 inst_7447 ( .QN(net_9293), .D(net_8243), .CK(net_15000) );
NAND2_X2 inst_3410 ( .ZN(net_9007), .A1(net_8489), .A2(net_8488) );
INV_X4 inst_4660 ( .ZN(net_6205), .A(net_5955) );
CLKBUF_X2 inst_14537 ( .A(net_12676), .Z(net_14456) );
OAI211_X2 inst_2120 ( .C2(net_6778), .ZN(net_6728), .A(net_6355), .B(net_6090), .C1(net_495) );
NOR2_X2 inst_2678 ( .ZN(net_5365), .A2(net_4758), .A1(net_2752) );
INV_X4 inst_5339 ( .A(net_4601), .ZN(net_1477) );
CLKBUF_X2 inst_13478 ( .A(net_13396), .Z(net_13397) );
CLKBUF_X2 inst_11506 ( .A(net_11424), .Z(net_11425) );
AOI22_X2 inst_9196 ( .A1(net_9886), .B1(net_9787), .B2(net_8041), .A2(net_6141), .ZN(net_6117) );
CLKBUF_X2 inst_15079 ( .A(net_14661), .Z(net_14998) );
CLKBUF_X2 inst_13216 ( .A(net_13134), .Z(net_13135) );
NOR2_X2 inst_2613 ( .A1(net_9073), .ZN(net_7280), .A2(net_6235) );
XOR2_X2 inst_17 ( .Z(net_2789), .B(net_2012), .A(net_1127) );
CLKBUF_X2 inst_15003 ( .A(net_14210), .Z(net_14922) );
AND2_X2 inst_10577 ( .A1(net_9618), .ZN(net_3308), .A2(net_2831) );
AOI21_X2 inst_10105 ( .B1(net_9979), .ZN(net_4875), .A(net_4505), .B2(net_2541) );
INV_X2 inst_7143 ( .A(net_1433), .ZN(net_811) );
XNOR2_X2 inst_249 ( .ZN(net_4121), .B(net_3967), .A(net_3966) );
DFF_X2 inst_7838 ( .Q(net_9923), .D(net_6457), .CK(net_14307) );
CLKBUF_X2 inst_12239 ( .A(net_12157), .Z(net_12158) );
NAND2_X2 inst_3866 ( .ZN(net_4367), .A2(net_4229), .A1(net_4083) );
CLKBUF_X2 inst_12407 ( .A(net_11043), .Z(net_12326) );
OAI211_X2 inst_2234 ( .C1(net_7229), .C2(net_6480), .ZN(net_6470), .B(net_5528), .A(net_3527) );
AND2_X4 inst_10460 ( .A1(net_10157), .ZN(net_1686), .A2(net_1225) );
INV_X4 inst_6251 ( .A(net_10226), .ZN(net_1208) );
DFF_X2 inst_8186 ( .QN(net_9168), .D(net_5007), .CK(net_13551) );
DFF_X2 inst_7976 ( .QN(net_10310), .D(net_5573), .CK(net_14212) );
CLKBUF_X2 inst_14509 ( .A(net_12895), .Z(net_14428) );
NAND2_X2 inst_4371 ( .A2(net_9933), .ZN(net_1137), .A1(net_777) );
INV_X4 inst_5204 ( .ZN(net_4265), .A(net_1530) );
INV_X4 inst_5253 ( .ZN(net_2693), .A(net_1681) );
OAI221_X2 inst_1649 ( .C1(net_10416), .B1(net_7124), .ZN(net_5539), .C2(net_4477), .B2(net_4455), .A(net_3507) );
DFF_X2 inst_7756 ( .Q(net_10405), .D(net_6451), .CK(net_15127) );
OAI221_X2 inst_1480 ( .C2(net_7671), .ZN(net_7604), .B1(net_7602), .A(net_7515), .B2(net_3881), .C1(net_3373) );
CLKBUF_X2 inst_12921 ( .A(net_12839), .Z(net_12840) );
CLKBUF_X2 inst_13594 ( .A(net_12371), .Z(net_13513) );
INV_X4 inst_5815 ( .ZN(net_678), .A(net_677) );
INV_X4 inst_5873 ( .ZN(net_633), .A(net_632) );
CLKBUF_X2 inst_15305 ( .A(net_10695), .Z(net_15224) );
CLKBUF_X2 inst_14121 ( .A(net_14039), .Z(net_14040) );
CLKBUF_X2 inst_10676 ( .A(net_10594), .Z(net_10595) );
CLKBUF_X2 inst_15708 ( .A(net_15626), .Z(net_15627) );
DFF_X1 inst_8697 ( .D(net_6739), .Q(net_148), .CK(net_12591) );
CLKBUF_X2 inst_12359 ( .A(net_11054), .Z(net_12278) );
AND2_X2 inst_10504 ( .A2(net_10378), .ZN(net_5970), .A1(net_1281) );
INV_X4 inst_6472 ( .ZN(net_370), .A(x715) );
DFF_X2 inst_7409 ( .QN(net_9401), .D(net_8364), .CK(net_14028) );
SDFF_X2 inst_669 ( .SI(net_9470), .Q(net_9470), .SE(net_3073), .CK(net_14643), .D(x3249) );
AOI22_X2 inst_9214 ( .A1(net_9907), .B1(net_9808), .A2(net_8042), .B2(net_6120), .ZN(net_6097) );
CLKBUF_X2 inst_13977 ( .A(net_11476), .Z(net_13896) );
CLKBUF_X2 inst_11638 ( .A(net_11556), .Z(net_11557) );
SDFF_X2 inst_664 ( .SI(net_9477), .Q(net_9477), .SE(net_3073), .CK(net_12400), .D(x2826) );
AOI21_X2 inst_10024 ( .B1(net_9364), .A(net_7916), .B2(net_7915), .ZN(net_7855) );
CLKBUF_X2 inst_12485 ( .A(net_12403), .Z(net_12404) );
AND2_X2 inst_10486 ( .A1(net_9560), .ZN(net_8396), .A2(net_8395) );
CLKBUF_X1 inst_8988 ( .A(x185142), .Z(x941) );
CLKBUF_X2 inst_14633 ( .A(net_14551), .Z(net_14552) );
CLKBUF_X2 inst_14262 ( .A(net_14180), .Z(net_14181) );
CLKBUF_X2 inst_14530 ( .A(net_14448), .Z(net_14449) );
AOI221_X2 inst_9911 ( .B1(net_9820), .C1(net_9721), .ZN(net_6448), .A(net_5716), .C2(net_3039), .B2(net_2556) );
AND2_X2 inst_10532 ( .A2(net_3928), .ZN(net_3925), .A1(net_3453) );
DFF_X2 inst_8236 ( .Q(net_10495), .D(net_4886), .CK(net_15212) );
OAI21_X2 inst_1918 ( .ZN(net_4569), .A(net_4148), .B2(net_4147), .B1(net_3984) );
CLKBUF_X2 inst_14500 ( .A(net_12922), .Z(net_14419) );
AOI22_X2 inst_9466 ( .B1(net_9907), .A1(net_9709), .B2(net_4969), .ZN(net_3861), .A2(net_3039) );
CLKBUF_X2 inst_15394 ( .A(net_12914), .Z(net_15313) );
NAND2_X2 inst_4064 ( .ZN(net_7502), .A1(net_2724), .A2(net_2723) );
CLKBUF_X2 inst_15806 ( .A(net_15724), .Z(net_15725) );
MUX2_X2 inst_4427 ( .A(net_9368), .S(net_7635), .Z(net_7596), .B(net_7595) );
CLKBUF_X2 inst_12543 ( .A(net_12461), .Z(net_12462) );
INV_X4 inst_4897 ( .ZN(net_4391), .A(net_2891) );
DFF_X2 inst_7603 ( .Q(net_9349), .D(net_7338), .CK(net_15296) );
INV_X4 inst_4635 ( .ZN(net_7161), .A(net_6589) );
OAI21_X2 inst_1844 ( .ZN(net_5989), .B2(net_5978), .A(net_2072), .B1(net_1368) );
NAND2_X2 inst_3839 ( .ZN(net_4679), .A2(net_4306), .A1(net_1512) );
OAI21_X2 inst_1913 ( .A(net_4680), .ZN(net_4610), .B2(net_4308), .B1(net_2232) );
INV_X4 inst_5209 ( .ZN(net_1822), .A(net_1524) );
DFF_X2 inst_7862 ( .Q(net_10000), .D(net_6269), .CK(net_15598) );
OAI21_X2 inst_1990 ( .ZN(net_2633), .A(net_1739), .B2(net_1570), .B1(net_222) );
NOR3_X2 inst_2368 ( .A3(net_10278), .A2(net_10277), .ZN(net_8260), .A1(net_1874) );
INV_X4 inst_5700 ( .A(net_1143), .ZN(net_791) );
XOR2_X2 inst_36 ( .B(net_9159), .A(net_9158), .Z(net_1726) );
NOR2_X2 inst_2735 ( .ZN(net_4200), .A1(net_3708), .A2(net_3707) );
NOR2_X2 inst_2767 ( .A2(net_3591), .ZN(net_3291), .A1(net_820) );
NOR2_X2 inst_2934 ( .A1(net_10356), .ZN(net_2237), .A2(net_1347) );
OAI222_X2 inst_1370 ( .B2(net_7660), .A2(net_7659), .C2(net_7658), .ZN(net_6273), .B1(net_4936), .A1(net_3523), .C1(net_1806) );
CLKBUF_X2 inst_15805 ( .A(net_15723), .Z(net_15724) );
NOR2_X2 inst_2512 ( .A2(net_8851), .ZN(net_8445), .A1(net_8266) );
CLKBUF_X2 inst_12770 ( .A(net_11359), .Z(net_12689) );
CLKBUF_X2 inst_14658 ( .A(net_14576), .Z(net_14577) );
CLKBUF_X2 inst_12093 ( .A(net_11784), .Z(net_12012) );
CLKBUF_X2 inst_13686 ( .A(net_13604), .Z(net_13605) );
AOI22_X2 inst_9039 ( .A2(net_7175), .ZN(net_7150), .B2(net_3931), .A1(net_3171), .B1(net_1643) );
CLKBUF_X2 inst_11948 ( .A(net_11866), .Z(net_11867) );
AOI22_X2 inst_9652 ( .B2(net_10351), .A2(net_10350), .ZN(net_3149), .B1(net_1285), .A1(net_804) );
CLKBUF_X2 inst_15175 ( .A(net_15093), .Z(net_15094) );
CLKBUF_X2 inst_11447 ( .A(net_11070), .Z(net_11366) );
CLKBUF_X2 inst_13040 ( .A(net_10811), .Z(net_12959) );
CLKBUF_X2 inst_12568 ( .A(net_12486), .Z(net_12487) );
CLKBUF_X2 inst_10721 ( .A(net_10639), .Z(net_10640) );
DFF_X2 inst_7998 ( .QN(net_10230), .D(net_5516), .CK(net_11743) );
NAND2_X2 inst_4124 ( .ZN(net_2328), .A2(net_2233), .A1(net_1619) );
DFF_X2 inst_7954 ( .QN(net_10215), .D(net_5636), .CK(net_15595) );
CLKBUF_X2 inst_13078 ( .A(net_12996), .Z(net_12997) );
CLKBUF_X2 inst_13284 ( .A(net_10686), .Z(net_13203) );
NAND4_X2 inst_3067 ( .ZN(net_5681), .A4(net_4761), .A2(net_3816), .A3(net_3776), .A1(net_3431) );
CLKBUF_X2 inst_13023 ( .A(net_12941), .Z(net_12942) );
CLKBUF_X2 inst_14456 ( .A(net_10656), .Z(net_14375) );
AOI221_X2 inst_9877 ( .B1(net_9784), .B2(net_9098), .A(net_6940), .C2(net_6939), .ZN(net_6824), .C1(net_6823) );
CLKBUF_X2 inst_14740 ( .A(net_11333), .Z(net_14659) );
AOI22_X2 inst_9142 ( .A1(net_9725), .A2(net_6402), .ZN(net_6343), .B2(net_5263), .B1(net_3246) );
CLKBUF_X2 inst_13737 ( .A(net_13655), .Z(net_13656) );
AOI21_X2 inst_10058 ( .ZN(net_7097), .B2(net_6661), .A(net_3201), .B1(net_2305) );
INV_X4 inst_5307 ( .ZN(net_5469), .A(net_1293) );
INV_X4 inst_5672 ( .ZN(net_1295), .A(net_812) );
CLKBUF_X2 inst_13188 ( .A(net_13106), .Z(net_13107) );
AOI211_X2 inst_10273 ( .A(net_7704), .ZN(net_7529), .C1(net_7165), .C2(net_6450), .B(x3390) );
SDFF_X2 inst_676 ( .SI(net_9490), .Q(net_9490), .SE(net_3073), .CK(net_11874), .D(x2027) );
AOI221_X2 inst_9755 ( .ZN(net_7751), .A(net_7749), .B2(net_7748), .C2(net_7747), .C1(net_7685), .B1(net_1993) );
NAND2_X4 inst_3348 ( .ZN(net_8906), .A1(net_8462), .A2(net_8460) );
DFF_X2 inst_7700 ( .Q(net_9803), .D(net_6281), .CK(net_13337) );
DFF_X2 inst_7888 ( .QN(net_10111), .D(net_6028), .CK(net_13268) );
NAND2_X2 inst_4222 ( .A2(net_3885), .ZN(net_1661), .A1(net_1060) );
INV_X4 inst_4848 ( .A(net_7503), .ZN(net_3698) );
CLKBUF_X2 inst_15139 ( .A(net_11729), .Z(net_15058) );
INV_X2 inst_7044 ( .A(net_2404), .ZN(net_1353) );
CLKBUF_X2 inst_11906 ( .A(net_10598), .Z(net_11825) );
INV_X2 inst_6669 ( .ZN(net_8359), .A(net_8302) );
OAI221_X2 inst_1684 ( .B1(net_7198), .ZN(net_5479), .C1(net_5478), .C2(net_4477), .B2(net_4455), .A(net_3527) );
INV_X4 inst_4820 ( .ZN(net_3984), .A(net_3527) );
INV_X4 inst_4859 ( .ZN(net_7649), .A(net_7620) );
CLKBUF_X2 inst_12588 ( .A(net_12506), .Z(net_12507) );
AOI21_X2 inst_10193 ( .ZN(net_3275), .A(net_2839), .B1(net_2629), .B2(net_2136) );
OAI222_X2 inst_1386 ( .B1(net_7665), .A2(net_7664), .C2(net_7663), .ZN(net_5959), .B2(net_5206), .A1(net_4130), .C1(net_1080) );
OAI211_X2 inst_2255 ( .C1(net_7234), .C2(net_6542), .ZN(net_6435), .B(net_5434), .A(net_3679) );
INV_X4 inst_4560 ( .ZN(net_8417), .A(net_8416) );
OAI22_X2 inst_1076 ( .B2(net_10483), .ZN(net_6654), .A2(net_6256), .A1(net_6255), .B1(net_4380) );
XNOR2_X2 inst_217 ( .ZN(net_4682), .B(net_4566), .A(net_4565) );
INV_X4 inst_6360 ( .ZN(net_4641), .A(net_133) );
INV_X4 inst_4852 ( .ZN(net_5370), .A(net_3286) );
INV_X4 inst_6078 ( .A(net_10104), .ZN(net_5825) );
CLKBUF_X2 inst_13292 ( .A(net_13210), .Z(net_13211) );
AOI22_X2 inst_9264 ( .A1(net_9076), .ZN(net_5810), .A2(net_5809), .B2(net_5808), .B1(net_807) );
OAI21_X2 inst_2000 ( .ZN(net_2297), .A(net_2296), .B1(net_2295), .B2(net_2294) );
INV_X4 inst_4616 ( .A(net_7506), .ZN(net_7489) );
NAND2_X2 inst_3748 ( .ZN(net_5302), .A2(net_5292), .A1(net_4476) );
AOI221_X2 inst_9816 ( .B1(net_9874), .B2(net_9101), .ZN(net_6947), .A(net_6945), .C1(net_6944), .C2(net_245) );
INV_X2 inst_6732 ( .ZN(net_7543), .A(net_7482) );
AOI21_X2 inst_10223 ( .ZN(net_2801), .B1(net_2299), .B2(net_2043), .A(net_1173) );
OAI211_X2 inst_2213 ( .C1(net_7219), .C2(net_6501), .ZN(net_6492), .B(net_5551), .A(net_3527) );
OAI22_X2 inst_1195 ( .A1(net_7136), .A2(net_5134), .B2(net_5133), .ZN(net_5058), .B1(net_1788) );
INV_X4 inst_6222 ( .A(net_10106), .ZN(net_5861) );
SDFF_X2 inst_672 ( .SI(net_9478), .Q(net_9478), .SE(net_3073), .CK(net_14639), .D(x2767) );
CLKBUF_X2 inst_15393 ( .A(net_14878), .Z(net_15312) );
OAI221_X2 inst_1471 ( .ZN(net_7800), .A(net_7797), .C2(net_6841), .B2(net_6619), .B1(net_5385), .C1(net_4799) );
AOI222_X1 inst_9699 ( .B1(net_9506), .A2(net_8295), .B2(net_8294), .C2(net_8293), .ZN(net_8279), .C1(net_8214), .A1(x3133) );
AOI22_X2 inst_9610 ( .A1(net_10073), .B1(net_10024), .A2(net_5319), .B2(net_5174), .ZN(net_3443) );
CLKBUF_X2 inst_12252 ( .A(net_12004), .Z(net_12171) );
NAND2_X2 inst_3826 ( .ZN(net_9074), .A2(net_4189), .A1(net_4030) );
CLKBUF_X2 inst_11829 ( .A(net_11075), .Z(net_11748) );
INV_X4 inst_6471 ( .ZN(net_578), .A(net_169) );
DFF_X2 inst_7523 ( .Q(net_9531), .D(net_7835), .CK(net_13985) );
OAI221_X2 inst_1525 ( .ZN(net_7279), .B2(net_7278), .C1(net_7277), .C2(net_7276), .A(net_6650), .B1(net_6228) );
INV_X2 inst_6839 ( .ZN(net_3871), .A(net_3870) );
NAND3_X2 inst_3230 ( .ZN(net_4952), .A1(net_4951), .A3(net_4950), .A2(net_2034) );
CLKBUF_X2 inst_11820 ( .A(net_11391), .Z(net_11739) );
OAI211_X2 inst_2248 ( .C1(net_7213), .C2(net_6480), .ZN(net_6456), .B(net_5647), .A(net_3679) );
NOR3_X2 inst_2453 ( .A3(net_9184), .A2(net_9182), .ZN(net_2151), .A1(net_2150) );
OAI22_X2 inst_1312 ( .B2(net_10043), .ZN(net_2286), .A1(net_2285), .A2(net_2284), .B1(net_2283) );
AOI22_X2 inst_9538 ( .B1(net_9781), .A1(net_9714), .ZN(net_3783), .A2(net_3039), .B2(net_2462) );
NAND3_X2 inst_3281 ( .A2(net_9111), .ZN(net_6669), .A1(net_3625), .A3(net_3624) );
OR3_X4 inst_703 ( .ZN(net_5375), .A2(net_4103), .A1(net_4097), .A3(net_3640) );
CLKBUF_X2 inst_11125 ( .A(net_11043), .Z(net_11044) );
AOI22_X2 inst_9474 ( .B1(net_9911), .A1(net_9713), .B2(net_4969), .ZN(net_3849), .A2(net_3039) );
NOR2_X2 inst_2546 ( .ZN(net_8108), .A2(net_8046), .A1(net_6192) );
CLKBUF_X2 inst_15145 ( .A(net_15063), .Z(net_15064) );
INV_X2 inst_7177 ( .A(net_9406), .ZN(net_8227) );
CLKBUF_X2 inst_11112 ( .A(net_11030), .Z(net_11031) );
AOI221_X2 inst_9882 ( .B1(net_9789), .B2(net_9098), .A(net_6940), .C2(net_6939), .ZN(net_6817), .C1(net_6816) );
INV_X4 inst_4693 ( .ZN(net_4834), .A(net_4650) );
CLKBUF_X2 inst_12504 ( .A(net_12422), .Z(net_12423) );
CLKBUF_X2 inst_15737 ( .A(net_11585), .Z(net_15656) );
AND2_X4 inst_10449 ( .A1(net_10262), .ZN(net_1530), .A2(net_1382) );
CLKBUF_X2 inst_14786 ( .A(net_14704), .Z(net_14705) );
CLKBUF_X2 inst_14289 ( .A(net_14207), .Z(net_14208) );
INV_X4 inst_5785 ( .ZN(net_813), .A(net_699) );
NAND2_X2 inst_3419 ( .ZN(net_9024), .A2(net_9023), .A1(net_9022) );
CLKBUF_X2 inst_12966 ( .A(net_11511), .Z(net_12885) );
OAI22_X2 inst_1067 ( .A2(net_7036), .B2(net_7035), .ZN(net_6962), .A1(net_3031), .B1(net_736) );
INV_X4 inst_6539 ( .A(net_9935), .ZN(net_338) );
CLKBUF_X2 inst_11970 ( .A(net_10652), .Z(net_11889) );
INV_X4 inst_4787 ( .ZN(net_4187), .A(net_4021) );
DFF_X2 inst_7411 ( .QN(net_9403), .D(net_8362), .CK(net_13956) );
CLKBUF_X2 inst_13749 ( .A(net_13667), .Z(net_13668) );
AOI222_X1 inst_9735 ( .B2(net_10401), .C2(net_10400), .A2(net_10399), .B1(net_10394), .C1(net_10393), .A1(net_10392), .ZN(net_1445) );
DFF_X1 inst_8406 ( .D(net_8815), .CK(net_14206), .Q(x637) );
AOI22_X2 inst_9231 ( .A1(net_9895), .B1(net_9796), .B2(net_6129), .A2(net_6109), .ZN(net_6080) );
INV_X4 inst_4951 ( .ZN(net_2561), .A(net_2560) );
CLKBUF_X2 inst_14954 ( .A(net_14815), .Z(net_14873) );
OAI21_X2 inst_1824 ( .B1(net_7157), .ZN(net_6569), .A(net_5925), .B2(net_5897) );
OAI22_X2 inst_1214 ( .A1(net_7190), .A2(net_5134), .B2(net_5133), .ZN(net_5035), .B1(net_3533) );
CLKBUF_X2 inst_15151 ( .A(net_15069), .Z(net_15070) );
DFF_X2 inst_8121 ( .Q(net_9742), .D(net_5145), .CK(net_12027) );
OAI22_X4 inst_971 ( .B2(net_8968), .ZN(net_8431), .A2(net_8430), .B1(net_8429), .A1(net_8429) );
OAI222_X2 inst_1417 ( .B2(net_7665), .A2(net_7664), .C2(net_7663), .ZN(net_5193), .B1(net_2978), .A1(net_2015), .C1(net_1257) );
OAI22_X2 inst_1219 ( .A1(net_7129), .A2(net_5139), .B2(net_5138), .ZN(net_5029), .B1(net_2574) );
CLKBUF_X2 inst_11103 ( .A(net_11021), .Z(net_11022) );
DFF_X2 inst_8018 ( .QN(net_10329), .D(net_5483), .CK(net_12128) );
NAND2_X2 inst_3459 ( .A1(net_9498), .A2(net_8473), .ZN(net_8465) );
CLKBUF_X2 inst_11887 ( .A(net_11805), .Z(net_11806) );
INV_X8 inst_4488 ( .ZN(net_8047), .A(net_7989) );
DFF_X2 inst_7633 ( .D(net_6760), .QN(net_123), .CK(net_12826) );
CLKBUF_X2 inst_15357 ( .A(net_15275), .Z(net_15276) );
NAND2_X4 inst_3335 ( .ZN(net_8941), .A2(net_8882), .A1(net_8881) );
NAND4_X2 inst_3073 ( .ZN(net_5197), .A4(net_4504), .A2(net_3841), .A1(net_3582), .A3(net_3439) );
CLKBUF_X2 inst_12716 ( .A(net_12634), .Z(net_12635) );
CLKBUF_X2 inst_11732 ( .A(net_11404), .Z(net_11651) );
CLKBUF_X2 inst_11741 ( .A(net_11659), .Z(net_11660) );
OAI21_X2 inst_1980 ( .ZN(net_2940), .A(net_2688), .B1(net_1850), .B2(net_680) );
AND2_X2 inst_10488 ( .ZN(net_8133), .A1(net_8132), .A2(net_8094) );
CLKBUF_X2 inst_15123 ( .A(net_13080), .Z(net_15042) );
INV_X4 inst_5868 ( .ZN(net_3739), .A(net_1507) );
AOI22_X2 inst_9454 ( .A1(net_6892), .B2(net_6625), .ZN(net_6433), .B1(net_3976), .A2(net_2817) );
AOI22_X2 inst_9325 ( .B1(net_9893), .A1(net_6828), .A2(net_5759), .B2(net_5758), .ZN(net_5651) );
NOR2_X2 inst_2885 ( .A1(net_2134), .ZN(net_1799), .A2(net_1798) );
INV_X2 inst_7222 ( .A(net_9324), .ZN(net_430) );
CLKBUF_X2 inst_12628 ( .A(net_12546), .Z(net_12547) );
AND2_X4 inst_10446 ( .A2(net_9195), .ZN(net_2445), .A1(net_1461) );
OAI211_X2 inst_2221 ( .C1(net_7190), .C2(net_6501), .ZN(net_6484), .B(net_5533), .A(net_3679) );
NOR2_X2 inst_2632 ( .A1(net_9219), .ZN(net_5928), .A2(net_5927) );
INV_X4 inst_4795 ( .ZN(net_3667), .A(net_3666) );
CLKBUF_X2 inst_12991 ( .A(net_12909), .Z(net_12910) );
OAI211_X2 inst_2082 ( .C2(net_6778), .ZN(net_6766), .A(net_6393), .B(net_6137), .C1(net_378) );
CLKBUF_X2 inst_12469 ( .A(net_12387), .Z(net_12388) );
INV_X4 inst_5842 ( .ZN(net_7562), .A(net_652) );
CLKBUF_X2 inst_15028 ( .A(net_14946), .Z(net_14947) );
AOI21_X2 inst_10135 ( .ZN(net_4251), .B2(net_3622), .B1(net_3283), .A(net_2104) );
NAND3_X2 inst_3286 ( .ZN(net_3110), .A3(net_2351), .A1(net_2052), .A2(net_1780) );
CLKBUF_X2 inst_15299 ( .A(net_15217), .Z(net_15218) );
CLKBUF_X2 inst_12907 ( .A(net_12825), .Z(net_12826) );
NAND2_X2 inst_4225 ( .A1(net_8687), .ZN(net_1655), .A2(net_115) );
INV_X4 inst_5625 ( .A(net_10435), .ZN(net_1637) );
CLKBUF_X2 inst_11371 ( .A(net_11097), .Z(net_11290) );
CLKBUF_X2 inst_11421 ( .A(net_11339), .Z(net_11340) );
AOI22_X2 inst_9533 ( .B1(net_10294), .A1(net_10189), .B2(net_4774), .A2(net_4217), .ZN(net_3788) );
NAND2_X2 inst_4141 ( .A1(net_4125), .ZN(net_2153), .A2(net_2150) );
CLKBUF_X2 inst_13004 ( .A(net_12922), .Z(net_12923) );
CLKBUF_X2 inst_14293 ( .A(net_14211), .Z(net_14212) );
OR3_X4 inst_692 ( .ZN(net_6501), .A1(net_5171), .A3(net_4789), .A2(net_4629) );
INV_X4 inst_4591 ( .A(net_8018), .ZN(net_8010) );
INV_X2 inst_6800 ( .ZN(net_5371), .A(net_5201) );
CLKBUF_X2 inst_14819 ( .A(net_14737), .Z(net_14738) );
INV_X2 inst_6897 ( .ZN(net_2584), .A(net_2583) );
OAI221_X2 inst_1517 ( .C1(net_10420), .B2(net_9063), .C2(net_9056), .ZN(net_7317), .B1(net_7127), .A(net_7063) );
INV_X4 inst_5318 ( .A(net_6311), .ZN(net_1278) );
AND2_X2 inst_10529 ( .ZN(net_3930), .A2(net_3928), .A1(net_3457) );
XNOR2_X2 inst_70 ( .ZN(net_8703), .A(net_8682), .B(net_2929) );
INV_X4 inst_5480 ( .A(net_7504), .ZN(net_1001) );
INV_X2 inst_6915 ( .A(net_2528), .ZN(net_2176) );
DFF_X2 inst_7587 ( .QN(net_9235), .D(net_7467), .CK(net_11256) );
DFF_X2 inst_7672 ( .D(net_6766), .QN(net_118), .CK(net_14319) );
CLKBUF_X2 inst_15662 ( .A(net_15580), .Z(net_15581) );
CLKBUF_X2 inst_12493 ( .A(net_11149), .Z(net_12412) );
AOI221_X2 inst_9865 ( .A(net_6889), .B2(net_6888), .C2(net_6887), .ZN(net_6851), .B1(net_2129), .C1(x4587) );
AOI22_X2 inst_9162 ( .A2(net_6402), .ZN(net_6312), .A1(net_6311), .B2(net_5263), .B1(net_1466) );
CLKBUF_X2 inst_14161 ( .A(net_14079), .Z(net_14080) );
CLKBUF_X2 inst_11290 ( .A(net_11208), .Z(net_11209) );
XNOR2_X2 inst_188 ( .ZN(net_5207), .A(net_4559), .B(net_2030) );
INV_X8 inst_4528 ( .A(net_9052), .ZN(net_9050) );
CLKBUF_X2 inst_13534 ( .A(net_13452), .Z(net_13453) );
NAND2_X2 inst_3768 ( .ZN(net_4972), .A2(net_4576), .A1(net_965) );
INV_X4 inst_6028 ( .ZN(net_7129), .A(x5548) );
INV_X4 inst_6093 ( .A(net_9565), .ZN(net_3365) );
CLKBUF_X2 inst_14586 ( .A(net_14504), .Z(net_14505) );
NAND2_X2 inst_4207 ( .A1(net_4017), .ZN(net_2904), .A2(net_1384) );
AOI22_X2 inst_9058 ( .B1(net_9679), .A2(net_6684), .B2(net_6683), .ZN(net_6608), .A1(net_248) );
CLKBUF_X2 inst_11308 ( .A(net_11226), .Z(net_11227) );
NOR2_X2 inst_3011 ( .ZN(net_1545), .A1(net_493), .A2(net_351) );
INV_X4 inst_6218 ( .ZN(net_4273), .A(net_270) );
CLKBUF_X2 inst_13306 ( .A(net_13100), .Z(net_13225) );
NOR2_X2 inst_2848 ( .A2(net_5983), .ZN(net_3720), .A1(net_2257) );
CLKBUF_X2 inst_15181 ( .A(net_11544), .Z(net_15100) );
CLKBUF_X2 inst_12686 ( .A(net_12604), .Z(net_12605) );
INV_X4 inst_4826 ( .ZN(net_7832), .A(net_5370) );
INV_X2 inst_6695 ( .ZN(net_8254), .A(net_8253) );
OAI221_X2 inst_1537 ( .B2(net_9047), .C2(net_7287), .ZN(net_7230), .C1(net_7229), .A(net_6795), .B1(net_5482) );
OAI211_X2 inst_2041 ( .C2(net_8102), .B(net_8098), .ZN(net_8045), .A(net_7944), .C1(net_5403) );
CLKBUF_X2 inst_13866 ( .A(net_13784), .Z(net_13785) );
INV_X4 inst_6323 ( .A(net_9984), .ZN(net_418) );
INV_X4 inst_5235 ( .ZN(net_1925), .A(net_1482) );
NAND2_X2 inst_3593 ( .ZN(net_7299), .A2(net_6861), .A1(net_6599) );
CLKBUF_X2 inst_15509 ( .A(net_15427), .Z(net_15428) );
DFF_X1 inst_8529 ( .Q(net_9969), .D(net_7317), .CK(net_13382) );
INV_X4 inst_4589 ( .ZN(net_8074), .A(net_8033) );
NAND3_X2 inst_3176 ( .A3(net_9560), .A2(net_9559), .ZN(net_8989), .A1(net_8386) );
DFF_X2 inst_7509 ( .QN(net_9376), .D(net_7938), .CK(net_14172) );
INV_X2 inst_6768 ( .ZN(net_6034), .A(net_5863) );
CLKBUF_X2 inst_11550 ( .A(net_11231), .Z(net_11469) );
CLKBUF_X2 inst_14830 ( .A(net_11168), .Z(net_14749) );
NAND2_X4 inst_3325 ( .ZN(net_9042), .A2(net_8608), .A1(net_8607) );
CLKBUF_X2 inst_13393 ( .A(net_13311), .Z(net_13312) );
CLKBUF_X2 inst_11145 ( .A(net_11063), .Z(net_11064) );
CLKBUF_X2 inst_11085 ( .A(net_11003), .Z(net_11004) );
AOI22_X2 inst_9083 ( .A2(net_6420), .ZN(net_6412), .B2(net_5263), .A1(net_1767), .B1(net_432) );
CLKBUF_X2 inst_13991 ( .A(net_13909), .Z(net_13910) );
CLKBUF_X2 inst_13889 ( .A(net_13807), .Z(net_13808) );
CLKBUF_X2 inst_12655 ( .A(net_12038), .Z(net_12574) );
NAND2_X2 inst_4168 ( .A1(net_9534), .ZN(net_7546), .A2(net_4788) );
XNOR2_X2 inst_195 ( .ZN(net_5192), .A(net_4546), .B(net_1808) );
CLKBUF_X2 inst_11835 ( .A(net_11714), .Z(net_11754) );
CLKBUF_X2 inst_12839 ( .A(net_12757), .Z(net_12758) );
OAI21_X2 inst_1987 ( .A(net_2792), .ZN(net_2740), .B2(net_2739), .B1(net_2719) );
CLKBUF_X2 inst_13730 ( .A(net_13648), .Z(net_13649) );
CLKBUF_X2 inst_10821 ( .A(net_10597), .Z(net_10740) );
CLKBUF_X2 inst_13418 ( .A(net_13336), .Z(net_13337) );
OAI22_X2 inst_1150 ( .A1(net_7229), .A2(net_5134), .B2(net_5133), .ZN(net_5123), .B1(net_453) );
DFF_X2 inst_7685 ( .Q(net_10069), .D(net_6567), .CK(net_10834) );
CLKBUF_X2 inst_14372 ( .A(net_14290), .Z(net_14291) );
INV_X4 inst_4914 ( .ZN(net_2799), .A(net_2798) );
CLKBUF_X2 inst_11355 ( .A(net_10658), .Z(net_11274) );
CLKBUF_X2 inst_11020 ( .A(net_10864), .Z(net_10939) );
INV_X4 inst_5605 ( .A(net_10473), .ZN(net_2625) );
INV_X2 inst_7070 ( .A(net_2005), .ZN(net_1237) );
INV_X2 inst_7106 ( .A(net_1817), .ZN(net_1022) );
INV_X4 inst_4780 ( .ZN(net_4135), .A(net_3298) );
CLKBUF_X2 inst_12981 ( .A(net_10557), .Z(net_12900) );
CLKBUF_X2 inst_15468 ( .A(net_15386), .Z(net_15387) );
CLKBUF_X2 inst_11770 ( .A(net_11688), .Z(net_11689) );
INV_X4 inst_4658 ( .A(net_9260), .ZN(net_6231) );
INV_X4 inst_5916 ( .A(net_606), .ZN(net_588) );
INV_X2 inst_7154 ( .A(net_2628), .ZN(net_713) );
DFF_X1 inst_8715 ( .QN(net_9207), .D(net_6580), .CK(net_11354) );
OAI221_X2 inst_1589 ( .B2(net_10271), .B1(net_6044), .ZN(net_5985), .A(net_5223), .C2(net_5218), .C1(net_4244) );
CLKBUF_X2 inst_11994 ( .A(net_11912), .Z(net_11913) );
INV_X4 inst_4535 ( .ZN(net_8749), .A(net_8746) );
CLKBUF_X2 inst_14114 ( .A(net_11106), .Z(net_14033) );
INV_X4 inst_5607 ( .ZN(net_2294), .A(net_2275) );
CLKBUF_X2 inst_14810 ( .A(net_14728), .Z(net_14729) );
CLKBUF_X2 inst_14095 ( .A(net_14013), .Z(net_14014) );
INV_X8 inst_4499 ( .ZN(net_6140), .A(net_5298) );
CLKBUF_X2 inst_12852 ( .A(net_12770), .Z(net_12771) );
CLKBUF_X2 inst_15263 ( .A(net_12872), .Z(net_15182) );
CLKBUF_X2 inst_10979 ( .A(net_10897), .Z(net_10898) );
INV_X2 inst_6825 ( .A(net_7602), .ZN(net_4186) );
DFF_X1 inst_8704 ( .Q(net_9148), .D(net_6782), .CK(net_10703) );
CLKBUF_X2 inst_15160 ( .A(net_15078), .Z(net_15079) );
XNOR2_X2 inst_335 ( .ZN(net_2979), .B(net_2491), .A(net_2327) );
CLKBUF_X2 inst_15244 ( .A(net_11993), .Z(net_15163) );
CLKBUF_X2 inst_12783 ( .A(net_11366), .Z(net_12702) );
CLKBUF_X2 inst_12827 ( .A(net_12745), .Z(net_12746) );
INV_X4 inst_5508 ( .ZN(net_3546), .A(net_1332) );
CLKBUF_X2 inst_12661 ( .A(net_12579), .Z(net_12580) );
CLKBUF_X2 inst_14406 ( .A(net_12872), .Z(net_14325) );
DFF_X1 inst_8611 ( .Q(net_9777), .D(net_7187), .CK(net_15463) );
SDFF_X2 inst_658 ( .SI(net_9491), .Q(net_9491), .SE(net_3073), .CK(net_12416), .D(x1974) );
INV_X4 inst_6190 ( .A(net_9738), .ZN(net_471) );
INV_X2 inst_6862 ( .A(net_3423), .ZN(net_3280) );
DFF_X1 inst_8420 ( .D(net_8774), .Q(net_247), .CK(net_14871) );
DFF_X2 inst_7779 ( .Q(net_9812), .D(net_6521), .CK(net_14231) );
CLKBUF_X2 inst_12192 ( .A(net_12110), .Z(net_12111) );
AOI22_X2 inst_9336 ( .B1(net_9812), .A2(net_5766), .B2(net_5765), .ZN(net_5616), .A1(net_250) );
INV_X8 inst_4520 ( .ZN(net_8924), .A(net_7608) );
CLKBUF_X2 inst_11562 ( .A(net_11480), .Z(net_11481) );
INV_X2 inst_7227 ( .A(net_9557), .ZN(net_8093) );
CLKBUF_X2 inst_14045 ( .A(net_10616), .Z(net_13964) );
CLKBUF_X2 inst_14276 ( .A(net_14194), .Z(net_14195) );
XNOR2_X2 inst_438 ( .B(net_9305), .ZN(net_1042), .A(net_213) );
CLKBUF_X2 inst_13311 ( .A(net_13229), .Z(net_13230) );
INV_X1 inst_7326 ( .A(net_9103), .ZN(net_9102) );
INV_X4 inst_6351 ( .ZN(net_1728), .A(x6401) );
CLKBUF_X2 inst_15090 ( .A(net_15008), .Z(net_15009) );
CLKBUF_X2 inst_10769 ( .A(net_10609), .Z(net_10688) );
AOI22_X2 inst_9626 ( .B1(net_9996), .A2(net_4694), .ZN(net_3421), .B2(net_2468), .A1(net_229) );
CLKBUF_X2 inst_14336 ( .A(net_14254), .Z(net_14255) );
AOI222_X1 inst_9692 ( .B1(net_9509), .A2(net_8301), .B2(net_8300), .C2(net_8299), .ZN(net_8289), .C1(net_8195), .A1(x1974) );
CLKBUF_X2 inst_11391 ( .A(net_11187), .Z(net_11310) );
XNOR2_X2 inst_324 ( .B(net_9618), .ZN(net_3029), .A(net_2831) );
CLKBUF_X2 inst_11640 ( .A(net_10555), .Z(net_11559) );
NAND2_X2 inst_3550 ( .A1(net_10509), .ZN(net_7874), .A2(net_7869) );
INV_X4 inst_6046 ( .ZN(net_7243), .A(x6028) );
NAND2_X2 inst_4083 ( .A1(net_5420), .ZN(net_3559), .A2(net_2871) );
CLKBUF_X2 inst_13581 ( .A(net_12242), .Z(net_13500) );
XOR2_X2 inst_43 ( .Z(net_2448), .B(net_666), .A(net_458) );
OAI211_X2 inst_2128 ( .C2(net_6778), .ZN(net_6720), .A(net_6419), .B(net_6139), .C1(net_548) );
INV_X4 inst_5936 ( .ZN(net_979), .A(net_851) );
OAI221_X2 inst_1707 ( .ZN(net_4379), .C1(net_4378), .B2(net_3597), .C2(net_3596), .B1(net_2851), .A(net_2550) );
INV_X2 inst_7213 ( .A(net_9391), .ZN(net_8214) );
INV_X2 inst_6715 ( .ZN(net_7941), .A(net_7917) );
AND2_X4 inst_10452 ( .A1(net_10367), .ZN(net_1674), .A2(net_1379) );
DFF_X2 inst_8115 ( .QN(net_9515), .D(net_5408), .CK(net_12729) );
XNOR2_X2 inst_375 ( .ZN(net_3955), .A(net_2473), .B(net_2472) );
CLKBUF_X2 inst_11241 ( .A(net_11159), .Z(net_11160) );
AOI221_X2 inst_9959 ( .C1(net_10500), .B1(net_10290), .C2(net_6415), .B2(net_4774), .ZN(net_4772), .A(net_4343) );
DFF_X1 inst_8606 ( .Q(net_9864), .D(net_7236), .CK(net_13466) );
NAND2_X2 inst_3490 ( .A1(net_8967), .ZN(net_8331), .A2(net_8239) );
CLKBUF_X2 inst_14472 ( .A(net_10669), .Z(net_14391) );
DFF_X2 inst_7384 ( .D(net_8655), .QN(net_271), .CK(net_12644) );
INV_X2 inst_7039 ( .A(net_2465), .ZN(net_1763) );
CLKBUF_X2 inst_15780 ( .A(net_15698), .Z(net_15699) );
CLKBUF_X2 inst_10933 ( .A(net_10851), .Z(net_10852) );
AOI21_X2 inst_10086 ( .B2(net_10094), .B1(net_10093), .ZN(net_5898), .A(net_5329) );
XNOR2_X2 inst_285 ( .ZN(net_3642), .B(net_3641), .A(net_2997) );
INV_X2 inst_7215 ( .A(net_9514), .ZN(net_448) );
OAI21_X2 inst_1830 ( .B1(net_7157), .ZN(net_6452), .B2(net_5693), .A(net_5537) );
AOI221_X2 inst_9887 ( .B1(net_9764), .B2(net_9098), .A(net_6940), .C2(net_6939), .ZN(net_6809), .C1(net_6808) );
CLKBUF_X2 inst_11780 ( .A(net_11141), .Z(net_11699) );
CLKBUF_X2 inst_11385 ( .A(net_11303), .Z(net_11304) );
AOI22_X2 inst_9313 ( .B1(net_9718), .A1(net_6821), .A2(net_5755), .B2(net_5754), .ZN(net_5664) );
DFF_X2 inst_8289 ( .Q(net_9753), .D(net_4738), .CK(net_14506) );
INV_X4 inst_5563 ( .ZN(net_1230), .A(net_936) );
OAI221_X2 inst_1563 ( .C1(net_10203), .C2(net_7295), .B2(net_7293), .ZN(net_7191), .B1(net_7190), .A(net_6809) );
INV_X4 inst_6363 ( .ZN(net_5798), .A(net_274) );
CLKBUF_X2 inst_10833 ( .A(net_10751), .Z(net_10752) );
CLKBUF_X2 inst_11402 ( .A(net_11227), .Z(net_11321) );
MUX2_X1 inst_4455 ( .S(net_6041), .A(net_291), .B(x5498), .Z(x198) );
DFF_X2 inst_7911 ( .Q(net_9223), .D(net_5942), .CK(net_13016) );
NAND3_X2 inst_3242 ( .ZN(net_4703), .A3(net_4584), .A1(net_4583), .A2(net_2701) );
DFF_X2 inst_7398 ( .D(net_8544), .Q(net_220), .CK(net_14614) );
CLKBUF_X2 inst_10638 ( .A(net_10556), .Z(net_10557) );
DFF_X2 inst_7907 ( .QN(net_10474), .D(net_5869), .CK(net_11393) );
AOI221_X2 inst_9895 ( .B1(net_9880), .B2(net_9101), .A(net_6945), .C2(net_6944), .ZN(net_6799), .C1(net_251) );
OR2_X2 inst_929 ( .A1(net_9105), .ZN(net_4077), .A2(net_2948) );
OAI22_X2 inst_982 ( .A2(net_8962), .B2(net_8659), .ZN(net_8658), .A1(net_6434), .B1(net_6230) );
NAND4_X2 inst_3138 ( .ZN(net_3450), .A3(net_2710), .A4(net_2709), .A1(net_2437), .A2(net_1519) );
OAI222_X2 inst_1397 ( .A2(net_7728), .C2(net_7727), .B2(net_7726), .ZN(net_5701), .A1(net_2885), .B1(net_1805), .C1(net_1490) );
CLKBUF_X2 inst_10864 ( .A(net_10604), .Z(net_10783) );
XNOR2_X2 inst_299 ( .B(net_9619), .ZN(net_3330), .A(net_3308) );
CLKBUF_X2 inst_13871 ( .A(net_13789), .Z(net_13790) );
AND2_X2 inst_10567 ( .A1(net_9205), .ZN(net_3513), .A2(net_3022) );
DFF_X2 inst_7656 ( .D(net_6694), .QN(net_188), .CK(net_12986) );
OAI21_X2 inst_1798 ( .B1(net_8012), .ZN(net_7444), .A(net_6979), .B2(net_6971) );
NOR2_X2 inst_2927 ( .A2(net_9062), .A1(net_8955), .ZN(net_8914) );
CLKBUF_X2 inst_13115 ( .A(net_13033), .Z(net_13034) );
NAND3_X2 inst_3303 ( .ZN(net_2175), .A2(net_2174), .A1(net_1699), .A3(net_1638) );
AND4_X4 inst_10336 ( .A2(net_10478), .ZN(net_2966), .A1(net_2715), .A4(net_1667), .A3(net_998) );
INV_X4 inst_6181 ( .A(net_10288), .ZN(net_474) );
CLKBUF_X2 inst_12938 ( .A(net_12033), .Z(net_12857) );
INV_X4 inst_5853 ( .A(net_739), .ZN(net_645) );
AND3_X2 inst_10383 ( .ZN(net_874), .A2(net_112), .A3(net_111), .A1(net_107) );
DFF_X1 inst_8727 ( .Q(net_9648), .D(net_5965), .CK(net_12830) );
NOR2_X2 inst_2760 ( .A1(net_9613), .ZN(net_3517), .A2(net_3029) );
OAI21_X2 inst_1938 ( .B2(net_5347), .A(net_4625), .ZN(net_4461), .B1(net_4360) );
INV_X4 inst_6478 ( .A(net_9988), .ZN(net_366) );
INV_X4 inst_6452 ( .A(net_10112), .ZN(net_5847) );
CLKBUF_X2 inst_11870 ( .A(net_11788), .Z(net_11789) );
CLKBUF_X2 inst_15213 ( .A(net_12321), .Z(net_15132) );
AOI22_X2 inst_9435 ( .A1(net_9853), .B1(net_6808), .ZN(net_4492), .A2(net_4491), .B2(net_4490) );
INV_X2 inst_7098 ( .A(net_2627), .ZN(net_1080) );
INV_X2 inst_6888 ( .A(net_3347), .ZN(net_2718) );
OAI211_X2 inst_2095 ( .C2(net_6778), .ZN(net_6753), .A(net_6410), .B(net_6074), .C1(net_5098) );
CLKBUF_X2 inst_15659 ( .A(net_15577), .Z(net_15578) );
INV_X4 inst_6288 ( .A(net_9652), .ZN(net_436) );
INV_X2 inst_7030 ( .A(net_10456), .ZN(net_1473) );
CLKBUF_X2 inst_15581 ( .A(net_15499), .Z(net_15500) );
INV_X4 inst_5129 ( .ZN(net_2527), .A(net_2131) );
CLKBUF_X2 inst_13524 ( .A(net_13442), .Z(net_13443) );
INV_X4 inst_5794 ( .ZN(net_3261), .A(net_2758) );
CLKBUF_X2 inst_14841 ( .A(net_14759), .Z(net_14760) );
CLKBUF_X2 inst_14103 ( .A(net_14021), .Z(net_14022) );
CLKBUF_X2 inst_10656 ( .A(net_10545), .Z(net_10575) );
INV_X4 inst_4995 ( .ZN(net_2569), .A(net_1584) );
INV_X4 inst_5652 ( .A(net_10514), .ZN(net_1498) );
NAND3_X2 inst_3260 ( .ZN(net_4437), .A1(net_4436), .A3(net_4435), .A2(net_2209) );
DFF_X2 inst_8262 ( .Q(net_10289), .D(net_4819), .CK(net_14516) );
NAND4_X2 inst_3158 ( .A4(net_1790), .ZN(net_1769), .A3(net_1029), .A1(net_1023), .A2(net_781) );
NAND2_X2 inst_4190 ( .ZN(net_1853), .A2(net_1852), .A1(net_1171) );
CLKBUF_X2 inst_13894 ( .A(net_11394), .Z(net_13813) );
CLKBUF_X2 inst_11248 ( .A(net_11166), .Z(net_11167) );
INV_X4 inst_5387 ( .A(net_5164), .ZN(net_1592) );
CLKBUF_X2 inst_14067 ( .A(net_13815), .Z(net_13986) );
CLKBUF_X2 inst_11813 ( .A(net_11731), .Z(net_11732) );
OR4_X4 inst_683 ( .A2(net_7583), .A1(net_4714), .ZN(net_4040), .A4(net_4039), .A3(net_3168) );
INV_X4 inst_5631 ( .A(net_10264), .ZN(net_3712) );
OAI211_X2 inst_2186 ( .C1(net_7184), .C2(net_6542), .ZN(net_6523), .B(net_5618), .A(net_3527) );
NAND3_X2 inst_3269 ( .ZN(net_4153), .A2(net_4152), .A3(net_3703), .A1(net_1581) );
CLKBUF_X2 inst_15745 ( .A(net_15663), .Z(net_15664) );
AOI22_X2 inst_9094 ( .A1(net_9675), .A2(net_6402), .ZN(net_6398), .B2(net_5263), .B1(net_113) );
OAI21_X2 inst_1944 ( .B2(net_10129), .A(net_10128), .ZN(net_4280), .B1(net_1588) );
AOI22_X2 inst_9079 ( .A1(net_9692), .ZN(net_6424), .B1(net_6423), .A2(net_6382), .B2(net_5263) );
XNOR2_X2 inst_210 ( .ZN(net_4936), .A(net_4392), .B(net_2337) );
CLKBUF_X2 inst_13763 ( .A(net_13681), .Z(net_13682) );
AOI22_X2 inst_9411 ( .A1(net_9952), .B1(net_6808), .ZN(net_4743), .A2(net_4742), .B2(net_4741) );
CLKBUF_X2 inst_11675 ( .A(net_11501), .Z(net_11594) );
NAND4_X2 inst_3101 ( .ZN(net_4342), .A2(net_3832), .A3(net_3831), .A1(net_3575), .A4(net_3574) );
DFF_X1 inst_8720 ( .QN(net_10171), .D(net_6267), .CK(net_12311) );
INV_X4 inst_4942 ( .A(net_6165), .ZN(net_4634) );
CLKBUF_X2 inst_14998 ( .A(net_14916), .Z(net_14917) );
CLKBUF_X2 inst_12103 ( .A(net_12021), .Z(net_12022) );
INV_X4 inst_5893 ( .A(net_677), .ZN(net_609) );
NAND2_X2 inst_3881 ( .A2(net_4027), .ZN(net_4025), .A1(net_4024) );
INV_X4 inst_5331 ( .ZN(net_3746), .A(net_1262) );
DFF_X2 inst_8164 ( .QN(net_10030), .D(net_5054), .CK(net_13700) );
INV_X2 inst_7123 ( .ZN(net_944), .A(net_943) );
CLKBUF_X2 inst_14580 ( .A(net_14498), .Z(net_14499) );
INV_X4 inst_4778 ( .ZN(net_4298), .A(net_3996) );
OAI22_X2 inst_1294 ( .B1(net_10041), .A1(net_9942), .A2(net_4274), .B2(net_3588), .ZN(net_3585) );
DFF_X2 inst_7663 ( .D(net_6726), .QN(net_159), .CK(net_12813) );
OAI221_X2 inst_1712 ( .B2(net_3910), .ZN(net_3740), .B1(net_3739), .A(net_2668), .C2(net_2443), .C1(net_1081) );
INV_X4 inst_5325 ( .ZN(net_5066), .A(net_3772) );
INV_X4 inst_5238 ( .A(net_1560), .ZN(net_1471) );
CLKBUF_X2 inst_15493 ( .A(net_15411), .Z(net_15412) );
CLKBUF_X2 inst_14605 ( .A(net_14523), .Z(net_14524) );
OR2_X4 inst_747 ( .ZN(net_7757), .A2(net_6184), .A1(net_5249) );
NAND4_X2 inst_3108 ( .ZN(net_4335), .A1(net_3858), .A3(net_3857), .A4(net_3676), .A2(net_3446) );
INV_X4 inst_4576 ( .A(net_8140), .ZN(net_8110) );
AOI22_X2 inst_9070 ( .B1(net_9690), .A1(net_6816), .A2(net_6684), .B2(net_6683), .ZN(net_6596) );
INV_X2 inst_6685 ( .ZN(net_8343), .A(net_8277) );
CLKBUF_X2 inst_12626 ( .A(net_12544), .Z(net_12545) );
NOR2_X2 inst_2853 ( .A2(net_10094), .A1(net_10093), .ZN(net_2180) );
NAND2_X2 inst_3806 ( .A1(net_10075), .A2(net_4534), .ZN(net_4532) );
INV_X8 inst_4486 ( .ZN(net_8479), .A(net_8415) );
CLKBUF_X2 inst_12893 ( .A(net_12811), .Z(net_12812) );
INV_X2 inst_7267 ( .A(net_8918), .ZN(net_8917) );
CLKBUF_X2 inst_15331 ( .A(net_13128), .Z(net_15250) );
AOI211_X2 inst_10291 ( .ZN(net_4669), .C2(net_4251), .A(net_3212), .C1(net_3197), .B(net_2416) );
CLKBUF_X2 inst_11362 ( .A(net_11280), .Z(net_11281) );
INV_X4 inst_6546 ( .A(net_10147), .ZN(net_898) );
CLKBUF_X2 inst_14946 ( .A(net_11893), .Z(net_14865) );
CLKBUF_X2 inst_12166 ( .A(net_11025), .Z(net_12085) );
NOR2_X2 inst_2775 ( .ZN(net_3180), .A2(net_3179), .A1(net_167) );
DFF_X2 inst_7855 ( .Q(net_9899), .D(net_6218), .CK(net_12783) );
CLKBUF_X2 inst_15055 ( .A(net_14973), .Z(net_14974) );
DFF_X1 inst_8553 ( .Q(net_8816), .D(net_7315), .CK(net_11778) );
INV_X4 inst_5589 ( .ZN(net_1289), .A(net_884) );
CLKBUF_X2 inst_15324 ( .A(net_15242), .Z(net_15243) );
CLKBUF_X2 inst_12334 ( .A(net_12252), .Z(net_12253) );
CLKBUF_X2 inst_11658 ( .A(net_11576), .Z(net_11577) );
XNOR2_X2 inst_305 ( .B(net_3985), .ZN(net_3252), .A(net_3010) );
INV_X2 inst_6795 ( .A(net_9267), .ZN(net_5416) );
CLKBUF_X2 inst_10853 ( .A(net_10771), .Z(net_10772) );
CLKBUF_X2 inst_13516 ( .A(net_11176), .Z(net_13435) );
OAI221_X2 inst_1595 ( .B1(net_10210), .C1(net_7127), .ZN(net_5643), .B2(net_5642), .C2(net_4905), .A(net_3731) );
DFF_X2 inst_7881 ( .QN(net_10095), .D(net_6037), .CK(net_15533) );
INV_X4 inst_5651 ( .A(net_10458), .ZN(net_1156) );
INV_X4 inst_6291 ( .A(net_10052), .ZN(net_4755) );
CLKBUF_X2 inst_14848 ( .A(net_14766), .Z(net_14767) );
DFF_X2 inst_7867 ( .QN(net_10155), .D(net_6005), .CK(net_13496) );
CLKBUF_X2 inst_12476 ( .A(net_12394), .Z(net_12395) );
CLKBUF_X2 inst_14547 ( .A(net_14465), .Z(net_14466) );
INV_X4 inst_5740 ( .ZN(net_936), .A(net_746) );
CLKBUF_X2 inst_13578 ( .A(net_11023), .Z(net_13497) );
CLKBUF_X2 inst_10926 ( .A(net_10569), .Z(net_10845) );
AND2_X2 inst_10602 ( .A1(net_3118), .ZN(net_2063), .A2(net_2062) );
CLKBUF_X2 inst_12319 ( .A(net_12237), .Z(net_12238) );
CLKBUF_X2 inst_10993 ( .A(net_10911), .Z(net_10912) );
INV_X4 inst_6227 ( .A(net_9831), .ZN(net_778) );
CLKBUF_X2 inst_13489 ( .A(net_13407), .Z(net_13408) );
CLKBUF_X2 inst_13069 ( .A(net_12987), .Z(net_12988) );
INV_X4 inst_6585 ( .A(net_9184), .ZN(net_5443) );
DFF_X2 inst_8079 ( .QN(net_10364), .D(net_5311), .CK(net_13614) );
CLKBUF_X2 inst_15595 ( .A(net_15513), .Z(net_15514) );
CLKBUF_X2 inst_14930 ( .A(net_14848), .Z(net_14849) );
CLKBUF_X2 inst_15511 ( .A(net_11491), .Z(net_15430) );
CLKBUF_X2 inst_14898 ( .A(net_13127), .Z(net_14817) );
DFF_X2 inst_7774 ( .Q(net_9725), .D(net_6528), .CK(net_15548) );
CLKBUF_X2 inst_11620 ( .A(net_11538), .Z(net_11539) );
CLKBUF_X2 inst_11605 ( .A(net_11523), .Z(net_11524) );
OAI33_X1 inst_963 ( .ZN(net_3635), .B3(net_3634), .A3(net_3634), .B2(net_3047), .A1(net_2722), .A2(net_2280), .B1(net_2120) );
OR2_X2 inst_907 ( .ZN(net_4948), .A2(net_4440), .A1(net_2755) );
OR2_X2 inst_922 ( .ZN(net_3386), .A1(net_3183), .A2(net_3182) );
OAI221_X2 inst_1614 ( .B1(net_10412), .C1(net_7192), .A(net_6546), .ZN(net_5599), .B2(net_4477), .C2(net_4455) );
CLKBUF_X2 inst_11323 ( .A(net_10654), .Z(net_11242) );
DFF_X2 inst_8225 ( .D(net_4869), .Q(net_226), .CK(net_10827) );
OAI221_X2 inst_1502 ( .C2(net_9063), .B2(net_9056), .ZN(net_7359), .C1(net_7209), .A(net_6991), .B1(net_5513) );
DFF_X1 inst_8773 ( .Q(net_10344), .D(net_4945), .CK(net_10623) );
CLKBUF_X2 inst_15072 ( .A(net_14990), .Z(net_14991) );
INV_X4 inst_5436 ( .ZN(net_1512), .A(net_1116) );
CLKBUF_X2 inst_12435 ( .A(net_12353), .Z(net_12354) );
CLKBUF_X2 inst_10693 ( .A(net_10611), .Z(net_10612) );
AOI22_X2 inst_9475 ( .B1(net_9893), .A1(net_9762), .B2(net_4969), .ZN(net_3848), .A2(net_2462) );
CLKBUF_X2 inst_14418 ( .A(net_14336), .Z(net_14337) );
INV_X4 inst_6115 ( .A(net_9931), .ZN(net_1339) );
DFF_X1 inst_8516 ( .QN(net_8819), .D(net_7484), .CK(net_12318) );
NAND2_X2 inst_4091 ( .A1(net_10156), .ZN(net_3015), .A2(net_2530) );
CLKBUF_X2 inst_12621 ( .A(net_12539), .Z(net_12540) );
DFF_X2 inst_7602 ( .Q(net_9348), .D(net_7339), .CK(net_15297) );
INV_X2 inst_6989 ( .ZN(net_1650), .A(net_1649) );
CLKBUF_X2 inst_13231 ( .A(net_13149), .Z(net_13150) );
NAND2_X2 inst_3907 ( .ZN(net_4361), .A2(net_4326), .A1(net_464) );
INV_X2 inst_6807 ( .ZN(net_5071), .A(net_4800) );
AOI22_X2 inst_9619 ( .B1(net_9787), .A2(net_6413), .ZN(net_3434), .A1(net_3433), .B2(net_2462) );
OAI221_X2 inst_1568 ( .C1(net_10218), .C2(net_7295), .B2(net_7293), .ZN(net_7183), .B1(net_7182), .A(net_6831) );
CLKBUF_X2 inst_11439 ( .A(net_10647), .Z(net_11358) );
CLKBUF_X2 inst_14752 ( .A(net_14670), .Z(net_14671) );
INV_X4 inst_6177 ( .ZN(net_5261), .A(net_177) );
CLKBUF_X2 inst_12383 ( .A(net_11905), .Z(net_12302) );
DFF_X1 inst_8487 ( .QN(net_9427), .D(net_7843), .CK(net_12667) );
CLKBUF_X2 inst_12223 ( .A(net_12141), .Z(net_12142) );
AOI22_X2 inst_9258 ( .B2(net_8041), .A2(net_6111), .ZN(net_6048), .A1(net_6047), .B1(net_1787) );
OR2_X2 inst_873 ( .A1(net_10503), .ZN(net_6977), .A2(net_6976) );
NAND2_X4 inst_3366 ( .ZN(net_4687), .A1(net_4031), .A2(net_3901) );
NAND2_X2 inst_3692 ( .A2(net_9257), .A1(net_8982), .ZN(net_6234) );
SDFF_X2 inst_653 ( .SI(net_9475), .Q(net_9475), .SE(net_3073), .CK(net_14651), .D(x2968) );
INV_X4 inst_6454 ( .ZN(net_4177), .A(net_156) );
CLKBUF_X2 inst_13439 ( .A(net_13357), .Z(net_13358) );
AOI21_X2 inst_10164 ( .A(net_5378), .ZN(net_3876), .B1(net_3875), .B2(net_3141) );
AOI21_X2 inst_10022 ( .B1(net_8595), .A(net_7916), .B2(net_7915), .ZN(net_7857) );
DFF_X1 inst_8563 ( .QN(net_9567), .D(net_7173), .CK(net_14265) );
DFF_X2 inst_8304 ( .QN(net_10244), .D(net_4568), .CK(net_11149) );
AOI211_X2 inst_10282 ( .ZN(net_5957), .C2(net_5338), .A(net_3613), .B(net_3306), .C1(net_3081) );
NAND2_X2 inst_3767 ( .ZN(net_4973), .A2(net_4577), .A1(net_954) );
OAI21_X2 inst_1746 ( .B1(net_8691), .ZN(net_8674), .B2(net_8646), .A(net_7853) );
CLKBUF_X2 inst_11099 ( .A(net_11017), .Z(net_11018) );
DFF_X1 inst_8839 ( .QN(net_9958), .D(net_2157), .CK(net_10755) );
DFF_X1 inst_8679 ( .D(net_6741), .Q(net_146), .CK(net_12598) );
MUX2_X2 inst_4431 ( .B(net_6854), .Z(net_6185), .S(net_6184), .A(net_1012) );
NAND2_X4 inst_3371 ( .ZN(net_3370), .A1(net_3285), .A2(net_3179) );
NAND4_X2 inst_3052 ( .ZN(net_5929), .A4(net_5184), .A3(net_3875), .A2(net_3344), .A1(net_2408) );
CLKBUF_X2 inst_13406 ( .A(net_13324), .Z(net_13325) );
DFF_X2 inst_8233 ( .Q(net_10491), .D(net_4892), .CK(net_15219) );
INV_X2 inst_6982 ( .ZN(net_3026), .A(net_2076) );
CLKBUF_X2 inst_15817 ( .A(net_15735), .Z(net_15736) );
NAND2_X2 inst_3649 ( .ZN(net_6782), .A2(net_6447), .A1(net_3847) );
CLKBUF_X2 inst_13548 ( .A(net_12133), .Z(net_13467) );
NOR2_X2 inst_2907 ( .ZN(net_2167), .A2(net_1425), .A1(net_199) );
INV_X4 inst_4609 ( .ZN(net_7588), .A(net_7556) );
NAND2_X2 inst_4072 ( .ZN(net_2656), .A1(net_2655), .A2(net_2654) );
INV_X4 inst_6526 ( .A(net_10511), .ZN(net_3686) );
CLKBUF_X2 inst_11843 ( .A(net_11761), .Z(net_11762) );
NOR2_X2 inst_2656 ( .A2(net_7615), .ZN(net_5402), .A1(net_5235) );
INV_X4 inst_5901 ( .A(net_2758), .ZN(net_2244) );
NOR2_X2 inst_3000 ( .A2(net_4641), .A1(net_4015), .ZN(net_2824) );
AOI22_X2 inst_9668 ( .B2(net_10080), .A2(net_10072), .B1(net_10071), .A1(net_10063), .ZN(net_954) );
OAI22_X2 inst_1163 ( .A1(net_7231), .A2(net_5151), .B2(net_5150), .ZN(net_5110), .B1(net_740) );
CLKBUF_X2 inst_10641 ( .A(net_10559), .Z(net_10560) );
DFF_X2 inst_8282 ( .Q(net_9754), .D(net_4737), .CK(net_14582) );
DFF_X2 inst_8301 ( .Q(net_9622), .D(net_4443), .CK(net_14086) );
OAI221_X2 inst_1604 ( .B1(net_10201), .C1(net_7243), .B2(net_5642), .ZN(net_5632), .C2(net_4905), .A(net_3731) );
NAND3_X2 inst_3239 ( .A1(net_7142), .ZN(net_4716), .A3(net_4713), .A2(net_1514) );
NOR4_X2 inst_2314 ( .A3(net_10304), .A1(net_10303), .ZN(net_7413), .A4(net_7065), .A2(net_544) );
AOI22_X2 inst_9426 ( .A1(net_9756), .B1(net_6828), .ZN(net_4623), .A2(net_4622), .B2(net_4621) );
CLKBUF_X2 inst_12885 ( .A(net_12803), .Z(net_12804) );
CLKBUF_X2 inst_13854 ( .A(net_13772), .Z(net_13773) );
NOR2_X2 inst_2812 ( .ZN(net_2647), .A1(net_2646), .A2(net_2645) );
CLKBUF_X2 inst_14441 ( .A(net_14359), .Z(net_14360) );
INV_X4 inst_4743 ( .A(net_4895), .ZN(net_4386) );
CLKBUF_X2 inst_15607 ( .A(net_15525), .Z(net_15526) );
DFF_X1 inst_8592 ( .Q(net_9667), .D(net_7098), .CK(net_11621) );
NAND3_X2 inst_3197 ( .ZN(net_7467), .A1(net_7383), .A3(net_5006), .A2(x813) );
INV_X4 inst_4651 ( .A(net_9255), .ZN(net_6233) );
AOI21_X2 inst_10126 ( .A(net_4460), .ZN(net_4318), .B2(net_3717), .B1(net_859) );
XOR2_X2 inst_7 ( .B(net_5374), .Z(net_4666), .A(net_4665) );
CLKBUF_X2 inst_13640 ( .A(net_13558), .Z(net_13559) );
AOI22_X2 inst_9672 ( .B2(net_10505), .A2(net_10504), .B1(net_10498), .A1(net_10497), .ZN(net_803) );
NAND2_X2 inst_3450 ( .A1(net_9495), .ZN(net_8474), .A2(net_8473) );
CLKBUF_X2 inst_14988 ( .A(net_14700), .Z(net_14907) );
DFF_X2 inst_8006 ( .QN(net_10121), .D(net_5502), .CK(net_12343) );
AOI222_X1 inst_9707 ( .B1(net_9504), .A2(net_8310), .B2(net_8309), .C2(net_8308), .ZN(net_8271), .C1(net_8209), .A1(x2767) );
CLKBUF_X2 inst_13742 ( .A(net_13660), .Z(net_13661) );
OAI22_X2 inst_1083 ( .ZN(net_6576), .A1(net_6575), .A2(net_5913), .B2(net_5912), .B1(net_534) );
INV_X4 inst_5408 ( .ZN(net_1962), .A(net_1157) );
NAND2_X2 inst_4073 ( .ZN(net_2652), .A2(net_2651), .A1(net_1955) );
INV_X4 inst_6123 ( .A(net_10225), .ZN(net_1088) );
CLKBUF_X2 inst_12036 ( .A(net_11954), .Z(net_11955) );
OAI22_X2 inst_1136 ( .A1(net_7229), .A2(net_5151), .B2(net_5150), .ZN(net_5141), .B1(net_394) );
NOR2_X4 inst_2466 ( .A2(net_9031), .A1(net_9030), .ZN(net_8562) );
CLKBUF_X2 inst_11979 ( .A(net_11897), .Z(net_11898) );
CLKBUF_X2 inst_11877 ( .A(net_11795), .Z(net_11796) );
CLKBUF_X2 inst_12070 ( .A(net_11988), .Z(net_11989) );
AND2_X4 inst_10402 ( .ZN(net_5390), .A1(net_5389), .A2(net_5388) );
CLKBUF_X2 inst_13615 ( .A(net_13533), .Z(net_13534) );
CLKBUF_X2 inst_13360 ( .A(net_13278), .Z(net_13279) );
CLKBUF_X2 inst_11262 ( .A(net_10679), .Z(net_11181) );
OR3_X4 inst_696 ( .A3(net_10199), .ZN(net_7660), .A1(net_4979), .A2(net_4978) );
AOI222_X1 inst_9719 ( .C1(net_10501), .B1(net_10396), .A1(net_9682), .C2(net_6415), .A2(net_5966), .ZN(net_4065), .B2(net_4062) );
AOI22_X2 inst_9621 ( .A1(net_10052), .B1(net_9823), .A2(net_5174), .ZN(net_3431), .B2(net_2556) );
CLKBUF_X2 inst_14474 ( .A(net_14392), .Z(net_14393) );
NAND3_X2 inst_3311 ( .A2(net_9226), .ZN(net_1766), .A1(net_1452), .A3(net_456) );
CLKBUF_X2 inst_13598 ( .A(net_13516), .Z(net_13517) );
CLKBUF_X2 inst_11890 ( .A(net_10690), .Z(net_11809) );
CLKBUF_X2 inst_15555 ( .A(net_15473), .Z(net_15474) );
CLKBUF_X2 inst_13339 ( .A(net_13257), .Z(net_13258) );
CLKBUF_X2 inst_12059 ( .A(net_10687), .Z(net_11978) );
CLKBUF_X2 inst_10755 ( .A(net_10673), .Z(net_10674) );
INV_X4 inst_5055 ( .ZN(net_2239), .A(net_1878) );
INV_X4 inst_5081 ( .ZN(net_2615), .A(net_1910) );
INV_X4 inst_5117 ( .ZN(net_2502), .A(net_1162) );
INV_X4 inst_4929 ( .A(net_8865), .ZN(net_2951) );
INV_X4 inst_5114 ( .A(net_2934), .ZN(net_1644) );
CLKBUF_X2 inst_13942 ( .A(net_13860), .Z(net_13861) );
INV_X4 inst_6128 ( .A(net_9555), .ZN(net_8179) );
CLKBUF_X2 inst_14885 ( .A(net_14803), .Z(net_14804) );
CLKBUF_X2 inst_10778 ( .A(net_10696), .Z(net_10697) );
CLKBUF_X2 inst_11712 ( .A(net_11630), .Z(net_11631) );
NAND2_X2 inst_3969 ( .A2(net_3378), .ZN(net_3377), .A1(net_578) );
AOI221_X2 inst_9909 ( .B1(net_9864), .B2(net_9101), .A(net_6945), .C2(net_6944), .ZN(net_6785), .C1(net_235) );
NOR3_X2 inst_2363 ( .ZN(net_8811), .A1(net_8809), .A3(net_8597), .A2(net_7901) );
INV_X4 inst_6014 ( .A(net_9998), .ZN(net_525) );
AND2_X4 inst_10423 ( .A2(net_10175), .ZN(net_4617), .A1(net_4006) );
INV_X4 inst_6257 ( .A(net_9848), .ZN(net_453) );
NAND2_X2 inst_4029 ( .A1(net_9046), .ZN(net_3147), .A2(net_2708) );
OAI221_X2 inst_1629 ( .B1(net_10336), .C1(net_7237), .B2(net_5591), .ZN(net_5578), .C2(net_4902), .A(net_3507) );
HA_X1 inst_7341 ( .S(net_6171), .CO(net_6170), .B(net_5236), .A(net_1241) );
CLKBUF_X2 inst_15583 ( .A(net_15501), .Z(net_15502) );
NAND2_X2 inst_3424 ( .A1(net_8967), .ZN(net_8506), .A2(net_8505) );
INV_X4 inst_6268 ( .A(net_10386), .ZN(net_446) );
CLKBUF_X2 inst_12138 ( .A(net_11084), .Z(net_12057) );
CLKBUF_X2 inst_13923 ( .A(net_11341), .Z(net_13842) );
NAND2_X2 inst_3713 ( .A1(net_5908), .ZN(net_5906), .A2(net_5905) );
NOR2_X2 inst_2580 ( .ZN(net_7310), .A2(net_7078), .A1(net_4603) );
INV_X4 inst_5681 ( .A(net_9243), .ZN(net_5268) );
NOR3_X2 inst_2394 ( .A1(net_7828), .ZN(net_7706), .A3(net_7568), .A2(x3390) );
CLKBUF_X2 inst_11342 ( .A(net_10725), .Z(net_11261) );
INV_X4 inst_4574 ( .ZN(net_8203), .A(net_8124) );
CLKBUF_X2 inst_14213 ( .A(net_11059), .Z(net_14132) );
DFF_X1 inst_8562 ( .QN(net_9564), .D(net_7174), .CK(net_14266) );
CLKBUF_X2 inst_12268 ( .A(net_12029), .Z(net_12187) );
AOI22_X2 inst_9404 ( .ZN(net_5201), .A2(net_4538), .B2(net_4537), .A1(net_4135), .B1(net_547) );
CLKBUF_X2 inst_15290 ( .A(net_15208), .Z(net_15209) );
CLKBUF_X2 inst_10681 ( .A(net_10549), .Z(net_10600) );
AND2_X2 inst_10612 ( .A1(net_9222), .ZN(net_2543), .A2(net_1845) );
INV_X4 inst_5840 ( .A(net_1351), .ZN(net_861) );
OAI211_X2 inst_2054 ( .C1(net_10134), .ZN(net_7796), .A(net_7795), .B(net_7304), .C2(net_6042) );
CLKBUF_X2 inst_12216 ( .A(net_11243), .Z(net_12135) );
CLKBUF_X2 inst_13448 ( .A(net_13366), .Z(net_13367) );
INV_X4 inst_5294 ( .A(net_1994), .ZN(net_1309) );
INV_X4 inst_5251 ( .A(net_7002), .ZN(net_1963) );
OAI22_X2 inst_1259 ( .B1(net_7201), .A2(net_4842), .B2(net_4841), .ZN(net_4814), .A1(net_4101) );
NAND2_X1 inst_4422 ( .ZN(net_4189), .A1(net_4188), .A2(net_4187) );
CLKBUF_X2 inst_12578 ( .A(net_12496), .Z(net_12497) );
CLKBUF_X2 inst_12219 ( .A(net_12137), .Z(net_12138) );
CLKBUF_X2 inst_14056 ( .A(net_12616), .Z(net_13975) );
CLKBUF_X2 inst_11905 ( .A(net_10755), .Z(net_11824) );
DFF_X1 inst_8623 ( .Q(net_9781), .D(net_7204), .CK(net_14395) );
DFF_X2 inst_7821 ( .Q(net_9179), .D(net_6297), .CK(net_13574) );
INV_X4 inst_5092 ( .ZN(net_5475), .A(net_1742) );
CLKBUF_X2 inst_10702 ( .A(net_10620), .Z(net_10621) );
OAI21_X2 inst_1796 ( .ZN(net_7446), .B1(net_7157), .A(net_6984), .B2(net_6977) );
CLKBUF_X2 inst_12318 ( .A(net_11228), .Z(net_12237) );
DFF_X2 inst_7649 ( .D(net_6753), .QN(net_179), .CK(net_14323) );
CLKBUF_X2 inst_11341 ( .A(net_11259), .Z(net_11260) );
SDFF_X2 inst_535 ( .D(net_9143), .SE(net_933), .CK(net_10997), .SI(x1792), .Q(x1153) );
CLKBUF_X2 inst_15330 ( .A(net_15248), .Z(net_15249) );
INV_X4 inst_5342 ( .ZN(net_1585), .A(net_1247) );
CLKBUF_X2 inst_12970 ( .A(net_12888), .Z(net_12889) );
OAI221_X2 inst_1670 ( .C1(net_7216), .A(net_6546), .B2(net_5642), .ZN(net_5499), .C2(net_4905), .B1(net_1350) );
CLKBUF_X2 inst_12932 ( .A(net_12736), .Z(net_12851) );
CLKBUF_X2 inst_11491 ( .A(net_11318), .Z(net_11410) );
AOI21_X2 inst_10059 ( .ZN(net_7096), .B2(net_7079), .A(net_3563), .B1(net_3399) );
DFF_X2 inst_7853 ( .Q(net_10399), .D(net_6213), .CK(net_15125) );
CLKBUF_X2 inst_11670 ( .A(net_10797), .Z(net_11589) );
AND3_X4 inst_10352 ( .ZN(net_7718), .A2(net_7574), .A3(net_7443), .A1(net_7421) );
DFF_X1 inst_8646 ( .Q(net_9791), .D(net_7208), .CK(net_13346) );
NOR3_X2 inst_2427 ( .ZN(net_4091), .A1(net_3632), .A3(net_1591), .A2(net_1392) );
AOI22_X2 inst_9028 ( .B1(net_9528), .A1(net_8002), .B2(net_8001), .ZN(net_7943), .A2(net_7899) );
AND2_X2 inst_10496 ( .A2(net_10345), .ZN(net_6667), .A1(net_1524) );
DFF_X1 inst_8603 ( .Q(net_9690), .D(net_7105), .CK(net_15244) );
CLKBUF_X2 inst_10677 ( .A(net_10595), .Z(net_10596) );
NAND2_X4 inst_3317 ( .ZN(net_8895), .A1(net_8741), .A2(net_7902) );
AND4_X4 inst_10327 ( .ZN(net_3323), .A4(net_3322), .A3(net_2860), .A1(net_1380), .A2(net_1127) );
INV_X4 inst_5027 ( .ZN(net_5459), .A(net_1938) );
INV_X4 inst_5883 ( .A(net_4172), .ZN(net_622) );
NAND4_X2 inst_3113 ( .ZN(net_4581), .A2(net_4265), .A4(net_4255), .A1(net_4114), .A3(net_2827) );
CLKBUF_X2 inst_13500 ( .A(net_13411), .Z(net_13419) );
CLKBUF_X2 inst_14616 ( .A(net_14534), .Z(net_14535) );
INV_X4 inst_6079 ( .ZN(net_1856), .A(net_119) );
CLKBUF_X2 inst_13245 ( .A(net_13163), .Z(net_13164) );
CLKBUF_X2 inst_11348 ( .A(net_11243), .Z(net_11267) );
NAND2_X2 inst_3695 ( .A2(net_9254), .A1(net_9082), .ZN(net_6226) );
CLKBUF_X2 inst_12309 ( .A(net_11802), .Z(net_12228) );
INV_X2 inst_7206 ( .A(net_9313), .ZN(net_468) );
NAND3_X4 inst_3168 ( .ZN(net_5520), .A2(net_4230), .A1(net_4226), .A3(x6599) );
INV_X2 inst_6687 ( .ZN(net_8339), .A(net_8275) );
NOR3_X2 inst_2385 ( .A1(net_7884), .ZN(net_7806), .A3(net_7805), .A2(net_5684) );
NOR4_X2 inst_2336 ( .ZN(net_4238), .A4(net_3284), .A3(net_2972), .A2(net_2791), .A1(net_1591) );
NAND2_X2 inst_3855 ( .ZN(net_8888), .A2(net_4187), .A1(net_1976) );
INV_X4 inst_5927 ( .ZN(net_1384), .A(net_578) );
DFF_X1 inst_8589 ( .Q(net_9865), .D(net_7107), .CK(net_14258) );
DFF_X1 inst_8574 ( .Q(net_9771), .D(net_7117), .CK(net_15633) );
CLKBUF_X2 inst_13549 ( .A(net_13467), .Z(net_13468) );
AND2_X2 inst_10594 ( .ZN(net_2372), .A2(net_2371), .A1(net_2208) );
AOI22_X2 inst_9482 ( .B1(net_9881), .A2(net_5173), .ZN(net_3841), .B2(net_2973), .A1(net_214) );
NAND2_X4 inst_3318 ( .A2(net_9004), .A1(net_9003), .ZN(net_8736) );
CLKBUF_X2 inst_12771 ( .A(net_12689), .Z(net_12690) );
XNOR2_X2 inst_223 ( .ZN(net_4567), .A(net_4123), .B(net_1784) );
AOI211_X2 inst_10299 ( .C1(net_3696), .ZN(net_3694), .B(net_3693), .C2(net_3692), .A(net_3088) );
INV_X2 inst_6814 ( .ZN(net_4727), .A(net_4726) );
INV_X4 inst_5278 ( .A(net_1570), .ZN(net_1329) );
INV_X4 inst_6042 ( .A(net_10437), .ZN(net_513) );
CLKBUF_X2 inst_13811 ( .A(net_13729), .Z(net_13730) );
NOR3_X2 inst_2420 ( .A2(net_9194), .ZN(net_5447), .A1(net_5101), .A3(net_459) );
NAND2_X2 inst_3564 ( .A2(net_7748), .ZN(net_7686), .A1(net_7685) );
INV_X4 inst_5176 ( .ZN(net_2886), .A(net_2279) );
CLKBUF_X2 inst_15453 ( .A(net_12886), .Z(net_15372) );
CLKBUF_X2 inst_12672 ( .A(net_12590), .Z(net_12591) );
NAND2_X2 inst_4205 ( .A1(net_10458), .A2(net_2049), .ZN(net_1778) );
OAI22_X2 inst_1322 ( .B2(net_2265), .ZN(net_1762), .A2(net_1761), .B1(net_1756), .A1(net_1755) );
CLKBUF_X2 inst_11862 ( .A(net_10892), .Z(net_11781) );
CLKBUF_X2 inst_11452 ( .A(net_11370), .Z(net_11371) );
AOI22_X2 inst_9633 ( .A1(net_10074), .A2(net_5319), .B2(net_5174), .ZN(net_3410), .B1(net_3409) );
CLKBUF_X2 inst_14891 ( .A(net_14809), .Z(net_14810) );
CLKBUF_X2 inst_10954 ( .A(net_10724), .Z(net_10873) );
CLKBUF_X2 inst_14004 ( .A(net_13296), .Z(net_13923) );
CLKBUF_X2 inst_10712 ( .A(net_10630), .Z(net_10631) );
CLKBUF_X2 inst_14237 ( .A(net_14155), .Z(net_14156) );
CLKBUF_X2 inst_15471 ( .A(net_13405), .Z(net_15390) );
AOI21_X2 inst_10248 ( .ZN(net_9115), .B1(net_9081), .A(net_5420), .B2(net_2554) );
CLKBUF_X2 inst_12027 ( .A(net_11945), .Z(net_11946) );
DFF_X2 inst_7668 ( .D(net_6689), .QN(net_173), .CK(net_15613) );
CLKBUF_X2 inst_11063 ( .A(net_10566), .Z(net_10982) );
AOI22_X2 inst_9408 ( .B1(net_9174), .A2(net_4802), .B2(net_4801), .ZN(net_4800), .A1(net_1730) );
AOI21_X2 inst_10156 ( .B1(net_4103), .ZN(net_4099), .A(net_4098), .B2(net_4097) );
DFF_X2 inst_8379 ( .D(net_1086), .Q(net_260), .CK(net_13863) );
NAND2_X2 inst_3493 ( .A1(net_8314), .ZN(net_8261), .A2(net_8147) );
INV_X4 inst_6156 ( .A(net_10265), .ZN(net_840) );
CLKBUF_X2 inst_13151 ( .A(net_10711), .Z(net_13070) );
AND2_X4 inst_10413 ( .ZN(net_4801), .A1(net_4376), .A2(net_4375) );
AOI221_X2 inst_9776 ( .B1(net_8982), .ZN(net_7422), .C2(net_7277), .A(net_7084), .B2(net_5997), .C1(net_2869) );
NOR2_X2 inst_3019 ( .A2(net_10198), .A1(net_10197), .ZN(net_661) );
INV_X4 inst_4622 ( .ZN(net_7131), .A(net_7011) );
NOR4_X2 inst_2327 ( .ZN(net_5379), .A3(net_5378), .A4(net_4672), .A1(net_3161), .A2(net_3160) );
CLKBUF_X2 inst_13430 ( .A(net_13348), .Z(net_13349) );
NAND2_X2 inst_3487 ( .ZN(net_8545), .A2(net_8377), .A1(net_3507) );
INV_X4 inst_5078 ( .ZN(net_2605), .A(net_1826) );
INV_X2 inst_6866 ( .A(net_3456), .ZN(net_3382) );
CLKBUF_X2 inst_14555 ( .A(net_14473), .Z(net_14474) );
CLKBUF_X2 inst_14421 ( .A(net_14339), .Z(net_14340) );
CLKBUF_X2 inst_11783 ( .A(net_11701), .Z(net_11702) );
NAND2_X2 inst_3597 ( .ZN(net_7269), .A2(net_6880), .A1(net_6608) );
DFF_X2 inst_8210 ( .Q(net_10085), .D(net_4850), .CK(net_10735) );
CLKBUF_X2 inst_10661 ( .A(net_10579), .Z(net_10580) );
CLKBUF_X2 inst_14976 ( .A(net_14894), .Z(net_14895) );
CLKBUF_X2 inst_11757 ( .A(net_11675), .Z(net_11676) );
CLKBUF_X2 inst_13422 ( .A(net_13296), .Z(net_13341) );
NOR2_X2 inst_2607 ( .ZN(net_6254), .A2(net_6253), .A1(net_5811) );
CLKBUF_X2 inst_11579 ( .A(net_11497), .Z(net_11498) );
XNOR2_X2 inst_113 ( .ZN(net_7891), .A(net_7817), .B(net_6893) );
CLKBUF_X2 inst_13893 ( .A(net_13811), .Z(net_13812) );
DFF_X2 inst_8133 ( .QN(net_9845), .D(net_5124), .CK(net_12492) );
CLKBUF_X2 inst_11395 ( .A(net_11313), .Z(net_11314) );
AND2_X4 inst_10433 ( .ZN(net_4694), .A2(net_3630), .A1(net_2763) );
DFF_X2 inst_7791 ( .Q(net_9796), .D(net_6505), .CK(net_13204) );
CLKBUF_X2 inst_14023 ( .A(net_12346), .Z(net_13942) );
NOR2_X2 inst_2690 ( .A2(net_10166), .ZN(net_4540), .A1(net_2258) );
AOI222_X1 inst_9680 ( .B1(net_9508), .A2(net_8310), .B2(net_8309), .C2(net_8308), .ZN(net_8307), .C1(net_8232), .A1(x2531) );
AOI22_X2 inst_9106 ( .A1(net_9686), .A2(net_6418), .ZN(net_6386), .B2(net_5263), .B1(net_4026) );
DFF_X1 inst_8479 ( .Q(net_9624), .D(net_7951), .CK(net_15027) );
DFF_X1 inst_8689 ( .D(net_6712), .Q(net_142), .CK(net_15099) );
CLKBUF_X2 inst_10849 ( .A(net_10767), .Z(net_10768) );
AND2_X4 inst_10467 ( .A2(net_10461), .ZN(net_2753), .A1(net_888) );
INV_X2 inst_7298 ( .ZN(net_9053), .A(net_3376) );
OAI221_X2 inst_1544 ( .B2(net_7295), .C2(net_7293), .C1(net_7221), .ZN(net_7218), .A(net_6825), .B1(net_5459) );
NAND2_X2 inst_4063 ( .A2(net_9199), .ZN(net_3891), .A1(net_2445) );
AOI21_X2 inst_10069 ( .B1(net_10280), .ZN(net_6972), .A(net_6678), .B2(net_264) );
DFF_X2 inst_8340 ( .QN(net_10165), .D(net_3007), .CK(net_12245) );
INV_X4 inst_6261 ( .A(net_9165), .ZN(net_1246) );
AOI22_X2 inst_9016 ( .A2(net_8030), .B2(net_8029), .ZN(net_8020), .B1(net_666), .A1(net_209) );
NOR2_X2 inst_2625 ( .ZN(net_6009), .A2(net_5428), .A1(net_5014) );
AOI221_X2 inst_9771 ( .B1(net_9529), .B2(net_8001), .ZN(net_7511), .C2(net_7474), .C1(net_5986), .A(net_3298) );
NAND4_X2 inst_3148 ( .ZN(net_2159), .A4(net_1136), .A2(net_975), .A1(net_650), .A3(net_634) );
CLKBUF_X2 inst_14088 ( .A(net_14006), .Z(net_14007) );
INV_X4 inst_6064 ( .ZN(net_6823), .A(net_254) );
CLKBUF_X2 inst_12652 ( .A(net_12570), .Z(net_12571) );
AOI22_X2 inst_9244 ( .A1(net_9948), .B1(net_9849), .A2(net_6141), .B2(net_6129), .ZN(net_6067) );
NAND2_X4 inst_3329 ( .A2(net_8938), .A1(net_8932), .ZN(net_8606) );
INV_X4 inst_4761 ( .ZN(net_4665), .A(net_3998) );
INV_X4 inst_5180 ( .ZN(net_7512), .A(net_1557) );
NOR2_X2 inst_3026 ( .ZN(net_580), .A2(net_276), .A1(net_275) );
INV_X4 inst_5769 ( .ZN(net_1349), .A(net_729) );
CLKBUF_X2 inst_13844 ( .A(net_13762), .Z(net_13763) );
NOR2_X2 inst_2847 ( .A2(net_3960), .ZN(net_3354), .A1(net_2258) );
OAI221_X2 inst_1442 ( .B1(net_8691), .ZN(net_8665), .B2(net_8610), .C2(net_7741), .A(net_7700), .C1(net_1306) );
DFF_X1 inst_8573 ( .Q(net_9675), .D(net_7099), .CK(net_14839) );
INV_X2 inst_6952 ( .A(net_6514), .ZN(net_1886) );
NAND2_X2 inst_3639 ( .ZN(net_6913), .A2(net_6912), .A1(net_2674) );
XNOR2_X2 inst_332 ( .ZN(net_2994), .B(net_2993), .A(net_2453) );
CLKBUF_X2 inst_14192 ( .A(net_12433), .Z(net_14111) );
NAND2_X2 inst_4013 ( .A1(net_4026), .ZN(net_3081), .A2(net_3080) );
OAI211_X2 inst_2132 ( .C2(net_6774), .ZN(net_6716), .A(net_6340), .B(net_6079), .C1(net_423) );
OAI22_X2 inst_1289 ( .A2(net_10232), .B2(net_8843), .ZN(net_3734), .A1(net_3546), .B1(net_1272) );
CLKBUF_X2 inst_13646 ( .A(net_10657), .Z(net_13565) );
INV_X4 inst_4979 ( .ZN(net_2604), .A(net_2291) );
AND2_X4 inst_10411 ( .ZN(net_5742), .A1(net_4788), .A2(net_4786) );
AOI22_X2 inst_9194 ( .A1(net_9884), .B1(net_9785), .A2(net_8042), .B2(net_8041), .ZN(net_6119) );
INV_X2 inst_7226 ( .ZN(net_416), .A(x3507) );
INV_X4 inst_4686 ( .ZN(net_5393), .A(net_4971) );
CLKBUF_X2 inst_14241 ( .A(net_11803), .Z(net_14160) );
CLKBUF_X2 inst_13130 ( .A(net_13048), .Z(net_13049) );
INV_X4 inst_4869 ( .A(net_8082), .ZN(net_8081) );
CLKBUF_X2 inst_12769 ( .A(net_12687), .Z(net_12688) );
NAND3_X2 inst_3245 ( .ZN(net_4700), .A3(net_4563), .A1(net_4562), .A2(net_2697) );
OR2_X4 inst_752 ( .ZN(net_5105), .A1(net_4475), .A2(net_4474) );
NAND3_X2 inst_3202 ( .ZN(net_7408), .A3(net_7407), .A2(net_6257), .A1(net_5815) );
NAND2_X2 inst_4279 ( .ZN(net_2950), .A2(net_952), .A1(net_690) );
OAI21_X2 inst_1951 ( .ZN(net_3924), .A(net_3561), .B1(net_2989), .B2(net_2985) );
XNOR2_X2 inst_378 ( .ZN(net_2452), .A(net_2451), .B(net_2450) );
DFF_X2 inst_7444 ( .QN(net_9297), .D(net_8207), .CK(net_11495) );
OAI222_X2 inst_1384 ( .B1(net_7665), .A2(net_7664), .C2(net_7663), .ZN(net_6001), .B2(net_5205), .A1(net_4203), .C1(net_1879) );
DFF_X2 inst_8151 ( .QN(net_9851), .D(net_5079), .CK(net_12122) );
OAI211_X2 inst_2118 ( .C2(net_6778), .ZN(net_6730), .A(net_6357), .B(net_6091), .C1(net_330) );
CLKBUF_X2 inst_11302 ( .A(net_11220), .Z(net_11221) );
DFF_X1 inst_8750 ( .Q(net_9170), .D(net_5788), .CK(net_11351) );
OAI211_X2 inst_2200 ( .C1(net_7294), .A(net_6546), .ZN(net_6507), .C2(net_6501), .B(net_5760) );
DFF_X2 inst_7749 ( .QN(net_10157), .D(net_6275), .CK(net_13499) );
DFF_X1 inst_8817 ( .QN(net_10234), .D(net_3253), .CK(net_10600) );
INV_X4 inst_4937 ( .ZN(net_3075), .A(net_3056) );
INV_X4 inst_5048 ( .A(net_5983), .ZN(net_1898) );
AND4_X4 inst_10320 ( .ZN(net_6850), .A4(net_5947), .A1(net_3772), .A3(net_1037), .A2(net_599) );
DFF_X2 inst_8284 ( .QN(net_10246), .D(net_4926), .CK(net_12177) );
DFF_X2 inst_8080 ( .Q(net_9574), .D(net_5264), .CK(net_11596) );
CLKBUF_X2 inst_11470 ( .A(net_11388), .Z(net_11389) );
AOI221_X2 inst_9948 ( .C2(net_10129), .B1(net_10128), .ZN(net_5274), .A(net_4591), .B2(net_4424), .C1(net_2876) );
CLKBUF_X2 inst_12693 ( .A(net_12611), .Z(net_12612) );
CLKBUF_X2 inst_14707 ( .A(net_14625), .Z(net_14626) );
XNOR2_X2 inst_250 ( .ZN(net_4118), .A(net_3959), .B(net_2046) );
NAND2_X2 inst_4356 ( .A2(net_9734), .ZN(net_1796), .A1(net_973) );
AOI22_X2 inst_9275 ( .B2(net_10131), .A1(net_10130), .ZN(net_5752), .A2(net_4932), .B1(net_4675) );
CLKBUF_X2 inst_11707 ( .A(net_11625), .Z(net_11626) );
DFF_X2 inst_7708 ( .Q(net_10004), .D(net_6263), .CK(net_12580) );
INV_X4 inst_5762 ( .A(net_1118), .ZN(net_950) );
CLKBUF_X2 inst_12250 ( .A(net_11730), .Z(net_12169) );
AOI221_X2 inst_9975 ( .B1(net_9913), .C1(net_9683), .C2(net_5966), .B2(net_4969), .ZN(net_4504), .A(net_4102) );
INV_X4 inst_6595 ( .ZN(net_767), .A(net_173) );
AOI22_X2 inst_9384 ( .B1(net_9705), .A1(net_5755), .B2(net_5754), .ZN(net_5440), .A2(net_242) );
INV_X4 inst_5329 ( .ZN(net_2276), .A(net_1265) );
NOR2_X2 inst_2539 ( .ZN(net_8285), .A2(net_8284), .A1(net_8082) );
OAI221_X2 inst_1523 ( .B1(net_10319), .B2(net_9047), .C1(net_7297), .ZN(net_7290), .C2(net_7287), .A(net_6947) );
AOI21_X2 inst_10141 ( .ZN(net_4244), .A(net_3935), .B2(net_3460), .B1(net_1594) );
AOI221_X2 inst_9941 ( .C1(net_10087), .B1(net_10065), .ZN(net_5394), .B2(net_5320), .C2(net_5319), .A(net_4660) );
OAI22_X2 inst_1048 ( .ZN(net_7537), .A1(net_7535), .A2(net_7393), .B2(net_7392), .B1(net_442) );
INV_X2 inst_7120 ( .A(net_1349), .ZN(net_1232) );
CLKBUF_X2 inst_13496 ( .A(net_13302), .Z(net_13415) );
NOR2_X2 inst_2797 ( .A2(net_3114), .ZN(net_2894), .A1(net_2253) );
NAND2_X2 inst_3431 ( .A1(net_9480), .A2(net_8490), .ZN(net_8485) );
CLKBUF_X2 inst_13537 ( .A(net_13455), .Z(net_13456) );
CLKBUF_X2 inst_13193 ( .A(net_12220), .Z(net_13112) );
OAI211_X2 inst_2270 ( .C1(net_7127), .C2(net_6480), .ZN(net_6274), .B(net_5687), .A(net_3679) );
OAI211_X2 inst_2085 ( .C2(net_6778), .ZN(net_6763), .A(net_6390), .B(net_6124), .C1(net_412) );
CLKBUF_X2 inst_11624 ( .A(net_11432), .Z(net_11543) );
NOR3_X2 inst_2401 ( .A3(net_7916), .ZN(net_7629), .A2(net_7502), .A1(net_3298) );
CLKBUF_X2 inst_11097 ( .A(net_11015), .Z(net_11016) );
CLKBUF_X2 inst_12979 ( .A(net_12897), .Z(net_12898) );
INV_X4 inst_5264 ( .ZN(net_2846), .A(net_1390) );
AOI21_X2 inst_10092 ( .B1(net_10280), .A(net_6678), .ZN(net_5770), .B2(net_5200) );
CLKBUF_X2 inst_14723 ( .A(net_14641), .Z(net_14642) );
CLKBUF_X2 inst_12649 ( .A(net_12567), .Z(net_12568) );
AOI22_X2 inst_9356 ( .B1(net_9911), .A2(net_5759), .B2(net_5758), .ZN(net_5566), .A1(net_250) );
DFF_X2 inst_8367 ( .QN(net_9176), .D(net_1746), .CK(net_11241) );
DFF_X2 inst_8015 ( .QN(net_10439), .D(net_5489), .CK(net_11382) );
CLKBUF_X2 inst_15564 ( .A(net_15482), .Z(net_15483) );
CLKBUF_X2 inst_12910 ( .A(net_12002), .Z(net_12829) );
INV_X4 inst_6150 ( .A(net_10476), .ZN(net_741) );
INV_X2 inst_7069 ( .ZN(net_2715), .A(net_1252) );
CLKBUF_X2 inst_14230 ( .A(net_14148), .Z(net_14149) );
DFF_X2 inst_8196 ( .QN(net_10032), .D(net_5028), .CK(net_12115) );
CLKBUF_X2 inst_11779 ( .A(net_11697), .Z(net_11698) );
SDFF_X2 inst_556 ( .D(net_9120), .SE(net_933), .CK(net_10566), .SI(x3194), .Q(x1384) );
INV_X4 inst_6050 ( .ZN(net_4304), .A(net_271) );
CLKBUF_X2 inst_14287 ( .A(net_12270), .Z(net_14206) );
NAND2_X2 inst_3632 ( .A1(net_10506), .ZN(net_6984), .A2(net_6976) );
INV_X4 inst_6204 ( .A(net_9384), .ZN(net_6949) );
DFF_X1 inst_8618 ( .Q(net_9663), .D(net_7266), .CK(net_13284) );
AOI222_X1 inst_9710 ( .A2(net_7930), .ZN(net_7888), .C1(net_7887), .B2(net_7807), .C2(net_5954), .A1(net_1964), .B1(net_685) );
XNOR2_X2 inst_420 ( .ZN(net_1402), .B(net_1401), .A(net_197) );
INV_X4 inst_5147 ( .ZN(net_6047), .A(net_1587) );
CLKBUF_X2 inst_13758 ( .A(net_13676), .Z(net_13677) );
NAND2_X2 inst_3992 ( .A2(net_10442), .ZN(net_3176), .A1(net_3175) );
CLKBUF_X2 inst_12522 ( .A(net_11890), .Z(net_12441) );
NAND3_X2 inst_3265 ( .A1(net_6203), .ZN(net_4825), .A2(net_4233), .A3(net_4229) );
CLKBUF_X2 inst_12573 ( .A(net_12491), .Z(net_12492) );
AOI22_X2 inst_9650 ( .B1(net_10433), .B2(net_3490), .A2(net_2686), .ZN(net_2414), .A1(net_1092) );
CLKBUF_X2 inst_15669 ( .A(net_15517), .Z(net_15588) );
CLKBUF_X2 inst_15641 ( .A(net_15559), .Z(net_15560) );
NAND3_X2 inst_3300 ( .A3(net_9108), .ZN(net_2420), .A2(net_638), .A1(net_620) );
DFF_X2 inst_7558 ( .QN(net_9384), .D(net_7674), .CK(net_13032) );
OAI22_X2 inst_1305 ( .B2(net_3531), .ZN(net_2708), .A1(net_2707), .B1(net_2706), .A2(net_2219) );
DFF_X2 inst_7997 ( .QN(net_10118), .D(net_5517), .CK(net_12362) );
XNOR2_X2 inst_314 ( .ZN(net_3221), .B(net_3004), .A(net_2342) );
CLKBUF_X2 inst_14813 ( .A(net_14731), .Z(net_14732) );
DFF_X1 inst_8713 ( .QN(net_10381), .D(net_6645), .CK(net_14493) );
NAND3_X2 inst_3225 ( .A2(net_9535), .A1(net_5353), .A3(net_5351), .ZN(net_5262) );
CLKBUF_X2 inst_13367 ( .A(net_13285), .Z(net_13286) );
DFF_X2 inst_7597 ( .Q(net_10401), .D(net_7444), .CK(net_15150) );
CLKBUF_X2 inst_12728 ( .A(net_12646), .Z(net_12647) );
CLKBUF_X2 inst_15342 ( .A(net_15260), .Z(net_15261) );
DFF_X1 inst_8757 ( .Q(net_10485), .D(net_5248), .CK(net_13733) );
NAND2_X2 inst_3822 ( .ZN(net_4901), .A1(net_4516), .A2(net_4181) );
AOI22_X2 inst_9603 ( .B1(net_9991), .A2(net_3500), .ZN(net_3465), .A1(net_3464), .B2(net_2468) );
SDFF_X2 inst_597 ( .QN(net_9266), .SE(net_4297), .SI(net_149), .D(net_115), .CK(net_13823) );
INV_X4 inst_6161 ( .A(net_9986), .ZN(net_478) );
DFF_X2 inst_7522 ( .QN(net_9532), .D(net_7824), .CK(net_12750) );
INV_X4 inst_4593 ( .A(net_9512), .ZN(net_7986) );
INV_X4 inst_5524 ( .A(net_10219), .ZN(net_1128) );
INV_X2 inst_7257 ( .A(net_9412), .ZN(net_8221) );
INV_X4 inst_6070 ( .ZN(net_505), .A(net_226) );
NAND3_X2 inst_3307 ( .A2(net_5096), .ZN(net_1841), .A1(net_1577), .A3(net_873) );
CLKBUF_X2 inst_11859 ( .A(net_11777), .Z(net_11778) );
INV_X2 inst_6927 ( .A(net_2754), .ZN(net_1955) );
CLKBUF_X2 inst_15115 ( .A(net_15033), .Z(net_15034) );
CLKBUF_X2 inst_12272 ( .A(net_12190), .Z(net_12191) );
OAI221_X2 inst_1587 ( .B1(net_10205), .B2(net_7295), .C2(net_7293), .ZN(net_7109), .C1(net_7108), .A(net_6929) );
OAI22_X2 inst_1185 ( .A1(net_7294), .A2(net_5151), .B2(net_5150), .ZN(net_5070), .B1(net_1768) );
INV_X4 inst_5452 ( .A(net_6054), .ZN(net_1079) );
DFF_X1 inst_8742 ( .Q(net_9145), .D(net_5725), .CK(net_11002) );
SDFF_X2 inst_472 ( .D(net_9577), .SI(net_2821), .SE(net_758), .Q(net_251), .CK(net_15046) );
XNOR2_X2 inst_447 ( .B(net_9307), .ZN(net_789), .A(net_215) );
INV_X4 inst_4533 ( .ZN(net_8798), .A(net_8797) );
CLKBUF_X2 inst_13715 ( .A(net_13516), .Z(net_13634) );
SDFF_X2 inst_457 ( .D(net_9583), .SI(net_5930), .SE(net_758), .Q(net_257), .CK(net_11582) );
INV_X4 inst_5987 ( .ZN(net_7231), .A(x4851) );
OAI21_X2 inst_1738 ( .ZN(net_8707), .B2(net_8706), .B1(net_8398), .A(net_8369) );
CLKBUF_X2 inst_12872 ( .A(net_12790), .Z(net_12791) );
NOR2_X2 inst_2802 ( .ZN(net_3230), .A2(net_2803), .A1(net_1798) );
NOR2_X2 inst_2623 ( .A1(net_9227), .ZN(net_6436), .A2(net_5707) );
OAI222_X2 inst_1391 ( .B1(net_7732), .A2(net_7731), .C2(net_7730), .ZN(net_5820), .B2(net_4937), .A1(net_3420), .C1(net_706) );
NAND2_X2 inst_4171 ( .ZN(net_2747), .A2(net_2205), .A1(net_1961) );
SDFF_X2 inst_665 ( .SI(net_9472), .Q(net_9472), .SE(net_3073), .CK(net_14646), .D(x3133) );
INV_X4 inst_4843 ( .A(net_4047), .ZN(net_3555) );
CLKBUF_X2 inst_15169 ( .A(net_15087), .Z(net_15088) );
CLKBUF_X2 inst_12929 ( .A(net_12847), .Z(net_12848) );
CLKBUF_X2 inst_12014 ( .A(net_11932), .Z(net_11933) );
CLKBUF_X2 inst_11276 ( .A(net_11194), .Z(net_11195) );
AOI21_X2 inst_10219 ( .ZN(net_2199), .B2(net_2198), .B1(net_2129), .A(net_668) );
NAND2_X2 inst_3538 ( .ZN(net_8246), .A2(net_8046), .A1(net_3287) );
CLKBUF_X2 inst_14984 ( .A(net_11433), .Z(net_14903) );
INV_X4 inst_5529 ( .A(net_9344), .ZN(net_1988) );
INV_X2 inst_7204 ( .A(net_9294), .ZN(net_470) );
AOI211_X2 inst_10250 ( .ZN(net_8810), .C2(net_8808), .C1(net_8803), .B(net_8628), .A(net_7907) );
INV_X4 inst_6103 ( .A(net_10001), .ZN(net_490) );
NAND2_X2 inst_3755 ( .ZN(net_5271), .A2(net_5266), .A1(net_2919) );
XNOR2_X2 inst_146 ( .ZN(net_7030), .B(net_7029), .A(net_6172) );
CLKBUF_X2 inst_15588 ( .A(net_15506), .Z(net_15507) );
DFF_X1 inst_8718 ( .QN(net_10241), .D(net_6291), .CK(net_10922) );
AOI221_X2 inst_9810 ( .B1(net_9961), .A(net_7090), .B2(net_7089), .C2(net_7088), .ZN(net_6992), .C1(net_6813) );
NAND2_X2 inst_3999 ( .ZN(net_4508), .A2(net_3390), .A1(net_1527) );
OAI22_X2 inst_1196 ( .A1(net_7249), .A2(net_5134), .B2(net_5133), .ZN(net_5057), .B1(net_1427) );
CLKBUF_X2 inst_12501 ( .A(net_11537), .Z(net_12420) );
CLKBUF_X2 inst_13815 ( .A(net_13191), .Z(net_13734) );
AND2_X2 inst_10589 ( .A2(net_4264), .A1(net_2417), .ZN(net_2390) );
OR2_X4 inst_817 ( .ZN(net_2142), .A2(net_947), .A1(net_780) );
XNOR2_X2 inst_326 ( .ZN(net_3008), .B(net_2806), .A(net_2063) );
CLKBUF_X2 inst_12550 ( .A(net_12468), .Z(net_12469) );
NAND2_X2 inst_3428 ( .A1(net_9479), .A2(net_8490), .ZN(net_8489) );
OAI211_X2 inst_2194 ( .C1(net_7229), .C2(net_6542), .ZN(net_6513), .B(net_5611), .A(net_3679) );
CLKBUF_X2 inst_10789 ( .A(net_10694), .Z(net_10708) );
AND2_X2 inst_10510 ( .ZN(net_4922), .A1(net_4921), .A2(net_4920) );
NAND2_X4 inst_3336 ( .A2(net_9027), .A1(net_9026), .ZN(net_8935) );
DFF_X2 inst_7963 ( .QN(net_10208), .D(net_5624), .CK(net_15589) );
AOI22_X2 inst_9034 ( .B2(net_10171), .ZN(net_7623), .A2(net_7491), .A1(net_7410), .B1(net_881) );
NAND3_X2 inst_3293 ( .A2(net_10070), .A3(net_4080), .A1(net_3630), .ZN(net_2746) );
CLKBUF_X2 inst_15825 ( .A(net_15743), .Z(net_15744) );
NAND2_X2 inst_3793 ( .A2(net_6319), .ZN(net_4731), .A1(net_922) );
NOR2_X2 inst_2837 ( .A2(net_2424), .ZN(net_2354), .A1(net_1513) );
INV_X2 inst_7115 ( .ZN(net_1256), .A(net_994) );
CLKBUF_X2 inst_11143 ( .A(net_10563), .Z(net_11062) );
OAI21_X2 inst_1845 ( .ZN(net_5988), .B2(net_5976), .A(net_2056), .B1(net_1372) );
XNOR2_X2 inst_108 ( .B(net_9429), .ZN(net_8115), .A(net_6293) );
NAND2_X2 inst_3778 ( .A2(net_9074), .ZN(net_4995), .A1(net_948) );
INV_X4 inst_4799 ( .A(net_3709), .ZN(net_3660) );
CLKBUF_X2 inst_14681 ( .A(net_11717), .Z(net_14600) );
AOI22_X2 inst_9296 ( .B1(net_10003), .A1(net_5743), .B2(net_5742), .ZN(net_5692), .A2(net_243) );
CLKBUF_X2 inst_15598 ( .A(net_15356), .Z(net_15517) );
INV_X2 inst_6905 ( .ZN(net_2253), .A(net_2252) );
NAND2_X2 inst_3940 ( .A1(net_9725), .ZN(net_3550), .A2(net_3039) );
INV_X4 inst_6503 ( .A(net_9615), .ZN(net_351) );
OAI222_X2 inst_1429 ( .ZN(net_3154), .C2(net_3153), .B2(net_3153), .A2(net_2317), .A1(net_2199), .B1(net_1006), .C1(net_788) );
DFF_X1 inst_8439 ( .D(net_8507), .CK(net_11108), .Q(x987) );
CLKBUF_X2 inst_11937 ( .A(net_11677), .Z(net_11856) );
SDFF_X2 inst_638 ( .Q(net_9440), .D(net_9440), .SE(net_3293), .CK(net_14159), .SI(x3133) );
DFF_X2 inst_7786 ( .Q(net_9820), .D(net_6510), .CK(net_13414) );
AOI211_X2 inst_10311 ( .C1(net_2984), .ZN(net_2566), .A(net_2565), .B(net_2564), .C2(net_1263) );
CLKBUF_X2 inst_12919 ( .A(net_12463), .Z(net_12838) );
SDFF_X2 inst_586 ( .Q(net_9254), .SE(net_4589), .D(net_137), .SI(net_103), .CK(net_13838) );
INV_X4 inst_5220 ( .ZN(net_2751), .A(net_1509) );
AOI221_X2 inst_9828 ( .B1(net_9872), .B2(net_9101), .A(net_6945), .C1(net_6944), .ZN(net_6917), .C2(net_243) );
INV_X2 inst_7176 ( .A(net_10267), .ZN(net_727) );
AND2_X2 inst_10563 ( .A1(net_4019), .ZN(net_3082), .A2(net_2225) );
NOR2_X2 inst_2591 ( .ZN(net_7386), .A2(net_7161), .A1(net_7018) );
AOI22_X2 inst_9237 ( .A1(net_9936), .B1(net_9837), .B2(net_6129), .A2(net_6111), .ZN(net_6074) );
NAND3_X2 inst_3275 ( .ZN(net_4094), .A1(net_3621), .A2(net_3450), .A3(net_2703) );
INV_X4 inst_5008 ( .A(net_2544), .ZN(net_2165) );
CLKBUF_X2 inst_15317 ( .A(net_14881), .Z(net_15236) );
OAI221_X2 inst_1466 ( .ZN(net_7885), .B1(net_7884), .B2(net_7710), .C2(net_7525), .A(net_5170), .C1(net_1314) );
NOR2_X2 inst_2841 ( .ZN(net_2331), .A2(net_2330), .A1(net_1335) );
OAI21_X2 inst_1726 ( .ZN(net_8797), .A(net_8796), .B1(net_7649), .B2(net_7605) );
INV_X2 inst_7157 ( .A(net_4157), .ZN(net_698) );
CLKBUF_X2 inst_15591 ( .A(net_15509), .Z(net_15510) );
NOR2_X2 inst_2652 ( .ZN(net_5892), .A2(net_5329), .A1(net_2107) );
INV_X4 inst_5221 ( .ZN(net_1811), .A(net_807) );
OAI22_X2 inst_1203 ( .A1(net_7241), .A2(net_5134), .B2(net_5133), .ZN(net_5048), .B1(net_1933) );
CLKBUF_X2 inst_14251 ( .A(net_14169), .Z(net_14170) );
OR2_X4 inst_802 ( .ZN(net_2145), .A2(net_1380), .A1(net_1364) );
XNOR2_X2 inst_296 ( .B(net_9107), .ZN(net_3561), .A(net_2948) );
INV_X2 inst_7118 ( .A(net_10352), .ZN(net_960) );
CLKBUF_X2 inst_14626 ( .A(net_14544), .Z(net_14545) );
CLKBUF_X2 inst_14576 ( .A(net_14494), .Z(net_14495) );
CLKBUF_X2 inst_10892 ( .A(net_10794), .Z(net_10811) );
OR2_X2 inst_905 ( .ZN(net_4636), .A1(net_4635), .A2(net_4454) );
CLKBUF_X2 inst_14677 ( .A(net_11729), .Z(net_14596) );
CLKBUF_X2 inst_11571 ( .A(net_11489), .Z(net_11490) );
NAND2_X2 inst_4370 ( .A2(net_2928), .ZN(net_2101), .A1(net_892) );
CLKBUF_X2 inst_14860 ( .A(net_14778), .Z(net_14779) );
CLKBUF_X2 inst_11218 ( .A(net_11136), .Z(net_11137) );
AOI22_X2 inst_9185 ( .A1(net_9875), .B1(net_9776), .A2(net_8042), .ZN(net_6130), .B2(net_6129) );
NAND2_X2 inst_4214 ( .ZN(net_2168), .A2(net_1719), .A1(net_1181) );
CLKBUF_X2 inst_12753 ( .A(net_12671), .Z(net_12672) );
CLKBUF_X2 inst_11047 ( .A(net_10965), .Z(net_10966) );
NAND2_X2 inst_3834 ( .ZN(net_4452), .A1(net_4328), .A2(net_4014) );
NAND2_X2 inst_3943 ( .A2(net_4071), .ZN(net_4016), .A1(net_2617) );
NAND2_X2 inst_3651 ( .ZN(net_6666), .A2(net_6665), .A1(net_2677) );
CLKBUF_X2 inst_14280 ( .A(net_14198), .Z(net_14199) );
OAI21_X2 inst_1759 ( .ZN(net_8453), .A(net_8374), .B2(net_8373), .B1(net_3984) );
CLKBUF_X2 inst_11792 ( .A(net_11550), .Z(net_11711) );
NOR2_X2 inst_2615 ( .A1(net_8117), .ZN(net_7048), .A2(net_6231) );
NOR2_X2 inst_2532 ( .A2(net_9592), .A1(net_9077), .ZN(net_8319) );
INV_X4 inst_5485 ( .A(net_10254), .ZN(net_4601) );
CLKBUF_X2 inst_13859 ( .A(net_12374), .Z(net_13778) );
CLKBUF_X2 inst_13263 ( .A(net_13181), .Z(net_13182) );
NAND2_X2 inst_3463 ( .A1(net_9491), .ZN(net_8460), .A2(net_8417) );
NOR2_X4 inst_2463 ( .A2(net_9009), .A1(net_9008), .ZN(net_8739) );
INV_X2 inst_7017 ( .ZN(net_1550), .A(net_1549) );
CLKBUF_X2 inst_11206 ( .A(net_10985), .Z(net_11125) );
CLKBUF_X2 inst_10907 ( .A(net_10825), .Z(net_10826) );
DFF_X2 inst_7617 ( .Q(net_10070), .D(net_6966), .CK(net_10844) );
CLKBUF_X2 inst_12492 ( .A(net_11710), .Z(net_12411) );
CLKBUF_X2 inst_11115 ( .A(net_10747), .Z(net_11034) );
INV_X4 inst_5610 ( .A(net_3261), .ZN(net_3065) );
INV_X4 inst_6375 ( .ZN(net_641), .A(net_171) );
NAND2_X2 inst_4055 ( .ZN(net_3236), .A2(net_2804), .A1(net_2666) );
OAI221_X2 inst_1464 ( .C1(net_8116), .B2(net_7974), .C2(net_7973), .ZN(net_7956), .A(net_7955), .B1(net_3053) );
OAI22_X2 inst_1247 ( .B1(net_7231), .ZN(net_4843), .A2(net_4842), .B2(net_4841), .A1(net_475) );
CLKBUF_X2 inst_15536 ( .A(net_15454), .Z(net_15455) );
CLKBUF_X2 inst_12778 ( .A(net_12696), .Z(net_12697) );
INV_X4 inst_5284 ( .A(net_6633), .ZN(net_3352) );
DFF_X1 inst_8490 ( .Q(net_9623), .D(net_7920), .CK(net_15116) );
INV_X4 inst_5031 ( .A(net_7583), .ZN(net_2173) );
CLKBUF_X2 inst_13275 ( .A(net_11068), .Z(net_13194) );
CLKBUF_X2 inst_14541 ( .A(net_14459), .Z(net_14460) );
CLKBUF_X2 inst_13498 ( .A(net_13416), .Z(net_13417) );
CLKBUF_X2 inst_13215 ( .A(net_11636), .Z(net_13134) );
OAI221_X2 inst_1493 ( .B1(net_10412), .C2(net_9063), .B2(net_9056), .ZN(net_7370), .C1(net_7192), .A(net_6992) );
INV_X4 inst_6441 ( .A(net_9977), .ZN(net_378) );
OAI22_X2 inst_1308 ( .ZN(net_2407), .A1(net_2406), .B2(net_2405), .B1(net_2205), .A2(net_1604) );
NAND4_X2 inst_3070 ( .ZN(net_5406), .A4(net_4970), .A1(net_4038), .A2(net_3812), .A3(net_3811) );
XNOR2_X2 inst_85 ( .ZN(net_8618), .A(net_8582), .B(net_8267) );
INV_X4 inst_4733 ( .ZN(net_4589), .A(net_4297) );
NOR2_X2 inst_2998 ( .A1(net_10116), .ZN(net_2134), .A2(net_631) );
CLKBUF_X2 inst_11734 ( .A(net_11652), .Z(net_11653) );
CLKBUF_X2 inst_15623 ( .A(net_15541), .Z(net_15542) );
CLKBUF_X2 inst_14116 ( .A(net_11553), .Z(net_14035) );
CLKBUF_X2 inst_13348 ( .A(net_13266), .Z(net_13267) );
NOR2_X2 inst_2612 ( .A1(net_8057), .ZN(net_7057), .A2(net_6241) );
INV_X4 inst_5963 ( .ZN(net_4033), .A(net_118) );
CLKBUF_X2 inst_14693 ( .A(net_14611), .Z(net_14612) );
AOI222_X1 inst_9681 ( .B1(net_9509), .A2(net_8310), .B2(net_8309), .C2(net_8308), .ZN(net_8306), .C1(net_8230), .A1(x2477) );
CLKBUF_X2 inst_11850 ( .A(net_11768), .Z(net_11769) );
CLKBUF_X2 inst_12598 ( .A(net_12516), .Z(net_12517) );
CLKBUF_X2 inst_11314 ( .A(net_11106), .Z(net_11233) );
NAND2_X2 inst_4022 ( .A1(net_7336), .ZN(net_7115), .A2(net_3071) );
OAI222_X2 inst_1362 ( .B1(net_7665), .A2(net_7664), .C2(net_7663), .ZN(net_6331), .B2(net_5398), .A1(net_4060), .C1(net_1920) );
CLKBUF_X2 inst_13798 ( .A(net_12118), .Z(net_13717) );
CLKBUF_X2 inst_12888 ( .A(net_12806), .Z(net_12807) );
DFF_X1 inst_8881 ( .Q(net_91), .CK(net_14108), .D(x3507) );
OAI21_X2 inst_1978 ( .ZN(net_2879), .A(net_2878), .B1(net_2243), .B2(net_1345) );
XNOR2_X2 inst_290 ( .B(net_4929), .ZN(net_3521), .A(net_3020) );
CLKBUF_X2 inst_15285 ( .A(net_11948), .Z(net_15204) );
CLKBUF_X2 inst_14311 ( .A(net_14229), .Z(net_14230) );
XNOR2_X2 inst_272 ( .ZN(net_3954), .A(net_3953), .B(net_1994) );
INV_X4 inst_4718 ( .ZN(net_5256), .A(net_4982) );
CLKBUF_X2 inst_14122 ( .A(net_14040), .Z(net_14041) );
OAI211_X2 inst_2112 ( .C2(net_6778), .ZN(net_6736), .A(net_6364), .B(net_6096), .C1(net_444) );
DFF_X2 inst_7743 ( .QN(net_10152), .D(net_6302), .CK(net_11250) );
CLKBUF_X2 inst_15431 ( .A(net_15349), .Z(net_15350) );
NAND4_X2 inst_3036 ( .A4(net_9581), .A2(net_9580), .ZN(net_8789), .A3(net_8780), .A1(net_8600) );
OR2_X4 inst_814 ( .A2(net_10369), .ZN(net_2381), .A1(net_1365) );
CLKBUF_X2 inst_13441 ( .A(net_13359), .Z(net_13360) );
AOI22_X2 inst_9465 ( .B1(net_10006), .A2(net_6442), .ZN(net_3862), .B2(net_2468), .A1(net_1262) );
AOI22_X2 inst_9213 ( .A1(net_9905), .B1(net_9806), .B2(net_6120), .A2(net_6111), .ZN(net_6098) );
INV_X4 inst_5203 ( .A(net_10351), .ZN(net_3177) );
NAND2_X2 inst_3471 ( .A1(net_9440), .A2(net_8952), .ZN(net_8436) );
OAI221_X2 inst_1458 ( .B2(net_7974), .C2(net_7973), .ZN(net_7968), .A(net_7967), .C1(net_7845), .B1(net_2584) );
NAND2_X2 inst_4133 ( .ZN(net_3722), .A1(net_1891), .A2(net_1011) );
CLKBUF_X2 inst_15177 ( .A(net_15095), .Z(net_15096) );
CLKBUF_X2 inst_11332 ( .A(net_10932), .Z(net_11251) );
OAI211_X2 inst_2275 ( .C1(net_7124), .C2(net_6548), .ZN(net_6236), .B(net_5757), .A(net_3507) );
OAI21_X2 inst_1860 ( .B2(net_10343), .ZN(net_5783), .A(net_2716), .B1(net_1523) );
OAI21_X2 inst_1810 ( .ZN(net_7033), .A(net_6892), .B1(net_6207), .B2(net_5962) );
OAI21_X2 inst_1806 ( .ZN(net_7394), .B2(net_7060), .A(net_5363), .B1(net_5362) );
OR2_X4 inst_789 ( .ZN(net_3073), .A2(net_1962), .A1(net_791) );
CLKBUF_X2 inst_15561 ( .A(net_15479), .Z(net_15480) );
CLKBUF_X2 inst_15727 ( .A(net_14291), .Z(net_15646) );
OAI21_X2 inst_1885 ( .ZN(net_4961), .B1(net_4959), .B2(net_4958), .A(net_1470) );
CLKBUF_X2 inst_13232 ( .A(net_13150), .Z(net_13151) );
AOI21_X2 inst_10212 ( .ZN(net_2433), .B1(net_2432), .B2(net_2186), .A(net_640) );
CLKBUF_X2 inst_11184 ( .A(net_11102), .Z(net_11103) );
DFF_X2 inst_7926 ( .QN(net_10330), .D(net_5494), .CK(net_14367) );
OR2_X4 inst_822 ( .A2(net_10355), .A1(net_10354), .ZN(net_1652) );
CLKBUF_X2 inst_14136 ( .A(net_14054), .Z(net_14055) );
CLKBUF_X2 inst_12053 ( .A(net_11971), .Z(net_11972) );
OAI22_X2 inst_1125 ( .A1(net_10534), .ZN(net_5156), .A2(net_5155), .B2(net_3984), .B1(net_354) );
NAND2_X2 inst_4341 ( .ZN(net_1743), .A2(net_1036), .A1(net_1035) );
INV_X4 inst_5996 ( .A(net_10116), .ZN(net_668) );
CLKBUF_X2 inst_13189 ( .A(net_13107), .Z(net_13108) );
INV_X4 inst_4885 ( .A(net_7586), .ZN(net_3910) );
CLKBUF_X2 inst_10984 ( .A(net_10902), .Z(net_10903) );
SDFF_X2 inst_609 ( .QN(net_10407), .D(net_4413), .SE(net_3673), .SI(net_750), .CK(net_10743) );
CLKBUF_X2 inst_11521 ( .A(net_11439), .Z(net_11440) );
DFF_X2 inst_8261 ( .Q(net_10288), .D(net_4820), .CK(net_14519) );
NOR2_X2 inst_2496 ( .ZN(net_8577), .A2(net_8568), .A1(net_8451) );
OR2_X4 inst_795 ( .A2(net_10258), .ZN(net_2147), .A1(net_1342) );
DFF_X2 inst_8393 ( .Q(net_9156), .CK(net_11804), .D(x3588) );
NOR2_X2 inst_2491 ( .ZN(net_8686), .A2(net_8685), .A1(net_3137) );
CLKBUF_X2 inst_13466 ( .A(net_13384), .Z(net_13385) );
CLKBUF_X2 inst_15158 ( .A(net_10564), .Z(net_15077) );
NAND2_X2 inst_4381 ( .A2(net_9233), .ZN(net_4328), .A1(net_463) );
INV_X2 inst_6668 ( .ZN(net_8360), .A(net_8303) );
CLKBUF_X2 inst_14127 ( .A(net_14045), .Z(net_14046) );
CLKBUF_X2 inst_11406 ( .A(net_11304), .Z(net_11325) );
CLKBUF_X2 inst_11179 ( .A(net_11097), .Z(net_11098) );
CLKBUF_X2 inst_12848 ( .A(net_12695), .Z(net_12767) );
CLKBUF_X2 inst_11280 ( .A(net_10971), .Z(net_11199) );
DFF_X2 inst_8215 ( .Q(net_10075), .D(net_4860), .CK(net_11096) );
DFF_X2 inst_8229 ( .Q(net_10287), .D(net_4804), .CK(net_14532) );
SDFF_X2 inst_619 ( .Q(net_9455), .D(net_9455), .SE(net_3293), .CK(net_11901), .SI(x2214) );
NOR2_X2 inst_2671 ( .ZN(net_4908), .A2(net_4907), .A1(net_2226) );
AOI22_X2 inst_9638 ( .A1(net_9840), .B1(net_9777), .A2(net_6413), .ZN(net_3404), .B2(net_2462) );
CLKBUF_X2 inst_14481 ( .A(net_14399), .Z(net_14400) );
CLKBUF_X2 inst_12139 ( .A(net_12057), .Z(net_12058) );
OAI221_X2 inst_1654 ( .C1(net_7216), .ZN(net_5521), .C2(net_5520), .B1(net_5009), .B2(net_4547), .A(net_3507) );
CLKBUF_X2 inst_14713 ( .A(net_14631), .Z(net_14632) );
CLKBUF_X2 inst_13068 ( .A(net_11368), .Z(net_12987) );
INV_X4 inst_4547 ( .A(net_8581), .ZN(net_8580) );
DFF_X2 inst_7831 ( .Q(net_9798), .D(net_6195), .CK(net_11961) );
OAI222_X2 inst_1355 ( .A1(net_7660), .B2(net_7659), .C2(net_7658), .ZN(net_7159), .A2(net_6649), .B1(net_4417), .C1(net_698) );
AND2_X2 inst_10545 ( .ZN(net_3963), .A2(net_3488), .A1(net_2366) );
OR2_X2 inst_877 ( .ZN(net_6613), .A1(net_6423), .A2(net_5957) );
INV_X4 inst_6612 ( .A(net_8924), .ZN(net_8923) );
AND2_X2 inst_10553 ( .ZN(net_3339), .A2(net_3338), .A1(net_3320) );
AOI211_X2 inst_10267 ( .ZN(net_7705), .A(net_7704), .C2(net_7599), .C1(net_4627), .B(x3390) );
CLKBUF_X2 inst_10704 ( .A(net_10622), .Z(net_10623) );
INV_X4 inst_6563 ( .A(net_10149), .ZN(net_683) );
CLKBUF_X2 inst_12698 ( .A(net_11486), .Z(net_12617) );
DFF_X2 inst_7372 ( .D(net_8688), .QN(net_255), .CK(net_15090) );
AOI211_X2 inst_10265 ( .ZN(net_7756), .B(net_7645), .C2(net_7621), .A(net_3298), .C1(net_2263) );
INV_X4 inst_6486 ( .A(net_10197), .ZN(net_359) );
OAI211_X2 inst_2076 ( .C2(net_6774), .ZN(net_6772), .A(net_6367), .B(net_6134), .C1(net_395) );
INV_X4 inst_5879 ( .ZN(net_2607), .A(net_625) );
INV_X4 inst_6384 ( .A(net_9749), .ZN(net_394) );
NOR2_X4 inst_2481 ( .A2(net_2139), .ZN(net_1786), .A1(net_959) );
DFF_X2 inst_7824 ( .Q(net_9651), .D(net_6179), .CK(net_14093) );
CLKBUF_X2 inst_14523 ( .A(net_14441), .Z(net_14442) );
CLKBUF_X2 inst_11474 ( .A(net_11392), .Z(net_11393) );
INV_X4 inst_5829 ( .ZN(net_909), .A(net_665) );
CLKBUF_X2 inst_13385 ( .A(net_10988), .Z(net_13304) );
NAND2_X2 inst_4285 ( .A1(net_9247), .ZN(net_1711), .A2(net_1340) );
CLKBUF_X2 inst_15386 ( .A(net_15304), .Z(net_15305) );
OAI22_X2 inst_1162 ( .A1(net_7211), .A2(net_5139), .B2(net_5138), .ZN(net_5111), .B1(net_401) );
AOI211_X2 inst_10274 ( .ZN(net_7528), .B(net_7251), .A(net_5172), .C1(net_4626), .C2(net_4209) );
INV_X4 inst_5904 ( .ZN(net_4978), .A(net_596) );
DFF_X2 inst_7485 ( .Q(net_9276), .D(net_8075), .CK(net_13129) );
CLKBUF_X2 inst_14384 ( .A(net_14302), .Z(net_14303) );
INV_X4 inst_6108 ( .A(net_10373), .ZN(net_7025) );
INV_X4 inst_6572 ( .A(net_10502), .ZN(net_4100) );
CLKBUF_X2 inst_13123 ( .A(net_13041), .Z(net_13042) );
DFF_X2 inst_7449 ( .QN(net_9295), .D(net_8248), .CK(net_14994) );
CLKBUF_X2 inst_10734 ( .A(net_10561), .Z(net_10653) );
NOR2_X2 inst_2973 ( .ZN(net_1564), .A1(net_484), .A2(net_433) );
CLKBUF_X2 inst_11013 ( .A(net_10931), .Z(net_10932) );
CLKBUF_X2 inst_11454 ( .A(net_11372), .Z(net_11373) );
OAI222_X2 inst_1433 ( .A1(net_2649), .ZN(net_2456), .C2(net_2455), .B2(net_2455), .A2(net_2028), .B1(net_992), .C1(net_586) );
OR2_X4 inst_793 ( .A1(net_10262), .ZN(net_2189), .A2(net_1382) );
AOI22_X2 inst_9206 ( .A1(net_9866), .B1(net_9767), .B2(net_6120), .A2(net_6109), .ZN(net_6105) );
OAI21_X2 inst_1894 ( .B1(net_7108), .B2(net_4862), .ZN(net_4858), .A(net_4530) );
CLKBUF_X2 inst_13960 ( .A(net_13878), .Z(net_13879) );
INV_X4 inst_4815 ( .ZN(net_4206), .A(net_3543) );
CLKBUF_X2 inst_15401 ( .A(net_10965), .Z(net_15320) );
INV_X2 inst_6707 ( .ZN(net_8147), .A(net_8146) );
OAI21_X2 inst_1999 ( .B1(net_10324), .ZN(net_2300), .A(net_2299), .B2(net_2298) );
INV_X4 inst_4643 ( .ZN(net_6025), .A(net_5844) );
CLKBUF_X2 inst_14379 ( .A(net_14297), .Z(net_14298) );
NOR2_X2 inst_2733 ( .ZN(net_4202), .A1(net_3712), .A2(net_3711) );
CLKBUF_X2 inst_12405 ( .A(net_11468), .Z(net_12324) );
CLKBUF_X2 inst_11750 ( .A(net_11668), .Z(net_11669) );
INV_X4 inst_6636 ( .A(net_9059), .ZN(net_9058) );
CLKBUF_X2 inst_15429 ( .A(net_15347), .Z(net_15348) );
CLKBUF_X2 inst_13677 ( .A(net_13595), .Z(net_13596) );
DFF_X1 inst_8808 ( .QN(net_9189), .D(net_3518), .CK(net_13608) );
SDFF_X2 inst_475 ( .SE(net_9540), .SI(net_8234), .Q(net_291), .D(net_291), .CK(net_11724) );
CLKBUF_X2 inst_13253 ( .A(net_11571), .Z(net_13172) );
AOI22_X2 inst_9436 ( .ZN(net_4638), .A2(net_4361), .B2(net_3604), .A1(net_1121), .B1(net_955) );
INV_X4 inst_4738 ( .ZN(net_4779), .A(net_4461) );
AOI22_X2 inst_9412 ( .A1(net_9953), .B1(net_6834), .ZN(net_4735), .A2(net_4734), .B2(net_4733) );
NOR2_X2 inst_2701 ( .A2(net_10481), .ZN(net_4389), .A1(net_2255) );
NAND2_X2 inst_4412 ( .A2(net_10226), .A1(net_10225), .ZN(net_2093) );
AOI22_X2 inst_9171 ( .A1(net_9911), .B1(net_9812), .A2(net_8042), .B2(net_8041), .ZN(net_6147) );
DFF_X2 inst_8321 ( .Q(net_10293), .D(net_3929), .CK(net_14500) );
CLKBUF_X2 inst_12595 ( .A(net_12513), .Z(net_12514) );
AND2_X4 inst_10385 ( .A2(net_9587), .ZN(net_8754), .A1(net_1320) );
NAND4_X2 inst_3165 ( .ZN(net_990), .A4(net_116), .A3(net_115), .A2(net_114), .A1(net_113) );
AOI22_X2 inst_9564 ( .B1(net_10035), .A1(net_9872), .B2(net_5174), .ZN(net_3755), .A2(net_2973) );
CLKBUF_X2 inst_12804 ( .A(net_12722), .Z(net_12723) );
CLKBUF_X2 inst_11222 ( .A(net_10999), .Z(net_11141) );
CLKBUF_X2 inst_15573 ( .A(net_15491), .Z(net_15492) );
SDFF_X2 inst_575 ( .D(net_9574), .SI(net_2569), .SE(net_758), .Q(net_248), .CK(net_11570) );
CLKBUF_X2 inst_11738 ( .A(net_11656), .Z(net_11657) );
INV_X4 inst_5724 ( .ZN(net_1094), .A(net_760) );
AOI21_X2 inst_10151 ( .ZN(net_4150), .B2(net_4149), .B1(net_4088), .A(net_3696) );
DFF_X2 inst_8276 ( .Q(net_9756), .D(net_4739), .CK(net_15415) );
NAND2_X2 inst_4331 ( .A2(net_10230), .ZN(net_2185), .A1(net_1115) );
CLKBUF_X2 inst_11054 ( .A(net_10972), .Z(net_10973) );
DFF_X2 inst_8049 ( .QN(net_9551), .D(net_9257), .CK(net_13754) );
INV_X4 inst_4705 ( .A(net_6678), .ZN(net_5345) );
CLKBUF_X2 inst_14606 ( .A(net_11261), .Z(net_14525) );
CLKBUF_X2 inst_10940 ( .A(net_10858), .Z(net_10859) );
SDFF_X2 inst_627 ( .Q(net_9458), .D(net_9458), .SE(net_3293), .CK(net_11899), .SI(x2027) );
INV_X4 inst_4725 ( .ZN(net_4613), .A(net_4492) );
INV_X2 inst_6831 ( .ZN(net_4012), .A(net_4011) );
NAND2_X4 inst_3352 ( .A2(net_9444), .A1(net_9016), .ZN(net_9013) );
XNOR2_X2 inst_344 ( .ZN(net_2864), .A(net_1872), .B(net_1491) );
CLKBUF_X2 inst_11543 ( .A(net_11461), .Z(net_11462) );
INV_X2 inst_6928 ( .A(net_2681), .ZN(net_1954) );
NAND2_X2 inst_3580 ( .ZN(net_7547), .A2(net_7119), .A1(net_2419) );
NAND2_X2 inst_3818 ( .A1(net_10087), .A2(net_4534), .ZN(net_4520) );
CLKBUF_X2 inst_15209 ( .A(net_14341), .Z(net_15128) );
CLKBUF_X2 inst_12321 ( .A(net_10575), .Z(net_12240) );
INV_X4 inst_5975 ( .A(net_10477), .ZN(net_694) );
OAI222_X2 inst_1338 ( .A1(net_7728), .B2(net_7727), .C2(net_7726), .ZN(net_7627), .A2(net_7471), .B1(net_4987), .C1(net_1896) );
CLKBUF_X2 inst_11531 ( .A(net_11351), .Z(net_11450) );
AOI21_X2 inst_10004 ( .B2(net_9570), .ZN(net_8793), .B1(net_4297), .A(net_3365) );
NOR3_X2 inst_2430 ( .ZN(net_4560), .A3(net_3382), .A1(net_3187), .A2(net_2963) );
NAND4_X2 inst_3080 ( .ZN(net_4704), .A4(net_4278), .A1(net_3846), .A2(net_3463), .A3(net_3402) );
INV_X2 inst_6857 ( .A(net_4460), .ZN(net_3335) );
CLKBUF_X2 inst_13093 ( .A(net_13011), .Z(net_13012) );
NOR3_X2 inst_2434 ( .A3(net_9622), .ZN(net_3504), .A1(net_3503), .A2(net_731) );
INV_X4 inst_4952 ( .A(net_4714), .ZN(net_2559) );
DFF_X2 inst_7432 ( .QN(net_9412), .D(net_8353), .CK(net_13930) );
NAND2_X2 inst_3731 ( .A1(net_10300), .ZN(net_5537), .A2(net_5536) );
OAI22_X2 inst_1107 ( .A1(net_7219), .ZN(net_6152), .B2(net_5879), .A2(net_5303), .B1(net_3945) );
CLKBUF_X2 inst_13932 ( .A(net_13850), .Z(net_13851) );
AOI21_X2 inst_10039 ( .ZN(net_7722), .B1(net_7640), .B2(net_7588), .A(net_4371) );
INV_X2 inst_6899 ( .A(net_7895), .ZN(net_2506) );
CLKBUF_X2 inst_15364 ( .A(net_13590), .Z(net_15283) );
OAI211_X2 inst_2028 ( .ZN(net_8374), .B(net_8373), .C2(net_8156), .C1(net_4515), .A(x962) );
INV_X4 inst_4839 ( .ZN(net_3526), .A(net_3378) );
CLKBUF_X2 inst_15335 ( .A(net_11853), .Z(net_15254) );
CLKBUF_X2 inst_12909 ( .A(net_12827), .Z(net_12828) );
INV_X4 inst_5930 ( .ZN(net_814), .A(net_576) );
AOI221_X2 inst_9916 ( .B1(net_10510), .ZN(net_6416), .B2(net_6415), .C1(net_6414), .C2(net_6413), .A(net_5688) );
DFF_X2 inst_8381 ( .QN(net_10094), .D(net_10093), .CK(net_11167) );
CLKBUF_X2 inst_15038 ( .A(net_14956), .Z(net_14957) );
CLKBUF_X2 inst_14904 ( .A(net_14822), .Z(net_14823) );
NAND2_X2 inst_4253 ( .A2(net_9172), .ZN(net_1836), .A1(net_911) );
NOR2_X2 inst_2776 ( .ZN(net_3595), .A2(net_3390), .A1(net_3172) );
OR2_X4 inst_722 ( .ZN(net_8427), .A2(net_8426), .A1(net_8405) );
AOI22_X2 inst_9646 ( .A1(net_2651), .ZN(net_2577), .B2(net_2576), .A2(net_1615), .B1(net_828) );
DFF_X1 inst_8612 ( .Q(net_9778), .D(net_7185), .CK(net_15564) );
OR2_X4 inst_746 ( .A1(net_9227), .ZN(net_5927), .A2(net_5361) );
INV_X4 inst_6019 ( .A(net_10157), .ZN(net_557) );
DFF_X2 inst_8093 ( .QN(net_10041), .D(net_5088), .CK(net_12507) );
CLKBUF_X2 inst_13016 ( .A(net_11968), .Z(net_12935) );
INV_X4 inst_6553 ( .A(net_9546), .ZN(net_8184) );
AOI22_X2 inst_9502 ( .B1(net_10390), .A1(net_9888), .B2(net_4062), .ZN(net_3821), .A2(net_2973) );
NAND2_X2 inst_4232 ( .A2(net_9039), .A1(net_6949), .ZN(net_2724) );
DFF_X1 inst_8660 ( .Q(net_9789), .D(net_7215), .CK(net_13341) );
OAI211_X2 inst_2267 ( .C1(net_7139), .C2(net_6501), .ZN(net_6278), .B(net_5698), .A(net_3679) );
NAND2_X2 inst_4270 ( .A2(net_10247), .ZN(net_1634), .A1(net_1015) );
NOR2_X2 inst_3010 ( .A2(net_9216), .ZN(net_837), .A1(net_836) );
DFF_X2 inst_8010 ( .QN(net_10433), .D(net_5497), .CK(net_13716) );
INV_X2 inst_7127 ( .A(net_1093), .ZN(net_893) );
CLKBUF_X2 inst_12282 ( .A(net_10585), .Z(net_12201) );
DFF_X2 inst_8207 ( .Q(net_10074), .D(net_4861), .CK(net_11098) );
NAND4_X2 inst_3133 ( .ZN(net_5335), .A4(net_5272), .A2(net_2918), .A3(net_2917), .A1(net_799) );
INV_X4 inst_5662 ( .A(net_10156), .ZN(net_2624) );
INV_X4 inst_6412 ( .A(net_10433), .ZN(net_643) );
DFF_X2 inst_7893 ( .QN(net_10099), .D(net_6021), .CK(net_15521) );
AOI21_X2 inst_10050 ( .ZN(net_7311), .A(net_7310), .B2(net_7078), .B1(net_1921) );
INV_X4 inst_5820 ( .A(net_2000), .ZN(net_673) );
DFF_X1 inst_8721 ( .QN(net_10486), .D(net_6268), .CK(net_13738) );
OAI221_X2 inst_1577 ( .B1(net_10212), .B2(net_7295), .C2(net_7293), .ZN(net_7140), .C1(net_7139), .A(net_6924) );
DFF_X2 inst_7722 ( .Q(net_9704), .D(net_6248), .CK(net_15607) );
NOR2_X2 inst_2588 ( .ZN(net_7051), .A1(net_7050), .A2(net_6614) );
OAI22_X2 inst_1110 ( .A1(net_7219), .ZN(net_6149), .B1(net_6148), .B2(net_5872), .A2(net_5301) );
INV_X4 inst_5778 ( .ZN(net_1708), .A(net_708) );
INV_X4 inst_6547 ( .A(net_9748), .ZN(net_3945) );
CLKBUF_X2 inst_14870 ( .A(net_11131), .Z(net_14789) );
NOR2_X2 inst_2873 ( .ZN(net_3594), .A2(net_3172), .A1(net_1949) );
DFF_X2 inst_7724 ( .Q(net_9805), .D(net_6280), .CK(net_12568) );
INV_X2 inst_6994 ( .A(net_2889), .ZN(net_1636) );
INV_X4 inst_4665 ( .A(net_6041), .ZN(net_5442) );
DFF_X1 inst_8468 ( .Q(net_9598), .D(net_7972), .CK(net_11520) );
NOR3_X2 inst_2442 ( .A3(net_9279), .A2(net_5331), .ZN(net_2890), .A1(net_2889) );
CLKBUF_X2 inst_15379 ( .A(net_13760), .Z(net_15298) );
AOI222_X1 inst_9676 ( .B2(net_9577), .A1(net_9576), .ZN(net_8624), .A2(net_8602), .C2(net_8601), .B1(net_1971), .C1(net_1384) );
OAI211_X2 inst_2066 ( .ZN(net_7753), .B(net_7509), .A(net_7441), .C1(net_7336), .C2(net_564) );
CLKBUF_X2 inst_12126 ( .A(net_12044), .Z(net_12045) );
INV_X4 inst_5712 ( .ZN(net_1050), .A(net_771) );
OAI21_X2 inst_1742 ( .ZN(net_8692), .B1(net_8691), .B2(net_8672), .A(net_7854) );
MUX2_X1 inst_4466 ( .S(net_6041), .A(net_6040), .B(x6198), .Z(x316) );
INV_X4 inst_5374 ( .ZN(net_1566), .A(net_1063) );
INV_X4 inst_5562 ( .ZN(net_3853), .A(net_919) );
CLKBUF_X2 inst_15543 ( .A(net_15461), .Z(net_15462) );
CLKBUF_X2 inst_12085 ( .A(net_12003), .Z(net_12004) );
CLKBUF_X2 inst_11058 ( .A(net_10976), .Z(net_10977) );
CLKBUF_X2 inst_13603 ( .A(net_11286), .Z(net_13522) );
CLKBUF_X2 inst_12091 ( .A(net_11880), .Z(net_12010) );
CLKBUF_X2 inst_11035 ( .A(net_10953), .Z(net_10954) );
INV_X4 inst_6236 ( .A(net_9742), .ZN(net_460) );
DFF_X1 inst_8447 ( .Q(net_9431), .D(net_8143), .CK(net_14930) );
NOR2_X2 inst_2875 ( .ZN(net_2648), .A2(net_1947), .A1(net_860) );
INV_X4 inst_4779 ( .ZN(net_8012), .A(net_4135) );
AOI22_X2 inst_9522 ( .A1(net_9868), .B2(net_5174), .ZN(net_3800), .B1(net_3799), .A2(net_2973) );
AOI22_X2 inst_9067 ( .B1(net_9687), .A2(net_6684), .B2(net_6683), .ZN(net_6599), .A1(net_256) );
CLKBUF_X2 inst_11084 ( .A(net_10769), .Z(net_11003) );
AND4_X2 inst_10341 ( .A2(net_9355), .A1(net_9354), .A4(net_7530), .ZN(net_6202), .A3(net_5786) );
INV_X2 inst_7162 ( .A(net_1774), .ZN(net_910) );
AOI22_X2 inst_9396 ( .B1(net_9708), .A1(net_5755), .B2(net_5754), .ZN(net_5404), .A2(net_245) );
NAND3_X2 inst_3175 ( .ZN(net_8495), .A1(net_8425), .A2(net_8423), .A3(net_8331) );
NOR4_X2 inst_2302 ( .A4(net_9583), .A3(net_9579), .ZN(net_8791), .A1(net_8789), .A2(net_8575) );
CLKBUF_X2 inst_11021 ( .A(net_10939), .Z(net_10940) );
NAND2_X2 inst_3389 ( .ZN(net_8751), .A2(net_8738), .A1(net_1671) );
INV_X4 inst_6248 ( .A(net_9225), .ZN(net_456) );
AOI221_X2 inst_9967 ( .C1(net_9989), .B1(net_9755), .B2(net_6442), .ZN(net_4761), .A(net_4351), .C2(net_2541) );
INV_X2 inst_7181 ( .ZN(net_521), .A(x3867) );
NOR3_X2 inst_2447 ( .ZN(net_2714), .A1(net_2713), .A2(net_711), .A3(net_462) );
OR2_X4 inst_782 ( .A1(net_2963), .ZN(net_2765), .A2(net_2540) );
INV_X4 inst_5744 ( .ZN(net_1362), .A(net_1209) );
CLKBUF_X2 inst_12043 ( .A(net_11014), .Z(net_11962) );
NOR2_X2 inst_2869 ( .A1(net_2049), .ZN(net_2027), .A2(net_1694) );
AND2_X2 inst_10546 ( .ZN(net_3964), .A1(net_3487), .A2(net_3486) );
AND2_X2 inst_10603 ( .A2(net_4115), .ZN(net_2061), .A1(net_2060) );
XOR2_X2 inst_6 ( .B(net_9525), .Z(net_5198), .A(net_4427) );
NOR2_X2 inst_2486 ( .A2(net_8765), .ZN(net_8763), .A1(net_8762) );
CLKBUF_X2 inst_11648 ( .A(net_11325), .Z(net_11567) );
INV_X4 inst_5461 ( .A(net_1364), .ZN(net_1275) );
NOR3_X2 inst_2410 ( .A1(net_10537), .A3(net_10535), .ZN(net_6426), .A2(x1074) );
CLKBUF_X2 inst_15408 ( .A(net_15326), .Z(net_15327) );
CLKBUF_X2 inst_11151 ( .A(net_11069), .Z(net_11070) );
CLKBUF_X2 inst_11832 ( .A(net_11750), .Z(net_11751) );
CLKBUF_X2 inst_10914 ( .A(net_10832), .Z(net_10833) );
AOI222_X1 inst_9695 ( .B1(net_9506), .A2(net_8286), .B2(net_8285), .C2(net_8284), .ZN(net_8283), .C1(net_8218), .A1(x1660) );
DFF_X2 inst_7622 ( .QN(net_10160), .D(net_6930), .CK(net_13515) );
DFF_X1 inst_8728 ( .Q(net_9141), .D(net_6155), .CK(net_10985) );
INV_X4 inst_6141 ( .A(net_10326), .ZN(net_1948) );
DFF_X2 inst_7921 ( .Q(net_9222), .D(net_5920), .CK(net_13007) );
CLKBUF_X2 inst_13303 ( .A(net_10685), .Z(net_13222) );
INV_X2 inst_7163 ( .A(net_3988), .ZN(net_598) );
CLKBUF_X2 inst_12760 ( .A(net_12678), .Z(net_12679) );
INV_X4 inst_4803 ( .ZN(net_7535), .A(net_5575) );
OR2_X2 inst_935 ( .A1(net_9172), .ZN(net_2444), .A2(net_2442) );
CLKBUF_X2 inst_14650 ( .A(net_12641), .Z(net_14569) );
INV_X4 inst_6619 ( .ZN(net_8945), .A(net_8668) );
CLKBUF_X2 inst_11726 ( .A(net_11644), .Z(net_11645) );
INV_X4 inst_5699 ( .A(net_1143), .ZN(net_782) );
CLKBUF_X2 inst_13030 ( .A(net_12948), .Z(net_12949) );
INV_X4 inst_4772 ( .ZN(net_4296), .A(net_4120) );
CLKBUF_X2 inst_12781 ( .A(net_12699), .Z(net_12700) );
INV_X4 inst_4634 ( .ZN(net_7046), .A(net_6225) );
DFF_X2 inst_8211 ( .Q(net_10389), .D(net_4805), .CK(net_15225) );
DFF_X2 inst_8108 ( .QN(net_10043), .D(net_5086), .CK(net_12497) );
INV_X4 inst_6031 ( .ZN(net_1143), .A(net_265) );
CLKBUF_X2 inst_11255 ( .A(net_11173), .Z(net_11174) );
DFF_X2 inst_7729 ( .Q(net_9702), .D(net_6438), .CK(net_15057) );
AOI22_X2 inst_9284 ( .B1(net_9798), .A1(net_5766), .B2(net_5765), .ZN(net_5721), .A2(net_236) );
CLKBUF_X2 inst_11587 ( .A(net_11505), .Z(net_11506) );
NOR2_X2 inst_2944 ( .A2(net_9202), .A1(net_9201), .ZN(net_1814) );
OAI22_X2 inst_1320 ( .B2(net_9743), .ZN(net_2001), .A2(net_2000), .A1(net_1254), .B1(net_193) );
OAI22_X2 inst_1026 ( .A2(net_8036), .B2(net_8018), .ZN(net_7992), .A1(net_5252), .B1(net_443) );
CLKBUF_X2 inst_15638 ( .A(net_15556), .Z(net_15557) );
INV_X4 inst_5011 ( .ZN(net_2128), .A(net_1760) );
CLKBUF_X2 inst_11289 ( .A(net_11207), .Z(net_11208) );
INV_X4 inst_6250 ( .ZN(net_4183), .A(net_161) );
CLKBUF_X2 inst_12826 ( .A(net_11846), .Z(net_12745) );
INV_X4 inst_5576 ( .A(net_9735), .ZN(net_900) );
NAND2_X4 inst_3376 ( .ZN(net_9052), .A1(net_1715), .A2(net_564) );
XNOR2_X2 inst_95 ( .ZN(net_8493), .A(net_8394), .B(net_8371) );
INV_X4 inst_5246 ( .A(net_3204), .ZN(net_1866) );
CLKBUF_X2 inst_15830 ( .A(net_15748), .Z(net_15749) );
CLKBUF_X2 inst_15186 ( .A(net_13989), .Z(net_15105) );
NOR2_X2 inst_2921 ( .A2(net_4309), .ZN(net_3613), .A1(net_1396) );
CLKBUF_X2 inst_13690 ( .A(net_13572), .Z(net_13609) );
CLKBUF_X2 inst_13058 ( .A(net_12976), .Z(net_12977) );
AND2_X2 inst_10622 ( .A1(net_9279), .ZN(net_7887), .A2(net_652) );
AND2_X2 inst_10499 ( .ZN(net_7023), .A1(net_6587), .A2(net_6168) );
DFF_X2 inst_8314 ( .D(net_4049), .QN(net_280), .CK(net_12845) );
NOR2_X2 inst_2862 ( .ZN(net_2059), .A1(net_2058), .A2(net_1432) );
DFF_X2 inst_7949 ( .QN(net_10200), .D(net_5646), .CK(net_12032) );
CLKBUF_X2 inst_14794 ( .A(net_14712), .Z(net_14713) );
DFF_X2 inst_8391 ( .Q(net_10304), .D(net_10303), .CK(net_12101) );
NAND2_X2 inst_4009 ( .A1(net_9521), .ZN(net_3482), .A2(net_3035) );
CLKBUF_X2 inst_13397 ( .A(net_13315), .Z(net_13316) );
CLKBUF_X2 inst_10870 ( .A(net_10788), .Z(net_10789) );
AOI221_X2 inst_9766 ( .ZN(net_7591), .A(net_7450), .C1(net_5353), .C2(net_4908), .B1(net_4294), .B2(net_3509) );
CLKBUF_X2 inst_15109 ( .A(net_12138), .Z(net_15028) );
DFF_X2 inst_8071 ( .QN(net_9658), .D(net_5334), .CK(net_14952) );
DFF_X2 inst_8297 ( .Q(net_9855), .D(net_4615), .CK(net_15410) );
INV_X4 inst_4900 ( .A(net_7823), .ZN(net_4294) );
INV_X4 inst_6510 ( .A(net_10143), .ZN(net_1755) );
CLKBUF_X2 inst_13325 ( .A(net_13243), .Z(net_13244) );
INV_X4 inst_5808 ( .ZN(net_1966), .A(net_684) );
INV_X4 inst_5394 ( .A(net_6628), .ZN(net_3718) );
INV_X4 inst_5837 ( .ZN(net_1010), .A(net_657) );
INV_X2 inst_7194 ( .A(net_9418), .ZN(net_8216) );
CLKBUF_X2 inst_13883 ( .A(net_13801), .Z(net_13802) );
CLKBUF_X2 inst_12181 ( .A(net_12099), .Z(net_12100) );
CLKBUF_X2 inst_13390 ( .A(net_11837), .Z(net_13309) );
CLKBUF_X2 inst_11268 ( .A(net_11186), .Z(net_11187) );
INV_X2 inst_6859 ( .ZN(net_3326), .A(net_3119) );
DFF_X2 inst_7439 ( .QN(net_9397), .D(net_8333), .CK(net_11754) );
DFF_X2 inst_7537 ( .QN(net_9352), .D(net_7787), .CK(net_11475) );
AND2_X4 inst_10407 ( .ZN(net_4903), .A1(net_4902), .A2(net_4901) );
MUX2_X1 inst_4454 ( .S(net_6041), .A(net_292), .B(x5427), .Z(x182) );
CLKBUF_X2 inst_12369 ( .A(net_12287), .Z(net_12288) );
CLKBUF_X2 inst_14758 ( .A(net_14676), .Z(net_14677) );
INV_X4 inst_4901 ( .A(net_3160), .ZN(net_2855) );
CLKBUF_X2 inst_12813 ( .A(net_12731), .Z(net_12732) );
NAND2_X2 inst_3590 ( .ZN(net_7352), .A1(net_7047), .A2(net_6652) );
DFF_X1 inst_8709 ( .Q(net_9125), .D(net_6935), .CK(net_10584) );
NAND2_X2 inst_4315 ( .A2(net_10245), .ZN(net_1184), .A1(net_732) );
XNOR2_X2 inst_365 ( .B(net_9653), .ZN(net_2523), .A(net_2166) );
XNOR2_X2 inst_67 ( .ZN(net_8718), .A(net_8717), .B(net_6161) );
OAI33_X1 inst_954 ( .B3(net_9087), .A2(net_9075), .A3(net_8990), .ZN(net_7084), .B1(net_7083), .A1(net_7083), .B2(net_3067) );
CLKBUF_X2 inst_13162 ( .A(net_13080), .Z(net_13081) );
AOI22_X2 inst_9252 ( .A2(net_8042), .B2(net_8041), .ZN(net_6058), .A1(net_6057), .B1(net_6056) );
DFF_X2 inst_8145 ( .Q(net_10035), .D(net_5099), .CK(net_14279) );
INV_X4 inst_4974 ( .ZN(net_2313), .A(net_2312) );
CLKBUF_X2 inst_10836 ( .A(net_10754), .Z(net_10755) );
DFF_X1 inst_8582 ( .Q(net_9671), .D(net_7101), .CK(net_11628) );
CLKBUF_X2 inst_14186 ( .A(net_14104), .Z(net_14105) );
CLKBUF_X2 inst_11216 ( .A(net_11134), .Z(net_11135) );
DFF_X1 inst_8569 ( .Q(net_9874), .D(net_7290), .CK(net_14847) );
NOR2_X4 inst_2476 ( .A2(net_8930), .ZN(net_8379), .A1(net_8235) );
CLKBUF_X2 inst_11685 ( .A(net_11603), .Z(net_11604) );
CLKBUF_X2 inst_12078 ( .A(net_11996), .Z(net_11997) );
OAI21_X2 inst_1823 ( .B1(net_7157), .ZN(net_6570), .A(net_5926), .B2(net_5899) );
INV_X4 inst_5084 ( .A(net_5265), .ZN(net_1795) );
XNOR2_X2 inst_202 ( .ZN(net_4956), .A(net_4402), .B(net_3955) );
DFF_X2 inst_8116 ( .Q(net_10036), .D(net_5157), .CK(net_14300) );
HA_X1 inst_7359 ( .CO(net_5378), .A(net_5261), .S(net_1731), .B(net_636) );
AOI22_X2 inst_9154 ( .A1(net_9753), .A2(net_6404), .ZN(net_6328), .B2(net_5263), .B1(net_3529) );
OAI211_X2 inst_2212 ( .C1(net_7221), .C2(net_6501), .ZN(net_6493), .B(net_5564), .A(net_3679) );
CLKBUF_X2 inst_13786 ( .A(net_13704), .Z(net_13705) );
OAI222_X2 inst_1401 ( .B2(net_7728), .A2(net_7727), .C2(net_7726), .ZN(net_5330), .B1(net_3217), .A1(net_2771), .C1(net_1274) );
INV_X8 inst_4502 ( .ZN(net_6141), .A(net_5296) );
INV_X4 inst_4830 ( .A(net_10280), .ZN(net_5344) );
CLKBUF_X2 inst_14258 ( .A(net_13771), .Z(net_14177) );
CLKBUF_X2 inst_13444 ( .A(net_13362), .Z(net_13363) );
OAI211_X2 inst_2030 ( .C1(net_10054), .ZN(net_8125), .B(net_8043), .A(net_7935), .C2(net_6778) );
DFF_X2 inst_8254 ( .Q(net_10184), .D(net_4833), .CK(net_12856) );
INV_X4 inst_5624 ( .A(net_1342), .ZN(net_1148) );
DFF_X2 inst_7451 ( .QN(net_8834), .D(net_8162), .CK(net_14769) );
CLKBUF_X2 inst_11172 ( .A(net_10865), .Z(net_11091) );
DFF_X2 inst_7458 ( .QN(net_9290), .D(net_8163), .CK(net_14985) );
CLKBUF_X2 inst_14072 ( .A(net_13990), .Z(net_13991) );
XOR2_X2 inst_30 ( .Z(net_2124), .A(net_1741), .B(net_1206) );
SDFF_X2 inst_610 ( .QN(net_10236), .SI(net_10224), .SE(net_3667), .D(net_1321), .CK(net_10929) );
OAI22_X2 inst_1036 ( .A2(net_8921), .B1(net_8918), .ZN(net_7945), .A1(net_7846), .B2(net_1396) );
INV_X4 inst_6271 ( .A(net_10295), .ZN(net_445) );
XNOR2_X2 inst_233 ( .ZN(net_4313), .A(net_4165), .B(net_1832) );
AOI222_X1 inst_9704 ( .B1(net_9509), .A2(net_8295), .B2(net_8294), .C2(net_8293), .ZN(net_8274), .C1(net_8212), .A1(x2968) );
DFF_X1 inst_8639 ( .Q(net_9693), .D(net_7256), .CK(net_15557) );
AOI21_X2 inst_10094 ( .B2(net_10175), .A(net_6679), .ZN(net_5431), .B1(net_627) );
DFF_X1 inst_8595 ( .Q(net_9681), .D(net_7267), .CK(net_12011) );
AND4_X4 inst_10334 ( .ZN(net_2788), .A4(net_2108), .A1(net_1409), .A3(net_1296), .A2(net_1045) );
CLKBUF_X2 inst_12296 ( .A(net_12214), .Z(net_12215) );
AOI22_X2 inst_9527 ( .B1(net_9901), .A1(net_9671), .A2(net_5966), .B2(net_4969), .ZN(net_3794) );
AOI22_X2 inst_9127 ( .A1(net_9712), .A2(net_6382), .ZN(net_6361), .B2(net_5263), .B1(net_3894) );
DFF_X1 inst_8653 ( .Q(net_9763), .D(net_7193), .CK(net_15453) );
XNOR2_X2 inst_60 ( .B(net_9309), .A(net_9308), .ZN(net_8808) );
INV_X4 inst_5694 ( .A(net_3598), .ZN(net_1155) );
INV_X2 inst_6651 ( .ZN(net_8772), .A(net_8764) );
CLKBUF_X2 inst_14700 ( .A(net_14403), .Z(net_14619) );
CLKBUF_X2 inst_13540 ( .A(net_13458), .Z(net_13459) );
CLKBUF_X2 inst_12141 ( .A(net_12059), .Z(net_12060) );
INV_X4 inst_4613 ( .ZN(net_7339), .A(net_7156) );
INV_X4 inst_5852 ( .A(net_2702), .ZN(net_646) );
DFF_X2 inst_7752 ( .Q(net_10504), .D(net_6217), .CK(net_12273) );
NOR3_X2 inst_2376 ( .A2(net_9274), .ZN(net_8035), .A3(net_8033), .A1(net_3984) );
CLKBUF_X2 inst_13285 ( .A(net_13203), .Z(net_13204) );
DFF_X2 inst_7496 ( .D(net_8019), .QN(net_198), .CK(net_15166) );
DFF_X2 inst_7925 ( .Q(net_9225), .D(net_5785), .CK(net_14168) );
CLKBUF_X2 inst_12862 ( .A(net_12780), .Z(net_12781) );
NAND2_X2 inst_4360 ( .ZN(net_2465), .A2(net_951), .A1(net_313) );
INV_X2 inst_7050 ( .A(net_1761), .ZN(net_1333) );
HA_X1 inst_7339 ( .S(net_6175), .CO(net_6174), .B(net_5238), .A(net_1541) );
CLKBUF_X2 inst_12189 ( .A(net_12107), .Z(net_12108) );
OR2_X2 inst_860 ( .A1(net_10503), .ZN(net_7870), .A2(net_7869) );
SDFF_X2 inst_563 ( .D(net_9130), .SE(net_933), .CK(net_10935), .SI(x2589), .Q(x1262) );
CLKBUF_X2 inst_14074 ( .A(net_13992), .Z(net_13993) );
NAND2_X2 inst_3962 ( .ZN(net_3606), .A1(net_3456), .A2(net_3453) );
AND2_X4 inst_10392 ( .ZN(net_8001), .A1(net_7095), .A2(net_7094) );
DFF_X2 inst_8389 ( .Q(net_10198), .D(net_847), .CK(net_13532) );
OR2_X2 inst_943 ( .A2(net_10325), .A1(net_10324), .ZN(net_1864) );
CLKBUF_X2 inst_14397 ( .A(net_14315), .Z(net_14316) );
NAND2_X2 inst_3478 ( .A1(net_9457), .A2(net_8951), .ZN(net_8434) );
CLKBUF_X2 inst_11252 ( .A(net_11170), .Z(net_11171) );
AOI21_X2 inst_10181 ( .B1(net_7620), .A(net_4294), .ZN(net_3520), .B2(net_3058) );
INV_X4 inst_5314 ( .ZN(net_1563), .A(net_1283) );
CLKBUF_X2 inst_15714 ( .A(net_15632), .Z(net_15633) );
INV_X2 inst_7147 ( .A(net_1071), .ZN(net_788) );
CLKBUF_X2 inst_15505 ( .A(net_15423), .Z(net_15424) );
NOR2_X2 inst_2782 ( .ZN(net_3703), .A1(net_3145), .A2(net_2999) );
INV_X4 inst_4711 ( .A(net_5178), .ZN(net_4998) );
INV_X2 inst_7248 ( .A(net_9554), .ZN(net_362) );
CLKBUF_X2 inst_12151 ( .A(net_12069), .Z(net_12070) );
OAI21_X2 inst_1964 ( .ZN(net_3366), .A(net_3365), .B1(net_3364), .B2(net_3139) );
OAI21_X2 inst_1765 ( .B1(net_9057), .ZN(net_8970), .B2(net_8927), .A(net_8153) );
DFF_X2 inst_7464 ( .QN(net_9516), .D(net_8105), .CK(net_14981) );
INV_X4 inst_5475 ( .ZN(net_1193), .A(net_1006) );
CLKBUF_X2 inst_13887 ( .A(net_13605), .Z(net_13806) );
CLKBUF_X2 inst_11191 ( .A(net_11109), .Z(net_11110) );
NAND2_X2 inst_3720 ( .A2(net_10484), .ZN(net_7072), .A1(net_2205) );
CLKBUF_X2 inst_14672 ( .A(net_14590), .Z(net_14591) );
CLKBUF_X2 inst_11964 ( .A(net_10892), .Z(net_11883) );
CLKBUF_X2 inst_12444 ( .A(net_11967), .Z(net_12363) );
OAI21_X2 inst_2005 ( .ZN(net_2807), .A(net_2143), .B1(net_2142), .B2(net_1649) );
CLKBUF_X2 inst_11988 ( .A(net_10936), .Z(net_11907) );
CLKBUF_X2 inst_13377 ( .A(net_13295), .Z(net_13296) );
OR2_X4 inst_736 ( .A2(net_7038), .ZN(net_6183), .A1(net_6182) );
SDFF_X2 inst_544 ( .Q(net_9307), .D(net_9307), .SI(net_9158), .SE(net_7553), .CK(net_14034) );
CLKBUF_X2 inst_13525 ( .A(net_13443), .Z(net_13444) );
INV_X4 inst_5865 ( .ZN(net_982), .A(net_639) );
DFF_X2 inst_8021 ( .QN(net_10437), .D(net_5479), .CK(net_13639) );
INV_X4 inst_5465 ( .A(net_10247), .ZN(net_1819) );
CLKBUF_X2 inst_11944 ( .A(net_11862), .Z(net_11863) );
INV_X4 inst_6357 ( .A(net_10478), .ZN(net_7021) );
DFF_X2 inst_8232 ( .Q(net_10492), .D(net_4891), .CK(net_12962) );
XNOR2_X2 inst_178 ( .B(net_5953), .ZN(net_5357), .A(net_5190) );
AOI22_X2 inst_9179 ( .A1(net_9878), .B1(net_9779), .A2(net_8042), .ZN(net_6137), .B2(net_6133) );
NAND2_X2 inst_4402 ( .A2(net_10300), .A1(net_10286), .ZN(net_650) );
OR2_X4 inst_734 ( .A1(net_9245), .A2(net_9170), .ZN(net_7167) );
HA_X1 inst_7352 ( .A(net_9181), .S(net_4293), .CO(net_4292), .B(net_4124) );
OAI22_X2 inst_1282 ( .ZN(net_4096), .A1(net_4095), .A2(net_4092), .B1(net_2595), .B2(net_2260) );
DFF_X1 inst_8528 ( .Q(net_9971), .D(net_7314), .CK(net_12609) );
DFF_X2 inst_8257 ( .Q(net_10282), .D(net_4824), .CK(net_12942) );
CLKBUF_X2 inst_14818 ( .A(net_14736), .Z(net_14737) );
INV_X4 inst_5941 ( .A(net_6958), .ZN(net_569) );
CLKBUF_X2 inst_15673 ( .A(net_15591), .Z(net_15592) );
CLKBUF_X2 inst_13562 ( .A(net_13480), .Z(net_13481) );
NAND2_X2 inst_3919 ( .A2(net_9055), .ZN(net_7967), .A1(net_568) );
OAI22_X2 inst_1148 ( .A1(net_7203), .A2(net_5134), .B2(net_5133), .ZN(net_5125), .B1(net_689) );
DFF_X2 inst_7661 ( .D(net_6692), .QN(net_170), .CK(net_12817) );
AND2_X4 inst_10425 ( .ZN(net_3723), .A1(net_3722), .A2(net_3334) );
AOI211_X2 inst_10292 ( .ZN(net_4348), .C2(net_4328), .B(net_4013), .C1(net_1958), .A(net_1600) );
DFF_X2 inst_8270 ( .Q(net_10396), .D(net_4845), .CK(net_12932) );
NAND2_X2 inst_4350 ( .A2(net_10121), .ZN(net_1855), .A1(net_973) );
INV_X4 inst_5634 ( .ZN(net_1098), .A(net_854) );
AOI22_X2 inst_9597 ( .B1(net_9959), .A2(net_4694), .ZN(net_3495), .B2(net_2541), .A1(net_224) );
NAND2_X2 inst_3587 ( .ZN(net_7391), .A2(net_7390), .A1(net_5908) );
DFF_X1 inst_8777 ( .QN(net_10168), .D(net_4685), .CK(net_12298) );
AOI21_X2 inst_10139 ( .ZN(net_4246), .A(net_3936), .B2(net_3458), .B1(net_1558) );
CLKBUF_X2 inst_13003 ( .A(net_12407), .Z(net_12922) );
AOI21_X2 inst_10147 ( .ZN(net_4201), .A(net_4200), .B1(net_3708), .B2(net_3707) );
AOI22_X2 inst_9659 ( .A2(net_10140), .ZN(net_3153), .B2(net_1071), .A1(net_749), .B1(net_696) );
INV_X4 inst_5543 ( .ZN(net_2554), .A(net_940) );
INV_X4 inst_6004 ( .ZN(net_3976), .A(net_268) );
INV_X4 inst_6392 ( .A(net_9321), .ZN(net_1993) );
OR2_X4 inst_842 ( .A2(net_10359), .A1(net_10358), .ZN(net_1433) );
INV_X4 inst_5588 ( .ZN(net_6628), .A(net_1093) );
CLKBUF_X2 inst_15465 ( .A(net_12372), .Z(net_15384) );
CLKBUF_X2 inst_11427 ( .A(net_11345), .Z(net_11346) );
OAI211_X2 inst_2068 ( .ZN(net_7436), .C1(net_7435), .C2(net_7434), .A(net_7143), .B(net_2990) );
AOI221_X2 inst_9897 ( .B1(net_9882), .B2(net_9101), .A(net_6945), .C2(net_6944), .ZN(net_6797), .C1(net_253) );
INV_X4 inst_6183 ( .A(net_9745), .ZN(net_709) );
AOI222_X1 inst_9697 ( .B1(net_9508), .A2(net_8286), .B2(net_8285), .C2(net_8284), .ZN(net_8281), .C1(net_8197), .A1(x1547) );
SDFF_X2 inst_551 ( .D(net_9153), .SE(net_7248), .SI(net_195), .Q(net_195), .CK(net_15266) );
OAI211_X2 inst_2101 ( .C2(net_6778), .ZN(net_6747), .A(net_6421), .B(net_6105), .C1(net_413) );
CLKBUF_X2 inst_11529 ( .A(net_11447), .Z(net_11448) );
DFF_X1 inst_8542 ( .Q(net_9976), .D(net_7349), .CK(net_15474) );
XNOR2_X2 inst_353 ( .ZN(net_2797), .B(net_2777), .A(net_1773) );
NAND2_X2 inst_3808 ( .A1(net_10077), .A2(net_4534), .ZN(net_4530) );
CLKBUF_X2 inst_15721 ( .A(net_14399), .Z(net_15640) );
OAI21_X2 inst_1940 ( .ZN(net_4286), .A(net_4119), .B2(net_3963), .B1(net_986) );
INV_X4 inst_6286 ( .A(net_10035), .ZN(net_5098) );
DFF_X1 inst_8492 ( .QN(net_9636), .D(net_7826), .CK(net_13796) );
INV_X4 inst_4632 ( .ZN(net_7304), .A(net_6329) );
AND2_X4 inst_10400 ( .A2(net_9100), .ZN(net_6939), .A1(net_4796) );
CLKBUF_X2 inst_15025 ( .A(net_14943), .Z(net_14944) );
CLKBUF_X2 inst_13456 ( .A(net_13374), .Z(net_13375) );
CLKBUF_X2 inst_13917 ( .A(net_13835), .Z(net_13836) );
INV_X4 inst_6212 ( .A(net_10505), .ZN(net_465) );
NAND2_X2 inst_4041 ( .ZN(net_4088), .A1(net_2854), .A2(net_2619) );
CLKBUF_X2 inst_13761 ( .A(net_11462), .Z(net_13680) );
NAND2_X2 inst_3701 ( .A2(net_9100), .A1(net_6165), .ZN(net_5935) );
NAND2_X4 inst_3357 ( .ZN(net_8416), .A2(net_8381), .A1(net_8380) );
AOI22_X2 inst_9559 ( .B1(net_9894), .A1(net_9763), .B2(net_4969), .ZN(net_3760), .A2(net_2462) );
CLKBUF_X2 inst_14184 ( .A(net_14102), .Z(net_14103) );
INV_X2 inst_7082 ( .ZN(net_1174), .A(net_1173) );
CLKBUF_X2 inst_11822 ( .A(net_11740), .Z(net_11741) );
XOR2_X2 inst_8 ( .Z(net_3949), .B(net_3231), .A(net_2879) );
CLKBUF_X2 inst_15559 ( .A(net_15477), .Z(net_15478) );
CLKBUF_X2 inst_15456 ( .A(net_15374), .Z(net_15375) );
CLKBUF_X2 inst_14588 ( .A(net_13631), .Z(net_14507) );
CLKBUF_X2 inst_13869 ( .A(net_13787), .Z(net_13788) );
CLKBUF_X2 inst_11321 ( .A(net_10848), .Z(net_11240) );
INV_X2 inst_6745 ( .ZN(net_6842), .A(net_6618) );
CLKBUF_X2 inst_14064 ( .A(net_13982), .Z(net_13983) );
INV_X2 inst_6984 ( .ZN(net_2371), .A(net_1669) );
OAI211_X2 inst_2090 ( .C2(net_6778), .ZN(net_6758), .A(net_6411), .B(net_6118), .C1(net_418) );
OAI33_X1 inst_965 ( .A1(net_7437), .ZN(net_3359), .A3(net_3075), .B1(net_2751), .B2(net_2613), .A2(net_2589), .B3(net_2279) );
CLKBUF_X2 inst_13980 ( .A(net_13526), .Z(net_13899) );
CLKBUF_X2 inst_12624 ( .A(net_11473), .Z(net_12543) );
DFF_X2 inst_8228 ( .D(net_4868), .Q(net_227), .CK(net_10824) );
NAND2_X4 inst_3370 ( .ZN(net_9082), .A1(net_4018), .A2(net_3886) );
INV_X2 inst_7134 ( .A(net_1385), .ZN(net_1316) );
AOI21_X2 inst_10168 ( .B2(net_10197), .ZN(net_8375), .A(net_4371), .B1(net_3683) );
CLKBUF_X2 inst_14583 ( .A(net_14466), .Z(net_14502) );
CLKBUF_X2 inst_15301 ( .A(net_11242), .Z(net_15220) );
CLKBUF_X2 inst_12267 ( .A(net_12185), .Z(net_12186) );
DFF_X1 inst_8677 ( .D(net_6743), .Q(net_134), .CK(net_12088) );
CLKBUF_X2 inst_11991 ( .A(net_11870), .Z(net_11910) );
AOI22_X2 inst_8993 ( .A2(net_8936), .ZN(net_8616), .A1(net_8614), .B2(net_7753), .B1(net_7656) );
CLKBUF_X2 inst_12284 ( .A(net_12202), .Z(net_12203) );
CLKBUF_X2 inst_11976 ( .A(net_11894), .Z(net_11895) );
INV_X4 inst_6579 ( .A(net_10397), .ZN(net_4101) );
INV_X4 inst_5392 ( .A(net_2216), .ZN(net_1573) );
INV_X2 inst_7210 ( .A(net_9407), .ZN(net_8226) );
OR2_X2 inst_901 ( .A1(net_10398), .ZN(net_5410), .A2(net_5409) );
INV_X4 inst_6179 ( .A(net_9363), .ZN(net_7856) );
CLKBUF_X2 inst_10992 ( .A(net_10685), .Z(net_10911) );
CLKBUF_X2 inst_15520 ( .A(net_15438), .Z(net_15439) );
INV_X4 inst_6094 ( .A(net_9521), .ZN(net_3565) );
INV_X2 inst_7261 ( .A(net_9167), .ZN(net_320) );
CLKBUF_X2 inst_13821 ( .A(net_13739), .Z(net_13740) );
DFF_X2 inst_7913 ( .Q(net_9219), .D(net_5928), .CK(net_13013) );
AOI221_X2 inst_9957 ( .C1(net_10498), .B1(net_10288), .C2(net_6415), .ZN(net_4775), .B2(net_4774), .A(net_4335) );
CLKBUF_X2 inst_13288 ( .A(net_13206), .Z(net_13207) );
CLKBUF_X2 inst_10863 ( .A(net_10781), .Z(net_10782) );
CLKBUF_X2 inst_14843 ( .A(net_14761), .Z(net_14762) );
CLKBUF_X2 inst_14013 ( .A(net_11084), .Z(net_13932) );
NOR3_X2 inst_2403 ( .ZN(net_7448), .A1(net_7148), .A3(net_5181), .A2(net_3697) );
INV_X4 inst_4948 ( .A(net_4041), .ZN(net_2769) );
AOI22_X2 inst_9104 ( .A1(net_9684), .A2(net_6420), .ZN(net_6388), .B2(net_5263), .B1(net_4019) );
CLKBUF_X2 inst_14545 ( .A(net_14097), .Z(net_14464) );
OAI21_X2 inst_1934 ( .A(net_4877), .ZN(net_4362), .B2(net_4361), .B1(net_3192) );
INV_X2 inst_6759 ( .A(net_6651), .ZN(net_6232) );
AOI22_X2 inst_9429 ( .ZN(net_4593), .A1(net_4421), .A2(net_4284), .B2(net_3734), .B1(net_3547) );
NAND4_X2 inst_3098 ( .ZN(net_4345), .A1(net_3781), .A3(net_3757), .A4(net_3567), .A2(net_3405) );
NAND2_X2 inst_3916 ( .A2(net_9053), .ZN(net_7971), .A1(net_637) );
INV_X4 inst_5739 ( .A(net_1029), .ZN(net_991) );
INV_X4 inst_5401 ( .A(net_4988), .ZN(net_1524) );
CLKBUF_X2 inst_13834 ( .A(net_13752), .Z(net_13753) );
CLKBUF_X2 inst_10679 ( .A(net_10577), .Z(net_10598) );
AOI221_X2 inst_9970 ( .C1(net_9961), .ZN(net_4696), .B2(net_4694), .A(net_4277), .C2(net_2541), .B1(net_226) );
DFF_X2 inst_8319 ( .Q(net_10188), .D(net_3930), .CK(net_12246) );
INV_X4 inst_6144 ( .A(net_10146), .ZN(net_973) );
DFF_X1 inst_8539 ( .Q(net_9961), .D(net_7370), .CK(net_14635) );
INV_X4 inst_5013 ( .ZN(net_2812), .A(net_2118) );
CLKBUF_X2 inst_13359 ( .A(net_11387), .Z(net_13278) );
CLKBUF_X2 inst_12034 ( .A(net_11952), .Z(net_11953) );
DFF_X1 inst_8464 ( .Q(net_9593), .D(net_7960), .CK(net_11530) );
CLKBUF_X2 inst_10968 ( .A(net_10886), .Z(net_10887) );
OAI211_X2 inst_2097 ( .C2(net_6774), .ZN(net_6751), .A(net_6424), .B(net_6112), .C1(net_375) );
CLKBUF_X2 inst_12943 ( .A(net_12861), .Z(net_12862) );
CLKBUF_X2 inst_15782 ( .A(net_15700), .Z(net_15701) );
OR2_X2 inst_928 ( .A1(net_2972), .A2(net_2955), .ZN(net_2954) );
INV_X8 inst_4484 ( .ZN(net_8475), .A(net_8384) );
INV_X4 inst_5910 ( .A(net_1843), .ZN(net_940) );
CLKBUF_X2 inst_10695 ( .A(net_10613), .Z(net_10614) );
CLKBUF_X2 inst_14948 ( .A(net_14866), .Z(net_14867) );
NOR2_X2 inst_2662 ( .ZN(net_5013), .A1(net_5012), .A2(net_4728) );
OAI221_X2 inst_1539 ( .B2(net_9047), .C2(net_7287), .ZN(net_7227), .C1(net_7226), .A(net_6794), .B1(net_5493) );
DFF_X2 inst_8053 ( .QN(net_9555), .D(net_9261), .CK(net_12616) );
INV_X4 inst_6215 ( .A(net_9207), .ZN(net_3967) );
OAI221_X2 inst_1718 ( .B2(net_3907), .ZN(net_3208), .B1(net_3207), .C1(net_3206), .A(net_2757), .C2(net_2439) );
CLKBUF_X2 inst_12225 ( .A(net_12143), .Z(net_12144) );
OAI22_X2 inst_1050 ( .ZN(net_7534), .A2(net_7391), .B2(net_7390), .A1(net_7157), .B1(net_445) );
INV_X4 inst_6476 ( .A(net_9382), .ZN(net_7336) );
AOI22_X2 inst_9424 ( .A1(net_10181), .A2(net_4656), .B2(net_4655), .ZN(net_4645), .B1(x4041) );
DFF_X1 inst_8549 ( .Q(net_9985), .D(net_7362), .CK(net_14777) );
CLKBUF_X2 inst_11126 ( .A(net_11044), .Z(net_11045) );
DFF_X2 inst_7654 ( .D(net_6704), .Q(net_186), .CK(net_12511) );
OAI22_X2 inst_1296 ( .B1(net_4749), .A2(net_4274), .B2(net_3588), .ZN(net_3569), .A1(net_479) );
INV_X4 inst_4661 ( .A(net_9269), .ZN(net_6581) );
CLKBUF_X2 inst_14443 ( .A(net_13490), .Z(net_14362) );
OAI21_X2 inst_1852 ( .ZN(net_5878), .B2(net_5877), .A(net_5293), .B1(net_4659) );
INV_X2 inst_6809 ( .ZN(net_8995), .A(net_4990) );
INV_X4 inst_6273 ( .A(net_9568), .ZN(net_2849) );
NAND2_X2 inst_3671 ( .A1(net_8057), .ZN(net_7281), .A2(net_6241) );
DFF_X2 inst_7978 ( .QN(net_10314), .D(net_5569), .CK(net_15581) );
NAND3_X2 inst_3282 ( .ZN(net_3632), .A1(net_3631), .A2(net_3630), .A3(net_3452) );
CLKBUF_X2 inst_12667 ( .A(net_12585), .Z(net_12586) );
CLKBUF_X2 inst_13121 ( .A(net_12832), .Z(net_13040) );
NAND2_X2 inst_4074 ( .A2(net_2963), .ZN(net_2891), .A1(net_2610) );
NAND2_X2 inst_3783 ( .A2(net_8986), .A1(net_7277), .ZN(net_4990) );
INV_X8 inst_4513 ( .ZN(net_1502), .A(net_771) );
CLKBUF_X2 inst_13613 ( .A(net_12877), .Z(net_13532) );
OAI221_X2 inst_1557 ( .C2(net_7295), .B2(net_7293), .ZN(net_7199), .B1(net_7198), .A(net_6818), .C1(net_5475) );
NOR3_X2 inst_2399 ( .ZN(net_7568), .A3(net_7455), .A1(net_4379), .A2(net_4317) );
CLKBUF_X2 inst_15078 ( .A(net_14996), .Z(net_14997) );
CLKBUF_X2 inst_12207 ( .A(net_10642), .Z(net_12126) );
NAND2_X2 inst_3412 ( .ZN(net_8524), .A2(net_8486), .A1(net_8485) );
INV_X4 inst_4698 ( .ZN(net_4829), .A(net_4645) );
CLKBUF_X2 inst_10855 ( .A(net_10689), .Z(net_10774) );
AOI22_X2 inst_9620 ( .A1(net_9852), .B1(net_9789), .A2(net_6413), .ZN(net_3432), .B2(net_2462) );
DFF_X1 inst_8485 ( .Q(net_9632), .D(net_7893), .CK(net_11516) );
INV_X4 inst_6290 ( .ZN(net_435), .A(net_222) );
MUX2_X1 inst_4452 ( .S(net_6041), .A(net_294), .B(x5289), .Z(x157) );
CLKBUF_X2 inst_11326 ( .A(net_11244), .Z(net_11245) );
CLKBUF_X2 inst_10633 ( .A(net_10545), .Z(net_10552) );
OAI221_X2 inst_1616 ( .C1(net_10411), .B1(net_7243), .ZN(net_5595), .C2(net_4477), .B2(net_4455), .A(net_3527) );
CLKBUF_X2 inst_14090 ( .A(net_13064), .Z(net_14009) );
DFF_X1 inst_8813 ( .QN(net_10445), .D(net_3499), .CK(net_11135) );
INV_X4 inst_5646 ( .ZN(net_1126), .A(net_841) );
CLKBUF_X2 inst_13167 ( .A(net_12310), .Z(net_13086) );
CLKBUF_X2 inst_11295 ( .A(net_11213), .Z(net_11214) );
CLKBUF_X2 inst_11403 ( .A(net_11321), .Z(net_11322) );
AOI221_X2 inst_9954 ( .C1(net_9971), .B1(net_9674), .B2(net_5966), .ZN(net_4778), .A(net_4336), .C2(net_2541) );
OAI21_X2 inst_1825 ( .B1(net_7785), .ZN(net_6568), .A(net_5924), .B2(net_5895) );
NAND2_X2 inst_4151 ( .ZN(net_2050), .A2(net_2049), .A1(net_805) );
NOR2_X2 inst_2851 ( .A2(net_6044), .ZN(net_3534), .A1(net_2249) );
OAI221_X2 inst_1606 ( .C1(net_10231), .B1(net_7237), .C2(net_5642), .ZN(net_5630), .B2(net_4905), .A(net_3527) );
INV_X4 inst_5356 ( .A(net_5405), .ZN(net_1229) );
CLKBUF_X2 inst_13110 ( .A(net_13028), .Z(net_13029) );
INV_X4 inst_5619 ( .ZN(net_5164), .A(net_865) );
INV_X4 inst_5126 ( .ZN(net_2247), .A(net_1971) );
XNOR2_X2 inst_410 ( .ZN(net_1536), .A(net_1535), .B(net_1534) );
XNOR2_X2 inst_316 ( .ZN(net_3219), .B(net_3002), .A(net_2033) );
DFF_X1 inst_8690 ( .D(net_6711), .Q(net_143), .CK(net_15098) );
CLKBUF_X2 inst_12860 ( .A(net_12778), .Z(net_12779) );
CLKBUF_X2 inst_11786 ( .A(net_11704), .Z(net_11705) );
CLKBUF_X2 inst_11621 ( .A(net_11533), .Z(net_11540) );
OAI22_X2 inst_1174 ( .A1(net_7203), .A2(net_5107), .B2(net_5105), .ZN(net_5087), .B1(net_721) );
OAI22_X2 inst_1023 ( .A2(net_8036), .B2(net_8018), .ZN(net_8015), .A1(net_3033), .B1(net_675) );
CLKBUF_X2 inst_15303 ( .A(net_15221), .Z(net_15222) );
NAND3_X2 inst_3186 ( .ZN(net_7818), .A1(net_7769), .A3(net_1046), .A2(net_1044) );
CLKBUF_X2 inst_15266 ( .A(net_15184), .Z(net_15185) );
DFF_X1 inst_8515 ( .QN(net_8821), .D(net_7485), .CK(net_11484) );
SDFF_X2 inst_678 ( .SI(net_9501), .Q(net_9501), .SE(net_3073), .CK(net_11358), .D(x1418) );
NAND2_X2 inst_3762 ( .ZN(net_5260), .A2(net_4985), .A1(net_1350) );
INV_X4 inst_5653 ( .A(net_10224), .ZN(net_1321) );
CLKBUF_X2 inst_10925 ( .A(net_10843), .Z(net_10844) );
NAND3_X2 inst_3259 ( .ZN(net_4450), .A3(net_4319), .A1(net_4186), .A2(net_3591) );
OR2_X2 inst_854 ( .A1(net_9272), .A2(net_9271), .ZN(net_8124) );
CLKBUF_X2 inst_12464 ( .A(net_11640), .Z(net_12383) );
CLKBUF_X2 inst_13293 ( .A(net_12303), .Z(net_13212) );
CLKBUF_X2 inst_13796 ( .A(net_13714), .Z(net_13715) );
CLKBUF_X2 inst_15369 ( .A(net_15287), .Z(net_15288) );
NAND2_X2 inst_4359 ( .A2(net_10160), .ZN(net_2655), .A1(net_614) );
INV_X2 inst_7310 ( .A(net_9088), .ZN(net_9087) );
CLKBUF_X2 inst_13177 ( .A(net_11368), .Z(net_13096) );
CLKBUF_X2 inst_15765 ( .A(net_15683), .Z(net_15684) );
NAND2_X2 inst_3678 ( .A1(net_9080), .A2(net_7043), .ZN(net_6225) );
NAND2_X2 inst_3979 ( .ZN(net_3262), .A2(net_3261), .A1(net_2887) );
INV_X4 inst_6297 ( .A(net_9651), .ZN(net_433) );
DFF_X2 inst_8033 ( .Q(net_9231), .D(net_5446), .CK(net_13568) );
CLKBUF_X2 inst_12191 ( .A(net_11867), .Z(net_12110) );
CLKBUF_X2 inst_15578 ( .A(net_13061), .Z(net_15497) );
OAI21_X2 inst_1946 ( .B2(net_4332), .ZN(net_4205), .B1(net_4204), .A(net_4175) );
DFF_X2 inst_7865 ( .QN(net_9378), .D(net_7505), .CK(net_13021) );
AND2_X2 inst_10478 ( .A2(net_9582), .ZN(net_8743), .A1(net_3121) );
AND2_X4 inst_10472 ( .A2(net_10363), .A1(net_10362), .ZN(net_2012) );
CLKBUF_X2 inst_12006 ( .A(net_11924), .Z(net_11925) );
DFF_X1 inst_8686 ( .D(net_6716), .Q(net_138), .CK(net_15730) );
AOI22_X2 inst_9226 ( .A1(net_9920), .B1(net_9821), .A2(net_6141), .B2(net_6129), .ZN(net_6085) );
INV_X4 inst_5322 ( .ZN(net_1562), .A(net_1272) );
DFF_X2 inst_8008 ( .QN(net_10228), .D(net_5499), .CK(net_11741) );
CLKBUF_X2 inst_13401 ( .A(net_13319), .Z(net_13320) );
AOI221_X2 inst_9786 ( .B1(net_9966), .A(net_7090), .B2(net_7089), .C1(net_7088), .ZN(net_7081), .C2(net_238) );
AOI22_X2 inst_9073 ( .B1(net_9692), .A1(net_6811), .A2(net_6684), .B2(net_6683), .ZN(net_6593) );
CLKBUF_X2 inst_10861 ( .A(net_10779), .Z(net_10780) );
NAND2_X2 inst_3457 ( .A2(net_9489), .A1(net_8476), .ZN(net_8467) );
CLKBUF_X2 inst_12996 ( .A(net_12914), .Z(net_12915) );
AOI22_X2 inst_9464 ( .B1(net_9708), .A1(net_9676), .A2(net_5966), .ZN(net_3863), .B2(net_3039) );
OR4_X2 inst_688 ( .A4(net_4914), .ZN(net_4911), .A3(net_3045), .A2(net_1263), .A1(net_1260) );
NOR2_X2 inst_2549 ( .ZN(net_8284), .A1(net_8082), .A2(net_7990) );
OAI21_X2 inst_1749 ( .ZN(net_8668), .A(net_8632), .B2(net_8589), .B1(net_8116) );
AOI222_X1 inst_9717 ( .A1(net_9070), .ZN(net_6320), .C2(net_6319), .A2(net_5994), .C1(net_5993), .B2(net_5973), .B1(net_4997) );
NAND2_X2 inst_3641 ( .ZN(net_7253), .A1(net_6903), .A2(net_6902) );
INV_X4 inst_6519 ( .A(net_10098), .ZN(net_5837) );
CLKBUF_X2 inst_14105 ( .A(net_11673), .Z(net_14024) );
INV_X4 inst_4894 ( .ZN(net_2897), .A(net_2896) );
INV_X4 inst_5514 ( .A(net_10354), .ZN(net_3668) );
CLKBUF_X2 inst_15372 ( .A(net_13300), .Z(net_15291) );
CLKBUF_X2 inst_12518 ( .A(net_12436), .Z(net_12437) );
AOI22_X2 inst_9071 ( .B1(net_9691), .A2(net_6684), .B2(net_6683), .ZN(net_6595), .A1(net_260) );
NOR3_X2 inst_2387 ( .A1(net_7884), .A3(net_7805), .ZN(net_7803), .A2(net_2607) );
CLKBUF_X2 inst_14416 ( .A(net_12124), .Z(net_14335) );
CLKBUF_X2 inst_13351 ( .A(net_11886), .Z(net_13270) );
CLKBUF_X2 inst_12980 ( .A(net_10925), .Z(net_12899) );
CLKBUF_X2 inst_12474 ( .A(net_12392), .Z(net_12393) );
CLKBUF_X2 inst_11872 ( .A(net_11790), .Z(net_11791) );
AOI22_X2 inst_9017 ( .B1(net_9526), .ZN(net_8004), .A1(net_8002), .B2(net_8001), .A2(net_7945) );
NAND2_X2 inst_4391 ( .A1(net_10158), .A2(net_9734), .ZN(net_2767) );
AOI21_X2 inst_10137 ( .ZN(net_4895), .A(net_4249), .B2(net_3635), .B1(net_3069) );
AOI21_X2 inst_10017 ( .B2(net_8947), .ZN(net_8051), .B1(net_7993), .A(net_7571) );
AOI21_X2 inst_10163 ( .B2(net_10444), .ZN(net_4136), .A(net_1676), .B1(net_1273) );
NAND4_X2 inst_3156 ( .ZN(net_3131), .A3(net_2105), .A1(net_1855), .A4(net_1854), .A2(net_899) );
INV_X4 inst_6423 ( .A(net_10071), .ZN(net_383) );
NOR2_X2 inst_2747 ( .ZN(net_4005), .A1(net_3988), .A2(net_3677) );
CLKBUF_X2 inst_13744 ( .A(net_13662), .Z(net_13663) );
OR2_X4 inst_840 ( .A2(net_10149), .A1(net_10148), .ZN(net_1437) );
OAI22_X2 inst_1220 ( .A1(net_7129), .A2(net_5107), .B2(net_5105), .ZN(net_5028), .B1(net_5027) );
DFF_X1 inst_8554 ( .Q(net_9987), .D(net_7354), .CK(net_12170) );
OAI211_X2 inst_2181 ( .C1(net_7237), .C2(net_6548), .ZN(net_6528), .B(net_5655), .A(net_3679) );
OAI221_X2 inst_1456 ( .B2(net_7974), .C2(net_7973), .ZN(net_7972), .A(net_7971), .C1(net_7846), .B1(net_1893) );
CLKBUF_X2 inst_11900 ( .A(net_11818), .Z(net_11819) );
CLKBUF_X2 inst_13523 ( .A(net_12046), .Z(net_13442) );
CLKBUF_X2 inst_12498 ( .A(net_12208), .Z(net_12417) );
INV_X4 inst_6117 ( .ZN(net_6813), .A(net_233) );
CLKBUF_X2 inst_10736 ( .A(net_10654), .Z(net_10655) );
INV_X4 inst_5154 ( .ZN(net_7495), .A(net_2281) );
INV_X4 inst_5876 ( .A(net_915), .ZN(net_908) );
DFF_X2 inst_7497 ( .D(net_8017), .QN(net_199), .CK(net_15162) );
AND2_X2 inst_10593 ( .A2(net_4265), .ZN(net_2373), .A1(net_2189) );
NAND2_X2 inst_4195 ( .ZN(net_7584), .A1(net_1836), .A2(net_1714) );
NAND2_X2 inst_4294 ( .A1(net_3102), .ZN(net_2426), .A2(net_1249) );
DFF_X1 inst_8473 ( .QN(net_9429), .D(net_7891), .CK(net_12672) );
AOI22_X2 inst_9305 ( .B1(net_9711), .A2(net_5755), .B2(net_5754), .ZN(net_5673), .A1(net_248) );
CLKBUF_X2 inst_13605 ( .A(net_13523), .Z(net_13524) );
DFF_X2 inst_7589 ( .QN(net_9301), .D(net_7498), .CK(net_14105) );
MUX2_X1 inst_4440 ( .S(net_6041), .A(net_306), .B(x4359), .Z(x73) );
CLKBUF_X2 inst_14302 ( .A(net_14220), .Z(net_14221) );
CLKBUF_X2 inst_10799 ( .A(net_10673), .Z(net_10718) );
INV_X4 inst_5710 ( .ZN(net_1101), .A(net_809) );
CLKBUF_X2 inst_11607 ( .A(net_11525), .Z(net_11526) );
INV_X4 inst_5959 ( .A(net_10512), .ZN(net_551) );
INV_X2 inst_7072 ( .A(net_2850), .ZN(net_1231) );
AOI22_X2 inst_9536 ( .B1(net_9871), .A1(net_9836), .A2(net_6413), .ZN(net_3785), .B2(net_2973) );
INV_X4 inst_5939 ( .A(net_1847), .ZN(net_943) );
AOI22_X2 inst_9149 ( .A1(net_9727), .A2(net_6418), .ZN(net_6336), .B2(net_5263), .B1(net_5161) );
CLKBUF_X2 inst_11846 ( .A(net_11764), .Z(net_11765) );
NAND2_X2 inst_4199 ( .A1(net_2952), .ZN(net_1797), .A2(net_1796) );
CLKBUF_X2 inst_13588 ( .A(net_13506), .Z(net_13507) );
INV_X4 inst_5679 ( .ZN(net_3270), .A(net_2212) );
INV_X2 inst_7272 ( .A(net_8944), .ZN(net_8943) );
CLKBUF_X2 inst_14370 ( .A(net_14288), .Z(net_14289) );
CLKBUF_X2 inst_11141 ( .A(net_11059), .Z(net_11060) );
AOI22_X2 inst_9200 ( .A1(net_9862), .B1(net_9763), .A2(net_8042), .B2(net_6140), .ZN(net_6113) );
CLKBUF_X2 inst_12718 ( .A(net_12636), .Z(net_12637) );
SDFF_X2 inst_617 ( .Q(net_9450), .D(net_9450), .SE(net_3293), .CK(net_14164), .SI(x2531) );
CLKBUF_X2 inst_14897 ( .A(net_14815), .Z(net_14816) );
AOI22_X2 inst_9167 ( .A2(net_6418), .ZN(net_6304), .B2(net_5263), .B1(net_2587), .A1(net_2567) );
INV_X4 inst_5734 ( .ZN(net_935), .A(net_749) );
INV_X4 inst_5749 ( .A(net_2545), .ZN(net_966) );
INV_X4 inst_6225 ( .ZN(net_3899), .A(net_151) );
CLKBUF_X2 inst_12754 ( .A(net_10917), .Z(net_12673) );
CLKBUF_X2 inst_10823 ( .A(net_10741), .Z(net_10742) );
CLKBUF_X2 inst_14209 ( .A(net_14127), .Z(net_14128) );
NAND2_X1 inst_4420 ( .ZN(net_8737), .A2(net_8736), .A1(net_8596) );
CLKBUF_X2 inst_13795 ( .A(net_13713), .Z(net_13714) );
OAI22_X2 inst_1057 ( .B2(net_10450), .A1(net_10449), .ZN(net_7307), .A2(net_7306), .B1(net_909) );
DFF_X2 inst_8123 ( .QN(net_9746), .D(net_5142), .CK(net_12494) );
CLKBUF_X2 inst_14097 ( .A(net_14015), .Z(net_14016) );
INV_X4 inst_6614 ( .ZN(net_8931), .A(net_8930) );
CLKBUF_X2 inst_15225 ( .A(net_15143), .Z(net_15144) );
AND3_X4 inst_10359 ( .ZN(net_5743), .A2(net_4788), .A3(net_4628), .A1(net_4466) );
DFF_X1 inst_8843 ( .Q(net_9198), .D(net_2501), .CK(net_11289) );
CLKBUF_X2 inst_14565 ( .A(net_14483), .Z(net_14484) );
INV_X4 inst_5191 ( .ZN(net_3807), .A(net_1546) );
CLKBUF_X2 inst_15749 ( .A(net_15667), .Z(net_15668) );
INV_X4 inst_6029 ( .ZN(net_1970), .A(net_121) );
INV_X4 inst_5602 ( .A(net_1379), .ZN(net_1281) );
CLKBUF_X2 inst_10743 ( .A(net_10661), .Z(net_10662) );
CLKBUF_X2 inst_11956 ( .A(net_11554), .Z(net_11875) );
AND2_X2 inst_10610 ( .A1(net_3897), .ZN(net_2671), .A2(net_1977) );
OR2_X4 inst_748 ( .ZN(net_5298), .A2(net_5178), .A1(net_4480) );
DFF_X1 inst_8609 ( .Q(net_9861), .D(net_7239), .CK(net_15469) );
NOR2_X2 inst_2839 ( .ZN(net_2341), .A2(net_2340), .A1(net_1607) );
INV_X2 inst_6730 ( .ZN(net_7569), .A(net_7532) );
CLKBUF_X2 inst_11373 ( .A(net_11291), .Z(net_11292) );
AOI22_X2 inst_9266 ( .ZN(net_6648), .A2(net_5228), .B1(net_3855), .B2(net_2897), .A1(net_2684) );
INV_X4 inst_4582 ( .ZN(net_8068), .A(net_8026) );
INV_X4 inst_5482 ( .ZN(net_2984), .A(net_187) );
INV_X2 inst_7159 ( .A(net_3104), .ZN(net_654) );
INV_X2 inst_6739 ( .ZN(net_7319), .A(net_7318) );
CLKBUF_X2 inst_15700 ( .A(net_15618), .Z(net_15619) );
INV_X8 inst_4526 ( .ZN(net_8975), .A(net_3370) );
INV_X4 inst_5532 ( .ZN(net_1665), .A(net_948) );
CLKBUF_X2 inst_14487 ( .A(net_12409), .Z(net_14406) );
CLKBUF_X2 inst_11070 ( .A(net_10988), .Z(net_10989) );
AOI221_X2 inst_9818 ( .B1(net_9767), .B2(net_9097), .ZN(net_6941), .A(net_6940), .C1(net_6939), .C2(net_237) );
DFF_X1 inst_8798 ( .QN(net_10272), .D(net_4116), .CK(net_14489) );
CLKBUF_X2 inst_15064 ( .A(net_14982), .Z(net_14983) );
NOR2_X2 inst_2909 ( .A1(net_10162), .ZN(net_3202), .A2(net_1543) );
OAI21_X2 inst_1986 ( .ZN(net_2793), .A(net_2792), .B1(net_2739), .B2(net_2102) );
INV_X4 inst_4587 ( .ZN(net_8063), .A(net_8021) );
OAI21_X2 inst_1949 ( .ZN(net_3980), .A(net_3666), .B2(net_3488), .B1(net_917) );
CLKBUF_X2 inst_12636 ( .A(net_12554), .Z(net_12555) );
INV_X4 inst_5726 ( .ZN(net_858), .A(net_757) );
INV_X4 inst_6170 ( .A(net_10395), .ZN(net_475) );
CLKBUF_X2 inst_12163 ( .A(net_10946), .Z(net_12082) );
CLKBUF_X2 inst_10644 ( .A(net_10553), .Z(net_10563) );
NAND4_X2 inst_3135 ( .ZN(net_2914), .A4(net_2913), .A3(net_2905), .A2(net_2904), .A1(net_1663) );
INV_X4 inst_5867 ( .A(net_2495), .ZN(net_1698) );
DFF_X2 inst_8243 ( .Q(net_10076), .D(net_4859), .CK(net_10680) );
OR3_X4 inst_701 ( .ZN(net_7664), .A3(net_4169), .A2(net_4160), .A1(net_1495) );
NOR2_X2 inst_2911 ( .A2(net_2824), .ZN(net_1499), .A1(net_1498) );
CLKBUF_X2 inst_13770 ( .A(net_13688), .Z(net_13689) );
NOR3_X2 inst_2380 ( .ZN(net_7897), .A3(net_7771), .A1(net_3984), .A2(x3390) );
CLKBUF_X2 inst_12337 ( .A(net_12255), .Z(net_12256) );
DFF_X2 inst_7583 ( .Q(net_10400), .D(net_7537), .CK(net_15151) );
INV_X4 inst_5261 ( .A(net_5166), .ZN(net_3142) );
DFF_X2 inst_7739 ( .Q(net_10071), .D(net_6199), .CK(net_11180) );
OAI21_X2 inst_1859 ( .B2(net_10238), .ZN(net_5784), .A(net_2103), .B1(net_1563) );
DFF_X2 inst_7734 ( .Q(net_9997), .D(net_6215), .CK(net_11978) );
DFF_X2 inst_8238 ( .Q(net_10500), .D(net_4881), .CK(net_15211) );
INV_X2 inst_6933 ( .A(net_3175), .ZN(net_1931) );
CLKBUF_X2 inst_15818 ( .A(net_15736), .Z(net_15737) );
NOR2_X2 inst_2815 ( .ZN(net_2618), .A2(net_2617), .A1(net_1940) );
OAI22_X2 inst_1007 ( .ZN(net_8589), .A1(net_8315), .B2(net_8314), .A2(net_8146), .B1(net_8104) );
CLKBUF_X2 inst_11011 ( .A(net_10630), .Z(net_10930) );
DFF_X2 inst_8267 ( .Q(net_10391), .D(net_4808), .CK(net_15206) );
INV_X4 inst_5754 ( .ZN(net_848), .A(net_734) );
CLKBUF_X2 inst_11674 ( .A(net_11592), .Z(net_11593) );
DFF_X1 inst_8426 ( .Q(net_9586), .D(net_8730), .CK(net_13817) );
NAND2_X2 inst_4208 ( .A2(net_2827), .A1(net_2204), .ZN(net_1764) );
NAND2_X2 inst_3605 ( .ZN(net_7261), .A2(net_6863), .A1(net_6601) );
CLKBUF_X2 inst_11932 ( .A(net_11850), .Z(net_11851) );
AOI22_X2 inst_9617 ( .B1(net_10281), .A1(net_9848), .A2(net_6413), .B2(net_4774), .ZN(net_3436) );
SDFF_X2 inst_651 ( .SI(net_9494), .Q(net_9494), .SE(net_3073), .CK(net_12428), .D(x1792) );
INV_X4 inst_5066 ( .A(net_4037), .ZN(net_1860) );
CLKBUF_X2 inst_11998 ( .A(net_10931), .Z(net_11917) );
CLKBUF_X2 inst_11392 ( .A(net_11112), .Z(net_11311) );
NOR2_X2 inst_2883 ( .A2(net_10351), .A1(net_10350), .ZN(net_2563) );
CLKBUF_X2 inst_11560 ( .A(net_11124), .Z(net_11479) );
CLKBUF_X2 inst_11313 ( .A(net_11191), .Z(net_11232) );
OAI22_X2 inst_1157 ( .A1(net_7184), .A2(net_5139), .B2(net_5138), .ZN(net_5116), .B1(net_3644) );
DFF_X2 inst_8065 ( .QN(net_10459), .D(net_5327), .CK(net_11381) );
AOI221_X2 inst_9993 ( .B2(net_10075), .C2(net_10074), .B1(net_10066), .C1(net_10065), .ZN(net_2114), .A(net_1253) );
CLKBUF_X2 inst_11108 ( .A(net_11026), .Z(net_11027) );
CLKBUF_X2 inst_13395 ( .A(net_13313), .Z(net_13314) );
DFF_X1 inst_8408 ( .D(net_8807), .CK(net_11934), .Q(x769) );
NAND2_X2 inst_3528 ( .ZN(net_9015), .A2(net_8087), .A1(net_8086) );
AOI21_X2 inst_10083 ( .B2(net_10448), .A(net_10447), .ZN(net_5396), .B1(net_1468) );
OAI211_X2 inst_2061 ( .B(net_7783), .C2(net_7782), .ZN(net_7742), .A(net_7686), .C1(net_2480) );
NAND2_X2 inst_3685 ( .ZN(net_6663), .A2(net_5991), .A1(net_2654) );
AND2_X2 inst_10527 ( .ZN(net_3968), .A1(net_3967), .A2(net_3966) );
CLKBUF_X2 inst_13486 ( .A(net_11870), .Z(net_13405) );
NAND2_X2 inst_4255 ( .ZN(net_2062), .A1(net_1387), .A2(net_1371) );
INV_X2 inst_6891 ( .A(net_3722), .ZN(net_2689) );
CLKBUF_X2 inst_11301 ( .A(net_11219), .Z(net_11220) );
OAI221_X2 inst_1472 ( .ZN(net_7799), .A(net_7795), .C2(net_6842), .B2(net_6617), .B1(net_5752), .C1(net_5274) );
NAND2_X2 inst_4261 ( .A1(net_10473), .ZN(net_2766), .A2(net_1961) );
DFF_X2 inst_7616 ( .QN(net_9214), .D(net_6962), .CK(net_11835) );
CLKBUF_X2 inst_12511 ( .A(net_12429), .Z(net_12430) );
INV_X4 inst_6138 ( .A(net_10122), .ZN(net_614) );
CLKBUF_X2 inst_14981 ( .A(net_14899), .Z(net_14900) );
CLKBUF_X2 inst_14784 ( .A(net_14702), .Z(net_14703) );
NAND2_X2 inst_3784 ( .A2(net_9590), .ZN(net_5388), .A1(net_4687) );
OAI22_X2 inst_1183 ( .A1(net_7224), .A2(net_5107), .B2(net_5105), .ZN(net_5076), .B1(net_5075) );
AOI22_X2 inst_9577 ( .B1(net_9976), .A2(net_5173), .ZN(net_3676), .B2(net_2541), .A1(net_210) );
OAI221_X2 inst_1489 ( .B1(net_10425), .C2(net_9063), .B2(net_9056), .ZN(net_7381), .C1(net_7294), .A(net_7091) );
NOR3_X2 inst_2415 ( .A3(net_9162), .ZN(net_5939), .A1(net_5370), .A2(x3683) );
INV_X4 inst_5272 ( .A(net_3529), .ZN(net_1356) );
CLKBUF_X2 inst_15242 ( .A(net_15160), .Z(net_15161) );
CLKBUF_X2 inst_12353 ( .A(net_10868), .Z(net_12272) );
NAND3_X2 inst_3288 ( .A1(net_5268), .A2(net_4717), .ZN(net_3087), .A3(net_2244) );
OAI211_X2 inst_2262 ( .C1(net_7139), .C2(net_6548), .ZN(net_6286), .B(net_5712), .A(net_3527) );
CLKBUF_X2 inst_14498 ( .A(net_14416), .Z(net_14417) );
INV_X4 inst_4981 ( .ZN(net_2582), .A(net_2243) );
DFF_X2 inst_8352 ( .Q(net_10280), .D(net_3191), .CK(net_12469) );
INV_X4 inst_5506 ( .ZN(net_7420), .A(net_980) );
AOI22_X2 inst_9131 ( .A1(net_9715), .A2(net_6404), .ZN(net_6357), .B2(net_5263), .B1(net_944) );
OAI222_X2 inst_1394 ( .A2(net_7728), .C2(net_7727), .B2(net_7726), .ZN(net_5704), .A1(net_2863), .C1(net_2016), .B1(net_1131) );
OAI22_X2 inst_1160 ( .A1(net_7201), .A2(net_5139), .B2(net_5138), .ZN(net_5113), .B1(net_744) );
CLKBUF_X2 inst_13724 ( .A(net_13642), .Z(net_13643) );
INV_X2 inst_7102 ( .ZN(net_1056), .A(net_1055) );
CLKBUF_X2 inst_10767 ( .A(net_10685), .Z(net_10686) );
OAI21_X2 inst_1808 ( .ZN(net_7396), .B2(net_7060), .A(net_5348), .B1(net_5347) );
DFF_X1 inst_8440 ( .D(net_8452), .CK(net_10846), .Q(x1029) );
OAI21_X2 inst_1876 ( .B2(net_9068), .A(net_8926), .ZN(net_5264), .B1(net_545) );
OAI22_X2 inst_988 ( .A2(net_8962), .B2(net_8659), .ZN(net_8652), .B1(net_6241), .A1(net_6209) );
AOI211_X2 inst_10288 ( .C1(net_10175), .C2(net_8832), .ZN(net_4979), .B(net_4667), .A(net_4222) );
CLKBUF_X2 inst_15668 ( .A(net_11208), .Z(net_15587) );
CLKBUF_X2 inst_14941 ( .A(net_14859), .Z(net_14860) );
AOI22_X2 inst_9333 ( .B1(net_9809), .A2(net_5766), .B2(net_5765), .ZN(net_5619), .A1(net_247) );
CLKBUF_X2 inst_12869 ( .A(net_11407), .Z(net_12788) );
OAI22_X2 inst_1315 ( .A2(net_2880), .B2(net_2646), .ZN(net_2152), .A1(net_2131), .B1(net_1061) );
INV_X4 inst_4954 ( .A(net_2854), .ZN(net_2553) );
INV_X4 inst_5035 ( .A(net_5930), .ZN(net_1934) );
NOR3_X2 inst_2392 ( .A3(net_9000), .ZN(net_7816), .A1(net_7715), .A2(net_7461) );
INV_X4 inst_4759 ( .ZN(net_4545), .A(net_4113) );
NAND2_X2 inst_4308 ( .A2(net_10352), .ZN(net_2031), .A1(net_902) );
INV_X4 inst_4678 ( .ZN(net_5694), .A(net_5361) );
CLKBUF_X2 inst_11026 ( .A(net_10579), .Z(net_10945) );
AOI22_X2 inst_9531 ( .B1(net_10022), .A1(net_9954), .A2(net_6443), .ZN(net_3790), .B2(net_2468) );
CLKBUF_X2 inst_13513 ( .A(net_11380), .Z(net_13432) );
NAND2_X2 inst_3667 ( .A2(net_10485), .A1(net_10484), .ZN(net_7071) );
DFF_X2 inst_7569 ( .QN(net_10267), .D(net_7580), .CK(net_11684) );
DFF_X2 inst_7972 ( .QN(net_10306), .D(net_5580), .CK(net_13242) );
MUX2_X1 inst_4434 ( .S(net_6041), .A(net_312), .B(x3889), .Z(x27) );
CLKBUF_X2 inst_14775 ( .A(net_14693), .Z(net_14694) );
INV_X4 inst_6380 ( .A(net_9616), .ZN(net_397) );
AOI21_X2 inst_10049 ( .ZN(net_7312), .B2(net_7291), .A(net_3562), .B1(net_3397) );
INV_X4 inst_4967 ( .ZN(net_2484), .A(net_2152) );
CLKBUF_X2 inst_15249 ( .A(net_15167), .Z(net_15168) );
CLKBUF_X2 inst_14953 ( .A(net_12937), .Z(net_14872) );
INV_X2 inst_7217 ( .A(net_9930), .ZN(net_441) );
AOI221_X2 inst_9808 ( .B1(net_9987), .A(net_7090), .B2(net_7089), .C2(net_7088), .ZN(net_6994), .C1(net_6816) );
INV_X2 inst_6785 ( .A(net_9261), .ZN(net_6238) );
CLKBUF_X2 inst_10792 ( .A(net_10710), .Z(net_10711) );
INV_X4 inst_5527 ( .A(net_10460), .ZN(net_4554) );
INV_X2 inst_7007 ( .A(net_2343), .ZN(net_1609) );
CLKBUF_X2 inst_13993 ( .A(net_13911), .Z(net_13912) );
CLKBUF_X2 inst_10866 ( .A(net_10784), .Z(net_10785) );
SDFF_X2 inst_656 ( .SI(net_9482), .Q(net_9482), .SE(net_3073), .CK(net_14138), .D(x2531) );
AOI222_X1 inst_9690 ( .B1(net_9510), .A2(net_8301), .B2(net_8300), .C2(net_8299), .ZN(net_8291), .C1(net_8223), .A1(x1911) );
INV_X2 inst_6718 ( .ZN(net_7938), .A(net_7912) );
INV_X2 inst_6900 ( .ZN(net_5963), .A(net_2408) );
CLKBUF_X2 inst_12562 ( .A(net_11145), .Z(net_12481) );
INV_X4 inst_5919 ( .ZN(net_1005), .A(net_586) );
XOR2_X2 inst_45 ( .A(net_7905), .B(net_7634), .Z(net_2446) );
CLKBUF_X2 inst_15351 ( .A(net_15269), .Z(net_15270) );
CLKBUF_X2 inst_13471 ( .A(net_12077), .Z(net_13390) );
AOI22_X2 inst_9551 ( .B1(net_9861), .A1(net_9695), .ZN(net_3769), .A2(net_3039), .B2(net_2973) );
CLKBUF_X2 inst_15125 ( .A(net_11990), .Z(net_15044) );
CLKBUF_X2 inst_12500 ( .A(net_12418), .Z(net_12419) );
NAND4_X2 inst_3093 ( .ZN(net_4377), .A4(net_3912), .A3(net_3808), .A1(net_3428), .A2(net_3427) );
SDFF_X2 inst_458 ( .SE(net_8747), .SI(net_8723), .Q(net_243), .D(net_112), .CK(net_12558) );
AOI221_X2 inst_9934 ( .B2(net_5867), .A(net_5862), .C2(net_5853), .ZN(net_5836), .C1(net_5835), .B1(x5850) );
OAI221_X2 inst_1562 ( .C1(net_10202), .C2(net_7295), .B2(net_7293), .ZN(net_7193), .B1(net_7192), .A(net_6814) );
NAND2_X2 inst_4148 ( .ZN(net_2073), .A1(net_2072), .A2(net_1369) );
CLKBUF_X2 inst_11814 ( .A(net_11732), .Z(net_11733) );
DFF_X1 inst_8644 ( .Q(net_9885), .D(net_7227), .CK(net_12154) );
INV_X4 inst_4618 ( .ZN(net_7553), .A(net_7016) );
INV_X4 inst_5539 ( .ZN(net_2257), .A(net_1366) );
INV_X2 inst_6827 ( .ZN(net_4137), .A(net_4136) );
OAI21_X2 inst_1922 ( .ZN(net_4551), .A(net_4263), .B1(net_3725), .B2(net_3724) );
NAND2_X4 inst_3361 ( .A2(net_8871), .A1(net_8870), .ZN(net_8164) );
NAND3_X2 inst_3170 ( .A3(net_8940), .ZN(net_8902), .A1(net_8591), .A2(net_8408) );
OR2_X4 inst_741 ( .ZN(net_7018), .A1(net_5955), .A2(net_4974) );
NAND3_X2 inst_3232 ( .ZN(net_4896), .A1(net_4895), .A3(net_4607), .A2(net_4606) );
DFF_X2 inst_8335 ( .Q(net_10385), .D(net_3555), .CK(net_12473) );
CLKBUF_X2 inst_13062 ( .A(net_12980), .Z(net_12981) );
AOI22_X2 inst_9377 ( .B1(net_10015), .A1(net_6821), .A2(net_5743), .B2(net_5742), .ZN(net_5528) );
AND2_X2 inst_10524 ( .ZN(net_4126), .A1(net_4125), .A2(net_4124) );
AND2_X4 inst_10444 ( .A1(net_10260), .ZN(net_3111), .A2(net_1394) );
INV_X2 inst_7195 ( .A(net_10528), .ZN(net_872) );
INV_X4 inst_5973 ( .A(net_9562), .ZN(net_3364) );
DFF_X1 inst_8700 ( .D(net_6776), .Q(net_110), .CK(net_15094) );
INV_X2 inst_6942 ( .A(net_3985), .ZN(net_1913) );
AOI22_X2 inst_9338 ( .B1(net_9814), .A2(net_5766), .B2(net_5765), .ZN(net_5614), .A1(net_252) );
OAI222_X2 inst_1350 ( .B1(net_7728), .A2(net_7727), .C2(net_7726), .ZN(net_7330), .B2(net_6914), .A1(net_5243), .C1(net_1304) );
CLKBUF_X2 inst_12156 ( .A(net_12074), .Z(net_12075) );
AOI21_X2 inst_10178 ( .ZN(net_3597), .A(net_3595), .B1(net_3594), .B2(net_3593) );
CLKBUF_X2 inst_12964 ( .A(net_12882), .Z(net_12883) );
NOR2_X2 inst_3012 ( .A1(net_5100), .A2(net_5011), .ZN(net_4125) );
CLKBUF_X2 inst_11369 ( .A(net_11287), .Z(net_11288) );
NOR2_X2 inst_2635 ( .A2(net_5927), .ZN(net_5920), .A1(net_2171) );
DFF_X2 inst_8124 ( .Q(net_9739), .D(net_5137), .CK(net_14294) );
NOR2_X2 inst_2828 ( .A2(net_3172), .ZN(net_3089), .A1(net_1959) );
CLKBUF_X2 inst_14014 ( .A(net_13932), .Z(net_13933) );
DFF_X1 inst_8673 ( .D(net_6748), .Q(net_105), .CK(net_14256) );
CLKBUF_X2 inst_13560 ( .A(net_13478), .Z(net_13479) );
DFF_X2 inst_7769 ( .Q(net_9719), .D(net_6535), .CK(net_12796) );
NAND2_X2 inst_3877 ( .ZN(net_4031), .A2(net_4027), .A1(net_1856) );
NAND2_X4 inst_3363 ( .A1(net_8976), .A2(net_8920), .ZN(net_7973) );
INV_X4 inst_4745 ( .A(net_10398), .ZN(net_5903) );
AOI221_X2 inst_9859 ( .A(net_6889), .B2(net_6888), .C2(net_6887), .ZN(net_6859), .B1(net_1215), .C1(x4851) );
NOR2_X2 inst_2666 ( .A2(net_9073), .A1(net_8117), .ZN(net_5812) );
INV_X2 inst_7320 ( .ZN(net_9111), .A(net_959) );
INV_X2 inst_7188 ( .A(net_9352), .ZN(net_7668) );
OAI22_X2 inst_1131 ( .A1(net_7226), .A2(net_5151), .B2(net_5150), .ZN(net_5147), .B1(net_409) );
CLKBUF_X2 inst_14617 ( .A(net_10741), .Z(net_14536) );
OAI222_X2 inst_1357 ( .B1(net_7665), .A2(net_7664), .C2(net_7663), .ZN(net_6932), .B2(net_5977), .A1(net_4426), .C1(net_1142) );
OR3_X4 inst_691 ( .ZN(net_6480), .A1(net_5171), .A3(net_4786), .A2(net_4628) );
CLKBUF_X2 inst_14538 ( .A(net_14456), .Z(net_14457) );
CLKBUF_X2 inst_11769 ( .A(net_11687), .Z(net_11688) );
CLKBUF_X2 inst_10938 ( .A(net_10545), .Z(net_10857) );
AOI22_X2 inst_9547 ( .B1(net_9902), .A1(net_9672), .A2(net_5966), .B2(net_4969), .ZN(net_3774) );
INV_X4 inst_6402 ( .A(net_9744), .ZN(net_1429) );
CLKBUF_X2 inst_12845 ( .A(net_12763), .Z(net_12764) );
OR2_X4 inst_770 ( .ZN(net_3188), .A2(net_3187), .A1(net_2318) );
SDFF_X2 inst_565 ( .D(net_9149), .SE(net_933), .CK(net_11048), .SI(x1459), .Q(x1104) );
OAI21_X2 inst_1971 ( .B1(net_3628), .B2(net_3558), .ZN(net_3159), .A(net_3158) );
SDFF_X2 inst_622 ( .Q(net_9444), .D(net_9444), .SE(net_3293), .CK(net_11366), .SI(x2890) );
INV_X4 inst_5302 ( .ZN(net_1533), .A(net_1299) );
DFF_X2 inst_7418 ( .QN(net_9418), .D(net_8346), .CK(net_11698) );
CLKBUF_X2 inst_14345 ( .A(net_14263), .Z(net_14264) );
CLKBUF_X2 inst_12342 ( .A(net_12260), .Z(net_12261) );
MUX2_X1 inst_4476 ( .S(net_6041), .A(net_3976), .B(x6445), .Z(x413) );
CLKBUF_X2 inst_14531 ( .A(net_14449), .Z(net_14450) );
CLKBUF_X2 inst_11307 ( .A(net_11225), .Z(net_11226) );
INV_X2 inst_6861 ( .A(net_3417), .ZN(net_3281) );
CLKBUF_X2 inst_11679 ( .A(net_11363), .Z(net_11598) );
XNOR2_X2 inst_409 ( .A(net_9371), .B(net_7632), .ZN(net_2995) );
CLKBUF_X2 inst_12323 ( .A(net_12241), .Z(net_12242) );
OAI211_X2 inst_2288 ( .C1(net_7294), .C2(net_6548), .ZN(net_6178), .B(net_5400), .A(net_3679) );
CLKBUF_X2 inst_13644 ( .A(net_11460), .Z(net_13563) );
CLKBUF_X2 inst_11505 ( .A(net_11423), .Z(net_11424) );
INV_X2 inst_6672 ( .ZN(net_8356), .A(net_8296) );
INV_X4 inst_5813 ( .ZN(net_2721), .A(net_681) );
INV_X4 inst_4841 ( .ZN(net_3325), .A(net_3116) );
CLKBUF_X2 inst_15611 ( .A(net_15529), .Z(net_15530) );
AOI22_X2 inst_9368 ( .B1(net_9913), .A2(net_5759), .B2(net_5758), .ZN(net_5554), .A1(net_252) );
OAI21_X2 inst_1834 ( .ZN(net_6291), .A(net_6013), .B2(net_5824), .B1(net_1589) );
CLKBUF_X2 inst_12933 ( .A(net_12851), .Z(net_12852) );
DFF_X2 inst_8013 ( .QN(net_10332), .D(net_5492), .CK(net_14468) );
NAND2_X2 inst_3506 ( .ZN(net_8967), .A2(net_8130), .A1(net_424) );
NAND2_X2 inst_3574 ( .ZN(net_8086), .A1(net_7572), .A2(net_7571) );
OAI211_X2 inst_2228 ( .C1(net_7243), .C2(net_6480), .ZN(net_6476), .B(net_5677), .A(net_3679) );
AOI22_X2 inst_9220 ( .A1(net_9913), .B1(net_9814), .B2(net_6140), .A2(net_6109), .ZN(net_6091) );
CLKBUF_X2 inst_11947 ( .A(net_11865), .Z(net_11866) );
INV_X2 inst_7092 ( .ZN(net_1106), .A(net_1105) );
DFF_X2 inst_7396 ( .D(net_8547), .Q(net_222), .CK(net_12380) );
CLKBUF_X2 inst_11389 ( .A(net_11307), .Z(net_11308) );
CLKBUF_X2 inst_15198 ( .A(net_10880), .Z(net_15117) );
OR2_X4 inst_768 ( .ZN(net_4491), .A1(net_4324), .A2(net_4073) );
DFF_X2 inst_7795 ( .Q(net_9910), .D(net_6498), .CK(net_12048) );
SDFF_X2 inst_663 ( .SI(net_9476), .Q(net_9476), .SE(net_3073), .CK(net_12405), .D(x2890) );
OAI211_X2 inst_2121 ( .C2(net_6778), .ZN(net_6727), .A(net_6354), .B(net_6089), .C1(net_526) );
INV_X4 inst_4850 ( .ZN(net_3685), .A(net_3297) );
NAND3_X2 inst_3227 ( .ZN(net_5222), .A3(net_4951), .A1(net_4950), .A2(net_2898) );
CLKBUF_X2 inst_12067 ( .A(net_11985), .Z(net_11986) );
INV_X4 inst_6639 ( .A(net_9077), .ZN(net_9076) );
CLKBUF_X2 inst_11001 ( .A(net_10919), .Z(net_10920) );
CLKBUF_X2 inst_13225 ( .A(net_11666), .Z(net_13144) );
INV_X2 inst_6774 ( .ZN(net_6027), .A(net_5848) );
NAND2_X2 inst_3494 ( .A2(net_8397), .ZN(net_8259), .A1(net_8173) );
NAND2_X2 inst_4224 ( .A1(net_8687), .ZN(net_1657), .A2(net_111) );
OAI21_X2 inst_1867 ( .ZN(net_5907), .A(net_5345), .B1(net_5344), .B2(net_5343) );
CLKBUF_X2 inst_13627 ( .A(net_13330), .Z(net_13546) );
INV_X4 inst_6314 ( .A(net_10024), .ZN(net_5096) );
DFF_X2 inst_7580 ( .Q(net_10505), .D(net_7538), .CK(net_14568) );
INV_X2 inst_7046 ( .ZN(net_2032), .A(net_1103) );
INV_X2 inst_7279 ( .A(net_8964), .ZN(net_8963) );
OAI211_X2 inst_2290 ( .B(net_10534), .ZN(net_5355), .C2(net_5155), .A(net_3679), .C1(net_1242) );
CLKBUF_X2 inst_13782 ( .A(net_12231), .Z(net_13701) );
DFF_X2 inst_7909 ( .QN(net_10472), .D(net_5822), .CK(net_11389) );
CLKBUF_X2 inst_11913 ( .A(net_11831), .Z(net_11832) );
INV_X4 inst_5670 ( .A(net_2410), .ZN(net_2378) );
CLKBUF_X2 inst_15222 ( .A(net_15140), .Z(net_15141) );
INV_X2 inst_6791 ( .ZN(net_5781), .A(net_5395) );
INV_X4 inst_5070 ( .ZN(net_2224), .A(net_1851) );
CLKBUF_X2 inst_13695 ( .A(net_11008), .Z(net_13614) );
CLKBUF_X2 inst_12575 ( .A(net_12493), .Z(net_12494) );
INV_X4 inst_5797 ( .ZN(net_1385), .A(net_793) );
CLKBUF_X2 inst_14143 ( .A(net_14061), .Z(net_14062) );
INV_X4 inst_4912 ( .ZN(net_3310), .A(net_2833) );
NAND2_X4 inst_3342 ( .ZN(net_9031), .A2(net_8910), .A1(net_8909) );
INV_X4 inst_4825 ( .A(net_7157), .ZN(net_6546) );
AOI221_X2 inst_9832 ( .A(net_6889), .B2(net_6888), .C2(net_6887), .ZN(net_6886), .B1(net_5861), .C1(x5427) );
CLKBUF_X2 inst_14640 ( .A(net_14558), .Z(net_14559) );
NOR2_X2 inst_2621 ( .ZN(net_6181), .A1(net_5764), .A2(net_3972) );
CLKBUF_X2 inst_14666 ( .A(net_14584), .Z(net_14585) );
CLKBUF_X2 inst_15743 ( .A(net_13042), .Z(net_15662) );
DFF_X2 inst_8175 ( .QN(net_9926), .D(net_5037), .CK(net_12118) );
AOI22_X2 inst_9159 ( .A2(net_6418), .ZN(net_6322), .A1(net_6321), .B2(net_5263), .B1(net_2988) );
CLKBUF_X2 inst_10815 ( .A(net_10733), .Z(net_10734) );
CLKBUF_X2 inst_14454 ( .A(net_14372), .Z(net_14373) );
NAND2_X2 inst_3895 ( .ZN(net_4119), .A2(net_3963), .A1(net_986) );
CLKBUF_X2 inst_11928 ( .A(net_11846), .Z(net_11847) );
AOI22_X2 inst_9358 ( .B1(net_9914), .A2(net_5759), .B2(net_5758), .ZN(net_5564), .A1(net_253) );
XNOR2_X2 inst_303 ( .ZN(net_3273), .B(net_3272), .A(net_3025) );
CLKBUF_X2 inst_13518 ( .A(net_13436), .Z(net_13437) );
CLKBUF_X2 inst_14324 ( .A(net_12728), .Z(net_14243) );
DFF_X2 inst_7699 ( .QN(net_9204), .D(net_6554), .CK(net_11324) );
NAND3_X2 inst_3263 ( .A2(net_5337), .ZN(net_4354), .A3(net_3868), .A1(net_2910) );
OAI221_X2 inst_1647 ( .C1(net_10414), .B1(net_7241), .ZN(net_5541), .C2(net_4477), .B2(net_4455), .A(net_3731) );
CLKBUF_X2 inst_12114 ( .A(net_10651), .Z(net_12033) );
OAI22_X2 inst_1275 ( .B1(net_8122), .ZN(net_4597), .A2(net_4159), .B2(net_4158), .A1(net_3701) );
XOR2_X2 inst_26 ( .A(net_10324), .B(net_5486), .Z(net_2267) );
CLKBUF_X2 inst_15326 ( .A(net_14895), .Z(net_15245) );
CLKBUF_X2 inst_13052 ( .A(net_12970), .Z(net_12971) );
AND2_X2 inst_10480 ( .A2(net_9579), .ZN(net_8685), .A1(net_807) );
DFF_X2 inst_8104 ( .QN(net_9842), .D(net_5127), .CK(net_12898) );
AOI21_X2 inst_10198 ( .ZN(net_2885), .B1(net_1804), .A(net_1625), .B2(net_1577) );
NOR2_X2 inst_2882 ( .ZN(net_2516), .A1(net_1815), .A2(net_1814) );
OAI222_X2 inst_1376 ( .B2(net_7660), .A2(net_7659), .C2(net_7658), .ZN(net_6010), .B1(net_4106), .A1(net_2816), .C1(net_1916) );
CLKBUF_X2 inst_12731 ( .A(net_12649), .Z(net_12650) );
CLKBUF_X2 inst_14038 ( .A(net_13652), .Z(net_13957) );
CLKBUF_X2 inst_12605 ( .A(net_12523), .Z(net_12524) );
AND2_X2 inst_10507 ( .ZN(net_5318), .A1(net_5317), .A2(net_5316) );
AOI21_X4 inst_10001 ( .B1(net_9019), .ZN(net_7040), .B2(net_6892), .A(net_3388) );
INV_X4 inst_6530 ( .ZN(net_7211), .A(x5289) );
DFF_X2 inst_7490 ( .D(net_8037), .Q(net_205), .CK(net_12521) );
CLKBUF_X2 inst_12895 ( .A(net_10549), .Z(net_12814) );
CLKBUF_X2 inst_11483 ( .A(net_11322), .Z(net_11402) );
DFF_X2 inst_8182 ( .Q(net_10532), .D(net_5026), .CK(net_14881) );
INV_X4 inst_4864 ( .ZN(net_5966), .A(net_2954) );
CLKBUF_X2 inst_10654 ( .A(net_10572), .Z(net_10573) );
INV_X4 inst_6188 ( .ZN(net_472), .A(x494) );
NAND2_X2 inst_3765 ( .ZN(net_4975), .A2(net_4974), .A1(net_4706) );
CLKBUF_X2 inst_10742 ( .A(net_10608), .Z(net_10661) );
OAI221_X2 inst_1659 ( .C1(net_7213), .C2(net_5520), .ZN(net_5512), .B1(net_5511), .B2(net_4547), .A(net_3507) );
NAND2_X2 inst_4218 ( .A2(net_3171), .ZN(net_1673), .A1(net_648) );
DFF_X2 inst_7718 ( .Q(net_9709), .D(net_6178), .CK(net_15072) );
CLKBUF_X2 inst_15808 ( .A(net_15726), .Z(net_15727) );
AOI21_X2 inst_10062 ( .ZN(net_7073), .B1(net_7068), .B2(net_7067), .A(net_6053) );
INV_X4 inst_6456 ( .A(net_10262), .ZN(net_2628) );
XNOR2_X2 inst_398 ( .ZN(net_1773), .A(net_1772), .B(net_787) );
INV_X4 inst_5702 ( .A(net_3884), .ZN(net_2246) );
DFF_X2 inst_8184 ( .Q(net_9953), .D(net_5000), .CK(net_13186) );
XNOR2_X2 inst_436 ( .B(net_9305), .ZN(net_1044), .A(net_228) );
INV_X2 inst_7064 ( .A(net_3546), .ZN(net_1266) );
CLKBUF_X2 inst_13265 ( .A(net_13183), .Z(net_13184) );
CLKBUF_X2 inst_11766 ( .A(net_11296), .Z(net_11685) );
AOI221_X2 inst_9852 ( .B1(net_9772), .B2(net_9097), .A(net_6940), .C1(net_6939), .ZN(net_6866), .C2(net_242) );
INV_X4 inst_6529 ( .A(net_9299), .ZN(net_608) );
CLKBUF_X2 inst_11636 ( .A(net_11554), .Z(net_11555) );
CLKBUF_X2 inst_13702 ( .A(net_13620), .Z(net_13621) );
NAND2_X2 inst_3705 ( .A1(net_10068), .ZN(net_5924), .A2(net_5894) );
DFF_X2 inst_7623 ( .D(net_6698), .QN(net_177), .CK(net_12744) );
CLKBUF_X2 inst_11469 ( .A(net_11387), .Z(net_11388) );
INV_X4 inst_5053 ( .ZN(net_5043), .A(net_1885) );
INV_X2 inst_6746 ( .ZN(net_6841), .A(net_6620) );
OAI211_X2 inst_2231 ( .A(net_8098), .C1(net_7221), .C2(net_6480), .ZN(net_6473), .B(net_5529) );
CLKBUF_X2 inst_15137 ( .A(net_15055), .Z(net_15056) );
XNOR2_X2 inst_144 ( .ZN(net_7138), .A(net_6986), .B(net_1923) );
OAI222_X1 inst_1438 ( .A1(net_7665), .B2(net_7664), .C2(net_7663), .ZN(net_7606), .A2(net_7463), .B1(net_5182), .C1(net_1082) );
AOI221_X2 inst_9750 ( .C1(net_9366), .C2(net_8783), .A(net_7916), .B2(net_7915), .ZN(net_7913), .B1(net_7905) );
AND2_X4 inst_10454 ( .A1(net_10365), .ZN(net_3114), .A2(net_908) );
AND2_X2 inst_10565 ( .ZN(net_3479), .A2(net_3027), .A1(net_2686) );
INV_X4 inst_6373 ( .A(net_10360), .ZN(net_1351) );
CLKBUF_X2 inst_13660 ( .A(net_13578), .Z(net_13579) );
CLKBUF_X2 inst_12681 ( .A(net_12599), .Z(net_12600) );
OR2_X2 inst_880 ( .A2(net_7038), .ZN(net_6428), .A1(net_6427) );
INV_X2 inst_6912 ( .A(net_2239), .ZN(net_2221) );
INV_X4 inst_4857 ( .ZN(net_4371), .A(net_3287) );
AOI221_X2 inst_9763 ( .ZN(net_7643), .B1(net_7642), .C2(net_7641), .A(net_7523), .C1(net_6854), .B2(net_6185) );
CLKBUF_X2 inst_12241 ( .A(net_12159), .Z(net_12160) );
CLKBUF_X2 inst_11437 ( .A(net_11355), .Z(net_11356) );
NOR2_X2 inst_2681 ( .ZN(net_5359), .A2(net_4640), .A1(net_4547) );
NAND2_X2 inst_3445 ( .A2(net_9451), .ZN(net_8908), .A1(net_8477) );
AOI21_X2 inst_10026 ( .B1(net_9366), .A(net_7916), .B2(net_7915), .ZN(net_7853) );
INV_X4 inst_5555 ( .A(net_10459), .ZN(net_1092) );
MUX2_X1 inst_4447 ( .S(net_6041), .A(net_299), .B(x4937), .Z(x116) );
AOI22_X2 inst_9118 ( .A1(net_9694), .A2(net_6418), .ZN(net_6371), .B2(net_5263), .B1(net_134) );
CLKBUF_X2 inst_12370 ( .A(net_11186), .Z(net_12289) );
INV_X4 inst_6194 ( .A(net_9362), .ZN(net_8595) );
DFF_X1 inst_8493 ( .QN(net_9635), .D(net_7899), .CK(net_13793) );
CLKBUF_X2 inst_15694 ( .A(net_15612), .Z(net_15613) );
AOI22_X2 inst_9044 ( .A1(net_9152), .A2(net_7155), .B2(net_7154), .ZN(net_7011), .B1(net_1990) );
NAND2_X2 inst_3972 ( .A1(net_4273), .ZN(net_3652), .A2(net_3040) );
INV_X2 inst_6670 ( .ZN(net_8358), .A(net_8298) );
CLKBUF_X2 inst_11633 ( .A(net_11551), .Z(net_11552) );
OAI222_X2 inst_1388 ( .B1(net_7728), .A2(net_7727), .C2(net_7726), .ZN(net_5869), .B2(net_5211), .A1(net_4195), .C1(net_1882) );
NOR2_X2 inst_2699 ( .A2(net_4552), .ZN(net_4392), .A1(net_2396) );
CLKBUF_X2 inst_12470 ( .A(net_10556), .Z(net_12389) );
INV_X4 inst_6329 ( .ZN(net_5374), .A(net_273) );
NAND2_X2 inst_3517 ( .A2(net_9594), .A1(net_8983), .ZN(net_8152) );
AOI22_X2 inst_9291 ( .B1(net_9805), .A1(net_5766), .B2(net_5765), .ZN(net_5706), .A2(net_243) );
CLKBUF_X2 inst_14937 ( .A(net_14855), .Z(net_14856) );
CLKBUF_X2 inst_14927 ( .A(net_14845), .Z(net_14846) );
DFF_X1 inst_8506 ( .QN(net_10268), .D(net_7666), .CK(net_11713) );
NAND2_X2 inst_3396 ( .A2(net_9084), .A1(net_9041), .ZN(net_8669) );
OAI222_X2 inst_1372 ( .B1(net_7665), .A2(net_7664), .C2(net_7663), .ZN(net_6038), .B2(net_5207), .A1(net_3674), .C1(net_1877) );
OAI222_X2 inst_1360 ( .B1(net_7728), .A2(net_7727), .C2(net_7726), .ZN(net_6922), .B2(net_5946), .A1(net_4314), .C1(net_1901) );
HA_X1 inst_7332 ( .S(net_7565), .CO(net_7564), .B(net_7468), .A(net_861) );
CLKBUF_X2 inst_12109 ( .A(net_11963), .Z(net_12028) );
CLKBUF_X2 inst_10631 ( .A(net_10549), .Z(net_10550) );
AOI221_X2 inst_9759 ( .A(net_7749), .B2(net_7748), .C2(net_7747), .ZN(net_7743), .C1(net_7677), .B1(net_393) );
SDFF_X2 inst_466 ( .SE(net_8756), .SI(net_8634), .Q(net_237), .D(net_106), .CK(net_13848) );
INV_X4 inst_6081 ( .ZN(net_7213), .A(x4041) );
NAND2_X2 inst_3981 ( .A1(net_10057), .A2(net_10056), .ZN(net_3257) );
NOR2_X2 inst_2761 ( .ZN(net_5353), .A1(net_5180), .A2(net_3263) );
OAI22_X2 inst_989 ( .A2(net_8962), .B2(net_8659), .ZN(net_8651), .B1(net_8326), .A1(net_6656) );
CLKBUF_X2 inst_14742 ( .A(net_14562), .Z(net_14661) );
INV_X4 inst_5205 ( .ZN(net_1894), .A(net_1528) );
CLKBUF_X2 inst_15087 ( .A(net_12210), .Z(net_15006) );
OAI211_X2 inst_2283 ( .C1(net_7108), .C2(net_6548), .ZN(net_6196), .B(net_5724), .A(net_3679) );
AOI21_X2 inst_10073 ( .B1(net_7928), .B2(net_7721), .ZN(net_6584), .A(net_6186) );
NAND4_X2 inst_3038 ( .ZN(net_8504), .A1(net_8410), .A2(net_8258), .A4(net_8111), .A3(net_8083) );
CLKBUF_X2 inst_14154 ( .A(net_14072), .Z(net_14073) );
OR2_X2 inst_858 ( .A2(net_9600), .A1(net_8965), .ZN(net_8538) );
DFF_X2 inst_7605 ( .Q(net_9310), .D(net_7327), .CK(net_14098) );
DFF_X2 inst_7542 ( .QN(net_9353), .D(net_7758), .CK(net_11851) );
NAND2_X2 inst_3864 ( .ZN(net_4915), .A1(net_4103), .A2(net_4098) );
AOI22_X2 inst_9111 ( .A1(net_9664), .A2(net_6402), .ZN(net_6378), .B2(net_5263), .B1(net_102) );
CLKBUF_X2 inst_15482 ( .A(net_15400), .Z(net_15401) );
CLKBUF_X2 inst_13779 ( .A(net_13697), .Z(net_13698) );
CLKBUF_X2 inst_12060 ( .A(net_11370), .Z(net_11979) );
CLKBUF_X2 inst_12735 ( .A(net_12653), .Z(net_12654) );
NOR2_X2 inst_2936 ( .A1(net_10460), .A2(net_2702), .ZN(net_1348) );
NOR2_X4 inst_2468 ( .ZN(net_8561), .A1(net_8523), .A2(net_8522) );
XOR2_X1 inst_54 ( .Z(net_2125), .A(net_1814), .B(net_984) );
CLKBUF_X2 inst_15596 ( .A(net_15514), .Z(net_15515) );
CLKBUF_X2 inst_12610 ( .A(net_10762), .Z(net_12529) );
AND2_X2 inst_10556 ( .A1(net_9619), .ZN(net_3653), .A2(net_3308) );
OAI221_X2 inst_1482 ( .ZN(net_7590), .B2(net_7589), .C2(net_7557), .A(net_7490), .C1(net_3691), .B1(net_3092) );
OAI222_X2 inst_1420 ( .B2(net_7665), .A2(net_7664), .C2(net_7663), .ZN(net_4924), .B1(net_4257), .A1(net_3271), .C1(net_1147) );
AOI221_X2 inst_9757 ( .A(net_7749), .B2(net_7748), .C2(net_7747), .ZN(net_7746), .C1(net_7681), .B1(net_1123) );
DFF_X2 inst_7406 ( .QN(net_9389), .D(net_8367), .CK(net_14032) );
CLKBUF_X2 inst_12177 ( .A(net_12095), .Z(net_12096) );
CLKBUF_X2 inst_12988 ( .A(net_12906), .Z(net_12907) );
INV_X4 inst_5214 ( .ZN(net_1982), .A(net_1521) );
INV_X2 inst_7283 ( .ZN(net_8973), .A(net_8972) );
INV_X4 inst_5337 ( .ZN(net_5032), .A(net_3429) );
CLKBUF_X2 inst_15170 ( .A(net_15088), .Z(net_15089) );
NAND2_X2 inst_4062 ( .ZN(net_7586), .A2(net_3347), .A1(net_2757) );
CLKBUF_X2 inst_13331 ( .A(net_13249), .Z(net_13250) );
INV_X4 inst_5730 ( .ZN(net_1146), .A(net_823) );
CLKBUF_X2 inst_15775 ( .A(net_15693), .Z(net_15694) );
CLKBUF_X2 inst_15685 ( .A(net_15603), .Z(net_15604) );
NAND2_X2 inst_4108 ( .ZN(net_2669), .A2(net_2368), .A1(net_1666) );
INV_X4 inst_4626 ( .ZN(net_7457), .A(net_6919) );
DFF_X1 inst_8780 ( .Q(net_10238), .D(net_4610), .CK(net_10915) );
CLKBUF_X2 inst_13838 ( .A(net_13756), .Z(net_13757) );
INV_X4 inst_4794 ( .ZN(net_7770), .A(net_4092) );
CLKBUF_X2 inst_13688 ( .A(net_13606), .Z(net_13607) );
CLKBUF_X2 inst_10804 ( .A(net_10722), .Z(net_10723) );
AOI22_X2 inst_9491 ( .B1(net_9818), .A1(net_9687), .A2(net_5966), .ZN(net_3832), .B2(net_2556) );
CLKBUF_X2 inst_11595 ( .A(net_11513), .Z(net_11514) );
NAND2_X2 inst_3829 ( .ZN(net_7730), .A2(net_4444), .A1(net_587) );
CLKBUF_X2 inst_14465 ( .A(net_14383), .Z(net_14384) );
DFF_X2 inst_7883 ( .QN(net_10106), .D(net_6034), .CK(net_14807) );
CLKBUF_X2 inst_15496 ( .A(net_15414), .Z(net_15415) );
CLKBUF_X2 inst_14621 ( .A(net_14539), .Z(net_14540) );
CLKBUF_X2 inst_13414 ( .A(net_12935), .Z(net_13333) );
AOI22_X2 inst_9012 ( .B1(net_9307), .A2(net_8030), .B2(net_8029), .ZN(net_8024), .A1(net_215) );
CLKBUF_X2 inst_15272 ( .A(net_15190), .Z(net_15191) );
SDFF_X2 inst_497 ( .SE(net_9540), .SI(net_8212), .Q(net_286), .D(net_286), .CK(net_12701) );
CLKBUF_X2 inst_10971 ( .A(net_10889), .Z(net_10890) );
AND4_X4 inst_10325 ( .ZN(net_3355), .A2(net_3354), .A3(net_3353), .A4(net_3352), .A1(net_2750) );
CLKBUF_X2 inst_15791 ( .A(net_15709), .Z(net_15710) );
CLKBUF_X2 inst_13918 ( .A(net_11396), .Z(net_13837) );
CLKBUF_X2 inst_13826 ( .A(net_11549), .Z(net_13745) );
DFF_X2 inst_7517 ( .QN(net_10466), .D(net_7844), .CK(net_11410) );
OAI211_X2 inst_2195 ( .C1(net_7226), .C2(net_6542), .ZN(net_6512), .B(net_5610), .A(net_3527) );
DFF_X2 inst_8161 ( .QN(net_9733), .D(net_5059), .CK(net_12265) );
DFF_X1 inst_8787 ( .Q(net_10449), .D(net_4572), .CK(net_11073) );
OAI211_X2 inst_2168 ( .C1(net_7243), .C2(net_6548), .ZN(net_6541), .B(net_5670), .A(net_3679) );
OAI222_X2 inst_1335 ( .ZN(net_7666), .A1(net_7665), .B2(net_7664), .C2(net_7663), .A2(net_7551), .B1(net_7032), .C1(net_628) );
CLKBUF_X2 inst_15197 ( .A(net_15115), .Z(net_15116) );
AOI221_X2 inst_9924 ( .B2(net_5867), .A(net_5862), .ZN(net_5857), .C1(net_5856), .C2(net_5853), .B1(x5289) );
NAND2_X2 inst_3845 ( .ZN(net_4517), .A1(net_4237), .A2(net_4081) );
INV_X2 inst_7173 ( .A(net_9394), .ZN(net_8212) );
AOI21_X2 inst_10124 ( .ZN(net_4418), .B1(net_4412), .B2(net_4411), .A(net_3133) );
INV_X4 inst_5168 ( .A(net_1568), .ZN(net_1565) );
INV_X2 inst_7241 ( .A(net_9313), .ZN(net_7685) );
NAND4_X2 inst_3128 ( .ZN(net_2936), .A4(net_2720), .A3(net_2487), .A1(net_2222), .A2(net_1967) );
CLKBUF_X2 inst_15060 ( .A(net_14978), .Z(net_14979) );
CLKBUF_X2 inst_10715 ( .A(net_10576), .Z(net_10634) );
OAI22_X2 inst_1078 ( .A2(net_9064), .ZN(net_6640), .B2(net_6639), .B1(net_4303), .A1(net_1505) );
NAND2_X2 inst_4322 ( .ZN(net_2674), .A2(net_1146), .A1(net_692) );
CLKBUF_X2 inst_14653 ( .A(net_14571), .Z(net_14572) );
NOR2_X2 inst_2517 ( .A2(net_8318), .ZN(net_8264), .A1(net_8263) );
INV_X4 inst_6497 ( .A(net_9298), .ZN(net_593) );
NAND2_X2 inst_4183 ( .A1(net_5268), .A2(net_2612), .ZN(net_1953) );
CLKBUF_X2 inst_10806 ( .A(net_10724), .Z(net_10725) );
NAND2_X2 inst_3557 ( .A1(net_8960), .A2(net_8916), .ZN(net_7861) );
OAI21_X2 inst_1992 ( .B1(net_5469), .ZN(net_2494), .A(net_2117), .B2(net_1745) );
OAI22_X2 inst_1039 ( .A1(net_8981), .B1(net_8919), .A2(net_8915), .ZN(net_7947), .B2(net_2875) );
OR3_X2 inst_714 ( .ZN(net_4358), .A1(net_4357), .A2(net_4356), .A3(net_4355) );
CLKBUF_X2 inst_15735 ( .A(net_15653), .Z(net_15654) );
CLKBUF_X2 inst_15518 ( .A(net_15436), .Z(net_15437) );
NOR2_X2 inst_3005 ( .A2(net_2818), .A1(net_2139), .ZN(net_855) );
NOR2_X2 inst_2895 ( .ZN(net_1967), .A2(net_1681), .A1(net_1129) );
INV_X4 inst_5449 ( .A(net_5268), .ZN(net_3068) );
AOI22_X2 inst_9005 ( .A2(net_9758), .ZN(net_8040), .A1(net_6420), .B2(net_5263), .B1(net_2706) );
NAND2_X2 inst_4048 ( .ZN(net_3266), .A2(net_2812), .A1(net_1315) );
DFF_X2 inst_7549 ( .QN(net_9240), .D(net_7707), .CK(net_11267) );
NAND2_X2 inst_4003 ( .ZN(net_7434), .A2(net_3390), .A1(net_1643) );
INV_X2 inst_6868 ( .ZN(net_3108), .A(net_3107) );
CLKBUF_X2 inst_15512 ( .A(net_11736), .Z(net_15431) );
DFF_X2 inst_8306 ( .QN(net_10454), .D(net_4571), .CK(net_11193) );
OAI22_X2 inst_1061 ( .A2(net_7167), .ZN(net_7017), .B1(net_3889), .B2(net_3361), .A1(net_3206) );
INV_X4 inst_5033 ( .ZN(net_5027), .A(net_1935) );
CLKBUF_X2 inst_13966 ( .A(net_13884), .Z(net_13885) );
CLKBUF_X2 inst_11201 ( .A(net_11119), .Z(net_11120) );
NOR4_X2 inst_2326 ( .ZN(net_5814), .A1(net_5813), .A4(net_5812), .A3(net_4996), .A2(net_4732) );
DFF_X1 inst_8846 ( .Q(net_8832), .D(net_1497), .CK(net_14574) );
INV_X4 inst_5363 ( .ZN(net_5484), .A(net_1219) );
INV_X2 inst_6657 ( .A(net_9433), .ZN(net_8491) );
XNOR2_X2 inst_72 ( .A(net_8943), .ZN(net_8694), .B(net_8265) );
INV_X2 inst_6967 ( .ZN(net_1823), .A(net_1822) );
CLKBUF_X2 inst_11703 ( .A(net_10601), .Z(net_11622) );
CLKBUF_X2 inst_15529 ( .A(net_12186), .Z(net_15448) );
NAND2_X2 inst_3542 ( .A2(net_9058), .ZN(net_8871), .A1(net_7989) );
OAI221_X2 inst_1634 ( .B1(net_10311), .C1(net_7124), .A(net_6546), .B2(net_5591), .ZN(net_5572), .C2(net_4902) );
AOI22_X2 inst_8998 ( .B1(net_9485), .A1(net_9477), .ZN(net_8500), .B2(net_8490), .A2(net_8487) );
INV_X4 inst_6300 ( .A(net_9238), .ZN(net_1643) );
XNOR2_X2 inst_115 ( .B(net_9426), .ZN(net_7889), .A(net_6219) );
DFF_X2 inst_7980 ( .QN(net_10422), .D(net_5574), .CK(net_15485) );
AND2_X2 inst_10619 ( .A1(net_9652), .ZN(net_2166), .A2(net_1564) );
INV_X2 inst_6729 ( .ZN(net_7695), .A(net_7646) );
INV_X2 inst_6650 ( .ZN(net_8773), .A(net_8768) );
CLKBUF_X2 inst_15609 ( .A(net_15527), .Z(net_15528) );
AOI22_X2 inst_9485 ( .B1(net_9915), .A1(net_9883), .B2(net_4969), .ZN(net_3838), .A2(net_2973) );
INV_X4 inst_4691 ( .ZN(net_4836), .A(net_4652) );
NAND2_X2 inst_3726 ( .A1(net_10294), .ZN(net_5773), .A2(net_5770) );
CLKBUF_X2 inst_12415 ( .A(net_12333), .Z(net_12334) );
CLKBUF_X2 inst_12357 ( .A(net_12275), .Z(net_12276) );
INV_X4 inst_4638 ( .ZN(net_7283), .A(net_6237) );
NAND4_X2 inst_3045 ( .ZN(net_7251), .A4(net_6566), .A3(net_4720), .A1(net_4042), .A2(net_3057) );
CLKBUF_X2 inst_11487 ( .A(net_10901), .Z(net_11406) );
AOI221_X2 inst_9801 ( .B1(net_9980), .A(net_7090), .B2(net_7089), .C2(net_7088), .ZN(net_7001), .C1(net_252) );
CLKBUF_X2 inst_13426 ( .A(net_13344), .Z(net_13345) );
OAI221_X2 inst_1582 ( .C1(net_10206), .C2(net_7295), .B2(net_7293), .ZN(net_7125), .B1(net_7124), .A(net_6941) );
CLKBUF_X2 inst_13202 ( .A(net_11633), .Z(net_13121) );
CLKBUF_X2 inst_12741 ( .A(net_12659), .Z(net_12660) );
INV_X4 inst_6334 ( .A(net_10362), .ZN(net_693) );
CLKBUF_X2 inst_13905 ( .A(net_13011), .Z(net_13824) );
INV_X4 inst_5846 ( .A(net_1036), .ZN(net_873) );
OAI21_X2 inst_1840 ( .B1(net_7157), .ZN(net_6214), .A(net_5773), .B2(net_5771) );
INV_X4 inst_6345 ( .A(net_10507), .ZN(net_410) );
XNOR2_X2 inst_133 ( .ZN(net_7417), .A(net_7323), .B(net_1904) );
OAI22_X2 inst_1263 ( .B1(net_7226), .A2(net_4842), .B2(net_4841), .ZN(net_4810), .A1(net_480) );
INV_X4 inst_6113 ( .A(net_9318), .ZN(net_2481) );
CLKBUF_X2 inst_14734 ( .A(net_14652), .Z(net_14653) );
CLKBUF_X2 inst_13847 ( .A(net_13692), .Z(net_13766) );
NAND2_X4 inst_3330 ( .A1(net_8939), .A2(net_8933), .ZN(net_8604) );
DFF_X2 inst_8047 ( .QN(net_10455), .D(net_5701), .CK(net_14706) );
AOI221_X2 inst_9988 ( .B1(net_4017), .B2(net_3602), .ZN(net_3601), .C2(net_2914), .A(net_2907), .C1(net_2217) );
AOI21_X2 inst_10225 ( .ZN(net_2104), .B1(net_2103), .B2(net_2094), .A(net_1088) );
CLKBUF_X2 inst_14688 ( .A(net_10960), .Z(net_14607) );
OAI221_X2 inst_1721 ( .B2(net_3496), .ZN(net_2835), .C1(net_2412), .A(net_2077), .B1(net_1510), .C2(net_1126) );
DFF_X2 inst_7374 ( .Q(net_9368), .D(net_8683), .CK(net_14191) );
OAI221_X2 inst_1445 ( .B1(net_8565), .ZN(net_8442), .C2(net_8441), .B2(net_8255), .A(net_3904), .C1(net_1404) );
CLKBUF_X2 inst_11907 ( .A(net_11825), .Z(net_11826) );
AOI221_X2 inst_9744 ( .ZN(net_7982), .C2(net_7932), .B2(net_7930), .C1(net_7910), .A(net_7885), .B1(net_2611) );
CLKBUF_X2 inst_10884 ( .A(net_10802), .Z(net_10803) );
NAND2_X2 inst_3990 ( .A1(net_10018), .ZN(net_3184), .A2(net_2468) );
CLKBUF_X2 inst_13156 ( .A(net_13074), .Z(net_13075) );
CLKBUF_X2 inst_12854 ( .A(net_10893), .Z(net_12773) );
CLKBUF_X2 inst_12115 ( .A(net_12033), .Z(net_12034) );
XNOR2_X2 inst_126 ( .ZN(net_7485), .A(net_7096), .B(net_1692) );
INV_X4 inst_5982 ( .ZN(net_2169), .A(x6445) );
DFF_X2 inst_7931 ( .QN(net_9548), .D(net_9254), .CK(net_13765) );
OAI221_X2 inst_1512 ( .C1(net_10428), .B2(net_9063), .C2(net_9056), .ZN(net_7348), .B1(net_7182), .A(net_7007) );
DFF_X2 inst_7932 ( .QN(net_10327), .D(net_5455), .CK(net_13649) );
NAND2_X2 inst_3887 ( .A2(net_10490), .ZN(net_4639), .A1(net_4015) );
AND3_X2 inst_10366 ( .A3(net_8074), .ZN(net_8073), .A1(net_3713), .A2(net_3328) );
CLKBUF_X2 inst_14163 ( .A(net_12963), .Z(net_14082) );
INV_X4 inst_5160 ( .ZN(net_5161), .A(net_1573) );
DFF_X1 inst_8733 ( .Q(net_9120), .D(net_5870), .CK(net_10583) );
OAI221_X2 inst_1631 ( .B1(net_10309), .C1(net_7241), .B2(net_5591), .ZN(net_5576), .A(net_5575), .C2(net_4902) );
CLKBUF_X2 inst_13209 ( .A(net_13118), .Z(net_13128) );
CLKBUF_X2 inst_12651 ( .A(net_12569), .Z(net_12570) );
DFF_X2 inst_7510 ( .QN(net_9373), .D(net_7941), .CK(net_11920) );
CLKBUF_X2 inst_14395 ( .A(net_14313), .Z(net_14314) );
CLKBUF_X2 inst_13106 ( .A(net_10818), .Z(net_13025) );
OAI22_X2 inst_1086 ( .A1(net_6575), .ZN(net_6572), .A2(net_5901), .B2(net_5900), .B1(net_492) );
CLKBUF_X2 inst_14360 ( .A(net_14278), .Z(net_14279) );
CLKBUF_X2 inst_10727 ( .A(net_10645), .Z(net_10646) );
NOR2_X2 inst_2643 ( .A2(net_5449), .ZN(net_5448), .A1(net_1713) );
CLKBUF_X2 inst_12088 ( .A(net_11217), .Z(net_12007) );
CLKBUF_X2 inst_13950 ( .A(net_13830), .Z(net_13869) );
CLKBUF_X2 inst_12615 ( .A(net_10971), .Z(net_12534) );
DFF_X2 inst_7692 ( .Q(net_10298), .D(net_6573), .CK(net_14550) );
CLKBUF_X2 inst_12713 ( .A(net_12631), .Z(net_12632) );
CLKBUF_X2 inst_14822 ( .A(net_14740), .Z(net_14741) );
OAI221_X2 inst_1688 ( .B1(net_7231), .C2(net_5642), .ZN(net_5472), .B2(net_4905), .A(net_3731), .C1(net_1492) );
CLKBUF_X2 inst_11691 ( .A(net_10683), .Z(net_11610) );
OAI211_X2 inst_2299 ( .ZN(net_3362), .B(net_2847), .C1(net_2074), .C2(net_1969), .A(net_802) );
CLKBUF_X2 inst_15621 ( .A(net_15539), .Z(net_15540) );
CLKBUF_X2 inst_13651 ( .A(net_11911), .Z(net_13570) );
CLKBUF_X2 inst_12441 ( .A(net_12359), .Z(net_12360) );
CLKBUF_X2 inst_13732 ( .A(net_13650), .Z(net_13651) );
CLKBUF_X2 inst_12146 ( .A(net_12064), .Z(net_12065) );
DFF_X2 inst_7504 ( .D(net_8016), .QN(net_200), .CK(net_15158) );
INV_X4 inst_5292 ( .ZN(net_1312), .A(net_1311) );
CLKBUF_X2 inst_14836 ( .A(net_14754), .Z(net_14755) );
CLKBUF_X2 inst_13084 ( .A(net_11970), .Z(net_13003) );
OR2_X2 inst_914 ( .A1(net_9522), .ZN(net_3727), .A2(net_3482) );
INV_X4 inst_6364 ( .A(net_9221), .ZN(net_1538) );
INV_X4 inst_5170 ( .ZN(net_1887), .A(net_1562) );
DFF_X2 inst_7578 ( .QN(net_10254), .D(net_7555), .CK(net_11674) );
INV_X4 inst_5182 ( .A(net_1975), .ZN(net_1556) );
CLKBUF_X2 inst_14963 ( .A(net_14438), .Z(net_14882) );
CLKBUF_X2 inst_12366 ( .A(net_12284), .Z(net_12285) );
CLKBUF_X2 inst_12198 ( .A(net_12116), .Z(net_12117) );
DFF_X2 inst_8166 ( .QN(net_9730), .D(net_5050), .CK(net_12261) );
CLKBUF_X2 inst_14962 ( .A(net_14880), .Z(net_14881) );
CLKBUF_X2 inst_11588 ( .A(net_11506), .Z(net_11507) );
OAI221_X2 inst_1642 ( .B1(net_10425), .C1(net_7294), .ZN(net_5546), .B2(net_4477), .C2(net_4455), .A(net_3731) );
XNOR2_X2 inst_384 ( .ZN(net_2278), .B(net_1562), .A(net_1227) );
OAI22_X2 inst_1252 ( .B1(net_7216), .A2(net_4826), .B2(net_4825), .ZN(net_4822), .A1(net_419) );
CLKBUF_X2 inst_12773 ( .A(net_11641), .Z(net_12692) );
NAND2_X2 inst_3800 ( .ZN(net_4791), .A2(net_4545), .A1(net_2399) );
CLKBUF_X2 inst_12703 ( .A(net_12621), .Z(net_12622) );
CLKBUF_X2 inst_13434 ( .A(net_13352), .Z(net_13353) );
XNOR2_X2 inst_199 ( .ZN(net_4989), .B(net_4988), .A(net_4708) );
INV_X4 inst_6086 ( .A(net_9991), .ZN(net_499) );
CLKBUF_X2 inst_12540 ( .A(net_12262), .Z(net_12459) );
CLKBUF_X2 inst_13259 ( .A(net_11164), .Z(net_13178) );
CLKBUF_X2 inst_12989 ( .A(net_11122), .Z(net_12908) );
AOI211_X2 inst_10271 ( .ZN(net_7598), .B(net_7597), .C1(net_7422), .C2(net_7401), .A(net_5995) );
OAI211_X2 inst_2209 ( .C1(net_7243), .C2(net_6501), .ZN(net_6496), .B(net_5651), .A(net_3679) );
NOR2_X2 inst_2722 ( .A1(net_7932), .A2(net_5885), .ZN(net_4173) );
CLKBUF_X2 inst_13034 ( .A(net_12952), .Z(net_12953) );
OAI22_X2 inst_1238 ( .B1(net_7201), .A2(net_4890), .B2(net_4889), .ZN(net_4879), .A1(net_4100) );
INV_X2 inst_6764 ( .ZN(net_6169), .A(net_5944) );
HA_X1 inst_7361 ( .B(net_9325), .S(net_2473), .CO(net_1458), .A(net_786) );
OAI211_X2 inst_2171 ( .C1(net_7221), .C2(net_6548), .ZN(net_6538), .B(net_5666), .A(net_3679) );
CLKBUF_X2 inst_15385 ( .A(net_10783), .Z(net_15304) );
CLKBUF_X2 inst_13313 ( .A(net_13231), .Z(net_13232) );
INV_X2 inst_6976 ( .ZN(net_1683), .A(net_1682) );
AOI22_X2 inst_9031 ( .A1(net_9369), .A2(net_7638), .B2(net_7635), .ZN(net_7631), .B1(net_623) );
DFF_X2 inst_7941 ( .QN(net_10423), .D(net_5547), .CK(net_14795) );
CLKBUF_X2 inst_14274 ( .A(net_13455), .Z(net_14193) );
DFF_X1 inst_8527 ( .Q(net_9974), .D(net_7381), .CK(net_15652) );
INV_X4 inst_4875 ( .ZN(net_7620), .A(net_3088) );
NAND2_X2 inst_3402 ( .ZN(net_8590), .A1(net_8589), .A2(net_8587) );
CLKBUF_X2 inst_14252 ( .A(net_14170), .Z(net_14171) );
CLKBUF_X2 inst_15412 ( .A(net_13989), .Z(net_15331) );
CLKBUF_X2 inst_14318 ( .A(net_13793), .Z(net_14237) );
OAI22_X2 inst_1011 ( .A2(net_8247), .B2(net_8246), .ZN(net_8244), .A1(net_3038), .B1(net_1911) );
SDFF_X2 inst_540 ( .D(net_9124), .SE(net_933), .CK(net_10567), .SI(x2968), .Q(x1329) );
NAND2_X2 inst_4114 ( .ZN(net_2353), .A1(net_2352), .A2(net_1623) );
NOR4_X2 inst_2356 ( .A3(net_1993), .ZN(net_1451), .A4(net_1450), .A2(net_590), .A1(net_563) );
XNOR2_X2 inst_404 ( .A(net_9157), .B(net_9156), .ZN(net_1723) );
OAI22_X2 inst_998 ( .A1(net_8627), .B2(net_8626), .ZN(net_8597), .A2(net_8596), .B1(net_8595) );
INV_X4 inst_6044 ( .A(net_10141), .ZN(net_717) );
DFF_X2 inst_7989 ( .QN(net_10415), .D(net_5540), .CK(net_15660) );
NAND3_X2 inst_3209 ( .ZN(net_6781), .A1(net_6444), .A2(net_3836), .A3(net_3835) );
INV_X4 inst_5952 ( .ZN(net_2174), .A(net_836) );
INV_X4 inst_5838 ( .ZN(net_882), .A(net_656) );
NAND2_X2 inst_3615 ( .A2(net_10137), .ZN(net_7118), .A1(net_1204) );
AOI22_X2 inst_9628 ( .B1(net_9998), .A1(net_9768), .ZN(net_3415), .B2(net_2468), .A2(net_2462) );
CLKBUF_X2 inst_13989 ( .A(net_13907), .Z(net_13908) );
CLKBUF_X2 inst_14042 ( .A(net_12611), .Z(net_13961) );
CLKBUF_X2 inst_12298 ( .A(net_12216), .Z(net_12217) );
AOI222_X1 inst_9730 ( .ZN(net_3201), .B2(net_3200), .A2(net_3200), .C2(net_3199), .C1(net_2639), .A1(net_1589), .B1(net_727) );
NAND3_X2 inst_3216 ( .ZN(net_5689), .A1(net_5176), .A2(net_3422), .A3(net_3421) );
DFF_X1 inst_8748 ( .Q(net_9123), .D(net_5406), .CK(net_10608) );
CLKBUF_X2 inst_15093 ( .A(net_15011), .Z(net_15012) );
AOI221_X2 inst_9792 ( .B1(net_9970), .A(net_7090), .B2(net_7089), .C1(net_7088), .ZN(net_7020), .C2(net_242) );
CLKBUF_X2 inst_11442 ( .A(net_11360), .Z(net_11361) );
AOI21_X2 inst_10205 ( .ZN(net_2632), .A(net_2631), .B2(net_2630), .B1(net_1887) );
AOI22_X2 inst_9242 ( .A1(net_9946), .B1(net_9847), .A2(net_8042), .B2(net_8041), .ZN(net_6069) );
INV_X4 inst_5090 ( .ZN(net_2619), .A(net_1749) );
CLKBUF_X2 inst_14400 ( .A(net_14318), .Z(net_14319) );
XNOR2_X2 inst_192 ( .ZN(net_5203), .A(net_4564), .B(net_2382) );
INV_X2 inst_6720 ( .A(net_7876), .ZN(net_7833) );
CLKBUF_X2 inst_15489 ( .A(net_15407), .Z(net_15408) );
NOR2_X2 inst_2715 ( .ZN(net_4557), .A2(net_4111), .A1(net_1809) );
CLKBUF_X2 inst_13059 ( .A(net_11050), .Z(net_12978) );
NAND2_X2 inst_4242 ( .A2(net_5166), .ZN(net_4635), .A1(net_1476) );
NAND2_X2 inst_3540 ( .A2(net_9623), .A1(net_8975), .ZN(net_8006) );
CLKBUF_X2 inst_15277 ( .A(net_15195), .Z(net_15196) );
DFF_X2 inst_7701 ( .Q(net_9706), .D(net_6286), .CK(net_12588) );
NAND2_X2 inst_4126 ( .A1(net_2394), .ZN(net_2324), .A2(net_1606) );
DFF_X2 inst_7434 ( .QN(net_9388), .D(net_8328), .CK(net_14479) );
CLKBUF_X2 inst_14005 ( .A(net_13923), .Z(net_13924) );
CLKBUF_X2 inst_10904 ( .A(net_10596), .Z(net_10823) );
DFF_X1 inst_8741 ( .Q(net_9147), .D(net_5727), .CK(net_11035) );
NAND2_X2 inst_3547 ( .A2(net_9272), .ZN(net_8033), .A1(net_7875) );
NAND2_X2 inst_4178 ( .A2(net_4788), .ZN(net_3692), .A1(net_1269) );
CLKBUF_X2 inst_12720 ( .A(net_10597), .Z(net_12639) );
NOR3_X2 inst_2413 ( .ZN(net_5381), .A3(net_4669), .A1(net_3213), .A2(net_2429) );
OAI221_X2 inst_1574 ( .B2(net_7437), .ZN(net_7169), .C2(net_7167), .A(net_4724), .B1(net_3292), .C1(net_3207) );
INV_X4 inst_6558 ( .A(net_9177), .ZN(net_618) );
DFF_X2 inst_7528 ( .QN(net_9321), .D(net_7781), .CK(net_13063) );
AOI222_X1 inst_9739 ( .B2(net_10297), .C2(net_10295), .A2(net_10294), .B1(net_10284), .C1(net_10282), .A1(net_10281), .ZN(net_1136) );
CLKBUF_X2 inst_14518 ( .A(net_14436), .Z(net_14437) );
XNOR2_X2 inst_228 ( .ZN(net_4404), .B(net_4403), .A(net_3956) );
SDFF_X2 inst_486 ( .SE(net_9540), .SI(net_8223), .Q(net_303), .D(net_303), .CK(net_13910) );
INV_X2 inst_7234 ( .A(net_9398), .ZN(net_8208) );
CLKBUF_X2 inst_12977 ( .A(net_12895), .Z(net_12896) );
CLKBUF_X2 inst_15117 ( .A(net_15035), .Z(net_15036) );
CLKBUF_X2 inst_14034 ( .A(net_13952), .Z(net_13953) );
INV_X2 inst_6872 ( .ZN(net_3041), .A(net_3040) );
CLKBUF_X2 inst_13365 ( .A(net_13283), .Z(net_13284) );
CLKBUF_X2 inst_12008 ( .A(net_11014), .Z(net_11927) );
OAI22_X2 inst_1240 ( .A1(net_7243), .ZN(net_4872), .A2(net_4871), .B2(net_4870), .B1(net_1415) );
INV_X4 inst_5445 ( .ZN(net_1544), .A(net_1092) );
INV_X4 inst_6597 ( .A(net_9729), .ZN(net_707) );
CLKBUF_X2 inst_12279 ( .A(net_12197), .Z(net_12198) );
DFF_X1 inst_8759 ( .QN(net_9603), .D(net_5377), .CK(net_15174) );
XNOR2_X2 inst_244 ( .B(net_9621), .ZN(net_4162), .A(net_3654) );
CLKBUF_X2 inst_13514 ( .A(net_13432), .Z(net_13433) );
INV_X4 inst_5262 ( .ZN(net_1394), .A(net_1393) );
CLKBUF_X2 inst_11472 ( .A(net_11390), .Z(net_11391) );
CLKBUF_X2 inst_13464 ( .A(net_12093), .Z(net_13383) );
CLKBUF_X2 inst_12136 ( .A(net_12054), .Z(net_12055) );
CLKBUF_X2 inst_11794 ( .A(net_11712), .Z(net_11713) );
INV_X4 inst_5537 ( .ZN(net_6057), .A(net_945) );
AOI22_X2 inst_9186 ( .A1(net_9876), .B1(net_9777), .A2(net_8042), .B2(net_6129), .ZN(net_6128) );
OAI221_X2 inst_1521 ( .B1(net_10214), .ZN(net_7298), .C1(net_7297), .B2(net_7295), .C2(net_7293), .A(net_6687) );
CLKBUF_X2 inst_11339 ( .A(net_11257), .Z(net_11258) );
INV_X4 inst_6620 ( .ZN(net_8952), .A(net_8378) );
CLKBUF_X2 inst_13692 ( .A(net_13610), .Z(net_13611) );
AOI222_X1 inst_9679 ( .B1(net_9507), .ZN(net_8311), .A2(net_8310), .B2(net_8309), .C2(net_8308), .C1(net_8233), .A1(x2589) );
NAND4_X2 inst_3079 ( .ZN(net_4705), .A4(net_4279), .A1(net_3983), .A3(net_3495), .A2(net_3465) );
CLKBUF_X2 inst_12976 ( .A(net_12894), .Z(net_12895) );
CLKBUF_X2 inst_11208 ( .A(net_11126), .Z(net_11127) );
CLKBUF_X2 inst_10766 ( .A(net_10684), .Z(net_10685) );
NOR2_X2 inst_2563 ( .ZN(net_7790), .A1(net_7719), .A2(net_7701) );
OAI22_X2 inst_1306 ( .B1(net_3496), .A2(net_3062), .ZN(net_2413), .A1(net_2412), .B2(net_2076) );
INV_X4 inst_4845 ( .ZN(net_7449), .A(net_3313) );
AOI21_X2 inst_10143 ( .A(net_4671), .ZN(net_4234), .B2(net_3560), .B1(net_3159) );
CLKBUF_X2 inst_12529 ( .A(net_12447), .Z(net_12448) );
CLKBUF_X2 inst_15640 ( .A(net_15558), .Z(net_15559) );
AOI221_X2 inst_9931 ( .B2(net_5867), .A(net_5862), .ZN(net_5842), .C1(net_5841), .C2(net_4725), .B1(x5961) );
CLKBUF_X2 inst_12916 ( .A(net_12834), .Z(net_12835) );
OAI222_X2 inst_1407 ( .B2(net_7728), .A2(net_7727), .C2(net_7726), .ZN(net_5312), .B1(net_3228), .A1(net_2790), .C1(net_1073) );
INV_X4 inst_5487 ( .ZN(net_1986), .A(net_1363) );
DFF_X2 inst_8096 ( .QN(net_9732), .D(net_5049), .CK(net_12271) );
CLKBUF_X2 inst_13803 ( .A(net_11210), .Z(net_13722) );
CLKBUF_X2 inst_13128 ( .A(net_13046), .Z(net_13047) );
DFF_X2 inst_7599 ( .QN(net_10476), .D(net_7330), .CK(net_11401) );
INV_X2 inst_7018 ( .A(net_4009), .ZN(net_1542) );
CLKBUF_X2 inst_11789 ( .A(net_10949), .Z(net_11708) );
AOI22_X2 inst_9132 ( .A1(net_9716), .A2(net_6402), .ZN(net_6356), .B2(net_5263), .B1(net_4177) );
INV_X4 inst_6052 ( .A(net_10496), .ZN(net_508) );
AOI211_X2 inst_10303 ( .C2(net_10073), .C1(net_10064), .B(net_9858), .A(net_9759), .ZN(net_3477) );
CLKBUF_X2 inst_11526 ( .A(net_11444), .Z(net_11445) );
NAND2_X2 inst_3606 ( .ZN(net_7260), .A2(net_6856), .A1(net_6600) );
XNOR2_X2 inst_93 ( .ZN(net_8536), .A(net_8444), .B(net_5384) );
INV_X4 inst_4832 ( .ZN(net_5004), .A(net_3375) );
INV_X2 inst_7026 ( .A(net_8677), .ZN(net_1511) );
CLKBUF_X2 inst_14631 ( .A(net_14549), .Z(net_14550) );
INV_X2 inst_6965 ( .ZN(net_1833), .A(net_1832) );
CLKBUF_X2 inst_11051 ( .A(net_10969), .Z(net_10970) );
CLKBUF_X2 inst_12105 ( .A(net_11627), .Z(net_12024) );
AOI21_X2 inst_10217 ( .ZN(net_2303), .B1(net_2302), .B2(net_2301), .A(net_1950) );
AOI222_X1 inst_9687 ( .B1(net_9507), .A2(net_8301), .B2(net_8300), .C2(net_8299), .ZN(net_8297), .C1(net_8225), .A1(x2098) );
DFF_X2 inst_7784 ( .Q(net_9817), .D(net_6513), .CK(net_13418) );
INV_X4 inst_4595 ( .A(net_7861), .ZN(net_7826) );
INV_X4 inst_5099 ( .ZN(net_8760), .A(net_1191) );
CLKBUF_X2 inst_11116 ( .A(net_11034), .Z(net_11035) );
INV_X4 inst_6134 ( .A(net_9237), .ZN(net_2085) );
OAI221_X2 inst_1675 ( .B1(net_7226), .C2(net_5591), .ZN(net_5494), .C1(net_5493), .B2(net_4902), .A(net_3507) );
AOI22_X2 inst_9561 ( .A1(net_9937), .B1(net_9806), .A2(net_6443), .ZN(net_3758), .B2(net_2556) );
SDFF_X2 inst_584 ( .Q(net_9259), .SE(net_4589), .D(net_142), .SI(net_108), .CK(net_13841) );
CLKBUF_X2 inst_11086 ( .A(net_10967), .Z(net_11005) );
NAND2_X2 inst_3433 ( .A1(net_9481), .A2(net_8490), .ZN(net_8483) );
DFF_X1 inst_8668 ( .D(net_6769), .Q(net_115), .CK(net_15110) );
SDFF_X2 inst_470 ( .D(net_8576), .SE(net_758), .Q(net_235), .SI(net_104), .CK(net_11575) );
CLKBUF_X2 inst_15566 ( .A(net_15484), .Z(net_15485) );
CLKBUF_X2 inst_11274 ( .A(net_11192), .Z(net_11193) );
INV_X4 inst_5149 ( .ZN(net_1827), .A(net_1365) );
CLKBUF_X2 inst_12917 ( .A(net_12835), .Z(net_12836) );
CLKBUF_X2 inst_13713 ( .A(net_10602), .Z(net_13632) );
NAND2_X2 inst_4237 ( .A2(net_10331), .ZN(net_2705), .A1(net_810) );
CLKBUF_X2 inst_10709 ( .A(net_10612), .Z(net_10628) );
DFF_X2 inst_8138 ( .Q(net_9925), .D(net_5119), .CK(net_13387) );
XNOR2_X2 inst_148 ( .ZN(net_7022), .B(net_7021), .A(net_6176) );
INV_X8 inst_4490 ( .ZN(net_6889), .A(net_5936) );
SDFF_X2 inst_554 ( .SI(net_9361), .Q(net_9361), .D(net_9159), .SE(net_7248), .CK(net_15341) );
OAI21_X2 inst_1752 ( .ZN(net_8632), .B2(net_8590), .B1(net_8445), .A(net_8314) );
CLKBUF_X2 inst_13675 ( .A(net_13593), .Z(net_13594) );
CLKBUF_X2 inst_13621 ( .A(net_13539), .Z(net_13540) );
OAI22_X2 inst_1187 ( .A1(net_7294), .A2(net_5139), .B2(net_5138), .ZN(net_5068), .B1(net_1929) );
INV_X4 inst_6000 ( .A(net_9388), .ZN(net_2369) );
NAND2_X2 inst_4333 ( .A1(net_4172), .ZN(net_2347), .A2(net_1108) );
INV_X2 inst_6816 ( .A(net_9160), .ZN(net_5235) );
OAI22_X2 inst_1063 ( .A1(net_7535), .ZN(net_6966), .A2(net_6431), .B2(net_6430), .B1(net_507) );
INV_X4 inst_5499 ( .ZN(net_1157), .A(net_987) );
NOR2_X2 inst_2700 ( .ZN(net_4890), .A1(net_4391), .A2(net_4079) );
CLKBUF_X2 inst_10740 ( .A(net_10658), .Z(net_10659) );
OAI21_X2 inst_1917 ( .ZN(net_4570), .A(net_4144), .B2(net_4143), .B1(net_3984) );
CLKBUF_X2 inst_14764 ( .A(net_14682), .Z(net_14683) );
NAND3_X2 inst_3252 ( .ZN(net_4564), .A1(net_4563), .A3(net_4562), .A2(net_2415) );
CLKBUF_X2 inst_13542 ( .A(net_13460), .Z(net_13461) );
INV_X4 inst_4565 ( .ZN(net_8382), .A(net_8165) );
CLKBUF_X2 inst_15302 ( .A(net_15220), .Z(net_15221) );
CLKBUF_X2 inst_15753 ( .A(net_12323), .Z(net_15672) );
CLKBUF_X2 inst_12695 ( .A(net_12613), .Z(net_12614) );
INV_X4 inst_4755 ( .ZN(net_4902), .A(net_4228) );
INV_X4 inst_4955 ( .ZN(net_2552), .A(net_2551) );
CLKBUF_X2 inst_11553 ( .A(net_11471), .Z(net_11472) );
CLKBUF_X2 inst_12386 ( .A(net_12304), .Z(net_12305) );
INV_X4 inst_5276 ( .ZN(net_1338), .A(net_1337) );
AOI22_X2 inst_9452 ( .B1(net_9863), .A1(net_9697), .ZN(net_3990), .A2(net_3039), .B2(net_2973) );
OAI22_X2 inst_1167 ( .A1(net_7139), .A2(net_5107), .B2(net_5105), .ZN(net_5099), .B1(net_5098) );
OAI211_X2 inst_2087 ( .C2(net_6774), .ZN(net_6761), .A(net_6388), .B(net_6122), .C1(net_461) );
INV_X2 inst_6879 ( .ZN(net_4626), .A(net_2851) );
CLKBUF_X2 inst_14595 ( .A(net_14513), .Z(net_14514) );
DFF_X1 inst_8767 ( .QN(net_9381), .D(net_5408), .CK(net_13152) );
CLKBUF_X2 inst_13891 ( .A(net_13809), .Z(net_13810) );
CLKBUF_X2 inst_15671 ( .A(net_12459), .Z(net_15590) );
AOI221_X2 inst_9881 ( .B1(net_9788), .B2(net_9097), .A(net_6940), .C2(net_6939), .ZN(net_6818), .C1(net_258) );
OAI22_X2 inst_1303 ( .ZN(net_2907), .A1(net_2906), .A2(net_2905), .B2(net_2904), .B1(net_852) );
OAI221_X2 inst_1623 ( .C1(net_10320), .B1(net_7294), .C2(net_5591), .ZN(net_5584), .B2(net_4902), .A(net_3507) );
DFF_X1 inst_8571 ( .Q(net_9875), .D(net_7288), .CK(net_13376) );
CLKBUF_X2 inst_12788 ( .A(net_12706), .Z(net_12707) );
NAND2_X2 inst_4088 ( .A1(net_2677), .ZN(net_2549), .A2(net_2548) );
INV_X4 inst_6163 ( .A(net_9741), .ZN(net_477) );
INV_X4 inst_4922 ( .ZN(net_2701), .A(net_2700) );
INV_X4 inst_6501 ( .ZN(net_7139), .A(x5364) );
OR2_X4 inst_819 ( .ZN(net_5954), .A1(net_1002), .A2(net_186) );
MUX2_X1 inst_4464 ( .S(net_6041), .A(net_282), .B(x6028), .Z(x293) );
NAND2_X4 inst_3320 ( .A2(net_8989), .A1(net_8988), .ZN(net_8727) );
DFF_X2 inst_8369 ( .QN(net_9421), .D(net_2713), .CK(net_12715) );
OAI221_X2 inst_1468 ( .ZN(net_7880), .A(net_7876), .C2(net_7163), .B2(net_7023), .B1(net_5932), .C1(net_5275) );
AOI21_X2 inst_10183 ( .ZN(net_3961), .B2(net_3232), .A(net_2730), .B1(net_2455) );
AOI22_X2 inst_9663 ( .B2(net_10299), .A2(net_10298), .B1(net_10285), .A1(net_10284), .ZN(net_975) );
NAND2_X2 inst_3452 ( .A1(net_9463), .ZN(net_8910), .A2(net_8475) );
NAND2_X2 inst_3776 ( .ZN(net_5875), .A1(net_4784), .A2(net_4781) );
OAI221_X2 inst_1516 ( .B1(net_10419), .C2(net_9063), .B2(net_9056), .ZN(net_7320), .C1(net_7129), .A(net_7061) );
CLKBUF_X2 inst_14695 ( .A(net_10789), .Z(net_14614) );
CLKBUF_X2 inst_14046 ( .A(net_13964), .Z(net_13965) );
XNOR2_X2 inst_386 ( .ZN(net_2274), .B(net_1568), .A(net_1325) );
CLKBUF_X2 inst_15110 ( .A(net_15028), .Z(net_15029) );
CLKBUF_X2 inst_12372 ( .A(net_10966), .Z(net_12291) );
DFF_X1 inst_8497 ( .QN(net_10055), .D(net_7840), .CK(net_13744) );
DFF_X1 inst_8857 ( .Q(net_10522), .D(net_94), .CK(net_10859) );
INV_X4 inst_5859 ( .ZN(net_3194), .A(net_1233) );
INV_X2 inst_7255 ( .A(net_9390), .ZN(net_8224) );
NOR2_X2 inst_2617 ( .ZN(net_6207), .A2(net_5797), .A1(net_454) );
AND2_X2 inst_10543 ( .ZN(net_3852), .A2(net_3491), .A1(net_1283) );
AOI221_X2 inst_9863 ( .A(net_6889), .B2(net_6888), .C2(net_6887), .ZN(net_6853), .B1(net_1442), .C1(x4285) );
DFF_X2 inst_8089 ( .Q(net_10024), .D(net_5097), .CK(net_12979) );
NAND2_X2 inst_3942 ( .A1(net_9724), .ZN(net_3548), .A2(net_3039) );
DFF_X2 inst_7826 ( .Q(net_10012), .D(net_6474), .CK(net_14755) );
CLKBUF_X2 inst_11040 ( .A(net_10958), .Z(net_10959) );
AOI22_X2 inst_9459 ( .A1(net_6892), .B2(net_6625), .ZN(net_6287), .B1(net_3933), .A2(net_1753) );
NAND4_X2 inst_3068 ( .ZN(net_5680), .A4(net_4760), .A3(net_3790), .A2(net_3780), .A1(net_3411) );
INV_X4 inst_5225 ( .ZN(net_4929), .A(net_1503) );
INV_X4 inst_5850 ( .ZN(net_8756), .A(net_758) );
AOI21_X2 inst_10173 ( .ZN(net_3633), .A(net_3392), .B2(net_3085), .B1(net_3065) );
AOI221_X2 inst_9826 ( .B1(net_9770), .B2(net_9097), .A(net_6940), .C1(net_6939), .ZN(net_6923), .C2(net_240) );
NOR2_X2 inst_2778 ( .ZN(net_3367), .A2(net_3168), .A1(net_2223) );
OAI211_X2 inst_2277 ( .C1(net_7124), .C2(net_6542), .ZN(net_6223), .B(net_5751), .A(net_3679) );
INV_X4 inst_5320 ( .A(net_3429), .ZN(net_1276) );
AOI22_X2 inst_9518 ( .A1(net_10194), .B1(net_9897), .B2(net_4969), .A2(net_4217), .ZN(net_3804) );
CLKBUF_X2 inst_11883 ( .A(net_11801), .Z(net_11802) );
DFF_X2 inst_8245 ( .Q(net_10078), .D(net_4857), .CK(net_11216) );
INV_X4 inst_5223 ( .ZN(net_1919), .A(net_1506) );
INV_X4 inst_5468 ( .A(net_1727), .ZN(net_1719) );
AOI22_X2 inst_9599 ( .ZN(net_3493), .B2(net_3492), .A2(net_2762), .A1(net_2435), .B1(net_1018) );
NOR2_X2 inst_2962 ( .ZN(net_1812), .A1(net_1374), .A2(net_677) );
AOI21_X2 inst_10060 ( .ZN(net_7075), .B1(net_7072), .B2(net_7071), .A(net_3799) );
DFF_X1 inst_8716 ( .QN(net_8826), .D(net_6562), .CK(net_14125) );
CLKBUF_X2 inst_11064 ( .A(net_10780), .Z(net_10983) );
CLKBUF_X2 inst_12375 ( .A(net_12293), .Z(net_12294) );
OR2_X4 inst_811 ( .A2(net_10250), .A1(net_10249), .ZN(net_1662) );
CLKBUF_X2 inst_13973 ( .A(net_13040), .Z(net_13892) );
AND2_X2 inst_10605 ( .ZN(net_2038), .A1(net_2037), .A2(net_2036) );
AOI221_X2 inst_9973 ( .C2(net_10079), .B2(net_10078), .C1(net_10070), .B1(net_10069), .ZN(net_4577), .A(net_4129) );
XNOR2_X2 inst_208 ( .ZN(net_4938), .A(net_4401), .B(net_2391) );
CLKBUF_X2 inst_13756 ( .A(net_10592), .Z(net_13675) );
CLKBUF_X2 inst_14272 ( .A(net_14190), .Z(net_14191) );
CLKBUF_X2 inst_15247 ( .A(net_15165), .Z(net_15166) );
NAND2_X2 inst_4202 ( .ZN(net_2555), .A1(net_2169), .A2(net_1779) );
AOI22_X2 inst_9591 ( .B1(net_9975), .A2(net_5173), .ZN(net_3567), .B2(net_2541), .A1(net_209) );
NAND2_X2 inst_3774 ( .ZN(net_5877), .A2(net_4785), .A1(net_4784) );
INV_X2 inst_7101 ( .ZN(net_1058), .A(net_1057) );
NAND2_X2 inst_3909 ( .A2(net_9055), .ZN(net_7975), .A1(net_593) );
INV_X4 inst_5282 ( .ZN(net_1560), .A(net_1326) );
OAI21_X2 inst_1869 ( .ZN(net_5917), .A(net_5363), .B1(net_5362), .B2(net_5343) );
OR2_X2 inst_897 ( .A1(net_10503), .ZN(net_5769), .A2(net_5768) );
CLKBUF_X2 inst_12751 ( .A(net_12669), .Z(net_12670) );
CLKBUF_X2 inst_11935 ( .A(net_11853), .Z(net_11854) );
CLKBUF_X2 inst_15592 ( .A(net_15510), .Z(net_15511) );
AOI211_X2 inst_10294 ( .ZN(net_3749), .B(net_3748), .C2(net_3319), .C1(net_2966), .A(net_871) );
NAND2_X2 inst_3945 ( .ZN(net_3510), .A2(net_3509), .A1(net_3508) );
CLKBUF_X2 inst_11656 ( .A(net_11574), .Z(net_11575) );
OAI22_X2 inst_1201 ( .A1(net_7241), .A2(net_5151), .B2(net_5150), .ZN(net_5050), .B1(net_1860) );
DFF_X1 inst_8760 ( .Q(net_9129), .D(net_5305), .CK(net_10941) );
INV_X4 inst_5899 ( .ZN(net_4160), .A(net_601) );
AOI22_X2 inst_9294 ( .B1(net_9904), .A1(net_5759), .B2(net_5758), .ZN(net_5698), .A2(net_243) );
SDFF_X2 inst_636 ( .Q(net_9457), .D(net_9457), .SE(net_3293), .CK(net_11892), .SI(x2098) );
CLKBUF_X2 inst_15823 ( .A(net_11571), .Z(net_15742) );
OAI21_X2 inst_1927 ( .B1(net_10533), .ZN(net_4471), .B2(net_4470), .A(net_4468) );
XNOR2_X2 inst_184 ( .ZN(net_5211), .A(net_4585), .B(net_2389) );
OAI21_X2 inst_1847 ( .ZN(net_5931), .B1(net_5930), .A(net_5709), .B2(net_5360) );
CLKBUF_X2 inst_12499 ( .A(net_12417), .Z(net_12418) );
DFF_X1 inst_8878 ( .Q(net_9509), .D(net_9285), .CK(net_12144) );
CLKBUF_X2 inst_12270 ( .A(net_12188), .Z(net_12189) );
CLKBUF_X2 inst_11777 ( .A(net_11695), .Z(net_11696) );
OAI21_X2 inst_1907 ( .B2(net_10174), .ZN(net_4764), .B1(net_4007), .A(x3828) );
INV_X2 inst_6921 ( .ZN(net_2089), .A(net_2088) );
INV_X2 inst_7015 ( .ZN(net_2264), .A(net_1569) );
DFF_X1 inst_8775 ( .Q(net_10169), .D(net_4955), .CK(net_12301) );
DFF_X2 inst_8384 ( .QN(net_10538), .D(net_583), .CK(net_14577) );
AOI211_X2 inst_10313 ( .ZN(net_2436), .A(net_2435), .B(net_2434), .C2(net_925), .C1(net_665) );
NAND2_X2 inst_3836 ( .A1(net_6381), .ZN(net_4312), .A2(net_4311) );
INV_X2 inst_6999 ( .ZN(net_1628), .A(net_1627) );
CLKBUF_X2 inst_13461 ( .A(net_13379), .Z(net_13380) );
AOI22_X2 inst_9409 ( .A1(net_9951), .B1(net_6813), .ZN(net_4757), .A2(net_4742), .B2(net_4741) );
DFF_X1 inst_8472 ( .QN(net_9428), .D(net_7890), .CK(net_12677) );
DFF_X2 inst_7742 ( .QN(net_10147), .D(net_6326), .CK(net_13508) );
AOI22_X2 inst_9125 ( .A1(net_9710), .A2(net_6404), .ZN(net_6364), .B2(net_5263), .B1(net_150) );
CLKBUF_X2 inst_10919 ( .A(net_10629), .Z(net_10838) );
OAI211_X2 inst_2192 ( .C1(net_7221), .C2(net_6542), .ZN(net_6517), .B(net_5613), .A(net_3679) );
INV_X4 inst_5980 ( .A(net_9645), .ZN(net_2850) );
DFF_X2 inst_7806 ( .Q(net_9895), .D(net_6484), .CK(net_13198) );
OAI211_X2 inst_2114 ( .C2(net_6778), .ZN(net_6734), .A(net_6361), .B(net_6136), .C1(net_429) );
CLKBUF_X2 inst_14675 ( .A(net_14080), .Z(net_14594) );
NOR2_X2 inst_2784 ( .ZN(net_3417), .A1(net_3104), .A2(net_3103) );
CLKBUF_X2 inst_13817 ( .A(net_13735), .Z(net_13736) );
NAND2_X2 inst_4216 ( .A1(net_1988), .ZN(net_1969), .A2(net_1383) );
INV_X4 inst_6330 ( .ZN(net_7297), .A(x5225) );
XNOR2_X2 inst_106 ( .ZN(net_8144), .A(net_8051), .B(net_6900) );
CLKBUF_X2 inst_13001 ( .A(net_12919), .Z(net_12920) );
NOR2_X2 inst_2583 ( .ZN(net_7065), .A2(net_6637), .A1(net_3743) );
CLKBUF_X2 inst_10753 ( .A(net_10671), .Z(net_10672) );
AOI22_X2 inst_9036 ( .ZN(net_7430), .A2(net_6959), .B1(net_6958), .B2(net_4307), .A1(net_4301) );
AND2_X2 inst_10538 ( .A1(net_9620), .ZN(net_3654), .A2(net_3653) );
INV_X2 inst_7149 ( .A(net_4446), .ZN(net_768) );
NAND2_X2 inst_3997 ( .A2(net_8565), .ZN(net_3372), .A1(net_758) );
CLKBUF_X2 inst_13458 ( .A(net_12417), .Z(net_13377) );
CLKBUF_X2 inst_13697 ( .A(net_13615), .Z(net_13616) );
CLKBUF_X2 inst_11344 ( .A(net_10839), .Z(net_11263) );
NAND2_X2 inst_4377 ( .A2(net_9751), .A1(net_6321), .ZN(net_4007) );
INV_X4 inst_5241 ( .A(net_9735), .ZN(net_1747) );
AOI221_X2 inst_9903 ( .B1(net_9888), .B2(net_9101), .A(net_6945), .C2(net_6944), .C1(net_6816), .ZN(net_6791) );
NAND2_X2 inst_4383 ( .A2(net_10357), .ZN(net_2236), .A1(net_674) );
NAND2_X2 inst_4301 ( .ZN(net_1839), .A2(net_1381), .A1(net_717) );
CLKBUF_X2 inst_13432 ( .A(net_13350), .Z(net_13351) );
DFF_X1 inst_8537 ( .Q(net_9959), .D(net_7372), .CK(net_15478) );
CLKBUF_X2 inst_15018 ( .A(net_14936), .Z(net_14937) );
CLKBUF_X2 inst_14507 ( .A(net_14425), .Z(net_14426) );
AOI22_X2 inst_9208 ( .A1(net_9868), .B1(net_9769), .A2(net_8042), .B2(net_6120), .ZN(net_6103) );
OAI222_X2 inst_1410 ( .B2(net_7728), .A2(net_7727), .C2(net_7726), .ZN(net_5309), .B1(net_2981), .A1(net_2018), .C1(net_1319) );
INV_X4 inst_5106 ( .ZN(net_5433), .A(net_2913) );
CLKBUF_X2 inst_14943 ( .A(net_14861), .Z(net_14862) );
CLKBUF_X2 inst_10675 ( .A(net_10593), .Z(net_10594) );
INV_X4 inst_5434 ( .ZN(net_1578), .A(net_1120) );
AND2_X4 inst_10418 ( .ZN(net_4400), .A2(net_4261), .A1(net_4115) );
NAND2_X2 inst_3756 ( .A2(net_7846), .ZN(net_5413), .A1(net_5261) );
INV_X4 inst_4991 ( .ZN(net_6165), .A(net_2615) );
CLKBUF_X2 inst_14993 ( .A(net_12973), .Z(net_14912) );
NAND2_X1 inst_4424 ( .A2(net_4319), .A1(net_4041), .ZN(net_3880) );
CLKBUF_X2 inst_10811 ( .A(net_10656), .Z(net_10730) );
OAI21_X2 inst_1733 ( .ZN(net_8752), .B2(net_8729), .B1(net_8687), .A(net_1657) );
AOI22_X2 inst_9489 ( .B1(net_9884), .A2(net_5173), .ZN(net_3834), .B2(net_2973), .A1(net_217) );
DFF_X1 inst_8832 ( .Q(net_10542), .D(net_2857), .CK(net_13597) );
CLKBUF_X2 inst_11714 ( .A(net_11389), .Z(net_11633) );
INV_X2 inst_7028 ( .A(net_2612), .ZN(net_1489) );
NAND2_X2 inst_3900 ( .ZN(net_4236), .A2(net_3618), .A1(x6599) );
OAI211_X2 inst_2199 ( .C1(net_7192), .C2(net_6542), .ZN(net_6508), .B(net_5605), .A(net_3679) );
OR2_X2 inst_918 ( .A2(net_9760), .A1(net_9759), .ZN(net_3260) );
INV_X4 inst_4751 ( .ZN(net_4547), .A(net_4365) );
INV_X4 inst_5994 ( .A(net_10491), .ZN(net_535) );
INV_X4 inst_6588 ( .A(net_10370), .ZN(net_823) );
DFF_X2 inst_7678 ( .D(net_6754), .QN(net_129), .CK(net_11990) );
AOI21_X2 inst_10210 ( .ZN(net_2503), .A(net_2502), .B2(net_2276), .B1(net_1880) );
CLKBUF_X2 inst_13921 ( .A(net_13784), .Z(net_13840) );
INV_X2 inst_6653 ( .ZN(net_8570), .A(net_8569) );
AOI22_X2 inst_9177 ( .A1(net_9894), .B1(net_9795), .A2(net_8042), .B2(net_8041), .ZN(net_6139) );
OAI211_X2 inst_2074 ( .ZN(net_6775), .C2(net_6774), .A(net_6401), .B(net_6135), .C1(net_335) );
NAND2_X2 inst_4035 ( .ZN(net_4950), .A1(net_2950), .A2(net_2949) );
CLKBUF_X2 inst_11330 ( .A(net_11248), .Z(net_11249) );
OAI21_X2 inst_1862 ( .ZN(net_5424), .A(net_5260), .B2(net_4985), .B1(net_1350) );
INV_X4 inst_4823 ( .A(net_7157), .ZN(net_4413) );
INV_X2 inst_7296 ( .A(net_9052), .ZN(net_9051) );
XNOR2_X2 inst_221 ( .ZN(net_4574), .B(net_4573), .A(net_4415) );
OAI22_X2 inst_1236 ( .B1(net_7231), .A2(net_4890), .B2(net_4889), .ZN(net_4881), .A1(net_425) );
CLKBUF_X2 inst_14108 ( .A(net_14026), .Z(net_14027) );
CLKBUF_X2 inst_12928 ( .A(net_12846), .Z(net_12847) );
INV_X4 inst_5112 ( .ZN(net_1648), .A(net_1647) );
CLKBUF_X2 inst_12640 ( .A(net_12385), .Z(net_12559) );
NAND3_X2 inst_3313 ( .A3(net_9521), .ZN(net_1696), .A1(net_855), .A2(net_814) );
INV_X4 inst_5929 ( .ZN(net_1364), .A(net_1212) );
AOI22_X2 inst_9545 ( .B1(net_10021), .A1(net_9953), .A2(net_6443), .ZN(net_3776), .B2(net_2468) );
NAND2_X2 inst_3562 ( .A2(net_7748), .ZN(net_7688), .A1(net_2524) );
CLKBUF_X2 inst_13502 ( .A(net_11928), .Z(net_13421) );
DFF_X2 inst_7466 ( .QN(net_9521), .D(net_8080), .CK(net_14975) );
CLKBUF_X2 inst_11967 ( .A(net_11885), .Z(net_11886) );
NOR4_X2 inst_2334 ( .ZN(net_4483), .A4(net_4035), .A1(net_3628), .A3(net_3345), .A2(net_2853) );
NOR3_X2 inst_2429 ( .A2(net_9638), .A3(net_4460), .A1(net_4332), .ZN(net_4004) );
CLKBUF_X2 inst_15292 ( .A(net_12063), .Z(net_15211) );
OAI211_X2 inst_2210 ( .C1(net_7203), .C2(net_6501), .ZN(net_6495), .B(net_5565), .A(net_3527) );
AND2_X2 inst_10596 ( .A1(net_9617), .ZN(net_2831), .A2(net_2197) );
AND2_X4 inst_10463 ( .A1(net_10472), .ZN(net_1646), .A2(net_1096) );
OR2_X4 inst_754 ( .ZN(net_5150), .A1(net_4475), .A2(net_4472) );
INV_X4 inst_6040 ( .ZN(net_1392), .A(x6531) );
AND2_X2 inst_10531 ( .A2(net_3928), .ZN(net_3926), .A1(net_3454) );
AOI21_X2 inst_10030 ( .A(net_7916), .B2(net_7915), .ZN(net_7849), .B1(net_7848) );
INV_X4 inst_5028 ( .ZN(net_5518), .A(net_1937) );
NOR2_X2 inst_2590 ( .A2(net_7046), .ZN(net_7045), .A1(net_6227) );
AND4_X4 inst_10332 ( .ZN(net_3191), .A4(net_2022), .A1(net_1693), .A2(net_1410), .A3(net_1355) );
NOR2_X2 inst_2913 ( .A2(net_2824), .ZN(net_1496), .A1(net_1495) );
DFF_X2 inst_7647 ( .D(net_6719), .QN(net_164), .CK(net_14243) );
CLKBUF_X2 inst_11577 ( .A(net_11012), .Z(net_11496) );
CLKBUF_X2 inst_10949 ( .A(net_10621), .Z(net_10868) );
AND2_X4 inst_10435 ( .ZN(net_3025), .A2(net_2510), .A1(net_1295) );
DFF_X1 inst_8783 ( .Q(net_9539), .D(net_4605), .CK(net_12760) );
INV_X4 inst_5025 ( .ZN(net_1940), .A(net_1939) );
NAND3_X2 inst_3295 ( .A1(net_3630), .A3(net_2744), .ZN(net_2743), .A2(net_223) );
DFF_X1 inst_8792 ( .QN(net_10535), .D(net_4362), .CK(net_10575) );
CLKBUF_X2 inst_13341 ( .A(net_12460), .Z(net_13260) );
INV_X4 inst_5057 ( .A(net_3289), .ZN(net_3206) );
DFF_X1 inst_8828 ( .QN(net_9609), .D(net_3106), .CK(net_15390) );
DFF_X2 inst_7394 ( .D(net_8556), .QN(net_232), .CK(net_14331) );
CLKBUF_X2 inst_13997 ( .A(net_13631), .Z(net_13916) );
CLKBUF_X2 inst_13140 ( .A(net_12721), .Z(net_13059) );
CLKBUF_X2 inst_12451 ( .A(net_12369), .Z(net_12370) );
CLKBUF_X2 inst_15261 ( .A(net_15179), .Z(net_15180) );
CLKBUF_X2 inst_12998 ( .A(net_11247), .Z(net_12917) );
MUX2_X1 inst_4459 ( .S(net_6041), .A(net_287), .B(x5722), .Z(x244) );
NOR2_X2 inst_2923 ( .A2(net_10460), .A1(net_10459), .ZN(net_3490) );
CLKBUF_X2 inst_14028 ( .A(net_13201), .Z(net_13947) );
DFF_X2 inst_7957 ( .QN(net_10201), .D(net_5632), .CK(net_13253) );
NOR2_X2 inst_2707 ( .ZN(net_4270), .A2(net_4269), .A1(net_2425) );
OAI22_X2 inst_1117 ( .ZN(net_5992), .A2(net_4963), .B2(net_4962), .B1(net_3710), .A1(net_2576) );
NAND2_X2 inst_4015 ( .A1(net_9534), .ZN(net_5889), .A2(net_2553) );
HA_X1 inst_7343 ( .S(net_5241), .CO(net_5240), .B(net_4429), .A(net_565) );
CLKBUF_X2 inst_13909 ( .A(net_13827), .Z(net_13828) );
CLKBUF_X2 inst_11374 ( .A(net_10969), .Z(net_11293) );
NAND2_X2 inst_3958 ( .ZN(net_3472), .A2(net_3471), .A1(net_2037) );
INV_X2 inst_6887 ( .ZN(net_4068), .A(net_2764) );
NOR2_X2 inst_2725 ( .A2(net_10490), .ZN(net_4325), .A1(net_3298) );
CLKBUF_X2 inst_14476 ( .A(net_14394), .Z(net_14395) );
INV_X4 inst_5141 ( .A(net_10456), .ZN(net_3175) );
INV_X2 inst_6681 ( .ZN(net_8347), .A(net_8281) );
DFF_X2 inst_8204 ( .Q(net_10292), .D(net_4815), .CK(net_12972) );
XNOR2_X2 inst_334 ( .ZN(net_2980), .A(net_2377), .B(net_2148) );
OAI221_X2 inst_1610 ( .C1(net_10206), .B1(net_7124), .C2(net_5642), .ZN(net_5626), .B2(net_4905), .A(net_3507) );
AND2_X4 inst_10465 ( .A1(net_9586), .A2(net_8756), .ZN(net_1086) );
AOI21_X2 inst_10166 ( .B2(net_10512), .ZN(net_8373), .A(net_4371), .B1(net_3686) );
INV_X4 inst_4620 ( .ZN(net_7133), .A(net_7013) );
CLKBUF_X2 inst_12674 ( .A(net_11228), .Z(net_12593) );
CLKBUF_X2 inst_15719 ( .A(net_15637), .Z(net_15638) );
AOI22_X2 inst_9277 ( .B1(net_9800), .A1(net_5766), .B2(net_5765), .ZN(net_5749), .A2(net_238) );
NAND2_X2 inst_3707 ( .A1(net_9227), .ZN(net_7036), .A2(net_5888) );
CLKBUF_X2 inst_13337 ( .A(net_13255), .Z(net_13256) );
CLKBUF_X2 inst_11869 ( .A(net_11596), .Z(net_11788) );
CLKBUF_X2 inst_14243 ( .A(net_14091), .Z(net_14162) );
OAI22_X2 inst_1042 ( .A2(net_9068), .B1(net_8923), .A1(net_8921), .ZN(net_7920), .B2(net_2201) );
CLKBUF_X2 inst_14190 ( .A(net_12510), .Z(net_14109) );
CLKBUF_X2 inst_12431 ( .A(net_11051), .Z(net_12350) );
AOI21_X2 inst_10158 ( .B2(net_9053), .ZN(net_4043), .A(net_3180), .B1(net_663) );
INV_X4 inst_5961 ( .ZN(net_550), .A(net_223) );
DFF_X2 inst_8131 ( .QN(net_9843), .D(net_5126), .CK(net_14733) );
CLKBUF_X2 inst_14767 ( .A(net_14685), .Z(net_14686) );
INV_X4 inst_5388 ( .A(net_6414), .ZN(net_3532) );
INV_X4 inst_5595 ( .ZN(net_2882), .A(net_2272) );
INV_X8 inst_4492 ( .ZN(net_6945), .A(net_5934) );
CLKBUF_X2 inst_13551 ( .A(net_13469), .Z(net_13470) );
DFF_X2 inst_8153 ( .QN(net_9950), .D(net_5077), .CK(net_13706) );
AOI221_X2 inst_9773 ( .B2(net_10275), .ZN(net_7492), .C2(net_7405), .A(net_7073), .C1(net_6908), .B1(net_2202) );
CLKBUF_X2 inst_14553 ( .A(net_14471), .Z(net_14472) );
NAND4_X2 inst_3056 ( .ZN(net_5730), .A4(net_4773), .A3(net_4218), .A1(net_3856), .A2(net_3445) );
CLKBUF_X2 inst_14550 ( .A(net_14214), .Z(net_14469) );
CLKBUF_X2 inst_12214 ( .A(net_12132), .Z(net_12133) );
DFF_X2 inst_8058 ( .QN(net_10322), .D(net_5582), .CK(net_13232) );
CLKBUF_X2 inst_13255 ( .A(net_13173), .Z(net_13174) );
SDFF_X2 inst_595 ( .Q(net_9263), .SE(net_4589), .D(net_146), .SI(net_112), .CK(net_12547) );
NOR2_X2 inst_2609 ( .ZN(net_8994), .A2(net_5814), .A1(net_5414) );
NOR2_X2 inst_2556 ( .ZN(net_7820), .A2(net_7734), .A1(net_3721) );
INV_X4 inst_5002 ( .A(net_2605), .ZN(net_2187) );
CLKBUF_X2 inst_15022 ( .A(net_14940), .Z(net_14941) );
INV_X4 inst_5371 ( .ZN(net_1957), .A(net_1393) );
DFF_X2 inst_8222 ( .Q(net_10177), .D(net_4838), .CK(net_12966) );
OAI221_X2 inst_1704 ( .B2(net_7157), .ZN(net_4878), .B1(net_4877), .C1(net_4876), .A(net_4471), .C2(net_4084) );
INV_X4 inst_6343 ( .A(net_9550), .ZN(net_603) );
CLKBUF_X2 inst_13554 ( .A(net_12176), .Z(net_13473) );
AOI22_X2 inst_9014 ( .A2(net_8030), .B2(net_8029), .ZN(net_8022), .A1(net_217), .B1(net_194) );
INV_X4 inst_4604 ( .A(net_7782), .ZN(net_7747) );
CLKBUF_X2 inst_15156 ( .A(net_15074), .Z(net_15075) );
CLKBUF_X2 inst_15766 ( .A(net_15684), .Z(net_15685) );
XNOR2_X2 inst_161 ( .ZN(net_5977), .A(net_5976), .B(net_2057) );
INV_X4 inst_4688 ( .ZN(net_4839), .A(net_4657) );
CLKBUF_X2 inst_12658 ( .A(net_11073), .Z(net_12577) );
CLKBUF_X2 inst_10956 ( .A(net_10874), .Z(net_10875) );
CLKBUF_X2 inst_15451 ( .A(net_15369), .Z(net_15370) );
INV_X4 inst_4798 ( .A(net_3711), .ZN(net_3661) );
NAND2_X2 inst_3849 ( .ZN(net_4516), .A1(net_4237), .A2(net_4074) );
INV_X4 inst_6118 ( .A(net_9950), .ZN(net_6060) );
CLKBUF_X2 inst_15575 ( .A(net_14950), .Z(net_15494) );
CLKBUF_X2 inst_12205 ( .A(net_12123), .Z(net_12124) );
CLKBUF_X2 inst_11287 ( .A(net_10888), .Z(net_11206) );
OAI22_X2 inst_1029 ( .ZN(net_7908), .A2(net_7906), .B2(net_7904), .A1(net_6582), .B1(net_700) );
AOI22_X2 inst_9624 ( .A1(net_10076), .B1(net_9765), .A2(net_5319), .ZN(net_3427), .B2(net_2462) );
INV_X4 inst_5413 ( .A(net_6057), .ZN(net_1152) );
CLKBUF_X2 inst_11764 ( .A(net_11682), .Z(net_11683) );
AOI22_X2 inst_9246 ( .A1(net_9952), .B1(net_9853), .A2(net_8042), .B2(net_6133), .ZN(net_6065) );
INV_X2 inst_6666 ( .ZN(net_8362), .A(net_8305) );
INV_X2 inst_6841 ( .ZN(net_3868), .A(net_3601) );
NOR3_X2 inst_2408 ( .ZN(net_6806), .A2(net_6408), .A1(net_6198), .A3(net_5378) );
AND2_X2 inst_10519 ( .ZN(net_4686), .A2(net_4390), .A1(net_205) );
AOI221_X2 inst_9778 ( .ZN(net_7176), .B2(net_7175), .C2(net_7142), .A(net_3599), .C1(net_2606), .B1(net_1155) );
OAI22_X2 inst_1324 ( .A1(net_2780), .B2(net_2643), .B1(net_2302), .A2(net_1759), .ZN(net_1758) );
CLKBUF_X2 inst_15585 ( .A(net_14147), .Z(net_15504) );
INV_X4 inst_6245 ( .A(net_9513), .ZN(net_8107) );
INV_X2 inst_7032 ( .A(net_1759), .ZN(net_1443) );
INV_X4 inst_6551 ( .A(net_10102), .ZN(net_5829) );
CLKBUF_X2 inst_11848 ( .A(net_11191), .Z(net_11767) );
CLKBUF_X2 inst_10646 ( .A(net_10564), .Z(net_10565) );
XNOR2_X2 inst_342 ( .B(net_9361), .ZN(net_2867), .A(net_2285) );
CLKBUF_X2 inst_13048 ( .A(net_11184), .Z(net_12967) );
INV_X4 inst_5767 ( .A(net_1204), .ZN(net_995) );
AOI21_X2 inst_10067 ( .B1(net_10490), .ZN(net_6976), .A(net_6680), .B2(net_264) );
INV_X4 inst_6443 ( .ZN(net_7219), .A(x4520) );
CLKBUF_X2 inst_14404 ( .A(net_14322), .Z(net_14323) );
SDFF_X2 inst_463 ( .D(net_9579), .SI(net_5265), .SE(net_758), .Q(net_253), .CK(net_15052) );
OAI221_X2 inst_1534 ( .B1(net_10309), .B2(net_9047), .C2(net_7287), .C1(net_7241), .ZN(net_7236), .A(net_6785) );
CLKBUF_X2 inst_10667 ( .A(net_10585), .Z(net_10586) );
AOI221_X2 inst_9985 ( .C1(net_10178), .B2(net_6442), .C2(net_4217), .ZN(net_4212), .B1(net_4211), .A(net_3564) );
CLKBUF_X2 inst_13571 ( .A(net_12965), .Z(net_13490) );
NAND2_X2 inst_3820 ( .A1(net_10089), .A2(net_4534), .ZN(net_4518) );
INV_X4 inst_4667 ( .A(net_9265), .ZN(net_8403) );
AOI22_X2 inst_9108 ( .A1(net_9689), .A2(net_6420), .ZN(net_6384), .B2(net_5263), .B1(net_4309) );
XNOR2_X2 inst_319 ( .B(net_8760), .ZN(net_3193), .A(net_2726) );
NOR3_X2 inst_2422 ( .ZN(net_4349), .A3(net_4249), .A1(net_4036), .A2(net_821) );
CLKBUF_X2 inst_12762 ( .A(net_12680), .Z(net_12681) );
INV_X2 inst_6992 ( .A(net_4412), .ZN(net_1641) );
CLKBUF_X2 inst_12745 ( .A(net_12663), .Z(net_12664) );
CLKBUF_X2 inst_10688 ( .A(net_10572), .Z(net_10607) );
INV_X4 inst_5923 ( .ZN(net_883), .A(net_582) );
SDFF_X2 inst_649 ( .SI(net_9474), .Q(net_9474), .SE(net_3073), .CK(net_14143), .D(x3022) );
OAI211_X2 inst_2158 ( .C2(net_6778), .ZN(net_6690), .A(net_6303), .B(net_6045), .C1(net_5021) );
INV_X4 inst_5790 ( .ZN(net_998), .A(net_694) );
CLKBUF_X2 inst_15702 ( .A(net_14909), .Z(net_15621) );
CLKBUF_X2 inst_15166 ( .A(net_15084), .Z(net_15085) );
INV_X4 inst_5560 ( .A(net_10250), .ZN(net_1287) );
OAI221_X2 inst_1711 ( .B2(net_4274), .ZN(net_3943), .C2(net_3942), .A(net_3415), .C1(net_1590), .B1(net_1587) );
CLKBUF_X2 inst_10660 ( .A(net_10548), .Z(net_10579) );
DFF_X1 inst_8504 ( .Q(net_9426), .D(net_7716), .CK(net_13788) );
NAND2_X2 inst_3426 ( .A2(net_9478), .ZN(net_8885), .A1(net_8490) );
NOR2_X2 inst_2597 ( .A1(net_9289), .A2(net_7505), .ZN(net_6951) );
CLKBUF_X2 inst_14269 ( .A(net_14187), .Z(net_14188) );
CLKBUF_X2 inst_12227 ( .A(net_12145), .Z(net_12146) );
INV_X4 inst_5185 ( .ZN(net_4927), .A(net_1555) );
INV_X4 inst_5569 ( .A(net_9243), .ZN(net_3169) );
OAI211_X2 inst_2052 ( .ZN(net_7812), .C2(net_7811), .B(net_7448), .A(net_4295), .C1(net_4087) );
OAI22_X2 inst_995 ( .B1(net_9367), .ZN(net_8629), .A1(net_8627), .B2(net_8626), .A2(net_8586) );
OAI221_X2 inst_1575 ( .B2(net_7437), .ZN(net_7168), .C2(net_7167), .A(net_4721), .C1(net_3739), .B1(net_1508) );
INV_X4 inst_6059 ( .A(net_9346), .ZN(net_554) );
AOI22_X2 inst_9644 ( .ZN(net_2784), .A2(net_2783), .B2(net_2782), .B1(net_2780), .A1(net_1189) );
DFF_X1 inst_8850 ( .Q(net_10521), .D(net_93), .CK(net_10894) );
DFF_X2 inst_7726 ( .Q(net_9904), .D(net_6278), .CK(net_12566) );
CLKBUF_X2 inst_13948 ( .A(net_13866), .Z(net_13867) );
CLKBUF_X2 inst_10697 ( .A(net_10615), .Z(net_10616) );
NOR2_X4 inst_2470 ( .ZN(net_8882), .A1(net_8519), .A2(net_8518) );
INV_X4 inst_6049 ( .A(net_9968), .ZN(net_509) );
INV_X4 inst_5522 ( .ZN(net_3429), .A(net_1362) );
OAI22_X2 inst_1258 ( .B1(net_7201), .A2(net_4826), .B2(net_4825), .ZN(net_4815), .A1(net_323) );
AOI21_X2 inst_10148 ( .ZN(net_4199), .A(net_4198), .B1(net_3706), .B2(net_3705) );
NAND4_X2 inst_3141 ( .ZN(net_2687), .A2(net_2686), .A4(net_2434), .A3(net_1648), .A1(net_1454) );
NAND2_X2 inst_3921 ( .A2(net_9053), .ZN(net_7957), .A1(net_608) );
OAI21_X2 inst_1957 ( .ZN(net_4255), .A(net_3324), .B2(net_3242), .B1(net_3111) );
NAND2_X2 inst_3857 ( .A2(net_4187), .ZN(net_4178), .A1(net_4177) );
INV_X4 inst_5151 ( .ZN(net_5983), .A(net_908) );
CLKBUF_X2 inst_13860 ( .A(net_13447), .Z(net_13779) );
AOI22_X2 inst_9524 ( .B1(net_9702), .A2(net_6413), .A1(net_6053), .ZN(net_3797), .B2(net_3039) );
OAI22_X2 inst_1060 ( .ZN(net_7037), .A2(net_7036), .B2(net_7035), .B1(net_5718), .A1(net_4163) );
INV_X4 inst_5920 ( .ZN(net_2786), .A(net_585) );
DFF_X2 inst_7446 ( .QN(net_9291), .D(net_8236), .CK(net_11607) );
AND2_X4 inst_10456 ( .A1(net_10369), .ZN(net_1516), .A2(net_1365) );
OR2_X2 inst_900 ( .A1(net_10503), .ZN(net_5439), .A2(net_5425) );
INV_X2 inst_6950 ( .ZN(net_1893), .A(net_1892) );
AND2_X2 inst_10568 ( .A1(net_3272), .A2(net_3025), .ZN(net_3021) );
CLKBUF_X2 inst_14511 ( .A(net_14429), .Z(net_14430) );
INV_X4 inst_4949 ( .A(net_2587), .ZN(net_2562) );
CLKBUF_X2 inst_13813 ( .A(net_13731), .Z(net_13732) );
CLKBUF_X2 inst_12677 ( .A(net_12595), .Z(net_12596) );
INV_X4 inst_4624 ( .ZN(net_7086), .A(net_7085) );
NOR2_X2 inst_2807 ( .A2(net_8864), .ZN(net_5367), .A1(net_2753) );
CLKBUF_X2 inst_12458 ( .A(net_12376), .Z(net_12377) );
DFF_X2 inst_7811 ( .Q(net_10013), .D(net_6473), .CK(net_13332) );
CLKBUF_X2 inst_11257 ( .A(net_11175), .Z(net_11176) );
CLKBUF_X2 inst_13608 ( .A(net_13526), .Z(net_13527) );
AOI22_X2 inst_9254 ( .A2(net_8042), .B2(net_6133), .ZN(net_6052), .A1(net_2592), .B1(net_1596) );
INV_X4 inst_6062 ( .ZN(net_6821), .A(net_255) );
DFF_X2 inst_7428 ( .QN(net_9405), .D(net_8360), .CK(net_13943) );
NOR2_X2 inst_2983 ( .A1(net_10247), .ZN(net_2731), .A2(net_1015) );
INV_X4 inst_5327 ( .ZN(net_1528), .A(net_1269) );
INV_X4 inst_6608 ( .A(net_9946), .ZN(net_3944) );
DFF_X2 inst_7778 ( .Q(net_9810), .D(net_6523), .CK(net_12051) );
INV_X4 inst_5423 ( .A(net_3853), .ZN(net_1506) );
AOI221_X1 inst_9995 ( .ZN(net_7145), .A(net_6583), .C2(net_6153), .B2(net_5891), .B1(net_4499), .C1(net_4356) );
DFF_X1 inst_8803 ( .QN(net_10131), .D(net_3702), .CK(net_10773) );
DFF_X1 inst_8651 ( .Q(net_9779), .D(net_7183), .CK(net_15458) );
DFF_X2 inst_7421 ( .QN(net_9392), .D(net_8342), .CK(net_14020) );
CLKBUF_X2 inst_13584 ( .A(net_13502), .Z(net_13503) );
CLKBUF_X2 inst_13233 ( .A(net_13151), .Z(net_13152) );
AOI221_X2 inst_9969 ( .B1(net_10034), .C1(net_9804), .B2(net_5174), .ZN(net_4736), .A(net_4352), .C2(net_2556) );
DFF_X1 inst_8862 ( .Q(net_9511), .D(net_9287), .CK(net_12146) );
CLKBUF_X2 inst_12881 ( .A(net_12322), .Z(net_12800) );
AND2_X4 inst_10470 ( .A2(net_9244), .A1(net_9242), .ZN(net_3914) );
OAI22_X2 inst_1120 ( .B2(net_7525), .A1(net_5685), .ZN(net_5332), .B1(net_5331), .A2(net_4636) );
CLKBUF_X2 inst_12986 ( .A(net_11966), .Z(net_12905) );
INV_X4 inst_6238 ( .A(net_9302), .ZN(net_458) );
DFF_X1 inst_8545 ( .Q(net_9979), .D(net_7357), .CK(net_13740) );
DFF_X2 inst_7882 ( .QN(net_10105), .D(net_6036), .CK(net_14911) );
CLKBUF_X2 inst_15029 ( .A(net_13529), .Z(net_14948) );
CLKBUF_X2 inst_11617 ( .A(net_11535), .Z(net_11536) );
CLKBUF_X2 inst_12161 ( .A(net_12079), .Z(net_12080) );
NAND3_X2 inst_3184 ( .A1(net_8949), .ZN(net_8087), .A3(net_7993), .A2(net_7572) );
INV_X2 inst_6767 ( .ZN(net_6036), .A(net_5865) );
AOI222_X1 inst_9715 ( .ZN(net_7582), .A2(net_7489), .C2(net_6981), .A1(net_6950), .B2(net_6203), .C1(net_3698), .B1(net_657) );
INV_X4 inst_6398 ( .A(net_10543), .ZN(net_3464) );
DFF_X2 inst_8084 ( .QN(net_9165), .D(net_5102), .CK(net_13557) );
CLKBUF_X2 inst_15381 ( .A(net_12158), .Z(net_15300) );
OR2_X4 inst_731 ( .ZN(net_7506), .A1(net_7115), .A2(net_7114) );
OAI33_X1 inst_947 ( .ZN(net_7650), .A3(net_7649), .B1(net_7648), .A1(net_7516), .B2(net_5331), .B3(net_4611), .A2(net_1314) );
OAI22_X2 inst_1225 ( .A1(net_7108), .A2(net_5107), .B2(net_5105), .ZN(net_5022), .B1(net_5021) );
CLKBUF_X2 inst_10909 ( .A(net_10574), .Z(net_10828) );
CLKBUF_X2 inst_13788 ( .A(net_13168), .Z(net_13707) );
CLKBUF_X2 inst_15005 ( .A(net_14923), .Z(net_14924) );
DFF_X2 inst_7535 ( .QN(net_9316), .D(net_7775), .CK(net_15321) );
CLKBUF_X2 inst_12411 ( .A(net_11966), .Z(net_12330) );
NOR3_X2 inst_2459 ( .A2(net_9184), .A1(net_9182), .A3(net_9181), .ZN(net_894) );
CLKBUF_X2 inst_14256 ( .A(net_14174), .Z(net_14175) );
XNOR2_X2 inst_363 ( .B(net_9154), .ZN(net_2558), .A(net_2476) );
XNOR2_X2 inst_301 ( .ZN(net_3296), .A(net_2201), .B(net_1584) );
INV_X4 inst_5316 ( .ZN(net_1587), .A(net_1281) );
INV_X2 inst_7165 ( .A(net_7025), .ZN(net_567) );
OAI211_X2 inst_2141 ( .C2(net_6778), .ZN(net_6707), .A(net_6334), .B(net_6070), .C1(net_5873) );
INV_X4 inst_5530 ( .ZN(net_1199), .A(net_949) );
CLKBUF_X2 inst_14427 ( .A(net_14345), .Z(net_14346) );
CLKBUF_X2 inst_14215 ( .A(net_14133), .Z(net_14134) );
CLKBUF_X2 inst_12041 ( .A(net_11959), .Z(net_11960) );
INV_X4 inst_4551 ( .ZN(net_8569), .A(net_8557) );
CLKBUF_X2 inst_11397 ( .A(net_11290), .Z(net_11316) );
NAND2_X2 inst_4313 ( .ZN(net_2677), .A2(net_1190), .A1(net_712) );
INV_X4 inst_6609 ( .A(net_10252), .ZN(net_1016) );
CLKBUF_X2 inst_13213 ( .A(net_10805), .Z(net_13132) );
INV_X2 inst_7079 ( .A(net_2626), .ZN(net_1192) );
CLKBUF_X2 inst_13153 ( .A(net_13071), .Z(net_13072) );
INV_X4 inst_4714 ( .ZN(net_5323), .A(net_4711) );
DFF_X2 inst_7870 ( .QN(net_10251), .D(net_6038), .CK(net_13921) );
CLKBUF_X2 inst_14021 ( .A(net_13939), .Z(net_13940) );
CLKBUF_X2 inst_12898 ( .A(net_12816), .Z(net_12817) );
NAND2_X2 inst_4348 ( .A2(net_10457), .ZN(net_2036), .A1(net_842) );
INV_X4 inst_4706 ( .A(net_6679), .ZN(net_5348) );
NOR2_X2 inst_2956 ( .A1(net_10456), .ZN(net_1549), .A2(net_1209) );
INV_X4 inst_4713 ( .ZN(net_5853), .A(net_4547) );
CLKBUF_X2 inst_14312 ( .A(net_14230), .Z(net_14231) );
NAND2_X2 inst_3729 ( .A1(net_10405), .ZN(net_5696), .A2(net_5409) );
DFF_X1 inst_8521 ( .QN(net_10301), .D(net_7413), .CK(net_10707) );
XNOR2_X2 inst_412 ( .A(net_9202), .B(net_9201), .ZN(net_1463) );
AND2_X4 inst_10430 ( .A1(net_4088), .ZN(net_3303), .A2(net_3302) );
DFF_X2 inst_7548 ( .QN(net_9248), .D(net_7705), .CK(net_11271) );
AOI22_X2 inst_9282 ( .B1(net_9998), .A1(net_5743), .B2(net_5742), .ZN(net_5736), .A2(net_238) );
DFF_X2 inst_8345 ( .Q(net_9612), .D(net_2788), .CK(net_14057) );
CLKBUF_X2 inst_14559 ( .A(net_14477), .Z(net_14478) );
CLKBUF_X2 inst_11687 ( .A(net_11605), .Z(net_11606) );
NOR2_X2 inst_2650 ( .A1(net_9218), .ZN(net_5888), .A2(net_5361) );
INV_X4 inst_5463 ( .A(net_10142), .ZN(net_2007) );
INV_X8 inst_4508 ( .ZN(net_6418), .A(net_5295) );
CLKBUF_X2 inst_14721 ( .A(net_12476), .Z(net_14640) );
DFF_X2 inst_7943 ( .QN(net_10421), .D(net_5548), .CK(net_15496) );
CLKBUF_X2 inst_13022 ( .A(net_11539), .Z(net_12941) );
CLKBUF_X2 inst_11626 ( .A(net_11544), .Z(net_11545) );
AOI22_X2 inst_9490 ( .B1(net_9917), .A1(net_9719), .B2(net_4969), .ZN(net_3833), .A2(net_3039) );
CLKBUF_X2 inst_11666 ( .A(net_11584), .Z(net_11585) );
DFF_X2 inst_8295 ( .Q(net_9853), .D(net_4613), .CK(net_12328) );
CLKBUF_X2 inst_13969 ( .A(net_12544), .Z(net_13888) );
NAND3_X2 inst_3189 ( .ZN(net_7717), .A1(net_7591), .A3(net_7576), .A2(net_7425) );
NAND4_X2 inst_3163 ( .A3(net_9194), .A4(net_2928), .ZN(net_2099), .A1(net_1246), .A2(net_519) );
NOR2_X2 inst_2504 ( .ZN(net_8530), .A2(net_8406), .A1(net_8401) );
CLKBUF_X2 inst_13511 ( .A(net_13429), .Z(net_13430) );
CLKBUF_X2 inst_12818 ( .A(net_12736), .Z(net_12737) );
INV_X4 inst_5548 ( .ZN(net_1215), .A(net_935) );
INV_X4 inst_5985 ( .A(net_9180), .ZN(net_2785) );
INV_X2 inst_6855 ( .A(net_7434), .ZN(net_3369) );
CLKBUF_X2 inst_14076 ( .A(net_13994), .Z(net_13995) );
CLKBUF_X2 inst_14188 ( .A(net_14106), .Z(net_14107) );
CLKBUF_X2 inst_14824 ( .A(net_14742), .Z(net_14743) );
CLKBUF_X2 inst_10902 ( .A(net_10820), .Z(net_10821) );
CLKBUF_X2 inst_15469 ( .A(net_15387), .Z(net_15388) );
OR4_X2 inst_684 ( .A4(net_9584), .A3(net_9582), .A1(net_9574), .ZN(net_8777), .A2(net_8776) );
INV_X4 inst_6263 ( .A(net_10464), .ZN(net_665) );
NAND2_X4 inst_3374 ( .A2(net_9046), .A1(net_8998), .ZN(net_3179) );
NAND2_X2 inst_4354 ( .A2(net_10460), .ZN(net_2399), .A1(net_921) );
NAND2_X2 inst_4400 ( .A2(net_10405), .A1(net_10397), .ZN(net_662) );
NAND2_X2 inst_3438 ( .A1(net_9476), .A2(net_8487), .ZN(net_8481) );
NAND3_X2 inst_3177 ( .ZN(net_8183), .A1(net_8054), .A3(net_7961), .A2(net_3381) );
CLKBUF_X2 inst_12187 ( .A(net_11353), .Z(net_12106) );
CLKBUF_X2 inst_12541 ( .A(net_11473), .Z(net_12460) );
AND2_X4 inst_10437 ( .ZN(net_2376), .A2(net_2375), .A1(net_1685) );
INV_X4 inst_4930 ( .ZN(net_4355), .A(net_2669) );
CLKBUF_X2 inst_14614 ( .A(net_12594), .Z(net_14533) );
DFF_X2 inst_7965 ( .QN(net_10315), .D(net_5592), .CK(net_15586) );
NAND2_X2 inst_3811 ( .A1(net_10080), .A2(net_4534), .ZN(net_4527) );
CLKBUF_X2 inst_11857 ( .A(net_11775), .Z(net_11776) );
NAND2_X2 inst_3653 ( .A2(net_6660), .ZN(net_6659), .A1(net_2513) );
INV_X2 inst_6959 ( .A(net_4927), .ZN(net_1873) );
CLKBUF_X2 inst_15652 ( .A(net_15570), .Z(net_15571) );
DFF_X2 inst_8213 ( .Q(net_10087), .D(net_4848), .CK(net_10750) );
CLKBUF_X2 inst_10700 ( .A(net_10590), .Z(net_10619) );
OAI22_X2 inst_1138 ( .A1(net_7211), .A2(net_5151), .B2(net_5150), .ZN(net_5137), .B1(net_358) );
CLKBUF_X2 inst_15438 ( .A(net_15356), .Z(net_15357) );
OAI22_X2 inst_1241 ( .A1(net_7192), .A2(net_4871), .B2(net_4870), .ZN(net_4869), .B1(net_505) );
OAI22_X2 inst_1038 ( .A1(net_9087), .A2(net_8922), .B1(net_8919), .ZN(net_7948), .B2(net_2225) );
CLKBUF_X2 inst_15418 ( .A(net_15336), .Z(net_15337) );
INV_X4 inst_6568 ( .A(net_9924), .ZN(net_327) );
OR2_X2 inst_940 ( .A2(net_2344), .ZN(net_1810), .A1(net_1809) );
OAI22_X2 inst_1004 ( .ZN(net_8414), .A1(net_8327), .B2(net_8325), .A2(net_8204), .B1(net_5805) );
AOI22_X2 inst_9417 ( .A1(net_10179), .A2(net_4656), .B2(net_4655), .ZN(net_4652), .B1(x4209) );
CLKBUF_X2 inst_11705 ( .A(net_11623), .Z(net_11624) );
CLKBUF_X2 inst_11641 ( .A(net_10912), .Z(net_11560) );
NAND2_X2 inst_3595 ( .ZN(net_7271), .A2(net_6891), .A1(net_6610) );
CLKBUF_X2 inst_11830 ( .A(net_11748), .Z(net_11749) );
AOI22_X2 inst_9316 ( .B1(net_9721), .A2(net_5755), .B2(net_5754), .ZN(net_5661), .A1(net_258) );
XNOR2_X2 inst_189 ( .ZN(net_5206), .A(net_4578), .B(net_1764) );
INV_X4 inst_4876 ( .ZN(net_3287), .A(net_3044) );
DFF_X2 inst_8103 ( .Q(net_9174), .D(net_5071), .CK(net_11247) );
DFF_X2 inst_7732 ( .Q(net_9799), .D(net_6223), .CK(net_11986) );
AOI22_X2 inst_9008 ( .B1(net_9303), .A2(net_8030), .B2(net_8029), .ZN(net_8028), .A1(net_211) );
NOR3_X2 inst_2450 ( .A3(net_9222), .ZN(net_2492), .A1(net_1766), .A2(net_1538) );
CLKBUF_X2 inst_13248 ( .A(net_13166), .Z(net_13167) );
DFF_X1 inst_8597 ( .Q(net_9686), .D(net_7260), .CK(net_15253) );
NAND2_X2 inst_4362 ( .ZN(net_930), .A1(net_929), .A2(net_928) );
DFF_X2 inst_7437 ( .QN(net_9408), .D(net_8357), .CK(net_13925) );
AOI22_X2 inst_9581 ( .A1(net_10064), .A2(net_5320), .B2(net_5174), .ZN(net_3582), .B1(net_2284) );
DFF_X2 inst_7430 ( .QN(net_9410), .D(net_8352), .CK(net_13936) );
CLKBUF_X2 inst_15761 ( .A(net_15679), .Z(net_15680) );
CLKBUF_X2 inst_11006 ( .A(net_10924), .Z(net_10925) );
AOI22_X2 inst_9529 ( .B1(net_10504), .A1(net_9662), .B2(net_6415), .A2(net_5966), .ZN(net_3792) );
XNOR2_X2 inst_62 ( .ZN(net_8732), .A(net_8720), .B(net_8096) );
CLKBUF_X2 inst_12608 ( .A(net_11584), .Z(net_12527) );
NAND2_X2 inst_4369 ( .A2(net_10120), .ZN(net_899), .A1(net_898) );
INV_X4 inst_4696 ( .ZN(net_4831), .A(net_4647) );
NAND2_X2 inst_3743 ( .ZN(net_5597), .A2(net_5323), .A1(net_3204) );
NOR2_X2 inst_2860 ( .A1(net_3490), .A2(net_2686), .ZN(net_2070) );
CLKBUF_X2 inst_11899 ( .A(net_11323), .Z(net_11818) );
INV_X4 inst_5194 ( .ZN(net_1981), .A(net_1850) );
CLKBUF_X2 inst_11236 ( .A(net_10590), .Z(net_11155) );
CLKBUF_X2 inst_14496 ( .A(net_14414), .Z(net_14415) );
CLKBUF_X2 inst_13076 ( .A(net_12994), .Z(net_12995) );
DFF_X2 inst_8387 ( .Q(net_10513), .D(net_866), .CK(net_13110) );
NAND2_X2 inst_4007 ( .A1(net_4481), .ZN(net_4480), .A2(net_3191) );
OR2_X2 inst_879 ( .A2(net_7038), .ZN(net_6434), .A1(net_6433) );
CLKBUF_X2 inst_11266 ( .A(net_11184), .Z(net_11185) );
INV_X4 inst_5888 ( .ZN(net_5684), .A(net_613) );
CLKBUF_X2 inst_13956 ( .A(net_13874), .Z(net_13875) );
CLKBUF_X2 inst_11162 ( .A(net_11080), .Z(net_11081) );
CLKBUF_X2 inst_12416 ( .A(net_12334), .Z(net_12335) );
DFF_X2 inst_8252 ( .Q(net_10182), .D(net_4840), .CK(net_12954) );
HA_X1 inst_7344 ( .S(net_5239), .CO(net_5238), .B(net_4425), .A(net_569) );
CLKBUF_X2 inst_15462 ( .A(net_12331), .Z(net_15381) );
INV_X8 inst_4482 ( .ZN(net_8490), .A(net_8420) );
NAND2_X2 inst_4291 ( .A2(net_10156), .A1(net_3496), .ZN(net_2682) );
INV_X4 inst_5692 ( .A(net_932), .ZN(net_790) );
SDFF_X2 inst_629 ( .Q(net_9447), .D(net_9447), .SE(net_3293), .CK(net_14160), .SI(x2707) );
INV_X4 inst_4903 ( .A(net_7095), .ZN(net_3044) );
OAI22_X2 inst_1100 ( .A1(net_9192), .A2(net_6299), .B2(net_6298), .ZN(net_6250), .B1(net_660) );
DFF_X2 inst_7903 ( .QN(net_10142), .D(net_6031), .CK(net_12368) );
CLKBUF_X2 inst_10872 ( .A(net_10790), .Z(net_10791) );
CLKBUF_X2 inst_15105 ( .A(net_10826), .Z(net_15024) );
OR2_X4 inst_791 ( .A1(net_10260), .ZN(net_2250), .A2(net_1957) );
CLKBUF_X2 inst_13371 ( .A(net_13289), .Z(net_13290) );
AND2_X4 inst_10427 ( .ZN(net_7589), .A2(net_3514), .A1(net_3512) );
OAI21_X2 inst_2021 ( .ZN(net_8862), .A(net_2417), .B2(net_2064), .B1(net_1674) );
AOI22_X2 inst_9631 ( .A1(net_9837), .B1(net_9773), .A2(net_6413), .ZN(net_3412), .B2(net_2462) );
NAND2_X2 inst_3383 ( .ZN(net_8775), .A2(net_8758), .A1(net_1654) );
NAND2_X2 inst_4379 ( .A2(net_10434), .A1(net_3104), .ZN(net_2404) );
CLKBUF_X2 inst_15682 ( .A(net_15600), .Z(net_15601) );
OAI22_X2 inst_1191 ( .A1(net_7127), .A2(net_5139), .B2(net_5138), .ZN(net_5063), .B1(net_1152) );
INV_X4 inst_5668 ( .ZN(net_3034), .A(net_814) );
CLKBUF_X2 inst_13326 ( .A(net_13244), .Z(net_13245) );
SDFF_X2 inst_533 ( .D(net_9121), .SE(net_933), .CK(net_10571), .SI(x3133), .Q(x1370) );
INV_X4 inst_5086 ( .ZN(net_1788), .A(net_1787) );
CLKBUF_X2 inst_15107 ( .A(net_14050), .Z(net_15026) );
CLKBUF_X2 inst_12811 ( .A(net_12604), .Z(net_12730) );
NOR2_X4 inst_2478 ( .A2(net_9523), .ZN(net_4268), .A1(net_3727) );
INV_X4 inst_4972 ( .A(net_5376), .ZN(net_3317) );
CLKBUF_X2 inst_14670 ( .A(net_14588), .Z(net_14589) );
NOR2_X2 inst_2751 ( .ZN(net_3981), .A2(net_3652), .A1(net_271) );
CLKBUF_X2 inst_14399 ( .A(net_14317), .Z(net_14318) );
DFF_X1 inst_8576 ( .Q(net_9870), .D(net_7128), .CK(net_15629) );
CLKBUF_X2 inst_13020 ( .A(net_12938), .Z(net_12939) );
CLKBUF_X2 inst_11924 ( .A(net_11842), .Z(net_11843) );
OAI21_X2 inst_1760 ( .ZN(net_8452), .A(net_8376), .B2(net_8375), .B1(net_7157) );
OAI21_X2 inst_1874 ( .ZN(net_5287), .A(net_5286), .B2(net_4363), .B1(x4587) );
CLKBUF_X2 inst_11888 ( .A(net_11806), .Z(net_11807) );
OAI21_X2 inst_2022 ( .ZN(net_8868), .A(net_2189), .B2(net_2078), .B1(net_1530) );
NAND2_X2 inst_3960 ( .ZN(net_3617), .A1(net_3456), .A2(net_3455) );
NOR2_X2 inst_2821 ( .A1(net_3908), .A2(net_3065), .ZN(net_2594) );
OAI22_X2 inst_1095 ( .A1(net_9186), .ZN(net_6300), .A2(net_6299), .B2(net_6298), .B1(net_2090) );
DFF_X2 inst_8042 ( .QN(net_9550), .D(net_9256), .CK(net_13764) );
AND2_X2 inst_10516 ( .ZN(net_4920), .A1(net_4603), .A2(net_4451) );
AOI21_X2 inst_10096 ( .B2(net_10385), .A(net_6677), .ZN(net_5409), .B1(net_627) );
AOI22_X2 inst_9052 ( .B1(net_9673), .A1(net_6684), .B2(net_6683), .ZN(net_6643), .A2(net_242) );
NOR3_X2 inst_2439 ( .ZN(net_3051), .A1(net_3050), .A3(net_3049), .A2(net_664) );
XNOR2_X2 inst_176 ( .ZN(net_5398), .A(net_4952), .B(net_2024) );
NOR2_X2 inst_2826 ( .ZN(net_3011), .A1(net_2505), .A2(net_2504) );
DFF_X2 inst_7848 ( .Q(net_9909), .D(net_6499), .CK(net_12038) );
INV_X4 inst_6143 ( .ZN(net_3885), .A(net_154) );
DFF_X2 inst_8142 ( .QN(net_9942), .D(net_5115), .CK(net_11443) );
INV_X2 inst_7304 ( .A(net_9073), .ZN(net_9072) );
AOI22_X2 inst_9069 ( .B1(net_9689), .A2(net_6684), .B2(net_6683), .ZN(net_6597), .A1(net_258) );
CLKBUF_X2 inst_10894 ( .A(net_10812), .Z(net_10813) );
CLKBUF_X2 inst_12864 ( .A(net_12782), .Z(net_12783) );
OAI222_X2 inst_1336 ( .A1(net_7732), .B2(net_7731), .C2(net_7730), .ZN(net_7662), .A2(net_7550), .B1(net_7026), .C1(net_567) );
INV_X4 inst_5472 ( .ZN(net_3699), .A(net_1010) );
AND2_X4 inst_10387 ( .A1(net_8961), .A2(net_8497), .ZN(net_8337) );
NAND2_X2 inst_4404 ( .A2(net_10510), .A1(net_10496), .ZN(net_630) );
OAI221_X2 inst_1665 ( .C1(net_7229), .C2(net_5520), .ZN(net_5504), .B2(net_4547), .A(net_3507), .B1(net_1838) );
INV_X8 inst_4500 ( .ZN(net_6129), .A(net_5298) );
CLKBUF_X2 inst_13962 ( .A(net_12544), .Z(net_13881) );
INV_X4 inst_4763 ( .ZN(net_4476), .A(net_4367) );
OR2_X4 inst_780 ( .ZN(net_4661), .A1(net_2956), .A2(net_2555) );
INV_X4 inst_5626 ( .ZN(net_3529), .A(net_2565) );
AOI22_X2 inst_9054 ( .B1(net_9670), .A1(net_6684), .B2(net_6683), .ZN(net_6641), .A2(net_239) );
INV_X4 inst_6581 ( .A(net_9179), .ZN(net_1729) );
DFF_X2 inst_8154 ( .QN(net_10049), .D(net_5074), .CK(net_14720) );
INV_X2 inst_6783 ( .ZN(net_6588), .A(net_5784) );
DFF_X2 inst_8255 ( .Q(net_10186), .D(net_4831), .CK(net_12853) );
CLKBUF_X2 inst_11261 ( .A(net_11179), .Z(net_11180) );
CLKBUF_X2 inst_15046 ( .A(net_14964), .Z(net_14965) );
CLKBUF_X2 inst_12016 ( .A(net_11687), .Z(net_11935) );
INV_X2 inst_6716 ( .ZN(net_7940), .A(net_7914) );
NAND2_X2 inst_3967 ( .ZN(net_3381), .A1(net_3380), .A2(net_3378) );
INV_X4 inst_5541 ( .A(net_10355), .ZN(net_1220) );
DFF_X1 inst_8722 ( .QN(net_10276), .D(net_6266), .CK(net_13960) );
NAND2_X2 inst_4018 ( .A2(net_7095), .A1(net_6949), .ZN(net_3512) );
NAND2_X2 inst_3669 ( .A1(net_8958), .A2(net_7378), .ZN(net_6905) );
OAI21_X2 inst_1767 ( .ZN(net_8085), .B2(net_8036), .A(net_8011), .B1(net_5807) );
INV_X4 inst_5636 ( .ZN(net_2761), .A(net_1074) );
OAI211_X2 inst_2219 ( .C1(net_7192), .C2(net_6501), .ZN(net_6486), .B(net_5561), .A(net_3679) );
DFF_X1 inst_8884 ( .D(net_10517), .CK(net_12650), .Q(x461) );
DFF_X2 inst_8331 ( .QN(net_10270), .D(net_3220), .CK(net_14432) );
SDFF_X2 inst_546 ( .D(net_9142), .SE(net_933), .CK(net_10657), .SI(x1865), .Q(x1161) );
OAI22_X2 inst_1284 ( .A1(net_4508), .A2(net_4092), .ZN(net_4090), .B1(net_2693), .B2(net_2248) );
CLKBUF_X2 inst_13564 ( .A(net_13482), .Z(net_13483) );
NOR2_X4 inst_2465 ( .ZN(net_9032), .A1(net_8528), .A2(net_8526) );
NOR3_X4 inst_2361 ( .ZN(net_6253), .A1(net_5273), .A3(net_4994), .A2(net_4992) );
OR3_X4 inst_704 ( .A3(net_2712), .ZN(net_2466), .A1(net_2465), .A2(net_185) );
CLKBUF_X2 inst_11497 ( .A(net_11055), .Z(net_11416) );
AOI21_X2 inst_10237 ( .ZN(net_8848), .A(net_8779), .B1(net_8771), .B2(net_8770) );
AOI22_X2 inst_9301 ( .B1(net_9992), .A1(net_6828), .A2(net_5743), .B2(net_5742), .ZN(net_5677) );
INV_X4 inst_6006 ( .A(net_9646), .ZN(net_625) );
CLKBUF_X2 inst_14652 ( .A(net_14570), .Z(net_14571) );
INV_X4 inst_4542 ( .ZN(net_8711), .A(net_8698) );
INV_X4 inst_5558 ( .ZN(net_2258), .A(net_1371) );
INV_X2 inst_7084 ( .ZN(net_1161), .A(net_1160) );
DFF_X2 inst_8285 ( .Q(net_10395), .D(net_4843), .CK(net_12928) );
INV_X2 inst_6802 ( .A(net_5258), .ZN(net_5232) );
CLKBUF_X2 inst_15538 ( .A(net_15456), .Z(net_15457) );
OAI211_X2 inst_2226 ( .C1(net_7182), .C2(net_6480), .ZN(net_6478), .B(net_5594), .A(net_3679) );
INV_X4 inst_5467 ( .ZN(net_2366), .A(net_2211) );
OR3_X4 inst_694 ( .ZN(net_6542), .A1(net_5171), .A3(net_4787), .A2(net_4630) );
CLKBUF_X2 inst_15689 ( .A(net_12971), .Z(net_15608) );
INV_X4 inst_5574 ( .ZN(net_1476), .A(net_905) );
INV_X4 inst_6382 ( .A(net_9249), .ZN(net_653) );
NOR2_X2 inst_2498 ( .A2(net_9007), .A1(net_9006), .ZN(net_8563) );
CLKBUF_X2 inst_12402 ( .A(net_10762), .Z(net_12321) );
NAND4_X2 inst_3154 ( .ZN(net_1909), .A2(net_1048), .A3(net_108), .A4(net_104), .A1(net_100) );
INV_X2 inst_6986 ( .ZN(net_1659), .A(net_1658) );
CLKBUF_X2 inst_11476 ( .A(net_11394), .Z(net_11395) );
CLKBUF_X2 inst_11523 ( .A(net_11231), .Z(net_11442) );
CLKBUF_X1 inst_8983 ( .A(x185142), .Z(x916) );
INV_X4 inst_5396 ( .ZN(net_1583), .A(net_1169) );
CLKBUF_X2 inst_13885 ( .A(net_13803), .Z(net_13804) );
CLKBUF_X2 inst_11467 ( .A(net_11385), .Z(net_11386) );
INV_X4 inst_5211 ( .ZN(net_2088), .A(net_1523) );
AOI22_X2 inst_9394 ( .B1(net_10002), .A1(net_5743), .B2(net_5742), .ZN(net_5415), .A2(net_242) );
NOR2_X2 inst_2971 ( .ZN(net_2375), .A1(net_1063), .A2(net_1062) );
OAI222_X2 inst_1342 ( .B1(net_7665), .A2(net_7664), .C2(net_7663), .ZN(net_7580), .B2(net_7418), .A1(net_6175), .C1(net_1862) );
CLKBUF_X2 inst_15531 ( .A(net_15449), .Z(net_15450) );
DFF_X2 inst_7814 ( .Q(net_10017), .D(net_6468), .CK(net_15691) );
CLKBUF_X2 inst_12071 ( .A(net_11989), .Z(net_11990) );
OR2_X4 inst_787 ( .ZN(net_5376), .A2(net_2074), .A1(net_2071) );
NAND2_X2 inst_4396 ( .A2(net_10401), .A1(net_10388), .ZN(net_716) );
CLKBUF_X2 inst_11211 ( .A(net_11129), .Z(net_11130) );
INV_X4 inst_4549 ( .ZN(net_8894), .A(net_8578) );
CLKBUF_X2 inst_12958 ( .A(net_11322), .Z(net_12877) );
CLKBUF_X2 inst_15541 ( .A(net_14859), .Z(net_15460) );
DFF_X2 inst_7483 ( .Q(net_9277), .D(net_8073), .CK(net_13133) );
CLKBUF_X2 inst_14439 ( .A(net_12142), .Z(net_14358) );
AND2_X2 inst_10551 ( .A2(net_6625), .A1(net_5972), .ZN(net_3388) );
INV_X4 inst_6012 ( .A(net_10467), .ZN(net_779) );
NAND2_X2 inst_3933 ( .ZN(net_3728), .A2(net_3378), .A1(net_642) );
OR2_X4 inst_825 ( .A2(net_10462), .A1(net_10461), .ZN(net_2710) );
NOR2_X2 inst_2586 ( .A1(net_7280), .ZN(net_7056), .A2(net_6621) );
OAI221_X2 inst_1656 ( .C1(net_7219), .C2(net_5520), .ZN(net_5517), .B2(net_4547), .A(net_3731), .B1(net_566) );
INV_X4 inst_5881 ( .ZN(net_2412), .A(net_677) );
DFF_X2 inst_7928 ( .QN(net_10213), .D(net_5639), .CK(net_15512) );
OAI21_X2 inst_1881 ( .ZN(net_5224), .B1(net_5220), .B2(net_5219), .A(net_1540) );
CLKBUF_X2 inst_15310 ( .A(net_15228), .Z(net_15229) );
CLKBUF_X2 inst_12886 ( .A(net_12386), .Z(net_12805) );
NOR2_X1 inst_3034 ( .ZN(net_1964), .A2(net_1963), .A1(net_1288) );
OAI21_X2 inst_1892 ( .B1(net_7190), .B2(net_4862), .ZN(net_4860), .A(net_4532) );
INV_X4 inst_5590 ( .ZN(net_4988), .A(net_3214) );
DFF_X2 inst_7860 ( .Q(net_9999), .D(net_6429), .CK(net_12779) );
CLKBUF_X2 inst_15507 ( .A(net_11162), .Z(net_15426) );
CLKBUF_X2 inst_11404 ( .A(net_11322), .Z(net_11323) );
XNOR2_X2 inst_295 ( .ZN(net_3389), .A(net_2931), .B(net_1054) );
OR2_X4 inst_726 ( .ZN(net_8691), .A1(net_7916), .A2(net_7699) );
AND2_X2 inst_10583 ( .A1(net_9223), .ZN(net_3098), .A2(net_2543) );
CLKBUF_X2 inst_13018 ( .A(net_12936), .Z(net_12937) );
INV_X4 inst_4726 ( .ZN(net_5178), .A(net_4482) );
DFF_X2 inst_8073 ( .D(net_5257), .QN(net_133), .CK(net_13193) );
XNOR2_X2 inst_320 ( .B(net_9224), .ZN(net_3126), .A(net_3098) );
SDFF_X2 inst_607 ( .QN(net_10302), .D(net_4413), .SE(net_3682), .SI(net_597), .CK(net_11046) );
INV_X4 inst_6484 ( .A(net_10063), .ZN(net_360) );
NOR3_X2 inst_2432 ( .A2(net_4876), .ZN(net_3870), .A3(net_3183), .A1(net_3182) );
CLKBUF_X2 inst_14698 ( .A(net_14616), .Z(net_14617) );
NAND2_X2 inst_4263 ( .ZN(net_2054), .A2(net_1370), .A1(net_860) );
DFF_X2 inst_8273 ( .Q(net_10053), .D(net_4754), .CK(net_14272) );
XOR2_X2 inst_1 ( .Z(net_6943), .A(net_6014), .B(net_1925) );
INV_X4 inst_5061 ( .A(net_3175), .ZN(net_1872) );
INV_X2 inst_6693 ( .ZN(net_8426), .A(net_8329) );
OAI21_X2 inst_1891 ( .B1(net_7192), .B2(net_4862), .ZN(net_4861), .A(net_4533) );
DFF_X2 inst_7614 ( .QN(net_9211), .D(net_6965), .CK(net_11845) );
AOI21_X2 inst_10130 ( .A(net_10409), .B1(net_10385), .ZN(net_4444), .B2(net_2823) );
DFF_X1 inst_8560 ( .Q(net_9770), .D(net_7130), .CK(net_15639) );
NAND2_X2 inst_4343 ( .A2(net_9174), .ZN(net_1034), .A1(net_1033) );
CLKBUF_X2 inst_15399 ( .A(net_15317), .Z(net_15318) );
CLKBUF_X2 inst_12794 ( .A(net_11717), .Z(net_12713) );
INV_X4 inst_5684 ( .ZN(net_3736), .A(net_1381) );
CLKBUF_X2 inst_11537 ( .A(net_11455), .Z(net_11456) );
INV_X4 inst_4558 ( .ZN(net_8482), .A(net_8419) );
INV_X4 inst_6627 ( .A(net_8975), .ZN(net_8972) );
CLKBUF_X2 inst_14862 ( .A(net_14780), .Z(net_14781) );
CLKBUF_X2 inst_14525 ( .A(net_12155), .Z(net_14444) );
CLKBUF_X2 inst_11841 ( .A(net_11759), .Z(net_11760) );
CLKBUF_X2 inst_11493 ( .A(net_11113), .Z(net_11412) );
XNOR2_X2 inst_235 ( .B(net_4910), .ZN(net_4302), .A(net_3982) );
NAND4_X2 inst_3063 ( .ZN(net_5722), .A4(net_4874), .A2(net_3834), .A1(net_3578), .A3(net_3437) );
CLKBUF_X2 inst_13881 ( .A(net_12267), .Z(net_13800) );
DFF_X1 inst_8610 ( .Q(net_9863), .D(net_7188), .CK(net_15468) );
OAI21_X2 inst_1812 ( .ZN(net_6927), .B2(net_6663), .A(net_3203), .B1(net_2322) );
DFF_X2 inst_7608 ( .QN(net_9343), .D(net_7131), .CK(net_15290) );
CLKBUF_X2 inst_12257 ( .A(net_11513), .Z(net_12176) );
INV_X4 inst_5643 ( .A(net_10455), .ZN(net_1117) );
INV_X2 inst_6750 ( .A(net_6902), .ZN(net_6615) );
CLKBUF_X2 inst_12555 ( .A(net_12127), .Z(net_12474) );
DFF_X2 inst_8217 ( .Q(net_10187), .D(net_4830), .CK(net_12869) );
CLKBUF_X2 inst_15036 ( .A(net_14954), .Z(net_14955) );
CLKBUF_X2 inst_14608 ( .A(net_14526), .Z(net_14527) );
DFF_X2 inst_8370 ( .Q(net_10540), .D(net_2264), .CK(net_12320) );
CLKBUF_X2 inst_12051 ( .A(net_10707), .Z(net_11970) );
NAND2_X2 inst_4338 ( .ZN(net_3047), .A2(net_1074), .A1(net_681) );
DFF_X1 inst_8806 ( .Q(net_10447), .D(net_3987), .CK(net_11067) );
CLKBUF_X2 inst_12726 ( .A(net_11908), .Z(net_12645) );
CLKBUF_X2 inst_13066 ( .A(net_12984), .Z(net_12985) );
INV_X4 inst_4721 ( .ZN(net_5351), .A(net_4907) );
CLKBUF_X2 inst_13601 ( .A(net_13519), .Z(net_13520) );
DFF_X2 inst_8194 ( .Q(net_9741), .D(net_5146), .CK(net_13180) );
CLKBUF_X2 inst_12846 ( .A(net_12764), .Z(net_12765) );
NOR2_X2 inst_2835 ( .A1(net_3024), .ZN(net_2367), .A2(net_2366) );
INV_X4 inst_6638 ( .A(net_9067), .ZN(net_9066) );
CLKBUF_X2 inst_11136 ( .A(net_10736), .Z(net_11055) );
AND2_X4 inst_10399 ( .ZN(net_6888), .A1(net_5937), .A2(net_5359) );
NOR2_X2 inst_2731 ( .A2(net_5344), .ZN(net_4494), .A1(net_4170) );
CLKBUF_X2 inst_13019 ( .A(net_12388), .Z(net_12938) );
DFF_X1 inst_8663 ( .D(net_6772), .Q(net_112), .CK(net_12608) );
OAI211_X2 inst_2207 ( .C1(net_7182), .C2(net_6501), .ZN(net_6498), .B(net_5652), .A(net_3679) );
DFF_X2 inst_7841 ( .Q(net_9720), .D(net_6534), .CK(net_15671) );
AOI21_X2 inst_10088 ( .A(net_5361), .ZN(net_5281), .B2(net_5280), .B1(net_2517) );
CLKBUF_X2 inst_15692 ( .A(net_15610), .Z(net_15611) );
INV_X4 inst_5902 ( .ZN(net_5075), .A(net_599) );
INV_X16 inst_7322 ( .ZN(net_8042), .A(net_5296) );
NAND2_X2 inst_3892 ( .ZN(net_3978), .A1(net_3977), .A2(net_3342) );
INV_X4 inst_4813 ( .A(net_7525), .ZN(net_5885) );
CLKBUF_X2 inst_14906 ( .A(net_12938), .Z(net_14825) );
DFF_X1 inst_8829 ( .QN(net_10233), .D(net_2494), .CK(net_10599) );
NAND2_X2 inst_3930 ( .ZN(net_4479), .A2(net_4046), .A1(net_3555) );
NOR2_X2 inst_2867 ( .A1(net_2752), .A2(net_2237), .ZN(net_2039) );
AOI222_X1 inst_9725 ( .A2(net_7586), .C2(net_7584), .ZN(net_4042), .A1(net_4041), .B2(net_3890), .B1(net_1230), .C1(net_827) );
AOI221_X2 inst_9768 ( .C2(net_7586), .ZN(net_7585), .B2(net_7584), .C1(net_7583), .B1(net_7583), .A(net_7440) );
CLKBUF_X2 inst_15348 ( .A(net_13562), .Z(net_15267) );
NAND2_X2 inst_3398 ( .ZN(net_8901), .A2(net_8662), .A1(net_8580) );
SDFF_X2 inst_477 ( .SE(net_9540), .SI(net_8232), .Q(net_293), .D(net_293), .CK(net_13974) );
DFF_X2 inst_7953 ( .QN(net_10214), .D(net_5638), .CK(net_14792) );
CLKBUF_X2 inst_14235 ( .A(net_14153), .Z(net_14154) );
NAND2_X2 inst_3576 ( .ZN(net_7611), .A2(net_7404), .A1(net_2428) );
AOI21_X2 inst_10006 ( .ZN(net_8719), .B1(net_8711), .A(net_8599), .B2(net_8395) );
XNOR2_X2 inst_423 ( .A(net_9618), .B(net_2928), .ZN(net_1391) );
OR2_X4 inst_835 ( .A2(net_10254), .A1(net_10253), .ZN(net_1702) );
NAND3_X2 inst_3305 ( .A3(net_2101), .A1(net_2099), .ZN(net_2086), .A2(net_2085) );
NAND4_X2 inst_3082 ( .A3(net_10280), .ZN(net_4795), .A4(net_4641), .A1(net_4517), .A2(net_3892) );
CLKBUF_X2 inst_14637 ( .A(net_14555), .Z(net_14556) );
NAND2_X2 inst_4137 ( .ZN(net_2188), .A1(net_2147), .A2(net_1683) );
OAI22_X2 inst_1112 ( .A2(net_6190), .B2(net_6184), .ZN(net_5951), .A1(net_5950), .B1(net_5949) );
INV_X2 inst_6852 ( .ZN(net_3383), .A(net_3382) );
AOI21_X2 inst_10153 ( .ZN(net_4132), .A(net_3659), .B2(net_3280), .B1(net_2623) );
AOI222_X1 inst_9678 ( .B1(net_9506), .ZN(net_8312), .A2(net_8310), .B2(net_8309), .C2(net_8308), .C1(net_8234), .A1(x2648) );
NAND2_X2 inst_4081 ( .A1(net_9535), .ZN(net_7823), .A2(net_2610) );
OR3_X2 inst_710 ( .A1(net_7531), .ZN(net_7522), .A3(net_7161), .A2(net_6189) );
OR2_X2 inst_941 ( .A1(net_9195), .ZN(net_1789), .A2(net_1461) );
CLKBUF_X2 inst_14571 ( .A(net_10730), .Z(net_14490) );
NAND2_X4 inst_3350 ( .A2(net_8908), .A1(net_8907), .ZN(net_8516) );
DFF_X1 inst_8869 ( .Q(net_9510), .D(net_9286), .CK(net_13727) );
DFF_X2 inst_8398 ( .Q(net_9157), .CK(net_11791), .D(x3574) );
AND3_X2 inst_10375 ( .A2(net_4230), .ZN(net_4228), .A3(net_4227), .A1(x6599) );
OAI21_X2 inst_1817 ( .ZN(net_7077), .B2(net_6646), .A(net_2347), .B1(net_1485) );
XOR2_X1 inst_56 ( .A(net_9348), .Z(net_1989), .B(net_1988) );
INV_X2 inst_6835 ( .ZN(net_3939), .A(net_3938) );
XNOR2_X2 inst_308 ( .ZN(net_3227), .B(net_2644), .A(net_2504) );
CLKBUF_X2 inst_11056 ( .A(net_10821), .Z(net_10975) );
OAI221_X2 inst_1546 ( .B2(net_7295), .C2(net_7293), .C1(net_7216), .ZN(net_7215), .A(net_6817), .B1(net_1350) );
INV_X2 inst_7208 ( .A(net_9167), .ZN(net_463) );
CLKBUF_X2 inst_11224 ( .A(net_11142), .Z(net_11143) );
AOI21_X2 inst_10081 ( .B2(net_9094), .ZN(net_8992), .A(net_4999), .B1(net_1732) );
XNOR2_X1 inst_455 ( .B(net_9651), .A(net_9650), .ZN(net_1040) );
DFF_X1 inst_8449 ( .Q(net_9430), .D(net_8084), .CK(net_12681) );
CLKBUF_X2 inst_14715 ( .A(net_14633), .Z(net_14634) );
AOI21_X2 inst_10015 ( .ZN(net_8172), .B2(net_8169), .A(net_7283), .B1(net_6904) );
NOR2_X2 inst_2871 ( .ZN(net_3690), .A1(net_1962), .A2(net_794) );
OAI221_X2 inst_1694 ( .B1(net_7201), .A(net_5637), .ZN(net_5463), .C1(net_5462), .C2(net_4477), .B2(net_4455) );
NOR2_X2 inst_2540 ( .ZN(net_8286), .A2(net_8284), .A1(net_8081) );
INV_X2 inst_6833 ( .ZN(net_3982), .A(net_3981) );
DFF_X2 inst_7475 ( .D(net_8071), .Q(net_219), .CK(net_15371) );
CLKBUF_X2 inst_13298 ( .A(net_13216), .Z(net_13217) );
NAND2_X2 inst_3629 ( .A1(net_9081), .ZN(net_7047), .A2(net_7046) );
CLKBUF_X2 inst_12593 ( .A(net_12165), .Z(net_12512) );
INV_X2 inst_7052 ( .A(net_2625), .ZN(net_1324) );
INV_X4 inst_6602 ( .ZN(net_7136), .A(x5647) );
DFF_X2 inst_8114 ( .QN(net_10257), .D(net_5195), .CK(net_12200) );
NOR2_X2 inst_3024 ( .A2(net_10303), .A1(net_10302), .ZN(net_597) );
CLKBUF_X2 inst_13370 ( .A(net_13288), .Z(net_13289) );
AOI221_X2 inst_9946 ( .C2(net_10234), .B1(net_10233), .ZN(net_5276), .A(net_4593), .B2(net_4422), .C1(net_4283) );
CLKBUF_X2 inst_15427 ( .A(net_12965), .Z(net_15346) );
DFF_X1 inst_8454 ( .QN(net_10278), .D(net_8061), .CK(net_10614) );
NAND2_X2 inst_4414 ( .ZN(net_577), .A2(net_188), .A1(net_187) );
INV_X2 inst_7129 ( .A(net_10142), .ZN(net_878) );
CLKBUF_X2 inst_11860 ( .A(net_11725), .Z(net_11779) );
AOI21_X2 inst_10052 ( .ZN(net_7289), .B1(net_7286), .B2(net_7285), .A(net_6054) );
NAND4_X2 inst_3085 ( .ZN(net_4502), .A4(net_4061), .A3(net_3549), .A1(net_3184), .A2(net_2746) );
CLKBUF_X2 inst_15337 ( .A(net_11802), .Z(net_15256) );
DFF_X1 inst_8648 ( .Q(net_8835), .D(net_7303), .CK(net_11412) );
DFF_X2 inst_7620 ( .QN(net_9217), .D(net_7037), .CK(net_11342) );
NAND2_X2 inst_3951 ( .ZN(net_3664), .A2(net_3485), .A1(net_938) );
DFF_X2 inst_8240 ( .D(net_4873), .Q(net_224), .CK(net_11120) );
NAND2_X2 inst_4282 ( .A2(net_10264), .ZN(net_2233), .A1(net_1208) );
INV_X4 inst_5428 ( .ZN(net_4788), .A(net_1240) );
NOR2_X2 inst_2943 ( .A1(net_10245), .ZN(net_1740), .A2(net_1332) );
OAI221_X2 inst_1593 ( .C1(net_10413), .B1(net_7190), .ZN(net_5650), .C2(net_4477), .B2(net_4455), .A(net_3731) );
CLKBUF_X2 inst_13768 ( .A(net_13686), .Z(net_13687) );
INV_X4 inst_5661 ( .A(net_4441), .ZN(net_1223) );
AOI221_X2 inst_9918 ( .B1(net_10507), .C1(net_9665), .B2(net_6415), .ZN(net_5967), .C2(net_5966), .A(net_5253) );
CLKBUF_X2 inst_11541 ( .A(net_11233), .Z(net_11460) );
CLKBUF_X2 inst_14120 ( .A(net_12870), .Z(net_14039) );
OR2_X4 inst_724 ( .ZN(net_8813), .A1(net_8647), .A2(net_7720) );
NAND2_X2 inst_4292 ( .A2(net_10327), .ZN(net_2880), .A1(net_773) );
CLKBUF_X2 inst_12083 ( .A(net_10545), .Z(net_12002) );
NOR3_X2 inst_2449 ( .A2(net_2711), .ZN(net_2580), .A1(net_2465), .A3(net_2083) );
CLKBUF_X2 inst_14869 ( .A(net_14787), .Z(net_14788) );
CLKBUF_X2 inst_14709 ( .A(net_13206), .Z(net_14628) );
INV_X4 inst_6570 ( .A(net_10532), .ZN(net_4877) );
OAI22_X2 inst_975 ( .A1(net_8813), .B2(net_8812), .ZN(net_8806), .A2(net_8804), .B1(net_408) );
CLKBUF_X2 inst_15546 ( .A(net_15464), .Z(net_15465) );
CLKBUF_X2 inst_13683 ( .A(net_13601), .Z(net_13602) );
CLKBUF_X2 inst_13096 ( .A(net_13014), .Z(net_13015) );
NAND3_X2 inst_3191 ( .A2(net_9385), .ZN(net_7655), .A1(net_7638), .A3(net_2724) );
NOR2_X2 inst_2789 ( .A1(net_3069), .ZN(net_3066), .A2(net_3065) );
DFF_X2 inst_7792 ( .Q(net_9797), .D(net_6504), .CK(net_15702) );
AOI22_X2 inst_9504 ( .B1(net_10296), .A1(net_10191), .B2(net_4774), .A2(net_4217), .ZN(net_3819) );
OAI222_X2 inst_1431 ( .B1(net_5486), .ZN(net_3150), .C2(net_3149), .B2(net_3149), .A2(net_2313), .A1(net_2307), .C1(net_1529) );
INV_X4 inst_5714 ( .ZN(net_1534), .A(net_769) );
NAND2_X2 inst_3760 ( .A1(net_9081), .A2(net_5383), .ZN(net_5229) );
CLKBUF_X2 inst_12841 ( .A(net_12759), .Z(net_12760) );
AOI21_X2 inst_10110 ( .ZN(net_4608), .A(net_4330), .B2(net_4068), .B1(net_955) );
OAI222_X2 inst_1398 ( .B2(net_7732), .A2(net_7731), .C2(net_7730), .ZN(net_5700), .B1(net_2977), .A1(net_2013), .C1(net_1179) );
DFF_X2 inst_7639 ( .D(net_6733), .QN(net_153), .CK(net_14248) );
CLKBUF_X2 inst_10783 ( .A(net_10701), .Z(net_10702) );
DFF_X1 inst_8477 ( .Q(net_9599), .D(net_7858), .CK(net_13799) );
INV_X2 inst_7122 ( .A(net_1177), .ZN(net_946) );
NOR2_X2 inst_2849 ( .A2(net_6960), .ZN(net_2256), .A1(net_1345) );
OAI21_X2 inst_1804 ( .ZN(net_7384), .B2(net_7041), .A(net_2349), .B1(net_1632) );
CLKBUF_X2 inst_13808 ( .A(net_13726), .Z(net_13727) );
NOR3_X2 inst_2440 ( .A2(net_9528), .A3(net_9527), .ZN(net_3624), .A1(net_2575) );
INV_X4 inst_6418 ( .A(net_10253), .ZN(net_4172) );
AOI22_X2 inst_9261 ( .A1(net_6892), .B2(net_6625), .ZN(net_6585), .B1(net_5953), .A2(net_5357) );
CLKBUF_X2 inst_15533 ( .A(net_15451), .Z(net_15452) );
CLKBUF_X2 inst_11037 ( .A(net_10799), .Z(net_10956) );
OAI211_X2 inst_2183 ( .C1(net_7241), .C2(net_6548), .ZN(net_6526), .B(net_5653), .A(net_3679) );
CLKBUF_X2 inst_11981 ( .A(net_10981), .Z(net_11900) );
NAND2_X4 inst_3327 ( .A1(net_9034), .A2(net_8942), .ZN(net_8875) );
INV_X4 inst_5068 ( .ZN(net_2201), .A(net_1857) );
AOI21_X2 inst_10241 ( .ZN(net_8856), .B1(net_4412), .B2(net_2680), .A(net_2679) );
NOR2_X2 inst_2659 ( .ZN(net_5179), .A2(net_4782), .A1(net_4353) );
INV_X4 inst_6545 ( .A(net_9205), .ZN(net_334) );
OAI211_X2 inst_2134 ( .C2(net_6774), .ZN(net_6714), .A(net_6339), .B(net_6077), .C1(net_481) );
OAI21_X2 inst_1744 ( .B1(net_8691), .ZN(net_8684), .B2(net_8664), .A(net_7855) );
CLKBUF_X2 inst_13878 ( .A(net_12608), .Z(net_13797) );
INV_X4 inst_4805 ( .ZN(net_4226), .A(net_3618) );
INV_X4 inst_5018 ( .A(net_4204), .ZN(net_2608) );
CLKBUF_X2 inst_11609 ( .A(net_11194), .Z(net_11528) );
INV_X4 inst_5628 ( .ZN(net_5314), .A(net_861) );
INV_X4 inst_5641 ( .A(net_10263), .ZN(net_2627) );
CLKBUF_X2 inst_11958 ( .A(net_11876), .Z(net_11877) );
CLKBUF_X2 inst_11134 ( .A(net_11052), .Z(net_11053) );
OAI22_X2 inst_1155 ( .A1(net_7226), .A2(net_5139), .B2(net_5138), .ZN(net_5118), .B1(net_3576) );
NAND2_X2 inst_4117 ( .ZN(net_2348), .A1(net_2347), .A2(net_1486) );
CLKBUF_X2 inst_11311 ( .A(net_11229), .Z(net_11230) );
XNOR2_X2 inst_207 ( .ZN(net_4945), .A(net_4679), .B(net_1917) );
AOI22_X2 inst_9329 ( .B1(net_9892), .A1(net_6834), .A2(net_5759), .B2(net_5758), .ZN(net_5644) );
DFF_X1 inst_8886 ( .Q(net_9504), .D(net_9280), .CK(net_14369) );
CLKBUF_X2 inst_14467 ( .A(net_14385), .Z(net_14386) );
CLKBUF_X2 inst_11198 ( .A(net_11116), .Z(net_11117) );
AOI21_X2 inst_10047 ( .ZN(net_7389), .A(net_7161), .B1(net_7018), .B2(net_6849) );
CLKBUF_X2 inst_11639 ( .A(net_11557), .Z(net_11558) );
CLKBUF_X2 inst_11954 ( .A(net_11872), .Z(net_11873) );
AND2_X2 inst_10490 ( .ZN(net_7669), .A1(net_7668), .A2(net_7588) );
INV_X2 inst_6940 ( .A(net_2876), .ZN(net_1916) );
AOI22_X2 inst_9615 ( .B1(net_10013), .A1(net_9783), .ZN(net_3438), .B2(net_2468), .A2(net_2462) );
OR3_X2 inst_712 ( .ZN(net_5746), .A2(net_5745), .A3(net_5368), .A1(net_5367) );
AOI221_X2 inst_9912 ( .B1(net_9822), .C1(net_9723), .ZN(net_6447), .A(net_5715), .C2(net_3039), .B2(net_2556) );
OAI22_X2 inst_1215 ( .A1(net_7192), .A2(net_5107), .B2(net_5105), .ZN(net_5034), .B1(net_1577) );
AOI22_X2 inst_9303 ( .B1(net_9694), .A1(net_6834), .A2(net_5755), .B2(net_5754), .ZN(net_5675) );
XNOR2_X2 inst_131 ( .ZN(net_7419), .A(net_7325), .B(net_1824) );
CLKBUF_X2 inst_14271 ( .A(net_13094), .Z(net_14190) );
CLKBUF_X2 inst_15353 ( .A(net_15271), .Z(net_15272) );
CLKBUF_X2 inst_12436 ( .A(net_12354), .Z(net_12355) );
INV_X4 inst_6104 ( .A(net_10298), .ZN(net_489) );
NAND4_X2 inst_3111 ( .ZN(net_4584), .A2(net_4267), .A4(net_4261), .A1(net_4115), .A3(net_2766) );
XOR2_X2 inst_47 ( .B(net_3733), .Z(net_1144), .A(net_1143) );
OAI211_X2 inst_2035 ( .C2(net_8102), .ZN(net_8099), .B(net_8098), .A(net_7997), .C1(net_3997) );
CLKBUF_X2 inst_12360 ( .A(net_12278), .Z(net_12279) );
CLKBUF_X2 inst_14958 ( .A(net_12001), .Z(net_14877) );
CLKBUF_X2 inst_13530 ( .A(net_11072), .Z(net_13449) );
OAI21_X2 inst_1984 ( .B1(net_5452), .ZN(net_2820), .A(net_2515), .B2(net_2184) );
INV_X4 inst_5231 ( .ZN(net_4041), .A(net_1487) );
CLKBUF_X2 inst_14567 ( .A(net_14485), .Z(net_14486) );
CLKBUF_X2 inst_11569 ( .A(net_11487), .Z(net_11488) );
AND2_X4 inst_10442 ( .A1(net_10470), .ZN(net_2783), .A2(net_1189) );
CLKBUF_X2 inst_14686 ( .A(net_14604), .Z(net_14605) );
CLKBUF_X2 inst_11121 ( .A(net_11039), .Z(net_11040) );
AOI22_X2 inst_9458 ( .A2(net_10374), .B2(net_8842), .ZN(net_3934), .B1(net_1327), .A1(net_1275) );
CLKBUF_X2 inst_15563 ( .A(net_15481), .Z(net_15482) );
INV_X4 inst_6520 ( .A(net_9836), .ZN(net_344) );
CLKBUF_X2 inst_14356 ( .A(net_14274), .Z(net_14275) );
CLKBUF_X2 inst_12564 ( .A(net_12482), .Z(net_12483) );
CLKBUF_X2 inst_12397 ( .A(net_12315), .Z(net_12316) );
NAND2_X2 inst_4101 ( .ZN(net_2756), .A2(net_2751), .A1(net_313) );
INV_X4 inst_6483 ( .A(net_10470), .ZN(net_364) );
AND4_X4 inst_10316 ( .ZN(net_8724), .A1(net_8705), .A4(net_8704), .A2(net_8679), .A3(net_5272) );
AOI22_X2 inst_9469 ( .B1(net_9810), .A1(net_9679), .A2(net_5966), .ZN(net_3858), .B2(net_2556) );
CLKBUF_X2 inst_12482 ( .A(net_10892), .Z(net_12401) );
INV_X4 inst_4792 ( .ZN(net_5859), .A(net_3678) );
DFF_X2 inst_7381 ( .D(net_8661), .QN(net_266), .CK(net_12645) );
CLKBUF_X2 inst_14027 ( .A(net_13945), .Z(net_13946) );
SDFF_X2 inst_525 ( .Q(net_9342), .D(net_9342), .SI(net_9334), .SE(net_7588), .CK(net_14677) );
CLKBUF_X2 inst_12738 ( .A(net_10860), .Z(net_12657) );
CLKBUF_X2 inst_15360 ( .A(net_15278), .Z(net_15279) );
XNOR2_X2 inst_434 ( .B(net_9306), .ZN(net_1046), .A(net_229) );
CLKBUF_X2 inst_12196 ( .A(net_12114), .Z(net_12115) );
CLKBUF_X2 inst_11774 ( .A(net_11692), .Z(net_11693) );
NAND2_X2 inst_3455 ( .A1(net_9464), .A2(net_8475), .ZN(net_8469) );
CLKBUF_X2 inst_12424 ( .A(net_12342), .Z(net_12343) );
OAI22_X2 inst_1032 ( .A1(net_9269), .A2(net_7906), .B2(net_7904), .ZN(net_7901), .B1(net_7848) );
CLKBUF_X1 inst_8985 ( .A(x185142), .Z(x926) );
CLKBUF_X2 inst_14099 ( .A(net_12384), .Z(net_14018) );
CLKBUF_X2 inst_12638 ( .A(net_12556), .Z(net_12557) );
INV_X2 inst_6711 ( .A(net_9595), .ZN(net_8104) );
OAI222_X2 inst_1392 ( .B1(net_7665), .A2(net_7664), .C2(net_7663), .ZN(net_5819), .B2(net_4934), .A1(net_3521), .C1(net_1914) );
INV_X4 inst_5932 ( .A(net_1976), .ZN(net_1055) );
DFF_X2 inst_7376 ( .Q(net_9366), .D(net_8674), .CK(net_14189) );
CLKBUF_X2 inst_11816 ( .A(net_10841), .Z(net_11735) );
NAND2_X2 inst_4044 ( .A2(net_8829), .ZN(net_2828), .A1(net_2824) );
DFF_X2 inst_7585 ( .QN(net_10477), .D(net_7497), .CK(net_11405) );
CLKBUF_X2 inst_11682 ( .A(net_11600), .Z(net_11601) );
OAI221_X2 inst_1476 ( .ZN(net_7675), .B1(net_7672), .C2(net_7671), .A(net_7585), .C1(net_7439), .B2(net_4208) );
DFF_X2 inst_8265 ( .Q(net_10388), .D(net_4807), .CK(net_12934) );
CLKBUF_X2 inst_11148 ( .A(net_11066), .Z(net_11067) );
OAI211_X2 inst_2249 ( .C1(net_7237), .C2(net_6480), .ZN(net_6455), .B(net_5524), .A(net_3679) );
CLKBUF_X2 inst_12339 ( .A(net_12257), .Z(net_12258) );
CLKBUF_X2 inst_11106 ( .A(net_10552), .Z(net_11025) );
CLKBUF_X2 inst_13773 ( .A(net_10764), .Z(net_13692) );
AOI22_X2 inst_8995 ( .A2(net_8935), .A1(net_8614), .ZN(net_8613), .B2(net_8612), .B1(net_7633) );
INV_X4 inst_5404 ( .A(net_3067), .ZN(net_1484) );
OAI211_X2 inst_2269 ( .C1(net_7129), .C2(net_6501), .ZN(net_6276), .B(net_5697), .A(net_3679) );
NOR3_X2 inst_2390 ( .A2(net_8838), .A1(net_8818), .ZN(net_7764), .A3(net_7623) );
OAI21_X2 inst_1780 ( .ZN(net_7759), .B2(net_7757), .A(net_7657), .B1(net_5949) );
CLKBUF_X2 inst_11839 ( .A(net_11757), .Z(net_11758) );
OAI222_X1 inst_1436 ( .ZN(net_7789), .A1(net_7660), .B2(net_7659), .C2(net_7658), .A2(net_7654), .B1(net_5763), .C1(net_1203) );
INV_X4 inst_6033 ( .A(net_9996), .ZN(net_517) );
CLKBUF_X2 inst_15149 ( .A(net_15067), .Z(net_15068) );
CLKBUF_X2 inst_14305 ( .A(net_14223), .Z(net_14224) );
OR2_X2 inst_852 ( .ZN(net_8497), .A1(net_8177), .A2(net_8176) );
CLKBUF_X2 inst_12792 ( .A(net_12710), .Z(net_12711) );
DFF_X1 inst_8424 ( .Q(net_9587), .D(net_8732), .CK(net_13821) );
NAND2_X2 inst_3871 ( .ZN(net_4628), .A2(net_4232), .A1(net_4080) );
AOI22_X2 inst_9268 ( .B1(net_9807), .ZN(net_5772), .A1(net_5766), .B2(net_5765), .A2(net_245) );
INV_X2 inst_6663 ( .ZN(net_8365), .A(net_8311) );
NAND2_X2 inst_4306 ( .A2(net_10439), .ZN(net_3399), .A1(net_542) );
CLKBUF_X2 inst_12528 ( .A(net_12446), .Z(net_12447) );
OAI221_X2 inst_1474 ( .A(net_7783), .C1(net_7782), .ZN(net_7691), .B2(net_7690), .C2(net_4404), .B1(net_1478) );
MUX2_X1 inst_4449 ( .S(net_6041), .A(net_297), .B(x5077), .Z(x126) );
INV_X4 inst_6077 ( .A(net_9343), .ZN(net_747) );
CLKBUF_X2 inst_11974 ( .A(net_11442), .Z(net_11893) );
DFF_X2 inst_7637 ( .D(net_6755), .QN(net_128), .CK(net_12000) );
OAI211_X2 inst_2045 ( .C1(net_10239), .ZN(net_7879), .A(net_7878), .B(net_7459), .C2(net_6668) );
OAI21_X2 inst_1920 ( .ZN(net_4561), .A(net_4153), .B2(net_4152), .B1(net_3984) );
CLKBUF_X2 inst_11746 ( .A(net_11444), .Z(net_11665) );
AOI22_X2 inst_9022 ( .B1(net_9522), .A1(net_8002), .B2(net_8001), .ZN(net_7997), .A2(net_7947) );
OAI22_X2 inst_1311 ( .B2(net_9944), .ZN(net_2288), .A2(net_2287), .A1(net_2285), .B1(net_2283) );
AOI22_X2 inst_9307 ( .B1(net_9713), .A2(net_5755), .B2(net_5754), .ZN(net_5671), .A1(net_250) );
INV_X2 inst_7185 ( .A(net_9558), .ZN(net_8091) );
NAND2_X2 inst_3415 ( .ZN(net_8521), .A1(net_8466), .A2(net_8434) );
CLKBUF_X2 inst_13269 ( .A(net_12306), .Z(net_13188) );
CLKBUF_X2 inst_12787 ( .A(net_12705), .Z(net_12706) );
AOI22_X2 inst_9534 ( .B1(net_10405), .A1(net_9866), .B2(net_4062), .ZN(net_3787), .A2(net_2973) );
CLKBUF_X2 inst_10780 ( .A(net_10698), .Z(net_10699) );
INV_X4 inst_4654 ( .A(net_9251), .ZN(net_6626) );
OAI221_X2 inst_1640 ( .B1(net_10421), .C1(net_7234), .ZN(net_5548), .B2(net_4477), .C2(net_4455), .A(net_3731) );
CLKBUF_X2 inst_11359 ( .A(net_11277), .Z(net_11278) );
CLKBUF_X2 inst_11194 ( .A(net_10842), .Z(net_11113) );
NAND3_X2 inst_3234 ( .A1(net_7142), .ZN(net_4724), .A3(net_4723), .A2(net_4719) );
NAND2_X2 inst_4143 ( .ZN(net_2120), .A1(net_2119), .A2(net_1863) );
CLKBUF_X2 inst_13928 ( .A(net_10789), .Z(net_13847) );
CLKBUF_X2 inst_15127 ( .A(net_15045), .Z(net_15046) );
NOR2_X2 inst_2639 ( .A2(net_5927), .ZN(net_5785), .A1(net_3663) );
INV_X4 inst_4747 ( .A(net_10503), .ZN(net_5918) );
DFF_X2 inst_7682 ( .QN(net_9118), .D(net_6611), .CK(net_10881) );
CLKBUF_X2 inst_11122 ( .A(net_10887), .Z(net_11041) );
DFF_X2 inst_7571 ( .QN(net_10162), .D(net_7578), .CK(net_13524) );
CLKBUF_X2 inst_15666 ( .A(net_15584), .Z(net_15585) );
INV_X4 inst_4630 ( .ZN(net_7175), .A(net_7167) );
NOR2_X2 inst_2509 ( .ZN(net_8400), .A1(net_8399), .A2(net_8398) );
INV_X4 inst_5971 ( .A(net_9322), .ZN(net_1450) );
INV_X4 inst_5897 ( .ZN(net_604), .A(net_603) );
NOR2_X2 inst_2542 ( .ZN(net_8310), .A2(net_8308), .A1(net_8081) );
INV_X4 inst_6632 ( .A(net_9037), .ZN(net_9036) );
NAND4_X2 inst_3091 ( .A3(net_9568), .A4(net_9566), .ZN(net_5346), .A2(net_4311), .A1(net_2850) );
NAND2_X2 inst_4197 ( .A1(net_2399), .ZN(net_1808), .A2(net_1336) );
CLKBUF_X2 inst_11791 ( .A(net_11709), .Z(net_11710) );
CLKBUF_X2 inst_15784 ( .A(net_13902), .Z(net_15703) );
AOI22_X2 inst_9506 ( .B1(net_10401), .A2(net_6413), .B2(net_4062), .ZN(net_3817), .A1(net_2945) );
INV_X2 inst_6829 ( .ZN(net_4079), .A(net_4078) );
DFF_X2 inst_7567 ( .QN(net_9382), .D(net_7628), .CK(net_13026) );
INV_X4 inst_6590 ( .A(net_10292), .ZN(net_323) );
CLKBUF_X2 inst_15354 ( .A(net_15272), .Z(net_15273) );
XNOR2_X2 inst_417 ( .ZN(net_1408), .B(net_1406), .A(net_194) );
SDFF_X2 inst_671 ( .SI(net_9486), .Q(net_9486), .SE(net_3073), .CK(net_12388), .D(x2278) );
DFF_X2 inst_7400 ( .D(net_8442), .QN(net_231), .CK(net_12071) );
CLKBUF_X2 inst_15812 ( .A(net_11259), .Z(net_15731) );
CLKBUF_X2 inst_13473 ( .A(net_13391), .Z(net_13392) );
CLKBUF_X2 inst_12733 ( .A(net_12651), .Z(net_12652) );
XOR2_X2 inst_21 ( .B(net_9369), .Z(net_2726), .A(net_2725) );
AOI22_X2 inst_9462 ( .B1(net_9905), .A1(net_9707), .B2(net_4969), .ZN(net_3865), .A2(net_3039) );
CLKBUF_X2 inst_14782 ( .A(net_11734), .Z(net_14701) );
CLKBUF_X2 inst_13745 ( .A(net_13663), .Z(net_13664) );
INV_X8 inst_4524 ( .A(net_8960), .ZN(net_8958) );
CLKBUF_X2 inst_11024 ( .A(net_10942), .Z(net_10943) );
INV_X4 inst_4871 ( .A(net_3298), .ZN(net_3297) );
AOI211_X2 inst_10286 ( .ZN(net_5181), .A(net_5180), .B(net_4907), .C2(net_4893), .C1(net_1070) );
INV_X4 inst_5520 ( .ZN(net_1326), .A(net_966) );
NAND2_X2 inst_3885 ( .ZN(net_7602), .A2(net_4016), .A1(net_2085) );
NOR4_X2 inst_2311 ( .A3(net_10514), .A1(net_10513), .ZN(net_7478), .A4(net_7273), .A2(net_551) );
NAND2_X2 inst_4257 ( .ZN(net_2913), .A2(net_1384), .A1(net_838) );
INV_X4 inst_4586 ( .ZN(net_8064), .A(net_8022) );
DFF_X2 inst_7703 ( .Q(net_10006), .D(net_6439), .CK(net_15075) );
CLKBUF_X2 inst_13722 ( .A(net_13640), .Z(net_13641) );
OAI22_X2 inst_1317 ( .A2(net_2880), .B2(net_2646), .ZN(net_2133), .A1(net_2132), .B1(net_2131) );
INV_X2 inst_6820 ( .A(net_5160), .ZN(net_4605) );
NAND2_X2 inst_3683 ( .A2(net_9115), .ZN(net_5999), .A1(net_5998) );
NOR2_X2 inst_2941 ( .ZN(net_1951), .A2(net_1733), .A1(net_1732) );
CLKBUF_X2 inst_13655 ( .A(net_10909), .Z(net_13574) );
AOI22_X2 inst_9623 ( .B1(net_9797), .A2(net_5174), .ZN(net_3428), .B2(net_2556), .A1(net_1885) );
CLKBUF_X2 inst_12603 ( .A(net_11210), .Z(net_12522) );
CLKBUF_X2 inst_13528 ( .A(net_13446), .Z(net_13447) );
CLKBUF_X2 inst_12351 ( .A(net_12269), .Z(net_12270) );
AOI221_X2 inst_9861 ( .A(net_6889), .B2(net_6888), .C2(net_6887), .ZN(net_6857), .B1(net_668), .C1(x4694) );
AOI22_X2 inst_9203 ( .A1(net_9863), .B1(net_9764), .A2(net_6141), .B2(net_6133), .ZN(net_6108) );
SDFF_X2 inst_624 ( .Q(net_9443), .D(net_9443), .SE(net_3293), .CK(net_14660), .SI(x2968) );
INV_X4 inst_6284 ( .A(net_9967), .ZN(net_437) );
INV_X4 inst_5728 ( .ZN(net_835), .A(net_755) );
DFF_X1 inst_8442 ( .Q(net_9433), .D(net_8402), .CK(net_14942) );
INV_X4 inst_6404 ( .A(net_9826), .ZN(net_390) );
CLKBUF_X2 inst_11930 ( .A(net_11324), .Z(net_11849) );
CLKBUF_X2 inst_10920 ( .A(net_10838), .Z(net_10839) );
INV_X4 inst_6419 ( .A(net_10006), .ZN(net_384) );
AOI221_X2 inst_9886 ( .B1(net_9792), .B2(net_9098), .A(net_6940), .C2(net_6939), .ZN(net_6810), .C1(net_262) );
CLKBUF_X2 inst_11247 ( .A(net_10919), .Z(net_11166) );
AOI22_X2 inst_9375 ( .B1(net_10011), .A2(net_5743), .B2(net_5742), .ZN(net_5530), .A1(net_251) );
NOR2_X2 inst_2637 ( .A2(net_5927), .ZN(net_5817), .A1(net_3126) );
AOI22_X2 inst_9604 ( .B1(net_9992), .A2(net_3500), .ZN(net_3463), .B2(net_2468), .A1(net_313) );
NAND2_X2 inst_3624 ( .ZN(net_7102), .A1(net_6886), .A2(net_6643) );
CLKBUF_X2 inst_13207 ( .A(net_11671), .Z(net_13126) );
XNOR2_X2 inst_236 ( .ZN(net_4262), .A(net_4261), .B(net_2061) );
CLKBUF_X2 inst_14598 ( .A(net_14028), .Z(net_14517) );
CLKBUF_X2 inst_11440 ( .A(net_11264), .Z(net_11359) );
INV_X4 inst_4539 ( .ZN(net_9010), .A(net_8727) );
CLKBUF_X2 inst_12389 ( .A(net_12307), .Z(net_12308) );
NAND2_X2 inst_3878 ( .ZN(net_4030), .A1(net_4029), .A2(net_4028) );
CLKBUF_X2 inst_13295 ( .A(net_13213), .Z(net_13214) );
CLKBUF_X2 inst_13262 ( .A(net_12958), .Z(net_13181) );
AOI221_X2 inst_9806 ( .B1(net_9985), .A(net_7090), .B2(net_7089), .C2(net_7088), .ZN(net_6996), .C1(net_257) );
CLKBUF_X2 inst_14805 ( .A(net_14723), .Z(net_14724) );
NAND3_X2 inst_3172 ( .A3(net_9005), .A1(net_8950), .ZN(net_8940), .A2(net_8497) );
OAI22_X2 inst_986 ( .A2(net_8962), .B2(net_8659), .ZN(net_8654), .A1(net_6294), .B1(net_6231) );
INV_X8 inst_4532 ( .A(net_9107), .ZN(net_9105) );
INV_X4 inst_4983 ( .ZN(net_2560), .A(net_2242) );
INV_X4 inst_6277 ( .ZN(net_443), .A(net_207) );
CLKBUF_X2 inst_12962 ( .A(net_12880), .Z(net_12881) );
OAI222_X2 inst_1422 ( .B2(net_7665), .A2(net_7664), .C2(net_7663), .ZN(net_4913), .B1(net_4256), .A1(net_3275), .C1(net_2097) );
INV_X4 inst_5600 ( .A(net_985), .ZN(net_881) );
AOI211_X2 inst_10263 ( .ZN(net_7892), .A(net_7809), .B(net_7563), .C2(net_5682), .C1(net_1636) );
DFF_X2 inst_8337 ( .QN(net_9565), .D(net_3247), .CK(net_14208) );
NAND2_X2 inst_3508 ( .A2(net_8930), .ZN(net_8165), .A1(net_8164) );
INV_X4 inst_5132 ( .ZN(net_1937), .A(net_1595) );
INV_X4 inst_6327 ( .A(net_10148), .ZN(net_4157) );
AOI222_X1 inst_9702 ( .B1(net_9507), .A2(net_8295), .B2(net_8294), .C2(net_8293), .ZN(net_8276), .C1(net_8211), .A1(x3071) );
INV_X2 inst_6893 ( .ZN(net_3106), .A(net_2927) );
CLKBUF_X2 inst_14955 ( .A(net_14873), .Z(net_14874) );
AND2_X2 inst_10522 ( .ZN(net_4445), .A1(net_4166), .A2(net_4165) );
OAI22_X2 inst_1221 ( .A2(net_5155), .ZN(net_5026), .A1(net_4877), .B1(net_4876), .B2(net_3387) );
DFF_X1 inst_8675 ( .D(net_6745), .Q(net_108), .CK(net_15615) );
OAI22_X2 inst_1133 ( .A1(net_7184), .A2(net_5151), .B2(net_5150), .ZN(net_5145), .B1(net_460) );
DFF_X2 inst_7750 ( .Q(net_9655), .D(net_6262), .CK(net_11824) );
CLKBUF_X2 inst_15000 ( .A(net_14918), .Z(net_14919) );
CLKBUF_X2 inst_12158 ( .A(net_11438), .Z(net_12077) );
INV_X4 inst_4580 ( .ZN(net_8070), .A(net_8028) );
AOI221_X2 inst_9990 ( .ZN(net_3451), .C2(net_3450), .B2(net_3450), .C1(net_2695), .A(net_2438), .B1(net_1348) );
OAI211_X2 inst_2103 ( .C2(net_6778), .ZN(net_6745), .A(net_6373), .B(net_6103), .C1(net_437) );
DFF_X2 inst_7951 ( .QN(net_10211), .D(net_5641), .CK(net_15493) );
DFF_X1 inst_8710 ( .Q(net_9379), .D(net_6954), .CK(net_13065) );
CLKBUF_X2 inst_14040 ( .A(net_13958), .Z(net_13959) );
CLKBUF_X2 inst_15121 ( .A(net_11382), .Z(net_15040) );
INV_X4 inst_5139 ( .ZN(net_3085), .A(net_3068) );
CLKBUF_X2 inst_10793 ( .A(net_10711), .Z(net_10712) );
NOR2_X2 inst_2664 ( .A2(net_9079), .ZN(net_5808), .A1(net_790) );
XNOR2_X2 inst_339 ( .ZN(net_2931), .B(net_1998), .A(net_1083) );
INV_X4 inst_4750 ( .A(net_4369), .ZN(net_4368) );
CLKBUF_X2 inst_13995 ( .A(net_13913), .Z(net_13914) );
XNOR2_X2 inst_351 ( .B(net_4283), .ZN(net_2815), .A(net_2509) );
INV_X4 inst_6615 ( .A(net_8935), .ZN(net_8934) );
CLKBUF_X2 inst_11615 ( .A(net_11533), .Z(net_11534) );
AOI211_X2 inst_10257 ( .A(net_8190), .ZN(net_8159), .C2(net_7929), .C1(net_7388), .B(net_3298) );
AOI22_X2 inst_9557 ( .B1(net_9726), .B2(net_6442), .A2(net_5173), .ZN(net_3763), .A1(net_197) );
DFF_X1 inst_8761 ( .Q(net_9134), .D(net_5299), .CK(net_10962) );
CLKBUF_X2 inst_15463 ( .A(net_13887), .Z(net_15382) );
DFF_X2 inst_7852 ( .Q(net_9800), .D(net_6222), .CK(net_13327) );
INV_X2 inst_6757 ( .ZN(net_6244), .A(net_6243) );
CLKBUF_X2 inst_12507 ( .A(net_12425), .Z(net_12426) );
DFF_X2 inst_8170 ( .QN(net_10027), .D(net_5044), .CK(net_13696) );
DFF_X2 inst_7915 ( .Q(net_9945), .D(net_5876), .CK(net_11944) );
INV_X4 inst_5862 ( .ZN(net_1352), .A(net_1036) );
DFF_X2 inst_7651 ( .D(net_6708), .QN(net_168), .CK(net_14242) );
CLKBUF_X2 inst_14007 ( .A(net_11630), .Z(net_13926) );
CLKBUF_X2 inst_10966 ( .A(net_10884), .Z(net_10885) );
OAI221_X2 inst_1560 ( .C2(net_9047), .B2(net_7287), .B1(net_7198), .ZN(net_7195), .A(net_6792), .C1(net_5491) );
DFF_X2 inst_7658 ( .D(net_6693), .QN(net_169), .CK(net_15076) );
CLKBUF_X2 inst_15253 ( .A(net_15171), .Z(net_15172) );
CLKBUF_X2 inst_11463 ( .A(net_11029), .Z(net_11382) );
CLKBUF_X2 inst_11381 ( .A(net_11299), .Z(net_11300) );
CLKBUF_X2 inst_12622 ( .A(net_12389), .Z(net_12541) );
CLKBUF_X2 inst_10868 ( .A(net_10786), .Z(net_10787) );
AND2_X2 inst_10570 ( .ZN(net_3467), .A2(net_3005), .A1(net_1500) );
CLKBUF_X2 inst_10994 ( .A(net_10912), .Z(net_10913) );
DFF_X2 inst_8051 ( .Q(net_9545), .D(net_9251), .CK(net_13864) );
CLKBUF_X2 inst_13915 ( .A(net_13833), .Z(net_13834) );
DFF_X1 inst_8413 ( .Q(net_9605), .D(net_8794), .CK(net_15191) );
CLKBUF_X2 inst_15811 ( .A(net_15729), .Z(net_15730) );
NAND2_X2 inst_3932 ( .ZN(net_3729), .A2(net_3378), .A1(net_726) );
AOI21_X2 inst_10203 ( .B1(net_5175), .A(net_2783), .ZN(net_2638), .B2(net_1145) );
INV_X2 inst_7035 ( .ZN(net_1422), .A(net_927) );
CLKBUF_X2 inst_13634 ( .A(net_13291), .Z(net_13553) );
AOI22_X2 inst_9224 ( .A1(net_9918), .B1(net_9819), .A2(net_8042), .B2(net_6140), .ZN(net_6087) );
CLKBUF_X2 inst_15205 ( .A(net_15123), .Z(net_15124) );
CLKBUF_X2 inst_11164 ( .A(net_11082), .Z(net_11083) );
AOI21_X2 inst_10161 ( .B1(net_9522), .ZN(net_3997), .A(net_3662), .B2(net_3482) );
INV_X4 inst_6295 ( .A(net_9734), .ZN(net_684) );
OR2_X2 inst_847 ( .A2(net_9581), .ZN(net_8704), .A1(net_767) );
NOR2_X2 inst_2720 ( .A1(net_5347), .ZN(net_4667), .A2(net_133) );
INV_X4 inst_6577 ( .A(net_9250), .ZN(net_558) );
OAI221_X2 inst_1716 ( .ZN(net_3621), .A(net_3152), .C1(net_2943), .C2(net_2315), .B2(net_2302), .B1(net_2301) );
OAI21_X2 inst_1942 ( .B2(net_10234), .A(net_10233), .ZN(net_4284), .B1(net_4283) );
CLKBUF_X2 inst_11433 ( .A(net_10842), .Z(net_11352) );
CLKBUF_X2 inst_10857 ( .A(net_10775), .Z(net_10776) );
AOI221_X2 inst_9788 ( .B1(net_9969), .A(net_7090), .B2(net_7089), .C1(net_7088), .ZN(net_7063), .C2(net_241) );
INV_X4 inst_5950 ( .A(net_5261), .ZN(net_1396) );
CLKBUF_X2 inst_13573 ( .A(net_13491), .Z(net_13492) );
AOI22_X2 inst_9136 ( .A1(net_9720), .A2(net_6418), .ZN(net_6352), .B2(net_5263), .B1(net_3897) );
CLKBUF_X2 inst_11429 ( .A(net_11016), .Z(net_11348) );
NOR2_X2 inst_2648 ( .ZN(net_5384), .A1(net_5383), .A2(net_4941) );
INV_X2 inst_7055 ( .ZN(net_1305), .A(net_610) );
CLKBUF_X2 inst_15470 ( .A(net_14812), .Z(net_15389) );
DFF_X2 inst_7919 ( .Q(net_9221), .D(net_5921), .CK(net_13009) );
DFF_X2 inst_8372 ( .QN(net_9117), .D(net_1511), .CK(net_11588) );
OAI22_X2 inst_1146 ( .A1(net_7182), .A2(net_5134), .B2(net_5133), .ZN(net_5127), .B1(net_633) );
CLKBUF_X2 inst_12947 ( .A(net_12865), .Z(net_12866) );
NAND2_X2 inst_3708 ( .ZN(net_5919), .A1(net_5918), .A2(net_5917) );
CLKBUF_X2 inst_13112 ( .A(net_13030), .Z(net_13031) );
INV_X4 inst_5512 ( .A(net_10327), .ZN(net_2132) );
CLKBUF_X2 inst_12265 ( .A(net_12183), .Z(net_12184) );
CLKBUF_X2 inst_11973 ( .A(net_10858), .Z(net_11892) );
NAND2_X2 inst_4023 ( .A2(net_7095), .ZN(net_6188), .A1(net_5938) );
NAND2_X2 inst_3781 ( .A2(net_7277), .ZN(net_4991), .A1(net_764) );
NAND2_X2 inst_3673 ( .A2(net_8326), .ZN(net_6894), .A1(net_5012) );
NAND4_X2 inst_3105 ( .ZN(net_4338), .A2(net_3795), .A3(net_3794), .A4(net_3793), .A1(net_3337) );
INV_X4 inst_5162 ( .ZN(net_1891), .A(net_1846) );
INV_X8 inst_4519 ( .A(net_8924), .ZN(net_8920) );
INV_X4 inst_5349 ( .ZN(net_1239), .A(net_668) );
INV_X4 inst_6210 ( .A(net_9302), .ZN(net_7499) );
AOI221_X2 inst_9899 ( .B1(net_9884), .B2(net_9101), .A(net_6945), .C2(net_6944), .C1(net_6821), .ZN(net_6795) );
AOI22_X2 inst_9081 ( .A1(net_9668), .ZN(net_6421), .A2(net_6420), .B2(net_5263), .B1(net_106) );
NAND2_X2 inst_3539 ( .ZN(net_8011), .A2(net_8010), .A1(net_208) );
NAND2_X2 inst_3552 ( .A1(net_10299), .ZN(net_7872), .A2(net_7865) );
NOR3_X2 inst_2457 ( .A3(net_4033), .A2(net_4022), .A1(net_1708), .ZN(net_1424) );
OAI221_X2 inst_1702 ( .ZN(net_5377), .B1(net_5376), .C2(net_5375), .B2(net_4915), .A(net_4911), .C1(net_3504) );
DFF_X2 inst_8307 ( .Q(net_9621), .D(net_4539), .CK(net_14084) );
AOI21_X2 inst_10188 ( .B2(net_4328), .ZN(net_3361), .A(net_3360), .B1(net_3170) );
XNOR2_X2 inst_274 ( .ZN(net_3951), .A(net_3243), .B(net_2893) );
CLKBUF_X2 inst_15076 ( .A(net_13168), .Z(net_14995) );
CLKBUF_X2 inst_14543 ( .A(net_14461), .Z(net_14462) );
OAI22_X2 inst_1277 ( .B2(net_7671), .A1(net_7602), .ZN(net_4459), .B1(net_3909), .A2(net_3882) );
HA_X1 inst_7329 ( .S(net_7654), .CO(net_7653), .B(net_7464), .A(net_5794) );
NOR2_X2 inst_2817 ( .ZN(net_3160), .A1(net_1977), .A2(net_593) );
CLKBUF_X2 inst_13135 ( .A(net_11986), .Z(net_13054) );
NAND2_X2 inst_4076 ( .A1(net_9538), .ZN(net_3302), .A2(net_2619) );
OAI211_X2 inst_2092 ( .C2(net_6774), .ZN(net_6756), .A(net_6384), .B(net_6116), .C1(net_478) );
CLKBUF_X2 inst_13436 ( .A(net_13354), .Z(net_13355) );
NAND3_X2 inst_3207 ( .ZN(net_6910), .A3(net_5967), .A1(net_3990), .A2(net_3814) );
NAND4_X2 inst_3143 ( .A3(net_9245), .ZN(net_2489), .A1(net_2488), .A4(net_2487), .A2(net_1459) );
INV_X2 inst_7112 ( .A(net_1386), .ZN(net_1318) );
CLKBUF_X2 inst_11387 ( .A(net_11305), .Z(net_11306) );
NOR2_X2 inst_2696 ( .ZN(net_4598), .A2(net_4414), .A1(net_1235) );
INV_X4 inst_5586 ( .ZN(net_6053), .A(net_1960) );
CLKBUF_X2 inst_14063 ( .A(net_13981), .Z(net_13982) );
CLKBUF_X2 inst_13784 ( .A(net_13702), .Z(net_13703) );
INV_X2 inst_7136 ( .ZN(net_832), .A(net_831) );
NOR2_X2 inst_2880 ( .ZN(net_2657), .A2(net_2210), .A1(net_1583) );
OAI21_X2 inst_1771 ( .ZN(net_8008), .A(net_7872), .B2(net_7866), .B1(net_7157) );
CLKBUF_X2 inst_14402 ( .A(net_14320), .Z(net_14321) );
OAI221_X4 inst_1440 ( .B2(net_9081), .C2(net_8992), .C1(net_8991), .ZN(net_6682), .A(net_5429), .B1(net_2247) );
CLKBUF_X2 inst_15522 ( .A(net_15440), .Z(net_15441) );
CLKBUF_X2 inst_13611 ( .A(net_13529), .Z(net_13530) );
AOI22_X2 inst_9415 ( .A1(net_10177), .A2(net_4656), .B2(net_4655), .ZN(net_4654), .B1(x4359) );
NOR2_X2 inst_2660 ( .ZN(net_5016), .A2(net_5015), .A1(net_2906) );
AOI221_X2 inst_9854 ( .A(net_6889), .B2(net_6888), .C2(net_6887), .ZN(net_6864), .B1(net_1232), .C1(x4117) );
CLKBUF_X2 inst_13734 ( .A(net_13171), .Z(net_13653) );
DFF_X2 inst_7859 ( .Q(net_10064), .D(net_6200), .CK(net_11176) );
CLKBUF_X2 inst_13729 ( .A(net_12281), .Z(net_13648) );
NAND2_X4 inst_3355 ( .A2(net_9012), .ZN(net_8384), .A1(net_8379) );
NOR3_X2 inst_2389 ( .A2(net_8835), .A1(net_8820), .ZN(net_7765), .A3(net_7625) );
INV_X4 inst_5912 ( .ZN(net_941), .A(net_590) );
CLKBUF_X2 inst_10802 ( .A(net_10720), .Z(net_10721) );
CLKBUF_X2 inst_12148 ( .A(net_11053), .Z(net_12067) );
INV_X4 inst_6199 ( .A(net_9377), .ZN(net_623) );
DFF_X2 inst_8179 ( .QN(net_9830), .D(net_5025), .CK(net_14438) );
INV_X4 inst_4946 ( .ZN(net_2570), .A(net_2569) );
OAI211_X2 inst_2148 ( .C2(net_6774), .ZN(net_6700), .A(net_6324), .B(net_6063), .C1(net_4753) );
INV_X4 inst_6213 ( .A(net_10108), .ZN(net_5856) );
INV_X4 inst_5784 ( .ZN(net_978), .A(net_701) );
CLKBUF_X2 inst_13488 ( .A(net_13406), .Z(net_13407) );
DFF_X2 inst_8354 ( .QN(net_10232), .D(net_2858), .CK(net_10983) );
NOR2_X2 inst_2900 ( .A2(net_6958), .ZN(net_1653), .A1(net_993) );
OAI221_X2 inst_1591 ( .B2(net_10166), .ZN(net_5982), .A(net_5224), .C2(net_5221), .C1(net_4246), .B1(net_3960) );
NAND2_X2 inst_3697 ( .ZN(net_7531), .A2(net_7015), .A1(net_2615) );
NAND3_X2 inst_3247 ( .ZN(net_5190), .A3(net_4665), .A1(net_621), .A2(net_580) );
CLKBUF_X2 inst_13544 ( .A(net_13325), .Z(net_13463) );
XNOR2_X2 inst_379 ( .B(net_9359), .ZN(net_2449), .A(net_1077) );
OR2_X2 inst_926 ( .A2(net_7521), .A1(net_6847), .ZN(net_2998) );
CLKBUF_X2 inst_12348 ( .A(net_11644), .Z(net_12267) );
INV_X4 inst_5470 ( .ZN(net_5407), .A(net_1382) );
CLKBUF_X2 inst_10997 ( .A(net_10688), .Z(net_10916) );
DFF_X2 inst_8312 ( .Q(net_9620), .D(net_4151), .CK(net_14081) );
DFF_X2 inst_7827 ( .Q(net_9992), .D(net_6476), .CK(net_14609) );
CLKBUF_X2 inst_12856 ( .A(net_12774), .Z(net_12775) );
NOR2_X2 inst_2570 ( .ZN(net_7815), .A1(net_7461), .A2(net_7376) );
NAND2_X2 inst_4153 ( .ZN(net_2044), .A2(net_2043), .A1(net_1174) );
CLKBUF_X2 inst_13586 ( .A(net_12172), .Z(net_13505) );
DFF_X1 inst_8684 ( .D(net_6720), .Q(net_136), .CK(net_15441) );
AND2_X2 inst_10624 ( .ZN(net_583), .A2(x3858), .A1(x3849) );
INV_X4 inst_4960 ( .A(net_3095), .ZN(net_2826) );
CLKBUF_X2 inst_15741 ( .A(net_15659), .Z(net_15660) );
CLKBUF_X2 inst_14205 ( .A(net_14123), .Z(net_14124) );
AOI22_X2 inst_9098 ( .A1(net_9679), .A2(net_6402), .ZN(net_6394), .B2(net_5263), .B1(net_4022) );
NAND2_X2 inst_3719 ( .A1(net_8107), .ZN(net_7038), .A2(net_5818) );
NAND2_X2 inst_3646 ( .A1(net_9502), .ZN(net_6838), .A2(net_6669) );
OR2_X2 inst_891 ( .A1(net_10058), .ZN(net_5897), .A2(net_5896) );
NAND2_X2 inst_4095 ( .ZN(net_2539), .A2(net_2538), .A1(net_1946) );
AOI22_X2 inst_9479 ( .B1(net_9880), .A2(net_5173), .ZN(net_3844), .B2(net_2973), .A1(net_213) );
XNOR2_X2 inst_74 ( .A(net_9042), .ZN(net_8672), .B(net_2995) );
CLKBUF_X2 inst_13357 ( .A(net_13275), .Z(net_13276) );
OAI211_X2 inst_2244 ( .C1(net_7213), .C2(net_6542), .ZN(net_6460), .B(net_5606), .A(net_3679) );
INV_X4 inst_5682 ( .ZN(net_2283), .A(net_1817) );
CLKBUF_X2 inst_14739 ( .A(net_14657), .Z(net_14658) );
XNOR2_X2 inst_288 ( .B(net_9206), .ZN(net_3524), .A(net_3513) );
CLKBUF_X2 inst_14414 ( .A(net_14332), .Z(net_14333) );
CLKBUF_X2 inst_11435 ( .A(net_11353), .Z(net_11354) );
NAND3_X2 inst_3284 ( .A1(net_4328), .A3(net_3891), .ZN(net_3449), .A2(net_757) );
CLKBUF_X2 inst_11729 ( .A(net_11647), .Z(net_11648) );
INV_X2 inst_7263 ( .ZN(net_315), .A(net_200) );
CLKBUF_X2 inst_14265 ( .A(net_14183), .Z(net_14184) );
OAI22_X2 inst_1298 ( .A2(net_10442), .B2(net_8839), .ZN(net_3396), .A1(net_3175), .B1(net_1117) );
INV_X8 inst_4512 ( .ZN(net_6892), .A(net_6625) );
INV_X4 inst_5648 ( .ZN(net_1166), .A(net_838) );
INV_X4 inst_5719 ( .A(net_1816), .ZN(net_763) );
CLKBUF_X2 inst_15059 ( .A(net_14977), .Z(net_14978) );
CLKBUF_X2 inst_14636 ( .A(net_10817), .Z(net_14555) );
AOI22_X2 inst_9147 ( .A1(net_9701), .A2(net_6382), .ZN(net_6338), .B2(net_5263), .B1(net_141) );
CLKBUF_X2 inst_14856 ( .A(net_14774), .Z(net_14775) );
CLKBUF_X2 inst_12032 ( .A(net_10841), .Z(net_11951) );
DFF_X2 inst_8241 ( .D(net_4872), .Q(net_225), .CK(net_10801) );
INV_X4 inst_6499 ( .A(net_9844), .ZN(net_688) );
DFF_X1 inst_8483 ( .QN(net_9629), .D(net_7947), .CK(net_15017) );
XNOR2_X2 inst_372 ( .ZN(net_2477), .B(net_2476), .A(net_2451) );
DFF_X2 inst_7388 ( .D(net_8653), .QN(net_273), .CK(net_14915) );
DFF_X2 inst_8031 ( .QN(net_10432), .D(net_5453), .CK(net_11459) );
CLKBUF_X2 inst_13619 ( .A(net_13537), .Z(net_13538) );
CLKBUF_X2 inst_11234 ( .A(net_11152), .Z(net_11153) );
INV_X4 inst_5991 ( .ZN(net_2928), .A(net_313) );
CLKBUF_X2 inst_15142 ( .A(net_15060), .Z(net_15061) );
CLKBUF_X2 inst_14623 ( .A(net_14541), .Z(net_14542) );
AOI22_X2 inst_9218 ( .A1(net_9893), .B1(net_9794), .B2(net_8041), .A2(net_6109), .ZN(net_6093) );
DFF_X1 inst_8512 ( .D(net_7594), .Q(net_263), .CK(net_15181) );
INV_X2 inst_6949 ( .ZN(net_1896), .A(net_1895) );
INV_X4 inst_5709 ( .A(net_1978), .ZN(net_831) );
CLKBUF_X2 inst_11401 ( .A(net_11319), .Z(net_11320) );
INV_X4 inst_5835 ( .A(net_4157), .ZN(net_658) );
CLKBUF_X2 inst_11128 ( .A(net_10633), .Z(net_11047) );
NOR3_X2 inst_2397 ( .A1(net_7828), .ZN(net_7613), .A3(net_7527), .A2(x3390) );
OAI21_X2 inst_1775 ( .ZN(net_7813), .A(net_7713), .B1(net_7644), .B2(net_7486) );
INV_X4 inst_5335 ( .A(net_2945), .ZN(net_2630) );
INV_X4 inst_6223 ( .A(net_10223), .ZN(net_2210) );
CLKBUF_X2 inst_12802 ( .A(net_10752), .Z(net_12721) );
CLKBUF_X2 inst_13539 ( .A(net_11882), .Z(net_13458) );
OAI22_X2 inst_1172 ( .B1(net_10040), .A1(net_7182), .A2(net_5107), .B2(net_5105), .ZN(net_5089) );
AOI222_X1 inst_9709 ( .ZN(net_7911), .A1(net_7910), .A2(net_7909), .B2(net_7801), .C2(net_5164), .C1(net_3088), .B1(net_685) );
OAI22_X2 inst_1090 ( .A1(net_9202), .A2(net_9064), .B2(net_6639), .ZN(net_6557), .B1(net_1463) );
AOI22_X2 inst_9088 ( .A1(net_9702), .A2(net_6420), .ZN(net_6406), .B2(net_5263), .B1(net_142) );
NAND2_X2 inst_3903 ( .A2(net_3903), .ZN(net_3902), .A1(net_102) );
NOR3_X2 inst_2372 ( .A3(net_10488), .A2(net_10487), .ZN(net_8156), .A1(net_1395) );
DFF_X2 inst_7467 ( .QN(net_9517), .D(net_8103), .CK(net_14972) );
CLKBUF_X2 inst_13454 ( .A(net_12308), .Z(net_13373) );
NOR2_X2 inst_2575 ( .A1(net_8858), .ZN(net_7292), .A2(net_7291) );
INV_X4 inst_5007 ( .A(net_2546), .ZN(net_2170) );
CLKBUF_X2 inst_10923 ( .A(net_10841), .Z(net_10842) );
OAI22_X2 inst_1239 ( .A1(net_7245), .ZN(net_4873), .A2(net_4871), .B2(net_4870), .B1(net_1995) );
CLKBUF_X2 inst_13521 ( .A(net_12534), .Z(net_13440) );
CLKBUF_X2 inst_12496 ( .A(net_12414), .Z(net_12415) );
INV_X4 inst_5655 ( .A(net_835), .ZN(net_827) );
CLKBUF_X2 inst_11874 ( .A(net_11792), .Z(net_11793) );
AOI22_X2 inst_8991 ( .A2(net_9583), .ZN(net_8744), .B2(net_8743), .A1(net_2601), .B1(net_1977) );
INV_X4 inst_5874 ( .ZN(net_1387), .A(net_631) );
CLKBUF_X2 inst_13832 ( .A(net_10870), .Z(net_13751) );
CLKBUF_X2 inst_14068 ( .A(net_13950), .Z(net_13987) );
NAND4_X2 inst_3126 ( .ZN(net_3316), .A1(net_2290), .A4(net_2286), .A2(net_1414), .A3(net_1097) );
INV_X2 inst_7094 ( .A(net_1193), .ZN(net_1089) );
CLKBUF_X2 inst_12547 ( .A(net_12465), .Z(net_12466) );
CLKBUF_X2 inst_11319 ( .A(net_11237), .Z(net_11238) );
SDFF_X2 inst_503 ( .SE(net_9540), .SI(net_8198), .Q(net_312), .D(net_312), .CK(net_11645) );
DFF_X2 inst_8028 ( .QN(net_10222), .D(net_5460), .CK(net_14452) );
CLKBUF_X2 inst_12107 ( .A(net_12025), .Z(net_12026) );
DFF_X1 inst_8770 ( .D(net_4973), .CK(net_11076), .Q(x1066) );
DFF_X1 inst_8556 ( .Q(net_9983), .D(net_7365), .CK(net_14773) );
CLKBUF_X2 inst_14445 ( .A(net_14363), .Z(net_14364) );
DFF_X1 inst_8724 ( .Q(net_9140), .D(net_6449), .CK(net_11009) );
DFF_X2 inst_8300 ( .QN(net_9514), .D(net_4542), .CK(net_12725) );
INV_X4 inst_5340 ( .A(net_5420), .ZN(net_1722) );
CLKBUF_X2 inst_13235 ( .A(net_13153), .Z(net_13154) );
AND2_X2 inst_10580 ( .A1(net_3115), .ZN(net_2667), .A2(net_2666) );
NAND3_X2 inst_3193 ( .A3(net_7575), .ZN(net_7574), .A1(net_7573), .A2(net_7420) );
OAI21_X2 inst_1936 ( .B2(net_5362), .A(net_4628), .ZN(net_4466), .B1(net_4360) );
INV_X4 inst_6458 ( .A(net_10050), .ZN(net_4749) );
INV_X4 inst_5088 ( .A(net_1919), .ZN(net_1776) );
OAI211_X2 inst_2099 ( .C2(net_6778), .ZN(net_6749), .A(net_6407), .B(net_6108), .C1(net_541) );
NAND2_X2 inst_4193 ( .ZN(net_2920), .A1(net_1847), .A2(net_1846) );
NAND2_X2 inst_4069 ( .ZN(net_2798), .A2(net_2668), .A1(net_2173) );
CLKBUF_X2 inst_13316 ( .A(net_13234), .Z(net_13235) );
INV_X2 inst_7074 ( .A(net_2624), .ZN(net_1226) );
CLKBUF_X2 inst_14200 ( .A(net_13383), .Z(net_14119) );
CLKBUF_X2 inst_12858 ( .A(net_12776), .Z(net_12777) );
OR4_X2 inst_686 ( .ZN(net_7883), .A2(net_7768), .A4(net_7149), .A1(net_5349), .A3(net_3694) );
OAI22_X2 inst_1097 ( .A1(net_9189), .A2(net_6299), .B2(net_6298), .ZN(net_6296), .B1(net_2785) );
INV_X4 inst_5433 ( .ZN(net_3192), .A(net_1121) );
AOI221_X2 inst_9871 ( .B1(net_9779), .B2(net_9097), .A(net_6940), .C2(net_6939), .ZN(net_6831), .C1(net_249) );
CLKBUF_X2 inst_14777 ( .A(net_13247), .Z(net_14696) );
CLKBUF_X2 inst_11079 ( .A(net_10745), .Z(net_10998) );
CLKBUF_X2 inst_15268 ( .A(net_15186), .Z(net_15187) );
INV_X4 inst_4892 ( .ZN(net_5226), .A(net_2572) );
NOR2_X2 inst_2888 ( .ZN(net_2530), .A2(net_1783), .A1(net_1345) );
AOI22_X2 inst_9382 ( .B1(net_9995), .A2(net_5743), .B2(net_5742), .ZN(net_5523), .A1(net_235) );
INV_X2 inst_6804 ( .ZN(net_5186), .A(net_5185) );
CLKBUF_X2 inst_12683 ( .A(net_11777), .Z(net_12602) );
CLKBUF_X2 inst_12633 ( .A(net_12551), .Z(net_12552) );
NAND2_X2 inst_3643 ( .A2(net_6905), .ZN(net_6901), .A1(net_6243) );
CLKBUF_X2 inst_12330 ( .A(net_12248), .Z(net_12249) );
AOI22_X2 inst_9235 ( .A1(net_9899), .B1(net_9800), .B2(net_6129), .A2(net_6109), .ZN(net_6076) );
OAI33_X1 inst_967 ( .B2(net_10254), .ZN(net_3213), .B1(net_3212), .A3(net_3212), .A1(net_1475), .A2(net_1063), .B3(net_1062) );
CLKBUF_X2 inst_13117 ( .A(net_12339), .Z(net_13036) );
CLKBUF_X2 inst_10635 ( .A(net_10553), .Z(net_10554) );
AOI22_X2 inst_9075 ( .B1(net_9665), .A1(net_6808), .A2(net_6684), .B2(net_6683), .ZN(net_6591) );
OAI211_X2 inst_2119 ( .C2(net_6778), .ZN(net_6729), .A(net_6356), .B(net_6144), .C1(net_374) );
OAI21_X2 inst_1929 ( .B1(net_7785), .ZN(net_4438), .A(net_4142), .B2(net_4141) );
CLKBUF_X2 inst_12665 ( .A(net_10834), .Z(net_12584) );
NAND2_X2 inst_3391 ( .A1(net_9371), .ZN(net_8896), .A2(net_8736) );
AOI22_X2 inst_9422 ( .A1(net_10186), .A2(net_4656), .B2(net_4655), .ZN(net_4647), .B1(x4781) );
DFF_X1 inst_8519 ( .QN(net_10406), .D(net_7412), .CK(net_11090) );
CLKBUF_X2 inst_11495 ( .A(net_11413), .Z(net_11414) );
DFF_X2 inst_7863 ( .Q(net_9995), .D(net_6461), .CK(net_13398) );
CLKBUF_X2 inst_12200 ( .A(net_11695), .Z(net_12119) );
AOI22_X2 inst_9025 ( .A1(net_8002), .B2(net_8001), .ZN(net_7978), .A2(net_7921), .B1(net_3034) );
CLKBUF_X2 inst_12472 ( .A(net_12390), .Z(net_12391) );
OAI21_X2 inst_1794 ( .ZN(net_7571), .B2(net_7472), .A(net_7284), .B1(net_7252) );
CLKBUF_X2 inst_12029 ( .A(net_10989), .Z(net_11948) );
OAI22_X2 inst_1227 ( .B1(net_7229), .ZN(net_4892), .A2(net_4890), .B2(net_4889), .A1(net_535) );
NOR4_X2 inst_2324 ( .ZN(net_6159), .A3(net_6158), .A1(net_5886), .A4(net_5332), .A2(net_2890) );
CLKBUF_X2 inst_15023 ( .A(net_14941), .Z(net_14942) );
AOI22_X2 inst_9443 ( .A1(net_10522), .B1(net_9795), .ZN(net_4058), .A2(net_4056), .B2(net_2556) );
INV_X4 inst_5856 ( .A(net_7481), .ZN(net_5792) );
INV_X4 inst_5732 ( .ZN(net_3448), .A(net_752) );
DFF_X2 inst_8126 ( .Q(net_9825), .D(net_5136), .CK(net_13389) );
NAND4_X2 inst_3047 ( .ZN(net_7409), .A1(net_7070), .A4(net_7069), .A2(net_6259), .A3(net_2749) );
INV_X4 inst_5957 ( .A(net_7031), .ZN(net_553) );
NAND2_X2 inst_3847 ( .ZN(net_4365), .A1(net_4237), .A2(net_4236) );
NOR2_X2 inst_2897 ( .A1(net_9059), .A2(net_8954), .ZN(net_7987) );
CLKBUF_X2 inst_15086 ( .A(net_15004), .Z(net_15005) );
CLKBUF_X2 inst_15687 ( .A(net_15605), .Z(net_15606) );
NOR2_X2 inst_2529 ( .ZN(net_8137), .A1(net_8136), .A2(net_8135) );
CLKBUF_X2 inst_11807 ( .A(net_11725), .Z(net_11726) );
OAI21_X2 inst_1787 ( .B2(net_7664), .ZN(net_7540), .A(net_7430), .B1(net_5239) );
CLKBUF_X2 inst_14494 ( .A(net_13262), .Z(net_14413) );
INV_X4 inst_5756 ( .A(net_3528), .ZN(net_731) );
CLKBUF_X2 inst_12581 ( .A(net_12499), .Z(net_12500) );
INV_X2 inst_7274 ( .A(net_8947), .ZN(net_8946) );
CLKBUF_X2 inst_11376 ( .A(net_11294), .Z(net_11295) );
CLKBUF_X2 inst_14290 ( .A(net_13033), .Z(net_14209) );
AOI221_X2 inst_9741 ( .B2(net_9584), .C1(net_9582), .ZN(net_8770), .C2(net_8769), .A(net_8748), .B1(net_1396) );
CLKBUF_X2 inst_14369 ( .A(net_10904), .Z(net_14288) );
INV_X4 inst_5943 ( .A(net_911), .ZN(net_907) );
AOI221_X2 inst_9891 ( .B1(net_9877), .B2(net_9101), .A(net_6945), .C2(net_6944), .ZN(net_6803), .C1(net_248) );
OAI221_X2 inst_1540 ( .B2(net_9047), .C2(net_7287), .ZN(net_7225), .C1(net_7224), .A(net_6793), .B1(net_1512) );
INV_X4 inst_6310 ( .ZN(net_3332), .A(net_202) );
AOI22_X2 inst_9493 ( .B1(net_9918), .A1(net_9720), .B2(net_4969), .ZN(net_3830), .A2(net_3039) );
AOI221_X2 inst_9748 ( .C1(net_9365), .C2(net_8783), .ZN(net_7917), .A(net_7916), .B2(net_7915), .B1(net_7634) );
NAND2_X2 inst_3536 ( .A2(net_9059), .ZN(net_8870), .A1(net_8047) );
NOR2_X2 inst_2742 ( .A2(net_9289), .ZN(net_4147), .A1(net_3685) );
OAI221_X2 inst_1660 ( .C1(net_7226), .C2(net_5520), .ZN(net_5510), .B2(net_4547), .A(net_3507), .B1(net_598) );
AOI21_X2 inst_10113 ( .A(net_8868), .ZN(net_4578), .B2(net_4396), .B1(net_4265) );
DFF_X2 inst_7515 ( .QN(net_9244), .D(net_7898), .CK(net_11282) );
NAND2_X2 inst_4375 ( .ZN(net_1425), .A2(net_1401), .A1(net_197) );
INV_X4 inst_5243 ( .ZN(net_1749), .A(net_797) );
CLKBUF_X2 inst_13416 ( .A(net_13334), .Z(net_13335) );
CLKBUF_X2 inst_12355 ( .A(net_11721), .Z(net_12274) );
SDFF_X2 inst_517 ( .Q(net_9332), .D(net_9332), .SI(net_9157), .SE(net_7588), .CK(net_13082) );
NOR4_X2 inst_2346 ( .A3(net_9726), .A4(net_6305), .ZN(net_2750), .A1(net_2749), .A2(net_1829) );
OAI22_X2 inst_1261 ( .B1(net_7229), .A2(net_4842), .B2(net_4841), .ZN(net_4812), .A1(net_446) );
INV_X4 inst_5368 ( .ZN(net_2295), .A(net_1215) );
CLKBUF_X2 inst_12486 ( .A(net_12404), .Z(net_12405) );
CLKBUF_X2 inst_12123 ( .A(net_12041), .Z(net_12042) );
AOI21_X2 inst_10220 ( .ZN(net_2140), .B1(net_2139), .A(net_1786), .B2(net_959) );
INV_X4 inst_6130 ( .A(net_10468), .ZN(net_879) );
INV_X4 inst_5382 ( .ZN(net_1194), .A(net_1193) );
CLKBUF_X2 inst_14661 ( .A(net_14579), .Z(net_14580) );
CLKBUF_X2 inst_15629 ( .A(net_15547), .Z(net_15548) );
CLKBUF_X2 inst_13653 ( .A(net_13571), .Z(net_13572) );
XNOR2_X2 inst_310 ( .ZN(net_3226), .B(net_2804), .A(net_2667) );
CLKBUF_X2 inst_15680 ( .A(net_14088), .Z(net_15599) );
CLKBUF_X2 inst_12291 ( .A(net_12209), .Z(net_12210) );
INV_X2 inst_7250 ( .A(net_9415), .ZN(net_8218) );
CLKBUF_X2 inst_15279 ( .A(net_15197), .Z(net_15198) );
AOI221_X2 inst_9746 ( .B2(net_7932), .ZN(net_7931), .C2(net_7930), .A(net_7803), .C1(net_2609), .B1(net_988) );
HA_X1 inst_7363 ( .A(net_9228), .S(net_1456), .CO(net_1455), .B(net_527) );
CLKBUF_X2 inst_15135 ( .A(net_15053), .Z(net_15054) );
INV_X2 inst_7171 ( .A(net_9213), .ZN(net_546) );
OAI22_X2 inst_1005 ( .A2(net_8931), .ZN(net_8328), .A1(net_8327), .B1(net_8326), .B2(net_8325) );
INV_X2 inst_6979 ( .ZN(net_3137), .A(net_2919) );
CLKBUF_X2 inst_14895 ( .A(net_14813), .Z(net_14814) );
OAI221_X2 inst_1580 ( .B1(net_10315), .B2(net_9047), .C2(net_7287), .ZN(net_7128), .C1(net_7127), .A(net_6918) );
NOR2_X2 inst_2688 ( .ZN(net_4546), .A2(net_4545), .A1(net_2398) );
OAI21_X2 inst_1842 ( .ZN(net_6198), .B1(net_5963), .A(net_5929), .B2(net_3162) );
INV_X4 inst_6172 ( .A(net_9517), .ZN(net_1704) );
INV_X4 inst_5592 ( .A(net_1250), .ZN(net_1135) );
NOR4_X2 inst_2351 ( .A4(net_3708), .ZN(net_3320), .A1(net_2624), .A3(net_2623), .A2(net_795) );
DFF_X2 inst_8067 ( .QN(net_10353), .D(net_5324), .CK(net_13623) );
CLKBUF_X2 inst_12302 ( .A(net_12220), .Z(net_12221) );
INV_X4 inst_5125 ( .ZN(net_1826), .A(net_1600) );
OAI21_X2 inst_1853 ( .ZN(net_5876), .B2(net_5875), .A(net_5289), .B1(net_452) );
DFF_X2 inst_7534 ( .QN(net_9315), .D(net_7776), .CK(net_15323) );
DFF_X2 inst_7576 ( .QN(net_10266), .D(net_7540), .CK(net_11679) );
CLKBUF_X2 inst_11101 ( .A(net_11019), .Z(net_11020) );
XNOR2_X2 inst_264 ( .B(net_9216), .ZN(net_3974), .A(net_3655) );
NAND2_X2 inst_3703 ( .A1(net_10066), .ZN(net_5926), .A2(net_5898) );
INV_X2 inst_6737 ( .A(net_8002), .ZN(net_7924) );
OAI222_X2 inst_1333 ( .ZN(net_7733), .A1(net_7732), .B2(net_7731), .C2(net_7730), .A2(net_7565), .B1(net_5645), .C1(net_1279) );
NAND2_X2 inst_3710 ( .A1(net_5915), .ZN(net_5913), .A2(net_5912) );
CLKBUF_X2 inst_12613 ( .A(net_12531), .Z(net_12532) );
NAND2_X2 inst_3953 ( .A1(net_10473), .ZN(net_3709), .A2(net_3417) );
INV_X2 inst_7315 ( .A(net_9096), .ZN(net_9095) );
CLKBUF_X2 inst_14505 ( .A(net_14423), .Z(net_14424) );
OAI221_X2 inst_1551 ( .C2(net_7295), .B2(net_7293), .B1(net_7224), .ZN(net_7207), .A(net_6819), .C1(net_2232) );
OAI22_X2 inst_1260 ( .B1(net_7182), .A2(net_4842), .B2(net_4841), .ZN(net_4813), .A1(net_352) );
AOI22_X2 inst_9579 ( .B1(net_9978), .A2(net_5173), .ZN(net_3584), .B2(net_2541), .A1(net_212) );
OAI22_X2 inst_1088 ( .A2(net_7721), .ZN(net_6565), .A1(net_6564), .B2(net_6563), .B1(net_865) );
INV_X4 inst_6490 ( .A(net_10044), .ZN(net_5873) );
CLKBUF_X2 inst_13200 ( .A(net_13118), .Z(net_13119) );
AOI21_X2 inst_10190 ( .ZN(net_3278), .A(net_2838), .B1(net_2626), .B2(net_2121) );
CLKBUF_X2 inst_15238 ( .A(net_12426), .Z(net_15157) );
DFF_X1 inst_8692 ( .D(net_6700), .Q(net_192), .CK(net_14337) );
CLKBUF_X2 inst_15498 ( .A(net_15416), .Z(net_15417) );
CLKBUF_X2 inst_11672 ( .A(net_11590), .Z(net_11591) );
NAND2_X4 inst_3332 ( .A2(net_9033), .A1(net_9032), .ZN(net_8605) );
DFF_X2 inst_7885 ( .QN(net_10108), .D(net_6032), .CK(net_14805) );
CLKBUF_X2 inst_13165 ( .A(net_13083), .Z(net_13084) );
INV_X4 inst_4898 ( .A(net_7644), .ZN(net_7618) );
NOR2_X2 inst_2717 ( .A2(net_10270), .A1(net_6044), .ZN(net_5217) );
INV_X4 inst_5844 ( .A(net_3332), .ZN(net_651) );
CLKBUF_X2 inst_13142 ( .A(net_13060), .Z(net_13061) );
DFF_X1 inst_8781 ( .Q(net_10343), .D(net_4609), .CK(net_10674) );
INV_X4 inst_6433 ( .A(net_10100), .ZN(net_5833) );
CLKBUF_X2 inst_13836 ( .A(net_12627), .Z(net_13755) );
NAND2_X2 inst_4176 ( .ZN(net_2666), .A2(net_1366), .A1(net_1127) );
XNOR2_X2 inst_129 ( .ZN(net_7473), .A(net_7292), .B(net_2341) );
NOR2_X2 inst_2740 ( .A2(net_10539), .ZN(net_4323), .A1(net_3872) );
OAI21_X2 inst_1754 ( .A(net_8851), .ZN(net_8582), .B2(net_8569), .B1(net_8263) );
CLKBUF_X2 inst_12941 ( .A(net_12859), .Z(net_12860) );
AOI221_X2 inst_9922 ( .B2(net_5867), .ZN(net_5863), .A(net_5862), .C1(net_5861), .C2(net_4725), .B1(x5427) );
INV_X2 inst_6974 ( .ZN(net_1690), .A(net_1689) );
CLKBUF_X2 inst_12955 ( .A(net_11300), .Z(net_12874) );
NOR2_X2 inst_2931 ( .ZN(net_2045), .A2(net_1354), .A1(net_655) );
CLKBUF_X2 inst_14483 ( .A(net_14401), .Z(net_14402) );
INV_X4 inst_4768 ( .A(net_4311), .ZN(net_4297) );
DFF_X2 inst_7789 ( .Q(net_9823), .D(net_6506), .CK(net_14228) );
NOR2_X2 inst_2727 ( .ZN(net_4411), .A2(net_3961), .A1(net_2657) );
NOR2_X2 inst_2530 ( .A2(net_9589), .A1(net_9096), .ZN(net_9057) );
DFF_X2 inst_7974 ( .QN(net_10308), .D(net_5577), .CK(net_13236) );
OAI221_X2 inst_1503 ( .B2(net_9063), .C2(net_9056), .ZN(net_7358), .B1(net_7213), .A(net_6993), .C1(net_5881) );
CLKBUF_X2 inst_12234 ( .A(net_12152), .Z(net_12153) );
DFF_X1 inst_8848 ( .D(net_1159), .QN(net_314), .CK(net_12755) );
INV_X4 inst_5656 ( .ZN(net_5420), .A(net_826) );
INV_X4 inst_6305 ( .A(net_9553), .ZN(net_8175) );
DFF_X2 inst_7874 ( .QN(net_10154), .D(net_6008), .CK(net_13484) );
OR2_X4 inst_777 ( .ZN(net_3143), .A2(net_2971), .A1(net_2963) );
DFF_X2 inst_8317 ( .QN(net_10376), .D(net_3948), .CK(net_12113) );
NAND2_X2 inst_3802 ( .A1(net_5374), .ZN(net_4939), .A2(net_4665) );
INV_X4 inst_6164 ( .A(net_10150), .ZN(net_1204) );
CLKBUF_X2 inst_14175 ( .A(net_12242), .Z(net_14094) );
CLKBUF_X2 inst_12926 ( .A(net_10942), .Z(net_12845) );
INV_X4 inst_5016 ( .ZN(net_3908), .A(net_2111) );
AOI211_X2 inst_10276 ( .ZN(net_7515), .C2(net_7514), .A(net_7168), .C1(net_4192), .B(net_3740) );
CLKBUF_X2 inst_11094 ( .A(net_11012), .Z(net_11013) );
CLKBUF_X2 inst_10718 ( .A(net_10636), .Z(net_10637) );
OR2_X2 inst_933 ( .ZN(net_2665), .A1(net_2664), .A2(net_2663) );
INV_X2 inst_7000 ( .A(net_2401), .ZN(net_2322) );
AOI221_X2 inst_9983 ( .C1(net_10180), .B1(net_9753), .B2(net_6442), .C2(net_4217), .ZN(net_4214), .A(net_3569) );
NAND2_X2 inst_3724 ( .A1(net_10399), .ZN(net_5778), .A2(net_5777) );
CLKBUF_X2 inst_14393 ( .A(net_12604), .Z(net_14312) );
CLKBUF_X2 inst_14138 ( .A(net_13647), .Z(net_14057) );
CLKBUF_X2 inst_13902 ( .A(net_13820), .Z(net_13821) );
CLKBUF_X2 inst_14362 ( .A(net_14280), .Z(net_14281) );
AND2_X2 inst_10509 ( .A2(net_10483), .ZN(net_5806), .A1(net_869) );
OAI22_X2 inst_1013 ( .A2(net_8247), .B2(net_8246), .ZN(net_8236), .A1(net_2866), .B1(net_1176) );
INV_X4 inst_6146 ( .ZN(net_6811), .A(net_261) );
CLKBUF_X2 inst_13978 ( .A(net_13896), .Z(net_13897) );
CLKBUF_X2 inst_11909 ( .A(net_11827), .Z(net_11828) );
NAND2_X2 inst_3613 ( .ZN(net_7233), .A1(net_6870), .A2(net_6641) );
INV_X4 inst_4965 ( .ZN(net_2486), .A(net_2135) );
CLKBUF_X2 inst_13039 ( .A(net_12957), .Z(net_12958) );
AOI22_X2 inst_9439 ( .A2(net_10059), .B1(net_9924), .B2(net_6443), .A1(net_5320), .ZN(net_4279) );
CLKBUF_X2 inst_11158 ( .A(net_11065), .Z(net_11077) );
NOR4_X2 inst_2354 ( .A3(net_9218), .A4(net_9210), .A2(net_2497), .ZN(net_1699), .A1(net_1698) );
AOI22_X2 inst_9447 ( .A1(net_10527), .B1(net_9966), .A2(net_4056), .ZN(net_4052), .B2(net_2541) );
DFF_X1 inst_8735 ( .QN(net_9502), .D(net_6563), .CK(net_12538) );
DFF_X2 inst_7790 ( .Q(net_9824), .D(net_6459), .CK(net_15544) );
CLKBUF_X2 inst_14054 ( .A(net_13258), .Z(net_13973) );
CLKBUF_X2 inst_12870 ( .A(net_12788), .Z(net_12789) );
DFF_X1 inst_8481 ( .QN(net_9630), .D(net_7949), .CK(net_15023) );
CLKBUF_X2 inst_10729 ( .A(net_10611), .Z(net_10648) );
NAND2_X2 inst_3515 ( .ZN(net_8120), .A1(net_8119), .A2(net_8118) );
XNOR2_X2 inst_124 ( .ZN(net_7550), .A(net_7324), .B(net_7025) );
CLKBUF_X2 inst_13315 ( .A(net_13233), .Z(net_13234) );
CLKBUF_X2 inst_15514 ( .A(net_15432), .Z(net_15433) );
CLKBUF_X2 inst_14965 ( .A(net_14883), .Z(net_14884) );
CLKBUF_X2 inst_12316 ( .A(net_12234), .Z(net_12235) );
CLKBUF_X2 inst_10883 ( .A(net_10787), .Z(net_10802) );
CLKBUF_X2 inst_10982 ( .A(net_10900), .Z(net_10901) );
NAND2_X2 inst_3869 ( .ZN(net_4625), .A2(net_4226), .A1(net_4080) );
NAND2_X2 inst_3488 ( .A2(net_8970), .ZN(net_8443), .A1(net_5389) );
CLKBUF_X2 inst_13849 ( .A(net_13767), .Z(net_13768) );
CLKBUF_X2 inst_12531 ( .A(net_12449), .Z(net_12450) );
CLKBUF_X2 inst_11593 ( .A(net_10593), .Z(net_11512) );
OAI22_X2 inst_1270 ( .ZN(net_4756), .A1(net_4755), .A2(net_4752), .B2(net_4751), .B1(net_1264) );
INV_X4 inst_6332 ( .ZN(net_414), .A(x637) );
NAND2_X2 inst_3448 ( .A1(net_9486), .ZN(net_9028), .A2(net_8476) );
DFF_X2 inst_8001 ( .QN(net_10122), .D(net_5508), .CK(net_12357) );
INV_X4 inst_6088 ( .ZN(net_4188), .A(net_159) );
CLKBUF_X2 inst_15801 ( .A(net_15719), .Z(net_15720) );
CLKBUF_X2 inst_12689 ( .A(net_12607), .Z(net_12608) );
INV_X4 inst_4563 ( .ZN(net_8391), .A(net_8252) );
AOI21_X2 inst_10123 ( .ZN(net_4465), .A(net_4464), .B2(net_4012), .B1(net_3891) );
CLKBUF_X2 inst_13032 ( .A(net_12950), .Z(net_12951) );
INV_X4 inst_5504 ( .ZN(net_3855), .A(net_981) );
CLKBUF_X2 inst_14561 ( .A(net_12089), .Z(net_14480) );
CLKBUF_X2 inst_15602 ( .A(net_11897), .Z(net_15521) );
INV_X4 inst_5361 ( .ZN(net_1958), .A(net_1221) );
CLKBUF_X2 inst_12489 ( .A(net_12407), .Z(net_12408) );
CLKBUF_X2 inst_13049 ( .A(net_12967), .Z(net_12968) );
DFF_X2 inst_7453 ( .QN(net_9644), .D(net_8159), .CK(net_13148) );
CLKBUF_X2 inst_15620 ( .A(net_15538), .Z(net_15539) );
OAI221_X2 inst_1519 ( .C1(net_10415), .B2(net_9063), .C2(net_9056), .ZN(net_7313), .B1(net_7108), .A(net_7076) );
INV_X2 inst_7243 ( .A(net_9314), .ZN(net_369) );
OAI211_X2 inst_2156 ( .C2(net_6778), .ZN(net_6692), .A(net_6313), .B(net_6051), .C1(net_5032) );
CLKBUF_X2 inst_13389 ( .A(net_13307), .Z(net_13308) );
AOI221_X2 inst_9936 ( .B2(net_5867), .A(net_5862), .ZN(net_5832), .C1(net_5831), .C2(net_4725), .B1(x5722) );
DFF_X1 inst_8461 ( .Q(net_9595), .D(net_7956), .CK(net_11542) );
INV_X4 inst_4989 ( .ZN(net_7423), .A(net_2226) );
CLKBUF_X2 inst_12142 ( .A(net_12060), .Z(net_12061) );
NAND2_X2 inst_4324 ( .ZN(net_1629), .A2(net_950), .A1(net_741) );
INV_X4 inst_5746 ( .ZN(net_742), .A(net_741) );
INV_X4 inst_5417 ( .ZN(net_1526), .A(net_614) );
INV_X4 inst_5597 ( .A(net_10261), .ZN(net_1169) );
INV_X2 inst_7009 ( .A(net_2392), .ZN(net_1606) );
CLKBUF_X2 inst_12705 ( .A(net_12623), .Z(net_12624) );
NOR2_X2 inst_2515 ( .A2(net_8319), .ZN(net_8269), .A1(net_8151) );
DFF_X1 inst_8531 ( .Q(net_9967), .D(net_7373), .CK(net_15645) );
CLKBUF_X2 inst_15798 ( .A(net_12137), .Z(net_15717) );
CLKBUF_X2 inst_12244 ( .A(net_12162), .Z(net_12163) );
OAI221_X2 inst_1491 ( .B1(net_10410), .C2(net_9063), .B2(net_9056), .ZN(net_7372), .C1(net_7245), .A(net_7010) );
DFF_X2 inst_8070 ( .QN(net_10365), .D(net_5306), .CK(net_13621) );
CLKBUF_X2 inst_12747 ( .A(net_12665), .Z(net_12666) );
DFF_X1 inst_8703 ( .Q(net_9146), .D(net_6783), .CK(net_11016) );
CLKBUF_X2 inst_15446 ( .A(net_13662), .Z(net_15365) );
CLKBUF_X2 inst_12900 ( .A(net_12818), .Z(net_12819) );
XNOR2_X2 inst_117 ( .B(net_9425), .ZN(net_7821), .A(net_6433) );
NOR2_X2 inst_2676 ( .ZN(net_5290), .A2(net_4780), .A1(net_3298) );
INV_X4 inst_5172 ( .ZN(net_3037), .A(net_1560) );
DFF_X1 inst_8566 ( .Q(net_9871), .D(net_7177), .CK(net_14857) );
XNOR2_X2 inst_154 ( .ZN(net_6267), .A(net_5991), .B(net_2656) );
CLKBUF_X2 inst_13104 ( .A(net_13022), .Z(net_13023) );
CLKBUF_X2 inst_15195 ( .A(net_15113), .Z(net_15114) );
NAND2_X2 inst_4106 ( .A2(net_9107), .A1(net_3364), .ZN(net_2374) );
AOI221_X2 inst_9794 ( .B1(net_9959), .A(net_7090), .B2(net_7089), .C2(net_7088), .ZN(net_7010), .C1(net_6834) );
SDFF_X2 inst_465 ( .SE(net_8812), .SI(net_8649), .CK(net_11909), .Q(x732), .D(x732) );
INV_X4 inst_6057 ( .A(net_9519), .ZN(net_2818) );
CLKBUF_X2 inst_11367 ( .A(net_11285), .Z(net_11286) );
NOR4_X2 inst_2304 ( .A3(net_9043), .ZN(net_8050), .A1(net_7889), .A4(net_7821), .A2(net_7400) );
CLKBUF_X2 inst_12325 ( .A(net_12243), .Z(net_12244) );
AOI21_X2 inst_10078 ( .ZN(net_9064), .A(net_5888), .B2(net_5694), .B1(net_2758) );
CLKBUF_X2 inst_13427 ( .A(net_13345), .Z(net_13346) );
AND3_X2 inst_10368 ( .ZN(net_5227), .A2(net_5226), .A3(net_4948), .A1(net_4947) );
NAND2_X2 inst_4240 ( .A1(net_2236), .ZN(net_1481), .A2(net_1137) );
CLKBUF_X2 inst_11701 ( .A(net_11619), .Z(net_11620) );
CLKBUF_X2 inst_10813 ( .A(net_10731), .Z(net_10732) );
OAI211_X2 inst_2173 ( .C1(net_7229), .C2(net_6548), .ZN(net_6536), .B(net_5664), .A(net_3507) );
CLKBUF_X2 inst_12570 ( .A(net_12488), .Z(net_12489) );
OAI21_X2 inst_1790 ( .B2(net_8827), .ZN(net_7592), .B1(net_6951), .A(net_3541) );
INV_X4 inst_6621 ( .ZN(net_8953), .A(net_8942) );
INV_X2 inst_7048 ( .A(net_2397), .ZN(net_1336) );
CLKBUF_X2 inst_15039 ( .A(net_13563), .Z(net_14958) );
NAND3_X2 inst_3214 ( .ZN(net_5787), .A3(net_5231), .A1(net_5230), .A2(net_5229) );
CLKBUF_X2 inst_10989 ( .A(net_10646), .Z(net_10908) );
CLKBUF_X2 inst_12940 ( .A(net_12858), .Z(net_12859) );
OAI21_X2 inst_1905 ( .B1(net_7219), .B2(net_4862), .ZN(net_4847), .A(net_4519) );
INV_X4 inst_6355 ( .A(net_9374), .ZN(net_405) );
CLKBUF_X2 inst_11917 ( .A(net_11700), .Z(net_11836) );
CLKBUF_X2 inst_13982 ( .A(net_13900), .Z(net_13901) );
OAI211_X2 inst_2264 ( .C1(net_7127), .C2(net_6542), .ZN(net_6281), .B(net_5708), .A(net_3507) );
CLKBUF_X2 inst_14925 ( .A(net_14843), .Z(net_14844) );
XNOR2_X2 inst_243 ( .ZN(net_4163), .A(net_3656), .B(net_2496) );
OAI222_X2 inst_1378 ( .B2(net_7660), .A2(net_7659), .C2(net_7658), .ZN(net_6007), .B1(net_2980), .A1(net_2011), .C1(net_1317) );
CLKBUF_X2 inst_14156 ( .A(net_14074), .Z(net_14075) );
CLKBUF_X2 inst_14049 ( .A(net_12196), .Z(net_13968) );
NOR2_X2 inst_2697 ( .ZN(net_4842), .A1(net_4391), .A2(net_4075) );
AOI21_X2 inst_10196 ( .ZN(net_3036), .A(net_3035), .B1(net_3034), .B2(net_2546) );
XOR2_X2 inst_15 ( .Z(net_2800), .A(net_2225), .B(net_1484) );
NAND2_X2 inst_3747 ( .ZN(net_5303), .A2(net_5286), .A1(net_4472) );
CLKBUF_X2 inst_15738 ( .A(net_15656), .Z(net_15657) );
DFF_X2 inst_8189 ( .QN(net_10534), .D(net_5156), .CK(net_14876) );
CLKBUF_X2 inst_11902 ( .A(net_11820), .Z(net_11821) );
INV_X2 inst_7281 ( .A(net_8970), .ZN(net_8969) );
NAND2_X2 inst_3496 ( .A1(net_9554), .ZN(net_8329), .A2(net_8250) );
INV_X2 inst_6704 ( .A(net_8186), .ZN(net_8149) );
AOI22_X2 inst_9501 ( .B1(net_9821), .A1(net_9690), .A2(net_5966), .ZN(net_3822), .B2(net_2556) );
CLKBUF_X2 inst_13082 ( .A(net_13000), .Z(net_13001) );
AOI221_X2 inst_9830 ( .ZN(net_6891), .A(net_6889), .B2(net_6888), .C2(net_6887), .B1(net_5866), .C1(x6102) );
CLKBUF_X2 inst_13642 ( .A(net_13560), .Z(net_13561) );
CLKBUF_X2 inst_12020 ( .A(net_10710), .Z(net_11939) );
DFF_X1 inst_8799 ( .QN(net_10167), .D(net_4117), .CK(net_12295) );
OAI211_X2 inst_2123 ( .C2(net_6778), .ZN(net_6725), .A(net_6352), .B(net_6087), .C1(net_400) );
NAND3_X2 inst_3229 ( .A2(net_10515), .A3(net_8511), .A1(net_7832), .ZN(net_5732) );
INV_X4 inst_4918 ( .ZN(net_5174), .A(net_3588) );
DFF_X1 inst_8615 ( .Q(net_9662), .D(net_7271), .CK(net_15561) );
NAND2_X2 inst_4135 ( .ZN(net_2927), .A1(net_2321), .A2(net_2235) );
CLKBUF_X2 inst_14459 ( .A(net_14377), .Z(net_14378) );
OAI222_X2 inst_1369 ( .B2(net_7660), .A2(net_7659), .C2(net_7658), .ZN(net_6275), .B1(net_4935), .A1(net_3424), .C1(net_1076) );
CLKBUF_X2 inst_14668 ( .A(net_13197), .Z(net_14587) );
NAND2_X2 inst_3988 ( .A1(net_9791), .ZN(net_3186), .A2(net_2462) );
XNOR2_X2 inst_349 ( .A(net_9085), .B(net_3976), .ZN(net_2817) );
CLKBUF_X2 inst_14145 ( .A(net_14063), .Z(net_14064) );
CLKBUF_X2 inst_10690 ( .A(net_10569), .Z(net_10609) );
INV_X4 inst_6548 ( .A(net_10020), .ZN(net_333) );
CLKBUF_X2 inst_14381 ( .A(net_11659), .Z(net_14300) );
CLKBUF_X2 inst_15172 ( .A(net_13929), .Z(net_15091) );
NAND2_X2 inst_4249 ( .ZN(net_2757), .A2(net_1004), .A1(net_723) );
CLKBUF_X2 inst_15280 ( .A(net_11137), .Z(net_15199) );
NAND2_X2 inst_4235 ( .A1(net_9109), .ZN(net_2218), .A2(net_1581) );
CLKBUF_X2 inst_13940 ( .A(net_13858), .Z(net_13859) );
NOR2_X2 inst_2561 ( .ZN(net_7745), .A2(net_7651), .A1(net_3535) );
DFF_X2 inst_7767 ( .Q(net_9717), .D(net_6537), .CK(net_12797) );
CLKBUF_X2 inst_13629 ( .A(net_10798), .Z(net_13548) );
CLKBUF_X2 inst_11507 ( .A(net_10966), .Z(net_11426) );
AOI22_X2 inst_9570 ( .B2(net_6442), .A2(net_5173), .ZN(net_3738), .B1(net_1265), .A1(net_572) );
INV_X4 inst_6024 ( .ZN(net_522), .A(net_203) );
DFF_X1 inst_8495 ( .Q(net_9955), .D(net_7820), .CK(net_14422) );
CLKBUF_X2 inst_14876 ( .A(net_14794), .Z(net_14795) );
DFF_X2 inst_8163 ( .QN(net_9931), .D(net_5056), .CK(net_14350) );
CLKBUF_X2 inst_13669 ( .A(net_10581), .Z(net_13588) );
CLKBUF_X2 inst_13257 ( .A(net_13175), .Z(net_13176) );
AOI22_X2 inst_9583 ( .B1(net_9982), .A2(net_5173), .ZN(net_3579), .B2(net_2541), .A1(net_216) );
CLKBUF_X2 inst_15725 ( .A(net_11072), .Z(net_15644) );
NAND2_X2 inst_4226 ( .A1(net_8687), .ZN(net_1654), .A2(net_113) );
OAI211_X2 inst_2252 ( .C1(net_7294), .A(net_6546), .C2(net_6480), .ZN(net_6439), .B(net_5744) );
CLKBUF_X2 inst_12289 ( .A(net_12207), .Z(net_12208) );
CLKBUF_X2 inst_12514 ( .A(net_11474), .Z(net_12433) );
AOI22_X2 inst_9222 ( .A1(net_9916), .B1(net_9817), .B2(net_6120), .A2(net_6111), .ZN(net_6089) );
NAND2_X2 inst_4229 ( .ZN(net_3134), .A1(net_2627), .A2(net_986) );
CLKBUF_X2 inst_12843 ( .A(net_12761), .Z(net_12762) );
INV_X4 inst_5795 ( .A(net_1016), .ZN(net_919) );
CLKBUF_X2 inst_12112 ( .A(net_11267), .Z(net_12031) );
CLKBUF_X2 inst_12065 ( .A(net_11983), .Z(net_11984) );
OAI211_X2 inst_2238 ( .C1(net_7297), .C2(net_6501), .ZN(net_6466), .B(net_5761), .A(net_3679) );
NOR2_X2 inst_2763 ( .A2(net_4070), .ZN(net_3890), .A1(net_835) );
INV_X4 inst_5207 ( .ZN(net_4573), .A(net_1526) );
INV_X4 inst_4543 ( .ZN(net_8883), .A(net_8662) );
INV_X4 inst_5072 ( .ZN(net_2200), .A(net_1848) );
CLKBUF_X2 inst_14334 ( .A(net_11166), .Z(net_14253) );
AOI211_X2 inst_10301 ( .B(net_6060), .ZN(net_3539), .A(net_3538), .C2(net_3094), .C1(net_2059) );
CLKBUF_X2 inst_14347 ( .A(net_13517), .Z(net_14266) );
NAND4_X2 inst_3151 ( .ZN(net_3196), .A3(net_2103), .A1(net_2094), .A4(net_2093), .A2(net_1017) );
AND2_X2 inst_10554 ( .ZN(net_3657), .A2(net_3312), .A1(net_363) );
INV_X2 inst_6798 ( .ZN(net_5960), .A(net_5244) );
CLKBUF_X2 inst_15312 ( .A(net_15230), .Z(net_15231) );
OR2_X4 inst_761 ( .A1(net_6165), .ZN(net_5139), .A2(net_4364) );
CLKBUF_X2 inst_13073 ( .A(net_12991), .Z(net_12992) );
CLKBUF_X2 inst_10764 ( .A(net_10682), .Z(net_10683) );
INV_X4 inst_4867 ( .A(net_4481), .ZN(net_3363) );
CLKBUF_X2 inst_13342 ( .A(net_13260), .Z(net_13261) );
MUX2_X1 inst_4436 ( .S(net_6041), .A(net_310), .B(x4041), .Z(x39) );
NOR2_X2 inst_2803 ( .ZN(net_3232), .A2(net_2802), .A1(net_2648) );
DFF_X2 inst_8180 ( .QN(net_10028), .D(net_5022), .CK(net_13691) );
CLKBUF_X2 inst_13042 ( .A(net_12960), .Z(net_12961) );
CLKBUF_X2 inst_14732 ( .A(net_14110), .Z(net_14651) );
NAND2_X2 inst_4120 ( .A1(net_4553), .ZN(net_2337), .A2(net_1610) );
INV_X4 inst_5801 ( .ZN(net_1956), .A(net_1347) );
AOI22_X2 inst_9363 ( .B1(net_9923), .A2(net_5759), .B2(net_5758), .ZN(net_5559), .A1(net_262) );
AOI22_X2 inst_9211 ( .A1(net_9902), .B1(net_9803), .A2(net_8042), .B2(net_6133), .ZN(net_6100) );
INV_X4 inst_5525 ( .A(net_10352), .ZN(net_2005) );
INV_X2 inst_6674 ( .ZN(net_8354), .A(net_8291) );
AOI21_X4 inst_10003 ( .ZN(net_9046), .B1(net_1502), .B2(net_187), .A(net_180) );
OAI211_X2 inst_2259 ( .C1(net_7211), .C2(net_6501), .ZN(net_6362), .B(net_5421), .A(net_3679) );
INV_X4 inst_5097 ( .ZN(net_1712), .A(net_1711) );
CLKBUF_X2 inst_12935 ( .A(net_12313), .Z(net_12854) );
NOR2_X2 inst_2641 ( .A1(net_9228), .ZN(net_5451), .A2(net_5449) );
INV_X4 inst_6196 ( .A(net_10043), .ZN(net_2284) );
CLKBUF_X2 inst_14314 ( .A(net_14232), .Z(net_14233) );
OAI221_X2 inst_1638 ( .B1(net_10410), .C1(net_7245), .ZN(net_5550), .B2(net_4477), .C2(net_4455), .A(net_3731) );
INV_X4 inst_6462 ( .ZN(net_6344), .A(net_164) );
CLKBUF_X2 inst_11450 ( .A(net_11368), .Z(net_11369) );
INV_X4 inst_5771 ( .A(net_749), .ZN(net_719) );
AOI221_X2 inst_9812 ( .B1(net_9990), .A(net_7090), .B2(net_7089), .C2(net_7088), .ZN(net_6990), .C1(net_262) );
NAND3_X2 inst_3220 ( .ZN(net_9100), .A2(net_5356), .A1(net_4906), .A3(net_4795) );
CLKBUF_X2 inst_14101 ( .A(net_14019), .Z(net_14020) );
CLKBUF_X2 inst_12824 ( .A(net_12742), .Z(net_12743) );
CLKBUF_X2 inst_11915 ( .A(net_11703), .Z(net_11834) );
DFF_X2 inst_8177 ( .QN(net_9735), .D(net_5031), .CK(net_12771) );
CLKBUF_X2 inst_12280 ( .A(net_10749), .Z(net_12199) );
CLKBUF_X2 inst_11072 ( .A(net_10975), .Z(net_10991) );
CLKBUF_X2 inst_11983 ( .A(net_11021), .Z(net_11902) );
INV_X4 inst_5354 ( .ZN(net_7435), .A(net_1230) );
INV_X4 inst_6428 ( .ZN(net_7186), .A(x5077) );
CLKBUF_X2 inst_14221 ( .A(net_14139), .Z(net_14140) );
INV_X2 inst_7312 ( .A(net_9091), .ZN(net_9090) );
INV_X4 inst_5373 ( .A(net_2007), .ZN(net_1206) );
DFF_X2 inst_7560 ( .QN(net_10150), .D(net_7607), .CK(net_12375) );
INV_X4 inst_4783 ( .A(net_6669), .ZN(net_3923) );
AOI22_X2 inst_9047 ( .B1(net_9669), .ZN(net_6685), .A1(net_6684), .B2(net_6683), .A2(net_238) );
NAND2_X2 inst_3862 ( .ZN(net_4113), .A2(net_3940), .A1(net_2334) );
INV_X4 inst_6556 ( .ZN(net_331), .A(net_206) );
INV_X4 inst_6532 ( .A(net_9315), .ZN(net_7681) );
CLKBUF_X2 inst_10749 ( .A(net_10667), .Z(net_10668) );
CLKBUF_X2 inst_10847 ( .A(net_10765), .Z(net_10766) );
INV_X4 inst_5304 ( .ZN(net_5457), .A(net_1297) );
CLKBUF_X2 inst_14326 ( .A(net_14244), .Z(net_14245) );
CLKBUF_X2 inst_12737 ( .A(net_12655), .Z(net_12656) );
AND2_X2 inst_10482 ( .A2(net_9577), .A1(net_9576), .ZN(net_8574) );
SDFF_X2 inst_633 ( .Q(net_9460), .D(net_9460), .SE(net_3293), .CK(net_12440), .SI(x1911) );
CLKBUF_X2 inst_12837 ( .A(net_12586), .Z(net_12756) );
SDFF_X2 inst_524 ( .Q(net_9341), .D(net_9341), .SI(net_9333), .SE(net_7588), .CK(net_14679) );
CLKBUF_X2 inst_15568 ( .A(net_15486), .Z(net_15487) );
CLKBUF_X2 inst_13027 ( .A(net_12945), .Z(net_12946) );
NAND2_X2 inst_4060 ( .ZN(net_4606), .A1(net_2761), .A2(net_2760) );
XNOR2_X2 inst_104 ( .ZN(net_8171), .A(net_8088), .B(net_6901) );
OAI211_X2 inst_2285 ( .C1(net_7108), .C2(net_6501), .ZN(net_6194), .B(net_5717), .A(net_3679) );
CLKBUF_X2 inst_14986 ( .A(net_14904), .Z(net_14905) );
AND2_X2 inst_10500 ( .A2(net_10450), .ZN(net_6043), .A1(net_1582) );
NOR4_X2 inst_2331 ( .ZN(net_5215), .A2(net_5214), .A4(net_5213), .A3(net_4575), .A1(net_3720) );
NAND2_X4 inst_3344 ( .ZN(net_8522), .A2(net_8484), .A1(net_8483) );
MUX2_X1 inst_4478 ( .S(net_6041), .A(net_3733), .B(x6531), .Z(x427) );
INV_X4 inst_6096 ( .ZN(net_3897), .A(net_160) );
CLKBUF_X2 inst_11878 ( .A(net_11545), .Z(net_11797) );
AOI221_X2 inst_9752 ( .B2(net_7932), .ZN(net_7896), .B1(net_7895), .A(net_7802), .C2(net_7526), .C1(net_4204) );
NAND2_X2 inst_3447 ( .A1(net_9494), .ZN(net_9029), .A2(net_8461) );
NOR3_X2 inst_2377 ( .ZN(net_8034), .A3(net_8033), .A2(net_4127), .A1(net_3984) );
NOR2_X2 inst_2522 ( .ZN(net_8253), .A1(net_8184), .A2(net_8183) );
CLKBUF_X2 inst_13793 ( .A(net_13711), .Z(net_13712) );
INV_X2 inst_7199 ( .A(net_9399), .ZN(net_8234) );
INV_X4 inst_4862 ( .ZN(net_4062), .A(net_3143) );
CLKBUF_X2 inst_15220 ( .A(net_15138), .Z(net_15139) );
CLKBUF_X2 inst_11910 ( .A(net_10814), .Z(net_11829) );
INV_X4 inst_4663 ( .ZN(net_5598), .A(net_5597) );
AND3_X4 inst_10360 ( .ZN(net_5755), .A2(net_4788), .A3(net_4625), .A1(net_4461) );
OR2_X2 inst_882 ( .A2(net_7038), .ZN(net_6294), .A1(net_6293) );
CLKBUF_X2 inst_10673 ( .A(net_10576), .Z(net_10592) );
CLKBUF_X2 inst_13935 ( .A(net_13853), .Z(net_13854) );
DFF_X2 inst_7967 ( .QN(net_10317), .D(net_5587), .CK(net_15487) );
AOI221_X2 inst_9848 ( .A(net_6889), .B2(net_6888), .C2(net_6887), .ZN(net_6870), .B1(net_5827), .C1(x5601) );
INV_X4 inst_5216 ( .A(net_2869), .ZN(net_1902) );
CLKBUF_X2 inst_13700 ( .A(net_13618), .Z(net_13619) );
NOR2_X2 inst_2938 ( .ZN(net_1809), .A1(net_1367), .A2(net_759) );
INV_X4 inst_5257 ( .A(net_6053), .ZN(net_1427) );
DFF_X2 inst_8011 ( .QN(net_10223), .D(net_5496), .CK(net_12204) );
AOI22_X2 inst_9116 ( .A1(net_9670), .A2(net_6404), .ZN(net_6373), .B2(net_5263), .B1(net_108) );
CLKBUF_X2 inst_15627 ( .A(net_15545), .Z(net_15546) );
CLKBUF_X2 inst_11226 ( .A(net_11144), .Z(net_11145) );
INV_X4 inst_5083 ( .ZN(net_1801), .A(net_1800) );
INV_X2 inst_6931 ( .ZN(net_3140), .A(net_2219) );
CLKBUF_X2 inst_15802 ( .A(net_15720), .Z(net_15721) );
OR3_X2 inst_708 ( .ZN(net_7817), .A1(net_7816), .A3(net_7815), .A2(net_7276) );
OAI222_X2 inst_1346 ( .A1(net_7660), .B2(net_7659), .C2(net_7658), .ZN(net_7554), .A2(net_7311), .B1(net_4604), .C1(net_1922) );
NAND2_X2 inst_3523 ( .ZN(net_8247), .A2(net_8108), .A1(net_8107) );
OAI222_X2 inst_1374 ( .B2(net_7660), .A2(net_7659), .C2(net_7658), .ZN(net_6031), .B1(net_3222), .A1(net_2124), .C1(net_1119) );
INV_X4 inst_4855 ( .ZN(net_7157), .A(net_3286) );
INV_X4 inst_5811 ( .ZN(net_2232), .A(net_1208) );
AOI22_X2 inst_9046 ( .B1(net_9668), .ZN(net_6686), .A1(net_6684), .B2(net_6683), .A2(net_237) );
NAND2_X2 inst_3510 ( .A1(net_9549), .ZN(net_8173), .A2(net_8145) );
NOR2_X2 inst_2510 ( .A2(net_8428), .ZN(net_8390), .A1(net_8389) );
INV_X4 inst_5108 ( .ZN(net_4080), .A(net_2964) );
INV_X2 inst_6723 ( .ZN(net_7779), .A(net_7746) );
OAI22_X2 inst_1071 ( .ZN(net_6855), .A1(net_6854), .A2(net_6848), .B2(net_6846), .B1(net_5405) );
NAND2_X2 inst_4277 ( .A1(net_4157), .ZN(net_2345), .A2(net_1244) );
INV_X4 inst_6421 ( .ZN(net_771), .A(net_188) );
INV_X4 inst_6316 ( .A(net_10357), .ZN(net_777) );
INV_X4 inst_5291 ( .A(net_6056), .ZN(net_1313) );
CLKBUF_X2 inst_11352 ( .A(net_11270), .Z(net_11271) );
CLKBUF_X2 inst_13211 ( .A(net_10673), .Z(net_13130) );
CLKBUF_X2 inst_11548 ( .A(net_11466), .Z(net_11467) );
CLKBUF_X2 inst_14199 ( .A(net_14117), .Z(net_14118) );
OAI21_X2 inst_1994 ( .ZN(net_3005), .B1(net_2502), .A(net_1839), .B2(net_1201) );
CLKBUF_X2 inst_15184 ( .A(net_15102), .Z(net_15103) );
CLKBUF_X2 inst_13132 ( .A(net_13050), .Z(net_13051) );
AOI22_X2 inst_9192 ( .A1(net_9882), .B1(net_9783), .A2(net_8042), .B2(net_6129), .ZN(net_6122) );
INV_X4 inst_5298 ( .ZN(net_1523), .A(net_1303) );
CLKBUF_X2 inst_14436 ( .A(net_14354), .Z(net_14355) );
AOI21_X2 inst_10108 ( .B2(net_10131), .ZN(net_4931), .B1(net_3272), .A(net_3026) );
CLKBUF_X2 inst_15179 ( .A(net_15097), .Z(net_15098) );
CLKBUF_X2 inst_14935 ( .A(net_14853), .Z(net_14854) );
CLKBUF_X2 inst_14744 ( .A(net_14662), .Z(net_14663) );
CLKBUF_X2 inst_13191 ( .A(net_11077), .Z(net_13110) );
OAI211_X2 inst_2162 ( .C1(net_7245), .ZN(net_6550), .C2(net_6548), .B(net_5675), .A(net_3679) );
XNOR2_X2 inst_392 ( .B(net_9231), .ZN(net_2156), .A(net_1441) );
XNOR2_X2 inst_120 ( .ZN(net_7622), .A(net_7493), .B(net_7045) );
CLKBUF_X2 inst_14533 ( .A(net_14451), .Z(net_14452) );
INV_X2 inst_6780 ( .ZN(net_6018), .A(net_5830) );
DFF_X2 inst_7747 ( .QN(net_10356), .D(net_6283), .CK(net_12212) );
CLKBUF_X2 inst_10917 ( .A(net_10835), .Z(net_10836) );
NAND2_X2 inst_4165 ( .ZN(net_2902), .A1(net_1972), .A2(net_1971) );
NAND2_X2 inst_4398 ( .A2(net_10123), .A1(net_10122), .ZN(net_1436) );
OAI221_X2 inst_1514 ( .B1(net_10416), .C2(net_9063), .B2(net_9056), .ZN(net_7335), .C1(net_7124), .A(net_7082) );
OAI211_X2 inst_2272 ( .C1(net_7129), .C2(net_6480), .ZN(net_6269), .B(net_5691), .A(net_3679) );
DFF_X2 inst_8361 ( .QN(net_8842), .D(net_2300), .CK(net_13679) );
SDFF_X2 inst_567 ( .D(net_9145), .SE(net_933), .CK(net_10990), .SI(x1660), .Q(x1134) );
OAI221_X2 inst_1608 ( .C1(net_10204), .B1(net_7241), .C2(net_5642), .ZN(net_5628), .B2(net_4905), .A(net_3731) );
NAND3_X2 inst_3200 ( .A3(net_9503), .A1(net_7424), .ZN(net_7421), .A2(net_7420) );
CLKBUF_X2 inst_11631 ( .A(net_11549), .Z(net_11550) );
AOI22_X2 inst_9134 ( .A1(net_9718), .A2(net_6420), .ZN(net_6354), .B2(net_5263), .B1(net_4190) );
OAI221_X2 inst_1484 ( .C2(net_7525), .ZN(net_7520), .B2(net_7519), .B1(net_7003), .A(net_5165), .C1(net_1310) );
OAI221_X2 inst_1601 ( .B1(net_10216), .C1(net_7186), .B2(net_5642), .ZN(net_5635), .C2(net_4905), .A(net_3731) );
NAND2_X2 inst_3526 ( .ZN(net_8237), .A1(net_8093), .A2(net_8092) );
AOI22_X2 inst_9010 ( .B1(net_9305), .A2(net_8030), .B2(net_8029), .ZN(net_8026), .A1(net_213) );
OR2_X2 inst_856 ( .ZN(net_8141), .A1(net_8093), .A2(net_8092) );
INV_X4 inst_5677 ( .ZN(net_1254), .A(net_193) );

endmodule
